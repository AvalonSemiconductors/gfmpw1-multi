magic
tech gf180mcuD
magscale 1 10
timestamp 1753968499
<< metal1 >>
rect 1344 46282 48608 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 48608 46282
rect 1344 46196 48608 46230
rect 19182 46114 19234 46126
rect 19182 46050 19234 46062
rect 22542 46114 22594 46126
rect 33182 46114 33234 46126
rect 25834 46062 25846 46114
rect 25898 46062 25910 46114
rect 22542 46050 22594 46062
rect 28814 46058 28866 46070
rect 33182 46050 33234 46062
rect 36990 46114 37042 46126
rect 36990 46050 37042 46062
rect 40798 46114 40850 46126
rect 40798 46050 40850 46062
rect 28814 45994 28866 46006
rect 44594 45950 44606 46002
rect 44658 45950 44670 46002
rect 7310 45890 7362 45902
rect 7310 45826 7362 45838
rect 10558 45890 10610 45902
rect 10558 45826 10610 45838
rect 12686 45890 12738 45902
rect 12686 45826 12738 45838
rect 13134 45890 13186 45902
rect 17502 45890 17554 45902
rect 13134 45826 13186 45838
rect 13906 45810 13918 45862
rect 13970 45810 13982 45862
rect 16146 45838 16158 45890
rect 16210 45838 16222 45890
rect 20750 45890 20802 45902
rect 17502 45826 17554 45838
rect 20066 45810 20078 45862
rect 20130 45810 20142 45862
rect 24446 45890 24498 45902
rect 20750 45826 20802 45838
rect 21522 45810 21534 45862
rect 21586 45810 21598 45862
rect 24446 45826 24498 45838
rect 24782 45890 24834 45902
rect 24782 45826 24834 45838
rect 26126 45890 26178 45902
rect 26126 45826 26178 45838
rect 26238 45890 26290 45902
rect 26238 45826 26290 45838
rect 26462 45890 26514 45902
rect 26462 45826 26514 45838
rect 27918 45890 27970 45902
rect 29486 45890 29538 45902
rect 28354 45838 28366 45890
rect 28418 45838 28430 45890
rect 28690 45838 28702 45890
rect 28754 45838 28766 45890
rect 27918 45826 27970 45838
rect 29486 45826 29538 45838
rect 29710 45890 29762 45902
rect 29710 45826 29762 45838
rect 30270 45890 30322 45902
rect 30270 45826 30322 45838
rect 30494 45890 30546 45902
rect 30494 45826 30546 45838
rect 30606 45890 30658 45902
rect 30606 45826 30658 45838
rect 30942 45890 30994 45902
rect 35310 45890 35362 45902
rect 30942 45826 30994 45838
rect 32162 45810 32174 45862
rect 32226 45810 32238 45862
rect 35018 45838 35030 45890
rect 35082 45838 35094 45890
rect 35310 45826 35362 45838
rect 35534 45890 35586 45902
rect 38670 45890 38722 45902
rect 35534 45826 35586 45838
rect 35970 45810 35982 45862
rect 36034 45810 36046 45862
rect 38670 45826 38722 45838
rect 38894 45890 38946 45902
rect 42478 45890 42530 45902
rect 38894 45826 38946 45838
rect 39778 45810 39790 45862
rect 39842 45810 39854 45862
rect 42478 45826 42530 45838
rect 42702 45890 42754 45902
rect 46286 45890 46338 45902
rect 42702 45826 42754 45838
rect 43586 45810 43598 45862
rect 43650 45810 43662 45862
rect 46286 45826 46338 45838
rect 46510 45890 46562 45902
rect 48078 45852 48130 45864
rect 46510 45826 46562 45838
rect 47350 45834 47402 45846
rect 21086 45778 21138 45790
rect 3894 45722 3946 45734
rect 3110 45666 3162 45678
rect 3110 45602 3162 45614
rect 3558 45666 3610 45678
rect 5574 45722 5626 45734
rect 3894 45658 3946 45670
rect 4566 45666 4618 45678
rect 3558 45602 3610 45614
rect 4566 45602 4618 45614
rect 5014 45666 5066 45678
rect 7030 45722 7082 45734
rect 5574 45658 5626 45670
rect 6246 45666 6298 45678
rect 5014 45602 5066 45614
rect 6246 45602 6298 45614
rect 6694 45666 6746 45678
rect 8598 45722 8650 45734
rect 7030 45658 7082 45670
rect 7646 45666 7698 45678
rect 6694 45602 6746 45614
rect 7646 45602 7698 45614
rect 8262 45666 8314 45678
rect 10166 45722 10218 45734
rect 8598 45658 8650 45670
rect 9830 45666 9882 45678
rect 8262 45602 8314 45614
rect 11398 45722 11450 45734
rect 10166 45658 10218 45670
rect 10894 45666 10946 45678
rect 9830 45602 9882 45614
rect 11398 45658 11450 45670
rect 11846 45722 11898 45734
rect 21086 45714 21138 45726
rect 25398 45722 25450 45734
rect 29194 45726 29206 45778
rect 29258 45726 29270 45778
rect 29978 45726 29990 45778
rect 30042 45726 30054 45778
rect 11846 45658 11898 45670
rect 12350 45666 12402 45678
rect 10894 45602 10946 45614
rect 12350 45602 12402 45614
rect 13470 45666 13522 45678
rect 13470 45602 13522 45614
rect 17166 45666 17218 45678
rect 31446 45722 31498 45734
rect 39162 45726 39174 45778
rect 39226 45726 39238 45778
rect 42970 45726 42982 45778
rect 43034 45726 43046 45778
rect 46778 45726 46790 45778
rect 46842 45726 46854 45778
rect 47350 45770 47402 45782
rect 47518 45778 47570 45790
rect 48078 45788 48130 45800
rect 48190 45834 48242 45846
rect 48190 45770 48242 45782
rect 25398 45658 25450 45670
rect 26798 45666 26850 45678
rect 17166 45602 17218 45614
rect 26798 45602 26850 45614
rect 27582 45666 27634 45678
rect 47518 45714 47570 45726
rect 31446 45658 31498 45670
rect 27582 45602 27634 45614
rect 1344 45498 48608 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 48608 45498
rect 1344 45412 48608 45446
rect 2662 45218 2714 45230
rect 2662 45154 2714 45166
rect 13022 45218 13074 45230
rect 13022 45154 13074 45166
rect 24446 45218 24498 45230
rect 24446 45154 24498 45166
rect 32398 45218 32450 45230
rect 32398 45154 32450 45166
rect 36262 45162 36314 45174
rect 40854 45162 40906 45174
rect 6190 45106 6242 45118
rect 5842 45054 5854 45106
rect 5906 45054 5918 45106
rect 6962 45054 6974 45106
rect 7026 45054 7038 45106
rect 9538 45054 9550 45106
rect 9602 45054 9614 45106
rect 9874 45069 9886 45121
rect 9938 45069 9950 45121
rect 10334 45106 10386 45118
rect 16270 45106 16322 45118
rect 11106 45054 11118 45106
rect 11170 45054 11182 45106
rect 15474 45054 15486 45106
rect 15538 45054 15550 45106
rect 6190 45042 6242 45054
rect 10334 45042 10386 45054
rect 16270 45042 16322 45054
rect 16942 45106 16994 45118
rect 16942 45042 16994 45054
rect 20750 45106 20802 45118
rect 20750 45042 20802 45054
rect 20974 45106 21026 45118
rect 20974 45042 21026 45054
rect 21198 45106 21250 45118
rect 21198 45042 21250 45054
rect 21758 45106 21810 45118
rect 21758 45042 21810 45054
rect 25230 45106 25282 45118
rect 28870 45106 28922 45118
rect 29150 45106 29202 45118
rect 26002 45054 26014 45106
rect 26066 45054 26078 45106
rect 29026 45054 29038 45106
rect 29090 45054 29102 45106
rect 25230 45042 25282 45054
rect 28870 45042 28922 45054
rect 29150 45042 29202 45054
rect 29710 45106 29762 45118
rect 29710 45042 29762 45054
rect 33070 45106 33122 45118
rect 36418 45110 36430 45162
rect 36482 45110 36494 45162
rect 36642 45110 36654 45162
rect 36706 45110 36718 45162
rect 36262 45098 36314 45110
rect 37550 45106 37602 45118
rect 33070 45042 33122 45054
rect 40854 45098 40906 45110
rect 41010 45084 41022 45136
rect 41074 45084 41086 45136
rect 41234 45093 41246 45145
rect 41298 45093 41310 45145
rect 42254 45106 42306 45118
rect 37550 45042 37602 45054
rect 42254 45042 42306 45054
rect 45390 45106 45442 45118
rect 46162 45054 46174 45106
rect 46226 45054 46238 45106
rect 45390 45042 45442 45054
rect 2214 44994 2266 45006
rect 2214 44930 2266 44942
rect 3110 44994 3162 45006
rect 3110 44930 3162 44942
rect 3558 44994 3610 45006
rect 3558 44930 3610 44942
rect 4006 44994 4058 45006
rect 4006 44930 4058 44942
rect 4454 44994 4506 45006
rect 4454 44930 4506 44942
rect 4902 44994 4954 45006
rect 4902 44930 4954 44942
rect 5350 44994 5402 45006
rect 17670 44994 17722 45006
rect 8866 44942 8878 44994
rect 8930 44942 8942 44994
rect 9986 44942 9998 44994
rect 10050 44942 10062 44994
rect 13570 44942 13582 44994
rect 13634 44942 13646 44994
rect 18050 44942 18062 44994
rect 18114 44942 18126 44994
rect 19954 44942 19966 44994
rect 20018 44942 20030 44994
rect 22530 44942 22542 44994
rect 22594 44942 22606 44994
rect 27906 44942 27918 44994
rect 27970 44942 27982 44994
rect 30482 44942 30494 44994
rect 30546 44942 30558 44994
rect 33842 44942 33854 44994
rect 33906 44942 33918 44994
rect 35746 44942 35758 44994
rect 35810 44942 35822 44994
rect 38322 44942 38334 44994
rect 38386 44942 38398 44994
rect 40226 44942 40238 44994
rect 40290 44942 40302 44994
rect 43026 44942 43038 44994
rect 43090 44942 43102 44994
rect 44930 44942 44942 44994
rect 44994 44942 45006 44994
rect 48066 44942 48078 44994
rect 48130 44942 48142 44994
rect 5350 44930 5402 44942
rect 17670 44930 17722 44942
rect 5686 44882 5738 44894
rect 5686 44818 5738 44830
rect 16606 44882 16658 44894
rect 28478 44882 28530 44894
rect 21466 44830 21478 44882
rect 21530 44830 21542 44882
rect 16606 44818 16658 44830
rect 28478 44818 28530 44830
rect 37214 44882 37266 44894
rect 37214 44818 37266 44830
rect 41806 44882 41858 44894
rect 41806 44818 41858 44830
rect 1344 44714 48608 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 48608 44714
rect 1344 44628 48608 44662
rect 12686 44546 12738 44558
rect 6794 44494 6806 44546
rect 6858 44494 6870 44546
rect 12686 44482 12738 44494
rect 22318 44546 22370 44558
rect 22318 44482 22370 44494
rect 25006 44546 25058 44558
rect 37998 44546 38050 44558
rect 26730 44494 26742 44546
rect 26794 44494 26806 44546
rect 29530 44494 29542 44546
rect 29594 44494 29606 44546
rect 25006 44482 25058 44494
rect 37998 44482 38050 44494
rect 40910 44546 40962 44558
rect 40910 44482 40962 44494
rect 45614 44546 45666 44558
rect 45614 44482 45666 44494
rect 25678 44434 25730 44446
rect 8262 44378 8314 44390
rect 10658 44382 10670 44434
rect 10722 44382 10734 44434
rect 14466 44382 14478 44434
rect 14530 44382 14542 44434
rect 18498 44382 18510 44434
rect 18562 44382 18574 44434
rect 2270 44322 2322 44334
rect 5966 44322 6018 44334
rect 3042 44270 3054 44322
rect 3106 44270 3118 44322
rect 2270 44258 2322 44270
rect 5966 44258 6018 44270
rect 6078 44322 6130 44334
rect 6078 44258 6130 44270
rect 7086 44322 7138 44334
rect 7086 44258 7138 44270
rect 7310 44322 7362 44334
rect 7870 44322 7922 44334
rect 7578 44270 7590 44322
rect 7642 44270 7654 44322
rect 7310 44258 7362 44270
rect 7870 44258 7922 44270
rect 8094 44322 8146 44334
rect 8262 44314 8314 44326
rect 8430 44322 8482 44334
rect 9090 44326 9102 44378
rect 9154 44326 9166 44378
rect 25678 44370 25730 44382
rect 8094 44258 8146 44270
rect 9662 44322 9714 44334
rect 11790 44322 11842 44334
rect 8430 44258 8482 44270
rect 8990 44266 9042 44278
rect 4958 44210 5010 44222
rect 9662 44258 9714 44270
rect 9986 44243 9998 44295
rect 10050 44243 10062 44295
rect 10210 44270 10222 44322
rect 10274 44270 10286 44322
rect 10770 44226 10782 44278
rect 10834 44226 10846 44278
rect 10994 44270 11006 44322
rect 11058 44270 11070 44322
rect 11790 44258 11842 44270
rect 13022 44322 13074 44334
rect 17614 44322 17666 44334
rect 14130 44270 14142 44322
rect 14194 44270 14206 44322
rect 13022 44258 13074 44270
rect 14354 44226 14366 44278
rect 14418 44226 14430 44278
rect 16818 44270 16830 44322
rect 16882 44270 16894 44322
rect 17614 44258 17666 44270
rect 17726 44322 17778 44334
rect 23998 44322 24050 44334
rect 17726 44258 17778 44270
rect 21298 44242 21310 44294
rect 21362 44242 21374 44294
rect 23998 44258 24050 44270
rect 24222 44322 24274 44334
rect 24222 44258 24274 44270
rect 25342 44322 25394 44334
rect 27022 44322 27074 44334
rect 25342 44258 25394 44270
rect 25510 44266 25562 44278
rect 25890 44270 25902 44322
rect 25954 44270 25966 44322
rect 6346 44158 6358 44210
rect 6410 44158 6422 44210
rect 8990 44202 9042 44214
rect 14926 44210 14978 44222
rect 4958 44146 5010 44158
rect 2102 44098 2154 44110
rect 9762 44102 9774 44154
rect 9826 44102 9838 44154
rect 14926 44146 14978 44158
rect 20414 44210 20466 44222
rect 24490 44158 24502 44210
rect 24554 44158 24566 44210
rect 25510 44202 25562 44214
rect 26238 44266 26290 44278
rect 27022 44258 27074 44270
rect 27246 44322 27298 44334
rect 27246 44258 27298 44270
rect 27918 44322 27970 44334
rect 28478 44322 28530 44334
rect 28186 44270 28198 44322
rect 28250 44270 28262 44322
rect 27918 44258 27970 44270
rect 28478 44258 28530 44270
rect 28590 44322 28642 44334
rect 28590 44258 28642 44270
rect 29150 44322 29202 44334
rect 29150 44258 29202 44270
rect 29262 44322 29314 44334
rect 29262 44258 29314 44270
rect 31614 44322 31666 44334
rect 36430 44322 36482 44334
rect 47518 44322 47570 44334
rect 32274 44270 32286 44322
rect 32338 44270 32350 44322
rect 26238 44202 26290 44214
rect 30494 44210 30546 44222
rect 30725 44214 30737 44266
rect 30789 44214 30801 44266
rect 31614 44258 31666 44270
rect 34178 44242 34190 44294
rect 34242 44242 34254 44294
rect 35541 44270 35553 44322
rect 35605 44270 35617 44322
rect 36430 44258 36482 44270
rect 36978 44242 36990 44294
rect 37042 44242 37054 44294
rect 39890 44242 39902 44294
rect 39954 44242 39966 44294
rect 43250 44240 43262 44292
rect 43314 44240 43326 44292
rect 43474 44231 43486 44283
rect 43538 44231 43550 44283
rect 43766 44266 43818 44278
rect 44258 44270 44270 44322
rect 44322 44270 44334 44322
rect 20414 44146 20466 44158
rect 29990 44154 30042 44166
rect 2102 44034 2154 44046
rect 11622 44098 11674 44110
rect 11622 44034 11674 44046
rect 12126 44098 12178 44110
rect 12126 44034 12178 44046
rect 13526 44098 13578 44110
rect 13526 44034 13578 44046
rect 27582 44098 27634 44110
rect 30494 44146 30546 44158
rect 35310 44210 35362 44222
rect 35310 44146 35362 44158
rect 42814 44210 42866 44222
rect 47170 44242 47182 44294
rect 47234 44242 47246 44294
rect 47518 44258 47570 44270
rect 47742 44322 47794 44334
rect 47742 44258 47794 44270
rect 43766 44202 43818 44214
rect 48010 44158 48022 44210
rect 48074 44158 48086 44210
rect 42814 44146 42866 44158
rect 29990 44090 30042 44102
rect 44102 44098 44154 44110
rect 27582 44034 27634 44046
rect 44102 44034 44154 44046
rect 1344 43930 48608 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 48608 43930
rect 1344 43844 48608 43878
rect 19294 43762 19346 43774
rect 4062 43650 4114 43662
rect 4062 43586 4114 43598
rect 6526 43650 6578 43662
rect 7074 43654 7086 43706
rect 7138 43654 7150 43706
rect 6526 43586 6578 43598
rect 8318 43650 8370 43662
rect 15586 43654 15598 43706
rect 15650 43654 15662 43706
rect 19294 43698 19346 43710
rect 38054 43706 38106 43718
rect 7422 43577 7474 43589
rect 8318 43586 8370 43598
rect 17670 43650 17722 43662
rect 4398 43538 4450 43550
rect 4722 43486 4734 43538
rect 4786 43486 4798 43538
rect 4946 43501 4958 43553
rect 5010 43501 5022 43553
rect 5406 43538 5458 43550
rect 7198 43538 7250 43550
rect 6270 43486 6282 43538
rect 6334 43486 6346 43538
rect 7422 43513 7474 43525
rect 7746 43486 7758 43538
rect 7810 43486 7822 43538
rect 4398 43474 4450 43486
rect 5406 43474 5458 43486
rect 7198 43474 7250 43486
rect 8150 43482 8202 43494
rect 8530 43486 8542 43538
rect 8594 43486 8606 43538
rect 8754 43514 8766 43566
rect 8818 43514 8830 43566
rect 9438 43538 9490 43550
rect 1878 43426 1930 43438
rect 1878 43362 1930 43374
rect 2326 43426 2378 43438
rect 2326 43362 2378 43374
rect 2774 43426 2826 43438
rect 2774 43362 2826 43374
rect 3222 43426 3274 43438
rect 3222 43362 3274 43374
rect 3670 43426 3722 43438
rect 9438 43474 9490 43486
rect 9662 43538 9714 43550
rect 9662 43474 9714 43486
rect 10222 43538 10274 43550
rect 10222 43474 10274 43486
rect 11006 43538 11058 43550
rect 12126 43538 12178 43550
rect 11870 43486 11882 43538
rect 11934 43486 11946 43538
rect 11006 43474 11058 43486
rect 12126 43474 12178 43486
rect 12574 43538 12626 43550
rect 13438 43486 13450 43538
rect 13502 43486 13514 43538
rect 14242 43516 14254 43568
rect 14306 43516 14318 43568
rect 14466 43525 14478 43577
rect 14530 43525 14542 43577
rect 15038 43538 15090 43550
rect 12574 43474 12626 43486
rect 14746 43430 14758 43482
rect 14810 43430 14822 43482
rect 15038 43474 15090 43486
rect 15710 43538 15762 43550
rect 15922 43542 15934 43594
rect 15986 43542 15998 43594
rect 17670 43586 17722 43598
rect 23102 43650 23154 43662
rect 23930 43598 23942 43650
rect 23994 43598 24006 43650
rect 38054 43642 38106 43654
rect 41022 43650 41074 43662
rect 23102 43586 23154 43598
rect 28086 43594 28138 43606
rect 16886 43538 16938 43550
rect 16370 43486 16382 43538
rect 16434 43486 16446 43538
rect 17938 43513 17950 43565
rect 18002 43513 18014 43565
rect 20862 43538 20914 43550
rect 15710 43474 15762 43486
rect 16886 43474 16938 43486
rect 21726 43486 21738 43538
rect 21790 43486 21802 43538
rect 22642 43514 22654 43566
rect 22706 43514 22718 43566
rect 23438 43538 23490 43550
rect 22866 43486 22878 43538
rect 22930 43486 22942 43538
rect 20862 43474 20914 43486
rect 23270 43482 23322 43494
rect 23438 43474 23490 43486
rect 23662 43538 23714 43550
rect 23662 43474 23714 43486
rect 24222 43538 24274 43550
rect 25902 43538 25954 43550
rect 27358 43538 27410 43550
rect 25442 43486 25454 43538
rect 25506 43486 25518 43538
rect 26766 43486 26778 43538
rect 26830 43486 26842 43538
rect 24222 43474 24274 43486
rect 25902 43474 25954 43486
rect 27358 43474 27410 43486
rect 27694 43538 27746 43550
rect 28086 43530 28138 43542
rect 28242 43516 28254 43568
rect 28306 43516 28318 43568
rect 28466 43525 28478 43577
rect 28530 43525 28542 43577
rect 31984 43575 32036 43587
rect 41022 43586 41074 43598
rect 45054 43650 45106 43662
rect 29934 43538 29986 43550
rect 27694 43474 27746 43486
rect 29934 43474 29986 43486
rect 30158 43538 30210 43550
rect 30482 43516 30494 43568
rect 30546 43516 30558 43568
rect 30818 43516 30830 43568
rect 30882 43516 30894 43568
rect 31278 43538 31330 43550
rect 30158 43474 30210 43486
rect 30986 43430 30998 43482
rect 31050 43430 31062 43482
rect 31278 43474 31330 43486
rect 31726 43538 31778 43550
rect 31826 43486 31838 43538
rect 31890 43486 31902 43538
rect 34414 43538 34466 43550
rect 31984 43511 32036 43523
rect 33058 43486 33070 43538
rect 33122 43486 33134 43538
rect 33730 43486 33742 43538
rect 33794 43486 33806 43538
rect 35522 43513 35534 43565
rect 35586 43513 35598 43565
rect 38558 43538 38610 43550
rect 39678 43538 39730 43550
rect 37874 43486 37886 43538
rect 37938 43486 37950 43538
rect 38789 43486 38801 43538
rect 38853 43486 38865 43538
rect 31726 43474 31778 43486
rect 34414 43474 34466 43486
rect 38558 43474 38610 43486
rect 39678 43474 39730 43486
rect 39902 43538 39954 43550
rect 41253 43542 41265 43594
rect 41317 43542 41329 43594
rect 45054 43586 45106 43598
rect 39902 43474 39954 43486
rect 42142 43538 42194 43550
rect 42690 43516 42702 43568
rect 42754 43516 42766 43568
rect 43026 43516 43038 43568
rect 43090 43516 43102 43568
rect 43486 43538 43538 43550
rect 42142 43474 42194 43486
rect 5058 43374 5070 43426
rect 5122 43374 5134 43426
rect 8150 43418 8202 43430
rect 9930 43374 9942 43426
rect 9994 43374 10006 43426
rect 23270 43418 23322 43430
rect 34078 43426 34130 43438
rect 43194 43430 43206 43482
rect 43258 43430 43270 43482
rect 43486 43474 43538 43486
rect 43934 43538 43986 43550
rect 45390 43538 45442 43550
rect 44798 43486 44810 43538
rect 44862 43486 44874 43538
rect 43934 43474 43986 43486
rect 45390 43474 45442 43486
rect 29642 43374 29654 43426
rect 29706 43374 29718 43426
rect 36194 43374 36206 43426
rect 36258 43374 36270 43426
rect 46162 43374 46174 43426
rect 46226 43374 46238 43426
rect 48066 43374 48078 43426
rect 48130 43374 48142 43426
rect 3670 43362 3722 43374
rect 34078 43362 34130 43374
rect 10558 43314 10610 43326
rect 10558 43250 10610 43262
rect 13694 43314 13746 43326
rect 13694 43250 13746 43262
rect 21982 43314 22034 43326
rect 21982 43250 22034 43262
rect 24558 43314 24610 43326
rect 24558 43250 24610 43262
rect 25286 43314 25338 43326
rect 25286 43250 25338 43262
rect 27022 43314 27074 43326
rect 27022 43250 27074 43262
rect 29038 43314 29090 43326
rect 29038 43250 29090 43262
rect 32398 43314 32450 43326
rect 32398 43250 32450 43262
rect 34750 43314 34802 43326
rect 34750 43250 34802 43262
rect 40238 43314 40290 43326
rect 40238 43250 40290 43262
rect 1344 43146 48608 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 48608 43146
rect 1344 43060 48608 43094
rect 7086 42978 7138 42990
rect 20638 42978 20690 42990
rect 5674 42926 5686 42978
rect 5738 42926 5750 42978
rect 14186 42926 14198 42978
rect 14250 42926 14262 42978
rect 7086 42914 7138 42926
rect 20638 42914 20690 42926
rect 26574 42978 26626 42990
rect 26574 42914 26626 42926
rect 28478 42978 28530 42990
rect 28478 42914 28530 42926
rect 32454 42978 32506 42990
rect 43038 42978 43090 42990
rect 32454 42914 32506 42926
rect 35870 42922 35922 42934
rect 15262 42866 15314 42878
rect 12450 42814 12462 42866
rect 12514 42814 12526 42866
rect 15262 42802 15314 42814
rect 21982 42866 22034 42878
rect 43038 42914 43090 42926
rect 45838 42978 45890 42990
rect 45838 42914 45890 42926
rect 23538 42814 23550 42866
rect 23602 42814 23614 42866
rect 25442 42814 25454 42866
rect 25506 42814 25518 42866
rect 32050 42814 32062 42866
rect 32114 42814 32126 42866
rect 35410 42814 35422 42866
rect 35474 42814 35486 42866
rect 35870 42858 35922 42870
rect 42254 42866 42306 42878
rect 21982 42802 22034 42814
rect 1598 42754 1650 42766
rect 4286 42754 4338 42766
rect 1598 42690 1650 42702
rect 3602 42687 3614 42739
rect 3666 42687 3678 42739
rect 3938 42702 3950 42754
rect 4002 42702 4014 42754
rect 4286 42690 4338 42702
rect 4398 42754 4450 42766
rect 4398 42690 4450 42702
rect 5966 42754 6018 42766
rect 5966 42690 6018 42702
rect 6190 42754 6242 42766
rect 6190 42690 6242 42702
rect 6414 42754 6466 42766
rect 6692 42754 6744 42766
rect 6514 42702 6526 42754
rect 6578 42702 6590 42754
rect 6414 42690 6466 42702
rect 6692 42690 6744 42702
rect 7646 42754 7698 42766
rect 7646 42690 7698 42702
rect 7870 42754 7922 42766
rect 7870 42690 7922 42702
rect 9102 42754 9154 42766
rect 13806 42754 13858 42766
rect 9874 42702 9886 42754
rect 9938 42702 9950 42754
rect 9102 42690 9154 42702
rect 12562 42687 12574 42739
rect 12626 42687 12638 42739
rect 12898 42702 12910 42754
rect 12962 42702 12974 42754
rect 13806 42690 13858 42702
rect 13918 42754 13970 42766
rect 16382 42754 16434 42766
rect 13918 42690 13970 42702
rect 14702 42698 14754 42710
rect 15026 42702 15038 42754
rect 15090 42702 15102 42754
rect 11790 42642 11842 42654
rect 3614 42586 3666 42598
rect 4666 42590 4678 42642
rect 4730 42590 4742 42642
rect 8138 42590 8150 42642
rect 8202 42590 8214 42642
rect 14702 42634 14754 42646
rect 15430 42698 15482 42710
rect 16146 42702 16158 42754
rect 16210 42702 16222 42754
rect 17166 42754 17218 42766
rect 15922 42646 15934 42698
rect 15986 42646 15998 42698
rect 16382 42690 16434 42702
rect 16550 42698 16602 42710
rect 17166 42690 17218 42702
rect 17390 42754 17442 42766
rect 17390 42690 17442 42702
rect 17502 42754 17554 42766
rect 17502 42690 17554 42702
rect 17726 42754 17778 42766
rect 19182 42754 19234 42766
rect 19966 42754 20018 42766
rect 20246 42754 20298 42766
rect 22150 42754 22202 42766
rect 22766 42754 22818 42766
rect 17994 42702 18006 42754
rect 18058 42702 18070 42754
rect 19730 42702 19742 42754
rect 19794 42702 19806 42754
rect 20066 42702 20078 42754
rect 20130 42702 20142 42754
rect 21746 42702 21758 42754
rect 21810 42702 21822 42754
rect 22306 42702 22318 42754
rect 22370 42702 22382 42754
rect 17726 42690 17778 42702
rect 19182 42690 19234 42702
rect 19966 42690 20018 42702
rect 20246 42690 20298 42702
rect 21522 42646 21534 42698
rect 21586 42646 21598 42698
rect 22150 42690 22202 42702
rect 22766 42690 22818 42702
rect 25902 42754 25954 42766
rect 27358 42754 27410 42766
rect 29710 42754 29762 42766
rect 26002 42702 26014 42754
rect 26066 42702 26078 42754
rect 28222 42702 28234 42754
rect 28286 42702 28298 42754
rect 25902 42690 25954 42702
rect 26168 42646 26180 42698
rect 26232 42646 26244 42698
rect 27358 42690 27410 42702
rect 29710 42690 29762 42702
rect 29934 42754 29986 42766
rect 32734 42754 32786 42766
rect 36878 42754 36930 42766
rect 31602 42702 31614 42754
rect 31666 42702 31678 42754
rect 29934 42690 29986 42702
rect 30798 42646 30810 42698
rect 30862 42646 30874 42698
rect 31938 42687 31950 42739
rect 32002 42687 32014 42739
rect 32274 42702 32286 42754
rect 32338 42702 32350 42754
rect 33506 42702 33518 42754
rect 33570 42702 33582 42754
rect 35970 42702 35982 42754
rect 36034 42702 36046 42754
rect 36194 42702 36206 42754
rect 36258 42702 36270 42754
rect 32734 42690 32786 42702
rect 36878 42690 36930 42702
rect 37102 42754 37154 42766
rect 40798 42754 40850 42766
rect 41570 42758 41582 42810
rect 41634 42758 41646 42810
rect 42254 42802 42306 42814
rect 42422 42810 42474 42822
rect 40002 42702 40014 42754
rect 40066 42702 40078 42754
rect 41010 42702 41022 42754
rect 41074 42702 41086 42754
rect 42422 42746 42474 42758
rect 47518 42754 47570 42766
rect 41694 42716 41746 42728
rect 37102 42690 37154 42702
rect 40798 42690 40850 42702
rect 43990 42698 44042 42710
rect 15430 42634 15482 42646
rect 16550 42634 16602 42646
rect 31054 42642 31106 42654
rect 38110 42642 38162 42654
rect 41694 42652 41746 42664
rect 43418 42646 43430 42698
rect 43482 42646 43494 42698
rect 43698 42646 43710 42698
rect 43762 42646 43774 42698
rect 45042 42674 45054 42726
rect 45106 42674 45118 42726
rect 47518 42690 47570 42702
rect 47742 42754 47794 42766
rect 47742 42690 47794 42702
rect 16874 42590 16886 42642
rect 16938 42590 16950 42642
rect 1934 42530 1986 42542
rect 1934 42466 1986 42478
rect 2774 42530 2826 42542
rect 2774 42466 2826 42478
rect 3222 42530 3274 42542
rect 11790 42578 11842 42590
rect 19574 42586 19626 42598
rect 3614 42522 3666 42534
rect 8934 42530 8986 42542
rect 3222 42466 3274 42478
rect 8934 42466 8986 42478
rect 18846 42530 18898 42542
rect 37370 42590 37382 42642
rect 37434 42590 37446 42642
rect 43990 42634 44042 42646
rect 48010 42590 48022 42642
rect 48074 42590 48086 42642
rect 31054 42578 31106 42590
rect 38110 42578 38162 42590
rect 19574 42522 19626 42534
rect 22486 42530 22538 42542
rect 18846 42466 18898 42478
rect 22486 42466 22538 42478
rect 29374 42530 29426 42542
rect 29374 42466 29426 42478
rect 41190 42530 41242 42542
rect 41190 42466 41242 42478
rect 1344 42362 48608 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 48608 42362
rect 1344 42276 48608 42310
rect 9662 42194 9714 42206
rect 9662 42130 9714 42142
rect 34582 42194 34634 42206
rect 4846 42082 4898 42094
rect 4846 42018 4898 42030
rect 7870 42082 7922 42094
rect 10322 42086 10334 42138
rect 10386 42086 10398 42138
rect 24546 42086 24558 42138
rect 24610 42086 24622 42138
rect 34582 42130 34634 42142
rect 40182 42194 40234 42206
rect 40182 42130 40234 42142
rect 43990 42194 44042 42206
rect 43990 42130 44042 42142
rect 28590 42082 28642 42094
rect 7870 42018 7922 42030
rect 27638 42026 27690 42038
rect 10670 42009 10722 42021
rect 1598 41970 1650 41982
rect 1598 41906 1650 41918
rect 4286 41970 4338 41982
rect 5966 41970 6018 41982
rect 5077 41918 5089 41970
rect 5141 41918 5153 41970
rect 4286 41906 4338 41918
rect 5966 41906 6018 41918
rect 6302 41970 6354 41982
rect 7702 41970 7754 41982
rect 6850 41918 6862 41970
rect 6914 41918 6926 41970
rect 8082 41918 8094 41970
rect 8146 41918 8158 41970
rect 8306 41946 8318 41998
rect 8370 41946 8382 41998
rect 9998 41970 10050 41982
rect 8754 41918 8766 41970
rect 8818 41918 8830 41970
rect 10322 41918 10334 41970
rect 10386 41918 10398 41970
rect 15896 42007 15948 42019
rect 10670 41945 10722 41957
rect 10894 41970 10946 41982
rect 6302 41906 6354 41918
rect 7702 41906 7754 41918
rect 9998 41906 10050 41918
rect 10894 41906 10946 41918
rect 11790 41970 11842 41982
rect 11790 41906 11842 41918
rect 12014 41970 12066 41982
rect 13022 41970 13074 41982
rect 15150 41970 15202 41982
rect 12450 41918 12462 41970
rect 12514 41918 12526 41970
rect 13886 41918 13898 41970
rect 13950 41918 13962 41970
rect 14858 41918 14870 41970
rect 14922 41918 14934 41970
rect 12014 41906 12066 41918
rect 13022 41906 13074 41918
rect 15150 41906 15202 41918
rect 15374 41970 15426 41982
rect 15374 41906 15426 41918
rect 15598 41970 15650 41982
rect 15698 41918 15710 41970
rect 15762 41918 15774 41970
rect 22430 42008 22482 42020
rect 15896 41943 15948 41955
rect 17614 41970 17666 41982
rect 20750 41970 20802 41982
rect 21870 41970 21922 41982
rect 18386 41918 18398 41970
rect 18450 41918 18462 41970
rect 21614 41918 21626 41970
rect 21678 41918 21690 41970
rect 24222 42009 24274 42021
rect 22430 41944 22482 41956
rect 22754 41918 22766 41970
rect 22818 41918 22830 41970
rect 15598 41906 15650 41918
rect 17614 41906 17666 41918
rect 20750 41906 20802 41918
rect 21870 41906 21922 41918
rect 23158 41914 23210 41926
rect 23762 41918 23774 41970
rect 23826 41918 23838 41970
rect 24222 41945 24274 41957
rect 24446 41970 24498 41982
rect 16270 41858 16322 41870
rect 2370 41806 2382 41858
rect 2434 41806 2446 41858
rect 7074 41750 7086 41802
rect 7138 41750 7150 41802
rect 16270 41794 16322 41806
rect 16886 41858 16938 41870
rect 22990 41858 23042 41870
rect 20290 41806 20302 41858
rect 20354 41806 20366 41858
rect 24446 41906 24498 41918
rect 25230 41970 25282 41982
rect 26686 41970 26738 41982
rect 26094 41918 26106 41970
rect 26158 41918 26170 41970
rect 25230 41906 25282 41918
rect 26686 41906 26738 41918
rect 26910 41970 26962 41982
rect 28590 42018 28642 42030
rect 37998 42082 38050 42094
rect 27178 41918 27190 41970
rect 27242 41918 27254 41970
rect 27638 41962 27690 41974
rect 27794 41948 27806 42000
rect 27858 41948 27870 42000
rect 28130 41948 28142 42000
rect 28194 41948 28206 42000
rect 30158 41970 30210 41982
rect 29138 41918 29150 41970
rect 29202 41918 29214 41970
rect 29474 41918 29486 41970
rect 29538 41918 29550 41970
rect 26910 41906 26962 41918
rect 30158 41906 30210 41918
rect 30942 41970 30994 41982
rect 31806 41974 31818 42026
rect 31870 41974 31882 42026
rect 30942 41906 30994 41918
rect 32062 41970 32114 41982
rect 32062 41906 32114 41918
rect 32958 41970 33010 41982
rect 32958 41906 33010 41918
rect 33294 41970 33346 41982
rect 33294 41906 33346 41918
rect 33966 41970 34018 41982
rect 33966 41906 34018 41918
rect 34302 41970 34354 41982
rect 34974 41970 35026 41982
rect 36642 41974 36654 42026
rect 36706 41974 36718 42026
rect 37998 42018 38050 42030
rect 39118 42026 39170 42038
rect 34738 41918 34750 41970
rect 34802 41918 34814 41970
rect 35838 41918 35850 41970
rect 35902 41918 35914 41970
rect 36978 41948 36990 42000
rect 37042 41948 37054 42000
rect 34302 41906 34354 41918
rect 34974 41906 35026 41918
rect 37830 41914 37882 41926
rect 38210 41918 38222 41970
rect 38274 41918 38286 41970
rect 38434 41946 38446 41998
rect 38498 41946 38510 41998
rect 44326 42026 44378 42038
rect 39118 41962 39170 41974
rect 40798 41970 40850 41982
rect 44482 41974 44494 42026
rect 44546 41974 44558 42026
rect 44818 41974 44830 42026
rect 44882 41974 44894 42026
rect 39442 41918 39454 41970
rect 39506 41918 39518 41970
rect 23158 41850 23210 41862
rect 36094 41858 36146 41870
rect 37146 41862 37158 41914
rect 37210 41862 37222 41914
rect 16886 41794 16938 41806
rect 22990 41794 23042 41806
rect 29598 41802 29650 41814
rect 8934 41746 8986 41758
rect 12294 41746 12346 41758
rect 11498 41694 11510 41746
rect 11562 41694 11574 41746
rect 8934 41682 8986 41694
rect 12294 41682 12346 41694
rect 14142 41746 14194 41758
rect 14142 41682 14194 41694
rect 26350 41746 26402 41758
rect 36094 41794 36146 41806
rect 37438 41858 37490 41870
rect 39846 41914 39898 41926
rect 40338 41918 40350 41970
rect 40402 41918 40414 41970
rect 44146 41918 44158 41970
rect 44210 41918 44222 41970
rect 44326 41962 44378 41974
rect 45714 41945 45726 41997
rect 45778 41945 45790 41997
rect 37830 41850 37882 41862
rect 39678 41858 39730 41870
rect 37438 41794 37490 41806
rect 40798 41906 40850 41918
rect 39846 41850 39898 41862
rect 41570 41806 41582 41858
rect 41634 41806 41646 41858
rect 43474 41806 43486 41858
rect 43538 41806 43550 41858
rect 46722 41806 46734 41858
rect 46786 41806 46798 41858
rect 39678 41794 39730 41806
rect 29598 41738 29650 41750
rect 30494 41746 30546 41758
rect 26350 41682 26402 41694
rect 30494 41682 30546 41694
rect 45278 41746 45330 41758
rect 45278 41682 45330 41694
rect 1344 41578 48608 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 48608 41578
rect 1344 41492 48608 41526
rect 2382 41410 2434 41422
rect 2382 41346 2434 41358
rect 12014 41410 12066 41422
rect 12014 41346 12066 41358
rect 14366 41410 14418 41422
rect 14366 41346 14418 41358
rect 16046 41410 16098 41422
rect 16046 41346 16098 41358
rect 19742 41410 19794 41422
rect 19742 41346 19794 41358
rect 22206 41410 22258 41422
rect 33070 41410 33122 41422
rect 22698 41358 22710 41410
rect 22762 41358 22774 41410
rect 35914 41358 35926 41410
rect 35978 41358 35990 41410
rect 1990 41298 2042 41310
rect 20402 41302 20414 41354
rect 20466 41302 20478 41354
rect 22206 41346 22258 41358
rect 33070 41346 33122 41358
rect 28646 41298 28698 41310
rect 12450 41246 12462 41298
rect 12514 41246 12526 41298
rect 24658 41246 24670 41298
rect 24722 41246 24734 41298
rect 25442 41246 25454 41298
rect 25506 41246 25518 41298
rect 1990 41234 2042 41246
rect 28646 41234 28698 41246
rect 37662 41298 37714 41310
rect 37662 41234 37714 41246
rect 37830 41242 37882 41254
rect 41346 41246 41358 41298
rect 41410 41246 41422 41298
rect 2718 41186 2770 41198
rect 3950 41186 4002 41198
rect 3266 41134 3278 41186
rect 3330 41134 3342 41186
rect 2718 41122 2770 41134
rect 3602 41107 3614 41159
rect 3666 41107 3678 41159
rect 3950 41122 4002 41134
rect 4510 41186 4562 41198
rect 4510 41122 4562 41134
rect 4622 41186 4674 41198
rect 4622 41122 4674 41134
rect 5518 41186 5570 41198
rect 9886 41186 9938 41198
rect 6290 41134 6302 41186
rect 6354 41134 6366 41186
rect 5518 41122 5570 41134
rect 8206 41074 8258 41086
rect 4890 41022 4902 41074
rect 4954 41022 4966 41074
rect 3378 40966 3390 41018
rect 3442 40966 3454 41018
rect 8206 41010 8258 41022
rect 8766 41074 8818 41086
rect 8997 41078 9009 41130
rect 9061 41078 9073 41130
rect 9886 41122 9938 41134
rect 10894 41186 10946 41198
rect 14926 41186 14978 41198
rect 10894 41122 10946 41134
rect 11758 41103 11770 41155
rect 11822 41103 11834 41155
rect 12562 41090 12574 41142
rect 12626 41090 12638 41142
rect 12786 41134 12798 41186
rect 12850 41134 12862 41186
rect 13414 41130 13466 41142
rect 8766 41010 8818 41022
rect 10614 41074 10666 41086
rect 13570 41104 13582 41156
rect 13634 41104 13646 41156
rect 13906 41078 13918 41130
rect 13970 41078 13982 41130
rect 14926 41122 14978 41134
rect 16718 41186 16770 41198
rect 19406 41186 19458 41198
rect 18610 41134 18622 41186
rect 18674 41134 18686 41186
rect 15790 41078 15802 41130
rect 15854 41078 15866 41130
rect 16718 41122 16770 41134
rect 19406 41122 19458 41134
rect 20078 41186 20130 41198
rect 22990 41186 23042 41198
rect 20402 41134 20414 41186
rect 20466 41134 20478 41186
rect 20626 41134 20638 41186
rect 20690 41134 20702 41186
rect 20078 41122 20130 41134
rect 21254 41130 21306 41142
rect 21522 41095 21534 41147
rect 21586 41095 21598 41147
rect 21802 41078 21814 41130
rect 21866 41078 21878 41130
rect 22990 41122 23042 41134
rect 23214 41186 23266 41198
rect 23214 41122 23266 41134
rect 23326 41186 23378 41198
rect 23326 41122 23378 41134
rect 23550 41186 23602 41198
rect 26574 41186 26626 41198
rect 23818 41134 23830 41186
rect 23882 41134 23894 41186
rect 23550 41122 23602 41134
rect 24770 41119 24782 41171
rect 24834 41119 24846 41171
rect 25106 41134 25118 41186
rect 25170 41134 25182 41186
rect 25554 41090 25566 41142
rect 25618 41090 25630 41142
rect 25890 41134 25902 41186
rect 25954 41134 25966 41186
rect 26574 41122 26626 41134
rect 29038 41186 29090 41198
rect 27438 41078 27450 41130
rect 27502 41078 27514 41130
rect 29038 41122 29090 41134
rect 29822 41186 29874 41198
rect 30942 41186 30994 41198
rect 30686 41134 30698 41186
rect 30750 41134 30762 41186
rect 29822 41122 29874 41134
rect 30942 41122 30994 41134
rect 31390 41186 31442 41198
rect 33406 41186 33458 41198
rect 32254 41134 32266 41186
rect 32318 41134 32330 41186
rect 31390 41122 31442 41134
rect 33406 41122 33458 41134
rect 34078 41186 34130 41198
rect 34078 41122 34130 41134
rect 34750 41186 34802 41198
rect 34750 41122 34802 41134
rect 35086 41186 35138 41198
rect 35086 41122 35138 41134
rect 36206 41186 36258 41198
rect 36206 41122 36258 41134
rect 36318 41186 36370 41198
rect 42758 41242 42810 41254
rect 36318 41122 36370 41134
rect 37202 41106 37214 41158
rect 37266 41106 37278 41158
rect 37426 41134 37438 41186
rect 37490 41134 37502 41186
rect 37830 41178 37882 41190
rect 38110 41186 38162 41198
rect 42198 41186 42250 41198
rect 38882 41134 38894 41186
rect 38946 41134 38958 41186
rect 38110 41122 38162 41134
rect 41458 41119 41470 41171
rect 41522 41119 41534 41171
rect 41794 41134 41806 41186
rect 41858 41134 41870 41186
rect 42198 41122 42250 41134
rect 42478 41186 42530 41198
rect 43206 41242 43258 41254
rect 48066 41246 48078 41298
rect 48130 41246 48142 41298
rect 42758 41178 42810 41190
rect 42926 41186 42978 41198
rect 42478 41122 42530 41134
rect 43206 41178 43258 41190
rect 45278 41186 45330 41198
rect 43586 41134 43598 41186
rect 43650 41134 43662 41186
rect 43934 41148 43986 41160
rect 42926 41122 42978 41134
rect 45278 41122 45330 41134
rect 45390 41186 45442 41198
rect 46162 41134 46174 41186
rect 46226 41134 46238 41186
rect 45390 41122 45442 41134
rect 13414 41066 13466 41078
rect 21254 41066 21306 41078
rect 27694 41074 27746 41086
rect 10614 41010 10666 41022
rect 24278 41018 24330 41030
rect 27694 41010 27746 41022
rect 32510 41074 32562 41086
rect 32510 41010 32562 41022
rect 40798 41074 40850 41086
rect 40798 41010 40850 41022
rect 42590 41074 42642 41086
rect 42590 41010 42642 41022
rect 43374 41074 43426 41086
rect 43934 41084 43986 41096
rect 43374 41010 43426 41022
rect 24278 40954 24330 40966
rect 29374 40962 29426 40974
rect 29374 40898 29426 40910
rect 33742 40962 33794 40974
rect 33742 40898 33794 40910
rect 34414 40962 34466 40974
rect 34414 40898 34466 40910
rect 35422 40962 35474 40974
rect 35422 40898 35474 40910
rect 44942 40962 44994 40974
rect 44942 40898 44994 40910
rect 1344 40794 48608 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 48608 40794
rect 1344 40708 48608 40742
rect 2886 40626 2938 40638
rect 2886 40562 2938 40574
rect 6638 40626 6690 40638
rect 6638 40562 6690 40574
rect 9718 40626 9770 40638
rect 9718 40562 9770 40574
rect 10166 40626 10218 40638
rect 10166 40562 10218 40574
rect 15318 40626 15370 40638
rect 15318 40562 15370 40574
rect 17614 40626 17666 40638
rect 1990 40514 2042 40526
rect 6246 40514 6298 40526
rect 8878 40514 8930 40526
rect 1990 40450 2042 40462
rect 3390 40458 3442 40470
rect 7242 40462 7254 40514
rect 7306 40462 7318 40514
rect 2438 40402 2490 40414
rect 3390 40394 3442 40406
rect 4162 40380 4174 40432
rect 4226 40380 4238 40432
rect 4386 40406 4398 40458
rect 4450 40406 4462 40458
rect 6246 40450 6298 40462
rect 7926 40458 7978 40470
rect 4846 40402 4898 40414
rect 2438 40338 2490 40350
rect 3994 40294 4006 40346
rect 4058 40294 4070 40346
rect 4846 40338 4898 40350
rect 5070 40402 5122 40414
rect 6974 40402 7026 40414
rect 5338 40350 5350 40402
rect 5402 40350 5414 40402
rect 5070 40338 5122 40350
rect 6974 40338 7026 40350
rect 7534 40402 7586 40414
rect 7534 40338 7586 40350
rect 7758 40402 7810 40414
rect 8082 40406 8094 40458
rect 8146 40406 8158 40458
rect 8306 40406 8318 40458
rect 8370 40406 8382 40458
rect 8878 40450 8930 40462
rect 14702 40514 14754 40526
rect 16482 40518 16494 40570
rect 16546 40518 16558 40570
rect 17614 40562 17666 40574
rect 19798 40626 19850 40638
rect 19798 40562 19850 40574
rect 24726 40626 24778 40638
rect 24726 40562 24778 40574
rect 32286 40626 32338 40638
rect 32286 40562 32338 40574
rect 7926 40394 7978 40406
rect 10614 40402 10666 40414
rect 7758 40338 7810 40350
rect 10882 40350 10894 40402
rect 10946 40350 10958 40402
rect 11218 40394 11230 40446
rect 11282 40394 11294 40446
rect 11976 40440 12028 40452
rect 11678 40402 11730 40414
rect 11778 40350 11790 40402
rect 11842 40350 11854 40402
rect 13582 40402 13634 40414
rect 14446 40406 14458 40458
rect 14510 40406 14522 40458
rect 14702 40450 14754 40462
rect 18230 40514 18282 40526
rect 28926 40514 28978 40526
rect 20906 40462 20918 40514
rect 20970 40462 20982 40514
rect 30942 40514 30994 40526
rect 16270 40441 16322 40453
rect 18230 40450 18282 40462
rect 16046 40402 16098 40414
rect 11976 40376 12028 40388
rect 12786 40350 12798 40402
rect 12850 40350 12862 40402
rect 13122 40350 13134 40402
rect 13186 40350 13198 40402
rect 15474 40350 15486 40402
rect 15538 40350 15550 40402
rect 25712 40439 25764 40451
rect 17278 40402 17330 40414
rect 16270 40377 16322 40389
rect 16594 40350 16606 40402
rect 16658 40350 16670 40402
rect 10614 40338 10666 40350
rect 11678 40338 11730 40350
rect 13582 40338 13634 40350
rect 16046 40338 16098 40350
rect 17278 40338 17330 40350
rect 19294 40402 19346 40414
rect 20414 40402 20466 40414
rect 20290 40350 20302 40402
rect 20354 40350 20366 40402
rect 19294 40338 19346 40350
rect 20414 40338 20466 40350
rect 20638 40402 20690 40414
rect 20638 40338 20690 40350
rect 21310 40402 21362 40414
rect 21590 40402 21642 40414
rect 21410 40350 21422 40402
rect 21474 40350 21486 40402
rect 21310 40338 21362 40350
rect 21590 40338 21642 40350
rect 22430 40402 22482 40414
rect 22430 40338 22482 40350
rect 22542 40402 22594 40414
rect 24222 40402 24274 40414
rect 22810 40350 22822 40402
rect 22874 40350 22886 40402
rect 22542 40338 22594 40350
rect 24222 40338 24274 40350
rect 25454 40402 25506 40414
rect 25554 40350 25566 40402
rect 25618 40350 25630 40402
rect 25712 40375 25764 40387
rect 26462 40402 26514 40414
rect 25454 40338 25506 40350
rect 26462 40338 26514 40350
rect 26686 40402 26738 40414
rect 26686 40338 26738 40350
rect 27526 40402 27578 40414
rect 27526 40338 27578 40350
rect 27806 40402 27858 40414
rect 28670 40406 28682 40458
rect 28734 40406 28746 40458
rect 28926 40450 28978 40462
rect 30662 40458 30714 40470
rect 27806 40338 27858 40350
rect 29766 40402 29818 40414
rect 30146 40406 30158 40458
rect 30210 40406 30222 40458
rect 30482 40380 30494 40432
rect 30546 40380 30558 40432
rect 36990 40514 37042 40526
rect 46398 40514 46450 40526
rect 30942 40450 30994 40462
rect 36710 40458 36762 40470
rect 30662 40394 30714 40406
rect 31278 40402 31330 40414
rect 29766 40338 29818 40350
rect 31278 40338 31330 40350
rect 31502 40402 31554 40414
rect 32622 40402 32674 40414
rect 31770 40350 31782 40402
rect 31834 40350 31846 40402
rect 31502 40338 31554 40350
rect 32622 40338 32674 40350
rect 32958 40402 33010 40414
rect 35646 40402 35698 40414
rect 36194 40406 36206 40458
rect 36258 40406 36270 40458
rect 33730 40350 33742 40402
rect 33794 40350 33806 40402
rect 36418 40389 36430 40441
rect 36482 40389 36494 40441
rect 42746 40462 42758 40514
rect 42810 40462 42822 40514
rect 36990 40450 37042 40462
rect 36710 40394 36762 40406
rect 37326 40402 37378 40414
rect 32958 40338 33010 40350
rect 35646 40338 35698 40350
rect 37326 40338 37378 40350
rect 37550 40402 37602 40414
rect 38334 40402 38386 40414
rect 37818 40350 37830 40402
rect 37882 40350 37894 40402
rect 37550 40338 37602 40350
rect 38334 40338 38386 40350
rect 38446 40402 38498 40414
rect 38446 40338 38498 40350
rect 39454 40402 39506 40414
rect 39454 40338 39506 40350
rect 39678 40402 39730 40414
rect 39678 40338 39730 40350
rect 40238 40402 40290 40414
rect 40238 40338 40290 40350
rect 40462 40402 40514 40414
rect 40462 40338 40514 40350
rect 41246 40402 41298 40414
rect 41526 40402 41578 40414
rect 41346 40350 41358 40402
rect 41410 40350 41422 40402
rect 41246 40338 41298 40350
rect 41526 40338 41578 40350
rect 42254 40402 42306 40414
rect 42254 40338 42306 40350
rect 42478 40402 42530 40414
rect 42478 40338 42530 40350
rect 43374 40402 43426 40414
rect 43642 40406 43654 40458
rect 43706 40406 43718 40458
rect 44494 40402 44546 40414
rect 45358 40406 45370 40458
rect 45422 40406 45434 40458
rect 46398 40450 46450 40462
rect 43474 40350 43486 40402
rect 43538 40350 43550 40402
rect 43374 40338 43426 40350
rect 44494 40338 44546 40350
rect 45614 40402 45666 40414
rect 45614 40338 45666 40350
rect 46062 40402 46114 40414
rect 46062 40338 46114 40350
rect 46230 40402 46282 40414
rect 46230 40338 46282 40350
rect 46510 40402 46562 40414
rect 46510 40338 46562 40350
rect 47126 40402 47178 40414
rect 47730 40406 47742 40458
rect 47794 40406 47806 40458
rect 47506 40350 47518 40402
rect 47570 40350 47582 40402
rect 47126 40338 47178 40350
rect 12350 40290 12402 40302
rect 11330 40238 11342 40290
rect 11394 40238 11406 40290
rect 21982 40290 22034 40302
rect 12350 40226 12402 40238
rect 13246 40234 13298 40246
rect 3222 40178 3274 40190
rect 3222 40114 3274 40126
rect 3726 40178 3778 40190
rect 21982 40226 22034 40238
rect 23494 40290 23546 40302
rect 23494 40226 23546 40238
rect 26126 40290 26178 40302
rect 41918 40290 41970 40302
rect 26954 40238 26966 40290
rect 27018 40238 27030 40290
rect 26126 40226 26178 40238
rect 41918 40226 41970 40238
rect 47294 40290 47346 40302
rect 47294 40226 47346 40238
rect 13246 40170 13298 40182
rect 18958 40178 19010 40190
rect 3726 40114 3778 40126
rect 18958 40114 19010 40126
rect 20134 40178 20186 40190
rect 20134 40114 20186 40126
rect 23886 40178 23938 40190
rect 44046 40178 44098 40190
rect 38714 40126 38726 40178
rect 38778 40126 38790 40178
rect 39162 40126 39174 40178
rect 39226 40126 39238 40178
rect 39946 40126 39958 40178
rect 40010 40126 40022 40178
rect 23886 40114 23938 40126
rect 44046 40114 44098 40126
rect 46790 40178 46842 40190
rect 46790 40114 46842 40126
rect 1344 40010 48608 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 48608 40010
rect 1344 39924 48608 39958
rect 8094 39842 8146 39854
rect 8094 39778 8146 39790
rect 10334 39842 10386 39854
rect 10334 39778 10386 39790
rect 12854 39842 12906 39854
rect 12854 39778 12906 39790
rect 16830 39842 16882 39854
rect 16830 39778 16882 39790
rect 36206 39842 36258 39854
rect 6302 39730 6354 39742
rect 17558 39730 17610 39742
rect 31390 39730 31442 39742
rect 32610 39734 32622 39786
rect 32674 39734 32686 39786
rect 36206 39778 36258 39790
rect 37718 39842 37770 39854
rect 37718 39778 37770 39790
rect 4274 39678 4286 39730
rect 4338 39678 4350 39730
rect 16258 39678 16270 39730
rect 16322 39678 16334 39730
rect 18610 39678 18622 39730
rect 18674 39678 18686 39730
rect 20514 39678 20526 39730
rect 20578 39678 20590 39730
rect 23538 39678 23550 39730
rect 23602 39678 23614 39730
rect 25442 39678 25454 39730
rect 25506 39678 25518 39730
rect 28522 39678 28534 39730
rect 28586 39678 28598 39730
rect 6302 39666 6354 39678
rect 17558 39666 17610 39678
rect 31390 39666 31442 39678
rect 37158 39674 37210 39686
rect 1598 39618 1650 39630
rect 12126 39618 12178 39630
rect 2370 39566 2382 39618
rect 2434 39566 2446 39618
rect 1598 39554 1650 39566
rect 5842 39538 5854 39590
rect 5906 39538 5918 39590
rect 6066 39566 6078 39618
rect 6130 39566 6142 39618
rect 6470 39562 6522 39574
rect 6962 39566 6974 39618
rect 7026 39566 7038 39618
rect 5126 39506 5178 39518
rect 6470 39498 6522 39510
rect 7142 39562 7194 39574
rect 9986 39566 9998 39618
rect 10050 39566 10062 39618
rect 11286 39562 11338 39574
rect 7410 39510 7422 39562
rect 7474 39510 7486 39562
rect 7690 39510 7702 39562
rect 7754 39510 7766 39562
rect 10770 39510 10782 39562
rect 10834 39510 10846 39562
rect 11106 39510 11118 39562
rect 11170 39510 11182 39562
rect 12126 39554 12178 39566
rect 12294 39618 12346 39630
rect 12294 39554 12346 39566
rect 12574 39618 12626 39630
rect 13806 39618 13858 39630
rect 13514 39566 13526 39618
rect 13578 39566 13590 39618
rect 12574 39554 12626 39566
rect 13806 39554 13858 39566
rect 13918 39618 13970 39630
rect 13918 39554 13970 39566
rect 14254 39618 14306 39630
rect 17166 39618 17218 39630
rect 15922 39566 15934 39618
rect 15986 39566 15998 39618
rect 14254 39554 14306 39566
rect 7142 39498 7194 39510
rect 11286 39498 11338 39510
rect 12462 39506 12514 39518
rect 15118 39510 15130 39562
rect 15182 39510 15194 39562
rect 5126 39442 5178 39454
rect 12462 39442 12514 39454
rect 15374 39506 15426 39518
rect 16090 39510 16102 39562
rect 16154 39510 16166 39562
rect 17166 39554 17218 39566
rect 17838 39618 17890 39630
rect 17838 39554 17890 39566
rect 21310 39618 21362 39630
rect 21310 39554 21362 39566
rect 22766 39618 22818 39630
rect 22174 39510 22186 39562
rect 22238 39510 22250 39562
rect 22766 39554 22818 39566
rect 26238 39618 26290 39630
rect 26238 39554 26290 39566
rect 27358 39618 27410 39630
rect 15374 39442 15426 39454
rect 22430 39506 22482 39518
rect 27102 39510 27114 39562
rect 27166 39510 27178 39562
rect 27358 39554 27410 39566
rect 28142 39618 28194 39630
rect 28142 39554 28194 39566
rect 28254 39618 28306 39630
rect 29710 39618 29762 39630
rect 29026 39566 29038 39618
rect 29090 39566 29102 39618
rect 28254 39554 28306 39566
rect 29710 39554 29762 39566
rect 30830 39618 30882 39630
rect 33070 39618 33122 39630
rect 30574 39510 30586 39562
rect 30638 39510 30650 39562
rect 30830 39554 30882 39566
rect 31222 39562 31274 39574
rect 31602 39566 31614 39618
rect 31666 39566 31678 39618
rect 32386 39566 32398 39618
rect 32450 39566 32462 39618
rect 32722 39566 32734 39618
rect 32786 39566 32798 39618
rect 31770 39510 31782 39562
rect 31834 39510 31846 39562
rect 33070 39554 33122 39566
rect 33294 39618 33346 39630
rect 34526 39618 34578 39630
rect 36542 39618 36594 39630
rect 33562 39566 33574 39618
rect 33626 39566 33638 39618
rect 34290 39566 34302 39618
rect 34354 39566 34366 39618
rect 35390 39566 35402 39618
rect 35454 39566 35466 39618
rect 33294 39554 33346 39566
rect 34526 39554 34578 39566
rect 36542 39554 36594 39566
rect 36990 39618 37042 39630
rect 37158 39610 37210 39622
rect 37438 39618 37490 39630
rect 37314 39566 37326 39618
rect 37378 39566 37390 39618
rect 36990 39554 37042 39566
rect 37438 39554 37490 39566
rect 38222 39618 38274 39630
rect 41358 39618 41410 39630
rect 45278 39618 45330 39630
rect 38994 39566 39006 39618
rect 39058 39566 39070 39618
rect 42130 39566 42142 39618
rect 42194 39566 42206 39618
rect 38222 39554 38274 39566
rect 41358 39554 41410 39566
rect 45278 39554 45330 39566
rect 45390 39618 45442 39630
rect 46162 39566 46174 39618
rect 46226 39566 46238 39618
rect 45390 39554 45442 39566
rect 31222 39498 31274 39510
rect 35646 39506 35698 39518
rect 22430 39442 22482 39454
rect 29206 39450 29258 39462
rect 6806 39394 6858 39406
rect 6806 39330 6858 39342
rect 9046 39394 9098 39406
rect 9046 39330 9098 39342
rect 9494 39394 9546 39406
rect 9494 39330 9546 39342
rect 9830 39394 9882 39406
rect 9830 39330 9882 39342
rect 11846 39394 11898 39406
rect 35646 39442 35698 39454
rect 40910 39506 40962 39518
rect 40910 39442 40962 39454
rect 44046 39506 44098 39518
rect 44046 39442 44098 39454
rect 48078 39506 48130 39518
rect 48078 39442 48130 39454
rect 29206 39386 29258 39398
rect 34134 39394 34186 39406
rect 11846 39330 11898 39342
rect 34134 39330 34186 39342
rect 44942 39394 44994 39406
rect 44942 39330 44994 39342
rect 1344 39226 48608 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 48608 39226
rect 1344 39140 48608 39174
rect 2270 39058 2322 39070
rect 2270 38994 2322 39006
rect 15598 39058 15650 39070
rect 15598 38994 15650 39006
rect 16606 39058 16658 39070
rect 16606 38994 16658 39006
rect 23494 39058 23546 39070
rect 4062 38946 4114 38958
rect 2606 38834 2658 38846
rect 2606 38770 2658 38782
rect 2942 38834 2994 38846
rect 3806 38838 3818 38890
rect 3870 38838 3882 38890
rect 4062 38882 4114 38894
rect 5182 38946 5234 38958
rect 14926 38946 14978 38958
rect 22306 38950 22318 39002
rect 22370 38950 22382 39002
rect 23494 38994 23546 39006
rect 27750 39058 27802 39070
rect 24546 38950 24558 39002
rect 24610 38950 24622 39002
rect 27750 38994 27802 39006
rect 37606 39058 37658 39070
rect 5182 38882 5234 38894
rect 8094 38890 8146 38902
rect 7870 38834 7922 38846
rect 7074 38782 7086 38834
rect 7138 38782 7150 38834
rect 8094 38826 8146 38838
rect 8206 38872 8258 38884
rect 14366 38872 14418 38884
rect 14926 38882 14978 38894
rect 26350 38946 26402 38958
rect 30706 38950 30718 39002
rect 30770 38950 30782 39002
rect 37606 38994 37658 39006
rect 39902 39058 39954 39070
rect 39902 38994 39954 39006
rect 41134 39058 41186 39070
rect 41134 38994 41186 39006
rect 8206 38808 8258 38820
rect 8766 38834 8818 38846
rect 2942 38770 2994 38782
rect 7870 38770 7922 38782
rect 9438 38834 9490 38846
rect 8766 38770 8818 38782
rect 8934 38778 8986 38790
rect 4678 38722 4730 38734
rect 12718 38820 12730 38872
rect 12782 38820 12794 38872
rect 13458 38782 13470 38834
rect 13522 38782 13534 38834
rect 15934 38834 15986 38846
rect 14366 38808 14418 38820
rect 14690 38782 14702 38834
rect 14754 38782 14766 38834
rect 9438 38770 9490 38782
rect 15094 38778 15146 38790
rect 8934 38714 8986 38726
rect 15934 38770 15986 38782
rect 16942 38834 16994 38846
rect 16942 38770 16994 38782
rect 17502 38834 17554 38846
rect 20850 38782 20862 38834
rect 20914 38782 20926 38834
rect 21074 38826 21086 38878
rect 21138 38826 21150 38878
rect 21982 38873 22034 38885
rect 21758 38834 21810 38846
rect 24042 38838 24054 38890
rect 24106 38838 24118 38890
rect 26350 38882 26402 38894
rect 31390 38946 31442 38958
rect 39230 38946 39282 38958
rect 24446 38834 24498 38846
rect 21982 38809 22034 38821
rect 22306 38782 22318 38834
rect 22370 38782 22382 38834
rect 23762 38782 23774 38834
rect 23826 38782 23838 38834
rect 17502 38770 17554 38782
rect 21758 38770 21810 38782
rect 24446 38770 24498 38782
rect 25230 38834 25282 38846
rect 26094 38813 26106 38865
rect 26158 38813 26170 38865
rect 28030 38834 28082 38846
rect 28894 38838 28906 38890
rect 28958 38838 28970 38890
rect 31390 38882 31442 38894
rect 32342 38890 32394 38902
rect 26786 38782 26798 38834
rect 26850 38782 26862 38834
rect 27122 38782 27134 38834
rect 27186 38782 27198 38834
rect 25230 38770 25282 38782
rect 28030 38770 28082 38782
rect 29150 38834 29202 38846
rect 29150 38770 29202 38782
rect 29934 38834 29986 38846
rect 31770 38838 31782 38890
rect 31834 38838 31846 38890
rect 30482 38782 30494 38834
rect 30546 38782 30558 38834
rect 32162 38812 32174 38864
rect 32226 38812 32238 38864
rect 35534 38890 35586 38902
rect 42422 38946 42474 38958
rect 32342 38826 32394 38838
rect 33070 38834 33122 38846
rect 35086 38834 35138 38846
rect 33934 38782 33946 38834
rect 33998 38782 34010 38834
rect 34794 38782 34806 38834
rect 34858 38782 34870 38834
rect 29934 38770 29986 38782
rect 33070 38770 33122 38782
rect 35086 38770 35138 38782
rect 35310 38834 35362 38846
rect 35802 38838 35814 38890
rect 35866 38838 35878 38890
rect 38144 38871 38196 38883
rect 39230 38882 39282 38894
rect 41507 38890 41559 38902
rect 45894 38946 45946 38958
rect 35534 38826 35586 38838
rect 36374 38834 36426 38846
rect 35310 38770 35362 38782
rect 36374 38770 36426 38782
rect 36542 38834 36594 38846
rect 36542 38770 36594 38782
rect 36766 38834 36818 38846
rect 36766 38770 36818 38782
rect 37886 38834 37938 38846
rect 37986 38782 37998 38834
rect 38050 38782 38062 38834
rect 38144 38807 38196 38819
rect 38894 38834 38946 38846
rect 37886 38770 37938 38782
rect 38894 38770 38946 38782
rect 39566 38834 39618 38846
rect 39566 38770 39618 38782
rect 40798 38834 40850 38846
rect 41682 38838 41694 38890
rect 41746 38838 41758 38890
rect 41918 38862 41970 38874
rect 41507 38826 41559 38838
rect 42130 38838 42142 38890
rect 42194 38838 42206 38890
rect 42422 38882 42474 38894
rect 44718 38890 44770 38902
rect 44158 38862 44210 38874
rect 43878 38834 43930 38846
rect 41918 38798 41970 38810
rect 43138 38782 43150 38834
rect 43202 38782 43214 38834
rect 43362 38782 43374 38834
rect 43426 38782 43438 38834
rect 44158 38798 44210 38810
rect 44382 38862 44434 38874
rect 44594 38838 44606 38890
rect 44658 38838 44670 38890
rect 44718 38826 44770 38838
rect 45054 38890 45106 38902
rect 47450 38894 47462 38946
rect 47514 38894 47526 38946
rect 45054 38826 45106 38838
rect 45166 38862 45218 38874
rect 44382 38798 44434 38810
rect 45166 38798 45218 38810
rect 45390 38862 45442 38874
rect 45602 38838 45614 38890
rect 45666 38838 45678 38890
rect 45894 38882 45946 38894
rect 45390 38798 45442 38810
rect 46286 38834 46338 38846
rect 46564 38834 46616 38846
rect 40798 38770 40850 38782
rect 43878 38770 43930 38782
rect 46386 38782 46398 38834
rect 46450 38782 46462 38834
rect 46286 38770 46338 38782
rect 46564 38770 46616 38782
rect 47742 38834 47794 38846
rect 47742 38770 47794 38782
rect 47854 38834 47906 38846
rect 47854 38770 47906 38782
rect 10210 38670 10222 38722
rect 10274 38670 10286 38722
rect 12114 38670 12126 38722
rect 12178 38670 12190 38722
rect 15094 38714 15146 38726
rect 22934 38722 22986 38734
rect 4678 38658 4730 38670
rect 13582 38666 13634 38678
rect 18274 38670 18286 38722
rect 18338 38670 18350 38722
rect 20178 38670 20190 38722
rect 20242 38670 20254 38722
rect 21186 38670 21198 38722
rect 21250 38670 21262 38722
rect 36206 38722 36258 38734
rect 22934 38658 22986 38670
rect 27246 38666 27298 38678
rect 13582 38602 13634 38614
rect 36206 38658 36258 38670
rect 38558 38722 38610 38734
rect 46958 38722 47010 38734
rect 38558 38658 38610 38670
rect 43486 38666 43538 38678
rect 27246 38602 27298 38614
rect 34190 38610 34242 38622
rect 46958 38658 47010 38670
rect 37034 38558 37046 38610
rect 37098 38558 37110 38610
rect 43486 38602 43538 38614
rect 34190 38546 34242 38558
rect 1344 38442 48608 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 48608 38442
rect 1344 38356 48608 38390
rect 7870 38274 7922 38286
rect 18622 38274 18674 38286
rect 7870 38210 7922 38222
rect 9774 38218 9826 38230
rect 2998 38162 3050 38174
rect 2998 38098 3050 38110
rect 3446 38162 3498 38174
rect 3446 38098 3498 38110
rect 6470 38162 6522 38174
rect 8642 38166 8654 38218
rect 8706 38166 8718 38218
rect 9774 38154 9826 38166
rect 12126 38218 12178 38230
rect 14590 38218 14642 38230
rect 12562 38166 12574 38218
rect 12626 38166 12638 38218
rect 12126 38154 12178 38166
rect 13862 38162 13914 38174
rect 6470 38098 6522 38110
rect 18622 38210 18674 38222
rect 22206 38274 22258 38286
rect 22206 38210 22258 38222
rect 28478 38274 28530 38286
rect 28478 38210 28530 38222
rect 31838 38274 31890 38286
rect 31838 38210 31890 38222
rect 32342 38274 32394 38286
rect 32342 38210 32394 38222
rect 34526 38274 34578 38286
rect 34526 38210 34578 38222
rect 35310 38274 35362 38286
rect 35310 38210 35362 38222
rect 35982 38274 36034 38286
rect 35982 38210 36034 38222
rect 39342 38274 39394 38286
rect 39342 38210 39394 38222
rect 39902 38274 39954 38286
rect 39902 38210 39954 38222
rect 42086 38274 42138 38286
rect 42086 38210 42138 38222
rect 43262 38218 43314 38230
rect 14590 38154 14642 38166
rect 22822 38162 22874 38174
rect 13862 38098 13914 38110
rect 22822 38098 22874 38110
rect 23214 38162 23266 38174
rect 23214 38098 23266 38110
rect 24614 38162 24666 38174
rect 24614 38098 24666 38110
rect 25174 38162 25226 38174
rect 43262 38154 43314 38166
rect 48066 38110 48078 38162
rect 48130 38110 48142 38162
rect 25174 38098 25226 38110
rect 2606 38050 2658 38062
rect 4062 38050 4114 38062
rect 3770 37998 3782 38050
rect 3834 37998 3846 38050
rect 2606 37986 2658 37998
rect 4062 37986 4114 37998
rect 4286 38050 4338 38062
rect 4846 38050 4898 38062
rect 4554 37998 4566 38050
rect 4618 37998 4630 38050
rect 4286 37986 4338 37998
rect 4846 37986 4898 37998
rect 4958 38050 5010 38062
rect 4958 37986 5010 37998
rect 6750 38050 6802 38062
rect 10110 38050 10162 38062
rect 14926 38050 14978 38062
rect 16046 38050 16098 38062
rect 6750 37986 6802 37998
rect 7614 37967 7626 38019
rect 7678 37967 7690 38019
rect 8418 37998 8430 38050
rect 8482 37998 8494 38050
rect 8754 37998 8766 38050
rect 8818 37998 8830 38050
rect 9426 37998 9438 38050
rect 9490 37998 9502 38050
rect 9650 37998 9662 38050
rect 9714 37998 9726 38050
rect 11666 37998 11678 38050
rect 11730 37998 11742 38050
rect 12002 37998 12014 38050
rect 12066 37998 12078 38050
rect 12562 37998 12574 38050
rect 12626 37998 12638 38050
rect 12786 37998 12798 38050
rect 12850 37998 12862 38050
rect 14242 37998 14254 38050
rect 14306 37998 14318 38050
rect 14466 37998 14478 38050
rect 14530 37998 14542 38050
rect 15790 37998 15802 38050
rect 15854 37998 15866 38050
rect 10110 37986 10162 37998
rect 10974 37942 10986 37994
rect 11038 37942 11050 37994
rect 14926 37986 14978 37998
rect 16046 37986 16098 37998
rect 16942 38050 16994 38062
rect 16942 37986 16994 37998
rect 18958 38050 19010 38062
rect 23550 38050 23602 38062
rect 18958 37986 19010 37998
rect 21254 37994 21306 38006
rect 11230 37938 11282 37950
rect 11230 37874 11282 37886
rect 19686 37938 19738 37950
rect 21466 37942 21478 37994
rect 21530 37942 21542 37994
rect 21634 37942 21646 37994
rect 21698 37942 21710 37994
rect 23550 37986 23602 37998
rect 23662 38050 23714 38062
rect 23662 37986 23714 37998
rect 26238 38050 26290 38062
rect 26238 37986 26290 37998
rect 26350 38050 26402 38062
rect 26350 37986 26402 37998
rect 26574 38050 26626 38062
rect 26574 37986 26626 37998
rect 26798 38050 26850 38062
rect 29150 38050 29202 38062
rect 30270 38050 30322 38062
rect 26798 37986 26850 37998
rect 27526 37994 27578 38006
rect 27794 37942 27806 37994
rect 27858 37942 27870 37994
rect 28018 37968 28030 38020
rect 28082 37968 28094 38020
rect 30014 37998 30026 38050
rect 30078 37998 30090 38050
rect 29150 37986 29202 37998
rect 30270 37986 30322 37998
rect 30718 38050 30770 38062
rect 34190 38050 34242 38062
rect 32162 37998 32174 38050
rect 32226 37998 32238 38050
rect 32610 37998 32622 38050
rect 32674 37998 32686 38050
rect 30718 37986 30770 37998
rect 31582 37942 31594 37994
rect 31646 37942 31658 37994
rect 34190 37986 34242 37998
rect 34862 38050 34914 38062
rect 34862 37986 34914 37998
rect 34974 38050 35026 38062
rect 34974 37986 35026 37998
rect 35646 38050 35698 38062
rect 35646 37986 35698 37998
rect 37438 38050 37490 38062
rect 37438 37986 37490 37998
rect 37998 38050 38050 38062
rect 37998 37986 38050 37998
rect 38110 38050 38162 38062
rect 39006 38050 39058 38062
rect 38110 37986 38162 37998
rect 38334 37994 38386 38006
rect 39006 37986 39058 37998
rect 40238 38050 40290 38062
rect 44214 38050 44266 38062
rect 40238 37986 40290 37998
rect 41134 38022 41186 38034
rect 41694 38015 41746 38027
rect 41134 37958 41186 37970
rect 21254 37930 21306 37942
rect 25946 37886 25958 37938
rect 26010 37886 26022 37938
rect 27066 37886 27078 37938
rect 27130 37886 27142 37938
rect 27526 37930 27578 37942
rect 19686 37874 19738 37886
rect 32790 37882 32842 37894
rect 37706 37886 37718 37938
rect 37770 37886 37782 37938
rect 38334 37930 38386 37942
rect 40854 37938 40906 37950
rect 41346 37942 41358 37994
rect 41410 37942 41422 37994
rect 41570 37942 41582 37994
rect 41634 37942 41646 37994
rect 41694 37951 41746 37963
rect 42366 38022 42418 38034
rect 42366 37958 42418 37970
rect 42590 38022 42642 38034
rect 42590 37958 42642 37970
rect 42814 38022 42866 38034
rect 42814 37958 42866 37970
rect 42926 37994 42978 38006
rect 43362 37998 43374 38050
rect 43426 37998 43438 38050
rect 43698 37998 43710 38050
rect 43762 37998 43774 38050
rect 44214 37986 44266 37998
rect 45278 38050 45330 38062
rect 45278 37986 45330 37998
rect 45390 38050 45442 38062
rect 46162 37998 46174 38050
rect 46226 37998 46238 38050
rect 45390 37986 45442 37998
rect 42926 37930 42978 37942
rect 2270 37826 2322 37838
rect 2270 37762 2322 37774
rect 5798 37826 5850 37838
rect 5798 37762 5850 37774
rect 16606 37826 16658 37838
rect 16606 37762 16658 37774
rect 17334 37826 17386 37838
rect 17334 37762 17386 37774
rect 17782 37826 17834 37838
rect 17782 37762 17834 37774
rect 18230 37826 18282 37838
rect 18230 37762 18282 37774
rect 20134 37826 20186 37838
rect 20134 37762 20186 37774
rect 20582 37826 20634 37838
rect 20582 37762 20634 37774
rect 23998 37826 24050 37838
rect 23998 37762 24050 37774
rect 25622 37826 25674 37838
rect 40854 37874 40906 37886
rect 32790 37818 32842 37830
rect 33462 37826 33514 37838
rect 25622 37762 25674 37774
rect 33462 37762 33514 37774
rect 33854 37826 33906 37838
rect 33854 37762 33906 37774
rect 37102 37826 37154 37838
rect 37102 37762 37154 37774
rect 38670 37826 38722 37838
rect 38670 37762 38722 37774
rect 44942 37826 44994 37838
rect 44942 37762 44994 37774
rect 1344 37658 48608 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 48608 37658
rect 1344 37572 48608 37606
rect 9046 37490 9098 37502
rect 9046 37426 9098 37438
rect 14646 37490 14698 37502
rect 14646 37426 14698 37438
rect 20246 37490 20298 37502
rect 20246 37426 20298 37438
rect 30662 37490 30714 37502
rect 30662 37426 30714 37438
rect 35646 37490 35698 37502
rect 35646 37426 35698 37438
rect 41246 37490 41298 37502
rect 41246 37426 41298 37438
rect 41918 37490 41970 37502
rect 41918 37426 41970 37438
rect 43374 37490 43426 37502
rect 43374 37426 43426 37438
rect 4846 37378 4898 37390
rect 7198 37378 7250 37390
rect 10110 37378 10162 37390
rect 13358 37378 13410 37390
rect 4846 37314 4898 37326
rect 6246 37322 6298 37334
rect 1598 37266 1650 37278
rect 4286 37266 4338 37278
rect 5966 37266 6018 37278
rect 2370 37214 2382 37266
rect 2434 37214 2446 37266
rect 5077 37214 5089 37266
rect 5141 37214 5153 37266
rect 8026 37326 8038 37378
rect 8090 37326 8102 37378
rect 7198 37314 7250 37326
rect 9942 37322 9994 37334
rect 6246 37258 6298 37270
rect 6402 37244 6414 37296
rect 6466 37244 6478 37296
rect 6738 37244 6750 37296
rect 6802 37244 6814 37296
rect 7646 37266 7698 37278
rect 1598 37202 1650 37214
rect 4286 37202 4338 37214
rect 5966 37202 6018 37214
rect 7646 37202 7698 37214
rect 7758 37266 7810 37278
rect 10110 37314 10162 37326
rect 10670 37322 10722 37334
rect 12842 37326 12854 37378
rect 12906 37326 12918 37378
rect 9942 37258 9994 37270
rect 13358 37314 13410 37326
rect 16382 37378 16434 37390
rect 25678 37378 25730 37390
rect 16382 37314 16434 37326
rect 22318 37322 22370 37334
rect 10322 37214 10334 37266
rect 10386 37214 10398 37266
rect 10670 37258 10722 37270
rect 11666 37214 11678 37266
rect 11730 37214 11742 37266
rect 12002 37229 12014 37281
rect 12066 37229 12078 37281
rect 12350 37266 12402 37278
rect 7758 37202 7810 37214
rect 12350 37202 12402 37214
rect 12574 37266 12626 37278
rect 12574 37202 12626 37214
rect 13190 37210 13242 37222
rect 13570 37214 13582 37266
rect 13634 37214 13646 37266
rect 13794 37242 13806 37294
rect 13858 37242 13870 37294
rect 16718 37266 16770 37278
rect 14466 37214 14478 37266
rect 14530 37214 14542 37266
rect 18274 37242 18286 37294
rect 18338 37242 18350 37294
rect 19070 37266 19122 37278
rect 18498 37214 18510 37266
rect 18562 37214 18574 37266
rect 8598 37154 8650 37166
rect 8598 37090 8650 37102
rect 9718 37154 9770 37166
rect 9718 37090 9770 37102
rect 11286 37154 11338 37166
rect 16718 37202 16770 37214
rect 18902 37210 18954 37222
rect 12114 37102 12126 37154
rect 12178 37102 12190 37154
rect 13190 37146 13242 37158
rect 15206 37154 15258 37166
rect 11286 37090 11338 37102
rect 15206 37090 15258 37102
rect 15990 37154 16042 37166
rect 15990 37090 16042 37102
rect 17782 37154 17834 37166
rect 17782 37090 17834 37102
rect 18734 37154 18786 37166
rect 19070 37202 19122 37214
rect 19294 37266 19346 37278
rect 20638 37266 20690 37278
rect 21502 37270 21514 37322
rect 21566 37270 21578 37322
rect 20402 37214 20414 37266
rect 20466 37214 20478 37266
rect 19294 37202 19346 37214
rect 20638 37202 20690 37214
rect 21758 37266 21810 37278
rect 25678 37314 25730 37326
rect 28366 37378 28418 37390
rect 40238 37378 40290 37390
rect 35018 37326 35030 37378
rect 35082 37326 35094 37378
rect 28366 37314 28418 37326
rect 40238 37314 40290 37326
rect 22318 37258 22370 37270
rect 24222 37266 24274 37278
rect 22642 37214 22654 37266
rect 22706 37214 22718 37266
rect 21758 37202 21810 37214
rect 23046 37210 23098 37222
rect 18902 37146 18954 37158
rect 22878 37154 22930 37166
rect 18734 37090 18786 37102
rect 26114 37244 26126 37296
rect 26178 37244 26190 37296
rect 26450 37244 26462 37296
rect 26514 37244 26526 37296
rect 27246 37266 27298 37278
rect 30214 37266 30266 37278
rect 24222 37202 24274 37214
rect 28110 37214 28122 37266
rect 28174 37214 28186 37266
rect 23046 37146 23098 37158
rect 23494 37154 23546 37166
rect 22878 37090 22930 37102
rect 23494 37090 23546 37102
rect 23886 37154 23938 37166
rect 23886 37090 23938 37102
rect 24726 37154 24778 37166
rect 25946 37158 25958 37210
rect 26010 37158 26022 37210
rect 27246 37202 27298 37214
rect 30214 37202 30266 37214
rect 31054 37266 31106 37278
rect 32174 37266 32226 37278
rect 31918 37214 31930 37266
rect 31982 37214 31994 37266
rect 31054 37202 31106 37214
rect 32174 37202 32226 37214
rect 33070 37266 33122 37278
rect 34190 37266 34242 37278
rect 33934 37214 33946 37266
rect 33998 37214 34010 37266
rect 33070 37202 33122 37214
rect 34190 37202 34242 37214
rect 34638 37266 34690 37278
rect 34638 37202 34690 37214
rect 34750 37266 34802 37278
rect 34750 37202 34802 37214
rect 35310 37266 35362 37278
rect 35310 37202 35362 37214
rect 37048 37266 37100 37278
rect 37326 37266 37378 37278
rect 37202 37214 37214 37266
rect 37266 37214 37278 37266
rect 37048 37202 37100 37214
rect 37326 37202 37378 37214
rect 37550 37266 37602 37278
rect 41582 37266 41634 37278
rect 38322 37214 38334 37266
rect 38386 37214 38398 37266
rect 37550 37202 37602 37214
rect 41582 37202 41634 37214
rect 42254 37266 42306 37278
rect 42254 37202 42306 37214
rect 42926 37266 42978 37278
rect 42926 37202 42978 37214
rect 43710 37266 43762 37278
rect 44258 37229 44270 37281
rect 44322 37229 44334 37281
rect 45166 37266 45218 37278
rect 44594 37214 44606 37266
rect 44658 37214 44670 37266
rect 43710 37202 43762 37214
rect 45166 37202 45218 37214
rect 45390 37266 45442 37278
rect 46218 37270 46230 37322
rect 46282 37270 46294 37322
rect 46734 37266 46786 37278
rect 46386 37214 46398 37266
rect 46450 37214 46462 37266
rect 45390 37202 45442 37214
rect 46734 37202 46786 37214
rect 46958 37266 47010 37278
rect 47518 37266 47570 37278
rect 47226 37214 47238 37266
rect 47290 37214 47302 37266
rect 46958 37202 47010 37214
rect 47518 37202 47570 37214
rect 47742 37266 47794 37278
rect 47742 37202 47794 37214
rect 24726 37090 24778 37102
rect 28982 37154 29034 37166
rect 28982 37090 29034 37102
rect 29766 37154 29818 37166
rect 29766 37090 29818 37102
rect 36262 37154 36314 37166
rect 36262 37090 36314 37102
rect 36654 37154 36706 37166
rect 44146 37102 44158 37154
rect 44210 37102 44222 37154
rect 46050 37102 46062 37154
rect 46114 37102 46126 37154
rect 36654 37090 36706 37102
rect 42590 37042 42642 37054
rect 19562 36990 19574 37042
rect 19626 36990 19638 37042
rect 45658 36990 45670 37042
rect 45722 36990 45734 37042
rect 48010 36990 48022 37042
rect 48074 36990 48086 37042
rect 42590 36978 42642 36990
rect 1344 36874 48608 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 48608 36874
rect 1344 36788 48608 36822
rect 18846 36706 18898 36718
rect 28478 36706 28530 36718
rect 10490 36654 10502 36706
rect 10554 36654 10566 36706
rect 4398 36594 4450 36606
rect 4398 36530 4450 36542
rect 5798 36594 5850 36606
rect 5798 36530 5850 36542
rect 6246 36594 6298 36606
rect 6246 36530 6298 36542
rect 8150 36594 8202 36606
rect 13570 36598 13582 36650
rect 13634 36598 13646 36650
rect 18846 36642 18898 36654
rect 20302 36650 20354 36662
rect 22474 36654 22486 36706
rect 22538 36654 22550 36706
rect 14422 36594 14474 36606
rect 28478 36642 28530 36654
rect 30382 36706 30434 36718
rect 30382 36642 30434 36654
rect 32286 36706 32338 36718
rect 40294 36706 40346 36718
rect 32286 36642 32338 36654
rect 34302 36650 34354 36662
rect 12674 36542 12686 36594
rect 12738 36542 12750 36594
rect 16370 36542 16382 36594
rect 16434 36542 16446 36594
rect 20302 36586 20354 36598
rect 32846 36594 32898 36606
rect 23650 36542 23662 36594
rect 23714 36542 23726 36594
rect 25554 36542 25566 36594
rect 25618 36542 25630 36594
rect 40294 36642 40346 36654
rect 41526 36706 41578 36718
rect 41526 36642 41578 36654
rect 34302 36586 34354 36598
rect 42870 36594 42922 36606
rect 8150 36530 8202 36542
rect 14422 36530 14474 36542
rect 2606 36482 2658 36494
rect 2606 36418 2658 36430
rect 3502 36482 3554 36494
rect 3502 36418 3554 36430
rect 3614 36482 3666 36494
rect 4230 36482 4282 36494
rect 6974 36482 7026 36494
rect 7534 36482 7586 36494
rect 3882 36430 3894 36482
rect 3946 36430 3958 36482
rect 4610 36430 4622 36482
rect 4674 36430 4686 36482
rect 3614 36418 3666 36430
rect 4230 36418 4282 36430
rect 4958 36426 5010 36438
rect 7242 36430 7254 36482
rect 7306 36430 7318 36482
rect 6974 36418 7026 36430
rect 7534 36418 7586 36430
rect 7758 36482 7810 36494
rect 7758 36418 7810 36430
rect 8430 36482 8482 36494
rect 8430 36418 8482 36430
rect 9550 36482 9602 36494
rect 10782 36482 10834 36494
rect 9874 36430 9886 36482
rect 9938 36430 9950 36482
rect 9294 36374 9306 36426
rect 9358 36374 9370 36426
rect 9550 36418 9602 36430
rect 10782 36418 10834 36430
rect 10894 36482 10946 36494
rect 12238 36482 12290 36494
rect 15486 36482 15538 36494
rect 11442 36430 11454 36482
rect 11506 36430 11518 36482
rect 11778 36430 11790 36482
rect 11842 36430 11854 36482
rect 12562 36430 12574 36482
rect 12626 36430 12638 36482
rect 13570 36430 13582 36482
rect 13634 36430 13646 36482
rect 13794 36430 13806 36482
rect 13858 36430 13870 36482
rect 10894 36418 10946 36430
rect 12238 36418 12290 36430
rect 15486 36418 15538 36430
rect 15598 36482 15650 36494
rect 15598 36418 15650 36430
rect 19966 36482 20018 36494
rect 21646 36482 21698 36494
rect 20402 36430 20414 36482
rect 20466 36430 20478 36482
rect 20738 36430 20750 36482
rect 20802 36430 20814 36482
rect 21354 36430 21366 36482
rect 21418 36430 21430 36482
rect 4958 36362 5010 36374
rect 18286 36370 18338 36382
rect 19077 36374 19089 36426
rect 19141 36374 19153 36426
rect 19966 36418 20018 36430
rect 21646 36418 21698 36430
rect 21870 36482 21922 36494
rect 21870 36418 21922 36430
rect 21982 36482 22034 36494
rect 21982 36418 22034 36430
rect 22206 36482 22258 36494
rect 22206 36418 22258 36430
rect 22878 36482 22930 36494
rect 22878 36418 22930 36430
rect 26014 36482 26066 36494
rect 29262 36482 29314 36494
rect 31994 36486 32006 36538
rect 32058 36486 32070 36538
rect 32846 36530 32898 36542
rect 35366 36538 35418 36550
rect 33518 36482 33570 36494
rect 35198 36482 35250 36494
rect 26878 36430 26890 36482
rect 26942 36430 26954 36482
rect 26014 36418 26066 36430
rect 28198 36426 28250 36438
rect 18286 36306 18338 36318
rect 27134 36370 27186 36382
rect 27682 36374 27694 36426
rect 27746 36374 27758 36426
rect 27906 36374 27918 36426
rect 27970 36374 27982 36426
rect 30126 36430 30138 36482
rect 30190 36430 30202 36482
rect 29262 36418 29314 36430
rect 31490 36400 31502 36452
rect 31554 36400 31566 36452
rect 33394 36430 33406 36482
rect 33458 36430 33470 36482
rect 33842 36430 33854 36482
rect 33906 36430 33918 36482
rect 34178 36430 34190 36482
rect 34242 36430 34254 36482
rect 46162 36542 46174 36594
rect 46226 36542 46238 36594
rect 42870 36530 42922 36542
rect 35366 36474 35418 36486
rect 35646 36482 35698 36494
rect 31714 36374 31726 36426
rect 31778 36374 31790 36426
rect 33228 36374 33240 36426
rect 33292 36374 33304 36426
rect 33518 36418 33570 36430
rect 35198 36418 35250 36430
rect 35646 36418 35698 36430
rect 36878 36482 36930 36494
rect 39566 36482 39618 36494
rect 37650 36430 37662 36482
rect 37714 36430 37726 36482
rect 44718 36482 44770 36494
rect 36878 36418 36930 36430
rect 39566 36418 39618 36430
rect 40574 36454 40626 36466
rect 41134 36447 41186 36459
rect 40574 36390 40626 36402
rect 28198 36362 28250 36374
rect 34918 36370 34970 36382
rect 27134 36306 27186 36318
rect 34918 36306 34970 36318
rect 35534 36370 35586 36382
rect 35534 36306 35586 36318
rect 35926 36370 35978 36382
rect 40786 36374 40798 36426
rect 40850 36374 40862 36426
rect 41010 36374 41022 36426
rect 41074 36374 41086 36426
rect 41134 36383 41186 36395
rect 41806 36454 41858 36466
rect 41806 36390 41858 36402
rect 42030 36454 42082 36466
rect 42030 36390 42082 36402
rect 42254 36454 42306 36466
rect 43486 36454 43538 36466
rect 42254 36390 42306 36402
rect 42366 36426 42418 36438
rect 44046 36447 44098 36459
rect 43486 36390 43538 36402
rect 42366 36362 42418 36374
rect 43206 36370 43258 36382
rect 43698 36374 43710 36426
rect 43762 36374 43774 36426
rect 43922 36374 43934 36426
rect 43986 36374 43998 36426
rect 44718 36418 44770 36430
rect 45390 36482 45442 36494
rect 45390 36418 45442 36430
rect 44046 36383 44098 36395
rect 35926 36306 35978 36318
rect 43206 36306 43258 36318
rect 48078 36370 48130 36382
rect 48078 36306 48130 36318
rect 2270 36258 2322 36270
rect 2270 36194 2322 36206
rect 6638 36258 6690 36270
rect 6638 36194 6690 36206
rect 10054 36258 10106 36270
rect 10054 36194 10106 36206
rect 15150 36258 15202 36270
rect 15150 36194 15202 36206
rect 31110 36258 31162 36270
rect 31110 36194 31162 36206
rect 36486 36258 36538 36270
rect 36486 36194 36538 36206
rect 45054 36258 45106 36270
rect 45054 36194 45106 36206
rect 1344 36090 48608 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 48608 36090
rect 1344 36004 48608 36038
rect 5910 35922 5962 35934
rect 5910 35858 5962 35870
rect 21030 35922 21082 35934
rect 21030 35858 21082 35870
rect 30438 35922 30490 35934
rect 30438 35858 30490 35870
rect 32566 35922 32618 35934
rect 32566 35858 32618 35870
rect 40294 35922 40346 35934
rect 5406 35810 5458 35822
rect 8878 35810 8930 35822
rect 4846 35736 4898 35748
rect 5406 35746 5458 35758
rect 5574 35754 5626 35766
rect 1598 35698 1650 35710
rect 2370 35646 2382 35698
rect 2434 35646 2446 35698
rect 10446 35810 10498 35822
rect 19742 35810 19794 35822
rect 8878 35746 8930 35758
rect 9494 35754 9546 35766
rect 4846 35672 4898 35684
rect 5170 35646 5182 35698
rect 5234 35646 5246 35698
rect 5574 35690 5626 35702
rect 6078 35718 6130 35730
rect 6234 35672 6246 35724
rect 6298 35672 6310 35724
rect 18442 35758 18454 35810
rect 18506 35758 18518 35810
rect 10446 35746 10498 35758
rect 18790 35754 18842 35766
rect 6078 35654 6130 35666
rect 6962 35646 6974 35698
rect 7026 35646 7038 35698
rect 9494 35690 9546 35702
rect 9650 35676 9662 35728
rect 9714 35676 9726 35728
rect 9874 35685 9886 35737
rect 9938 35685 9950 35737
rect 11006 35698 11058 35710
rect 12126 35698 12178 35710
rect 11870 35646 11882 35698
rect 11934 35646 11946 35698
rect 1598 35634 1650 35646
rect 11006 35634 11058 35646
rect 12126 35634 12178 35646
rect 12574 35698 12626 35710
rect 14030 35698 14082 35710
rect 17838 35698 17890 35710
rect 13438 35646 13450 35698
rect 13502 35646 13514 35698
rect 14802 35646 14814 35698
rect 14866 35646 14878 35698
rect 12574 35634 12626 35646
rect 14030 35634 14082 35646
rect 17838 35634 17890 35646
rect 17950 35698 18002 35710
rect 17950 35634 18002 35646
rect 18174 35698 18226 35710
rect 19002 35702 19014 35754
rect 19066 35702 19078 35754
rect 19742 35746 19794 35758
rect 26686 35810 26738 35822
rect 26686 35746 26738 35758
rect 29038 35810 29090 35822
rect 29038 35746 29090 35758
rect 31838 35810 31890 35822
rect 33394 35814 33406 35866
rect 33458 35814 33470 35866
rect 40294 35858 40346 35870
rect 41806 35922 41858 35934
rect 41806 35858 41858 35870
rect 42478 35922 42530 35934
rect 42478 35858 42530 35870
rect 35422 35810 35474 35822
rect 46274 35814 46286 35866
rect 46338 35814 46350 35866
rect 34570 35758 34582 35810
rect 34634 35758 34646 35810
rect 31838 35746 31890 35758
rect 35422 35746 35474 35758
rect 36374 35754 36426 35766
rect 38602 35758 38614 35810
rect 38666 35758 38678 35810
rect 44426 35758 44438 35810
rect 44490 35758 44502 35810
rect 18790 35690 18842 35702
rect 19170 35685 19182 35737
rect 19234 35685 19246 35737
rect 20470 35727 20522 35739
rect 20178 35646 20190 35698
rect 20242 35646 20254 35698
rect 21758 35698 21810 35710
rect 20470 35663 20522 35675
rect 20850 35646 20862 35698
rect 20914 35646 20926 35698
rect 25330 35676 25342 35728
rect 25394 35676 25406 35728
rect 25666 35676 25678 35728
rect 25730 35676 25742 35728
rect 26126 35698 26178 35710
rect 18174 35634 18226 35646
rect 21758 35634 21810 35646
rect 13694 35586 13746 35598
rect 21590 35586 21642 35598
rect 25834 35590 25846 35642
rect 25898 35590 25910 35642
rect 26126 35634 26178 35646
rect 26518 35642 26570 35654
rect 26898 35646 26910 35698
rect 26962 35646 26974 35698
rect 27122 35674 27134 35726
rect 27186 35674 27198 35726
rect 27918 35698 27970 35710
rect 30718 35698 30770 35710
rect 33854 35698 33906 35710
rect 28782 35646 28794 35698
rect 28846 35646 28858 35698
rect 31582 35646 31594 35698
rect 31646 35646 31658 35698
rect 33170 35646 33182 35698
rect 33234 35646 33246 35698
rect 27918 35634 27970 35646
rect 30718 35634 30770 35646
rect 33854 35634 33906 35646
rect 34078 35698 34130 35710
rect 34078 35634 34130 35646
rect 34302 35698 34354 35710
rect 35858 35676 35870 35728
rect 35922 35676 35934 35728
rect 36082 35684 36094 35736
rect 36146 35684 36158 35736
rect 36374 35690 36426 35702
rect 36654 35698 36706 35710
rect 34302 35634 34354 35646
rect 36654 35634 36706 35646
rect 36766 35698 36818 35710
rect 36766 35634 36818 35646
rect 37438 35698 37490 35710
rect 37718 35698 37770 35710
rect 37538 35646 37550 35698
rect 37602 35646 37614 35698
rect 37438 35634 37490 35646
rect 37718 35634 37770 35646
rect 38894 35698 38946 35710
rect 38894 35634 38946 35646
rect 39118 35698 39170 35710
rect 39118 35634 39170 35646
rect 39342 35698 39394 35710
rect 39342 35634 39394 35646
rect 39454 35698 39506 35710
rect 40798 35698 40850 35710
rect 39722 35646 39734 35698
rect 39786 35646 39798 35698
rect 39454 35634 39506 35646
rect 40798 35634 40850 35646
rect 41470 35698 41522 35710
rect 41470 35634 41522 35646
rect 42142 35698 42194 35710
rect 42142 35634 42194 35646
rect 43374 35698 43426 35710
rect 43374 35634 43426 35646
rect 44046 35698 44098 35710
rect 44046 35634 44098 35646
rect 44718 35698 44770 35710
rect 44718 35634 44770 35646
rect 44830 35698 44882 35710
rect 44830 35634 44882 35646
rect 45166 35698 45218 35710
rect 45378 35702 45390 35754
rect 45442 35702 45454 35754
rect 46622 35737 46674 35749
rect 46274 35646 46286 35698
rect 46338 35646 46350 35698
rect 46622 35673 46674 35685
rect 46846 35698 46898 35710
rect 47394 35646 47406 35698
rect 47458 35646 47470 35698
rect 47730 35690 47742 35742
rect 47794 35690 47806 35742
rect 45166 35634 45218 35646
rect 46846 35634 46898 35646
rect 4274 35534 4286 35586
rect 4338 35534 4350 35586
rect 16706 35534 16718 35586
rect 16770 35534 16782 35586
rect 20626 35534 20638 35586
rect 20690 35534 20702 35586
rect 22530 35534 22542 35586
rect 22594 35534 22606 35586
rect 24434 35534 24446 35586
rect 24498 35534 24510 35586
rect 26518 35578 26570 35590
rect 29990 35586 30042 35598
rect 13694 35522 13746 35534
rect 21590 35522 21642 35534
rect 29990 35522 30042 35534
rect 38110 35586 38162 35598
rect 38110 35522 38162 35534
rect 43710 35586 43762 35598
rect 47842 35534 47854 35586
rect 47906 35534 47918 35586
rect 43710 35522 43762 35534
rect 17502 35474 17554 35486
rect 41134 35474 41186 35486
rect 37034 35422 37046 35474
rect 37098 35422 37110 35474
rect 17502 35410 17554 35422
rect 41134 35410 41186 35422
rect 43038 35474 43090 35486
rect 45658 35422 45670 35474
rect 45722 35422 45734 35474
rect 43038 35410 43090 35422
rect 1344 35306 48608 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 48608 35306
rect 1344 35220 48608 35254
rect 12798 35138 12850 35150
rect 2650 35086 2662 35138
rect 2714 35086 2726 35138
rect 8138 35086 8150 35138
rect 8202 35086 8214 35138
rect 12798 35074 12850 35086
rect 15150 35138 15202 35150
rect 15150 35074 15202 35086
rect 19630 35138 19682 35150
rect 23326 35138 23378 35150
rect 19630 35074 19682 35086
rect 21646 35082 21698 35094
rect 6694 35026 6746 35038
rect 6694 34962 6746 34974
rect 7086 35026 7138 35038
rect 23326 35074 23378 35086
rect 28478 35138 28530 35150
rect 28478 35074 28530 35086
rect 30270 35138 30322 35150
rect 30270 35074 30322 35086
rect 32734 35138 32786 35150
rect 32734 35074 32786 35086
rect 42422 35138 42474 35150
rect 42422 35074 42474 35086
rect 45726 35138 45778 35150
rect 45726 35074 45778 35086
rect 46398 35138 46450 35150
rect 48122 35086 48134 35138
rect 48186 35086 48198 35138
rect 46398 35074 46450 35086
rect 21646 35018 21698 35030
rect 37662 35026 37714 35038
rect 7086 34962 7138 34974
rect 38278 35026 38330 35038
rect 44942 35026 44994 35038
rect 2942 34914 2994 34926
rect 2942 34850 2994 34862
rect 3166 34914 3218 34926
rect 3166 34850 3218 34862
rect 3390 34914 3442 34926
rect 4510 34914 4562 34926
rect 5966 34914 6018 34926
rect 4254 34862 4266 34914
rect 4318 34862 4330 34914
rect 5170 34862 5182 34914
rect 5234 34862 5246 34914
rect 3390 34850 3442 34862
rect 4510 34850 4562 34862
rect 5966 34850 6018 34862
rect 6190 34914 6242 34926
rect 8430 34914 8482 34926
rect 6190 34850 6242 34862
rect 6918 34858 6970 34870
rect 7298 34862 7310 34914
rect 7362 34862 7374 34914
rect 7522 34806 7534 34858
rect 7586 34806 7598 34858
rect 8430 34850 8482 34862
rect 8654 34914 8706 34926
rect 8654 34850 8706 34862
rect 9214 34914 9266 34926
rect 10334 34914 10386 34926
rect 9445 34862 9457 34914
rect 9509 34862 9521 34914
rect 9214 34850 9266 34862
rect 10334 34850 10386 34862
rect 10782 34914 10834 34926
rect 10782 34850 10834 34862
rect 11006 34914 11058 34926
rect 12506 34918 12518 34970
rect 12570 34918 12582 34970
rect 11006 34850 11058 34862
rect 14030 34914 14082 34926
rect 12002 34806 12014 34858
rect 12066 34806 12078 34858
rect 12338 34806 12350 34858
rect 12402 34806 12414 34858
rect 14030 34850 14082 34862
rect 16046 34914 16098 34926
rect 14894 34806 14906 34858
rect 14958 34806 14970 34858
rect 16046 34850 16098 34862
rect 16270 34914 16322 34926
rect 16270 34850 16322 34862
rect 16494 34914 16546 34926
rect 19070 34914 19122 34926
rect 16494 34850 16546 34862
rect 17222 34858 17274 34870
rect 17490 34806 17502 34858
rect 17554 34806 17566 34858
rect 17770 34806 17782 34858
rect 17834 34806 17846 34858
rect 19070 34850 19122 34862
rect 19294 34914 19346 34926
rect 19294 34850 19346 34862
rect 20750 34914 20802 34926
rect 22878 34914 22930 34926
rect 21746 34862 21758 34914
rect 21810 34862 21822 34914
rect 21970 34862 21982 34914
rect 22034 34862 22046 34914
rect 5674 34750 5686 34802
rect 5738 34750 5750 34802
rect 6918 34794 6970 34806
rect 11274 34750 11286 34802
rect 11338 34750 11350 34802
rect 16762 34750 16774 34802
rect 16826 34750 16838 34802
rect 17222 34794 17274 34806
rect 18174 34802 18226 34814
rect 19861 34806 19873 34858
rect 19925 34806 19937 34858
rect 20750 34850 20802 34862
rect 22878 34850 22930 34862
rect 22990 34914 23042 34926
rect 24558 34914 24610 34926
rect 26898 34918 26910 34970
rect 26962 34918 26974 34970
rect 37662 34962 37714 34974
rect 37830 34970 37882 34982
rect 24322 34862 24334 34914
rect 24386 34862 24398 34914
rect 29150 34914 29202 34926
rect 33070 34914 33122 34926
rect 35758 34914 35810 34926
rect 39218 34974 39230 35026
rect 39282 34974 39294 35026
rect 41122 34974 41134 35026
rect 41186 34974 41198 35026
rect 38278 34962 38330 34974
rect 44942 34962 44994 34974
rect 22990 34850 23042 34862
rect 24558 34850 24610 34862
rect 25422 34831 25434 34883
rect 25486 34831 25498 34883
rect 26070 34858 26122 34870
rect 25678 34802 25730 34814
rect 18778 34750 18790 34802
rect 18842 34750 18854 34802
rect 26798 34858 26850 34870
rect 26070 34794 26122 34806
rect 26238 34802 26290 34814
rect 18174 34738 18226 34750
rect 25678 34738 25730 34750
rect 26798 34794 26850 34806
rect 27526 34858 27578 34870
rect 27794 34806 27806 34858
rect 27858 34806 27870 34858
rect 28018 34832 28030 34884
rect 28082 34832 28094 34884
rect 30014 34862 30026 34914
rect 30078 34862 30090 34914
rect 29150 34850 29202 34862
rect 31782 34858 31834 34870
rect 33842 34862 33854 34914
rect 33906 34862 33918 34914
rect 36082 34862 36094 34914
rect 36146 34862 36158 34914
rect 37830 34906 37882 34918
rect 38446 34914 38498 34926
rect 27526 34794 27578 34806
rect 31558 34802 31610 34814
rect 26238 34738 26290 34750
rect 31938 34806 31950 34858
rect 32002 34806 32014 34858
rect 32274 34806 32286 34858
rect 32338 34806 32350 34858
rect 33070 34850 33122 34862
rect 35758 34850 35810 34862
rect 36990 34858 37042 34870
rect 31782 34794 31834 34806
rect 36990 34794 37042 34806
rect 37102 34858 37154 34870
rect 42926 34914 42978 34926
rect 38446 34850 38498 34862
rect 41514 34846 41526 34898
rect 41578 34846 41590 34898
rect 41694 34886 41746 34898
rect 41694 34822 41746 34834
rect 41918 34886 41970 34898
rect 41918 34822 41970 34834
rect 42142 34886 42194 34898
rect 42926 34850 42978 34862
rect 43150 34914 43202 34926
rect 43710 34914 43762 34926
rect 43418 34862 43430 34914
rect 43482 34862 43494 34914
rect 43150 34850 43202 34862
rect 43710 34850 43762 34862
rect 45278 34914 45330 34926
rect 45278 34850 45330 34862
rect 45390 34914 45442 34926
rect 45390 34850 45442 34862
rect 46062 34914 46114 34926
rect 46062 34850 46114 34862
rect 47294 34914 47346 34926
rect 47294 34850 47346 34862
rect 47518 34914 47570 34926
rect 47518 34850 47570 34862
rect 47630 34914 47682 34926
rect 47630 34850 47682 34862
rect 47854 34914 47906 34926
rect 47854 34850 47906 34862
rect 42142 34822 42194 34834
rect 37102 34794 37154 34806
rect 47002 34750 47014 34802
rect 47066 34750 47078 34802
rect 31558 34738 31610 34750
rect 5014 34690 5066 34702
rect 5014 34626 5066 34638
rect 13750 34690 13802 34702
rect 13750 34626 13802 34638
rect 15710 34690 15762 34702
rect 15710 34626 15762 34638
rect 22542 34690 22594 34702
rect 22542 34626 22594 34638
rect 24166 34690 24218 34702
rect 24166 34626 24218 34638
rect 31110 34690 31162 34702
rect 31110 34626 31162 34638
rect 36262 34690 36314 34702
rect 36262 34626 36314 34638
rect 44046 34690 44098 34702
rect 44046 34626 44098 34638
rect 1344 34522 48608 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 48608 34522
rect 1344 34436 48608 34470
rect 8094 34354 8146 34366
rect 8094 34290 8146 34302
rect 9662 34354 9714 34366
rect 9662 34290 9714 34302
rect 36990 34354 37042 34366
rect 36990 34290 37042 34302
rect 41806 34354 41858 34366
rect 41806 34290 41858 34302
rect 4846 34242 4898 34254
rect 3894 34186 3946 34198
rect 5742 34242 5794 34254
rect 10894 34242 10946 34254
rect 14646 34242 14698 34254
rect 4050 34134 4062 34186
rect 4114 34134 4126 34186
rect 4274 34134 4286 34186
rect 4338 34134 4350 34186
rect 4846 34178 4898 34190
rect 5574 34186 5626 34198
rect 5742 34178 5794 34190
rect 6302 34186 6354 34198
rect 7130 34190 7142 34242
rect 7194 34190 7206 34242
rect 12954 34190 12966 34242
rect 13018 34190 13030 34242
rect 3894 34122 3946 34134
rect 5574 34122 5626 34134
rect 10334 34168 10386 34180
rect 10894 34178 10946 34190
rect 14646 34178 14698 34190
rect 22598 34242 22650 34254
rect 5954 34078 5966 34130
rect 6018 34078 6030 34130
rect 6302 34122 6354 34134
rect 6638 34130 6690 34142
rect 6638 34066 6690 34078
rect 6862 34130 6914 34142
rect 6862 34066 6914 34078
rect 8430 34130 8482 34142
rect 8430 34066 8482 34078
rect 9102 34130 9154 34142
rect 9102 34066 9154 34078
rect 9998 34130 10050 34142
rect 12462 34130 12514 34142
rect 10334 34104 10386 34116
rect 9998 34066 10050 34078
rect 11062 34074 11114 34086
rect 11330 34078 11342 34130
rect 11394 34078 11406 34130
rect 3670 34018 3722 34030
rect 3670 33954 3722 33966
rect 7702 34018 7754 34030
rect 10210 34022 10222 34074
rect 10274 34022 10286 34074
rect 12462 34066 12514 34078
rect 12686 34130 12738 34142
rect 12686 34066 12738 34078
rect 13918 34130 13970 34142
rect 14366 34130 14418 34142
rect 13918 34066 13970 34078
rect 14086 34074 14138 34086
rect 14242 34078 14254 34130
rect 14306 34078 14318 34130
rect 11062 34010 11114 34022
rect 13638 34018 13690 34030
rect 7702 33954 7754 33966
rect 14366 34066 14418 34078
rect 14926 34130 14978 34142
rect 14926 34066 14978 34078
rect 15150 34130 15202 34142
rect 16930 34078 16942 34130
rect 16994 34078 17006 34130
rect 17266 34078 17278 34130
rect 17330 34078 17342 34130
rect 18050 34078 18062 34130
rect 18114 34078 18126 34130
rect 19954 34105 19966 34157
rect 20018 34105 20030 34157
rect 20570 34094 20582 34146
rect 20634 34094 20646 34146
rect 20738 34134 20750 34186
rect 20802 34134 20814 34186
rect 20974 34158 21026 34170
rect 21186 34134 21198 34186
rect 21250 34134 21262 34186
rect 22598 34178 22650 34190
rect 28366 34242 28418 34254
rect 28366 34178 28418 34190
rect 30326 34242 30378 34254
rect 30326 34178 30378 34190
rect 45278 34242 45330 34254
rect 46386 34246 46398 34298
rect 46450 34246 46462 34298
rect 20974 34094 21026 34106
rect 21478 34130 21530 34142
rect 15150 34066 15202 34078
rect 21478 34066 21530 34078
rect 21870 34130 21922 34142
rect 22318 34130 22370 34142
rect 21870 34066 21922 34078
rect 22038 34074 22090 34086
rect 22194 34078 22206 34130
rect 22258 34078 22270 34130
rect 14086 34010 14138 34022
rect 22318 34066 22370 34078
rect 23662 34130 23714 34142
rect 23662 34066 23714 34078
rect 23774 34130 23826 34142
rect 23774 34066 23826 34078
rect 23998 34130 24050 34142
rect 26798 34130 26850 34142
rect 25666 34078 25678 34130
rect 25730 34078 25742 34130
rect 26002 34078 26014 34130
rect 26066 34078 26078 34130
rect 26506 34078 26518 34130
rect 26570 34078 26582 34130
rect 23998 34066 24050 34078
rect 26798 34066 26850 34078
rect 26910 34130 26962 34142
rect 26910 34066 26962 34078
rect 27246 34130 27298 34142
rect 29598 34130 29650 34142
rect 28110 34078 28122 34130
rect 28174 34078 28186 34130
rect 27246 34066 27298 34078
rect 29598 34066 29650 34078
rect 29766 34130 29818 34142
rect 30046 34130 30098 34142
rect 29922 34078 29934 34130
rect 29986 34078 29998 34130
rect 29766 34066 29818 34078
rect 30046 34066 30098 34078
rect 30718 34130 30770 34142
rect 31838 34130 31890 34142
rect 31582 34078 31594 34130
rect 31646 34078 31658 34130
rect 30718 34066 30770 34078
rect 31838 34066 31890 34078
rect 33070 34130 33122 34142
rect 33934 34134 33946 34186
rect 33998 34134 34010 34186
rect 45278 34178 45330 34190
rect 33070 34066 33122 34078
rect 34526 34130 34578 34142
rect 36542 34130 36594 34142
rect 35653 34078 35665 34130
rect 35717 34078 35729 34130
rect 34526 34066 34578 34078
rect 36542 34066 36594 34078
rect 37326 34130 37378 34142
rect 39230 34130 39282 34142
rect 37426 34078 37438 34130
rect 37490 34078 37502 34130
rect 38938 34078 38950 34130
rect 39002 34078 39014 34130
rect 37326 34066 37378 34078
rect 39230 34066 39282 34078
rect 39454 34130 39506 34142
rect 39454 34066 39506 34078
rect 39678 34130 39730 34142
rect 39678 34066 39730 34078
rect 39790 34130 39842 34142
rect 40798 34130 40850 34142
rect 40058 34078 40070 34130
rect 40122 34078 40134 34130
rect 39790 34066 39842 34078
rect 40798 34066 40850 34078
rect 41470 34130 41522 34142
rect 41470 34066 41522 34078
rect 42590 34130 42642 34142
rect 46510 34130 46562 34142
rect 43362 34078 43374 34130
rect 43426 34078 43438 34130
rect 46834 34105 46846 34157
rect 46898 34105 46910 34157
rect 47170 34078 47182 34130
rect 47234 34078 47246 34130
rect 47618 34122 47630 34174
rect 47682 34122 47694 34174
rect 47842 34078 47854 34130
rect 47906 34078 47918 34130
rect 42590 34066 42642 34078
rect 46510 34066 46562 34078
rect 22038 34010 22090 34022
rect 25398 34018 25450 34030
rect 13638 33954 13690 33966
rect 25398 33954 25450 33966
rect 28982 34018 29034 34030
rect 8766 33906 8818 33918
rect 17446 33906 17498 33918
rect 15418 33854 15430 33906
rect 15482 33854 15494 33906
rect 8766 33842 8818 33854
rect 17446 33842 17498 33854
rect 23326 33906 23378 33918
rect 25890 33910 25902 33962
rect 25954 33910 25966 33962
rect 28982 33954 29034 33966
rect 32566 34018 32618 34030
rect 32566 33954 32618 33966
rect 42422 34018 42474 34030
rect 42422 33954 42474 33966
rect 45894 34018 45946 34030
rect 47506 33966 47518 34018
rect 47570 33966 47582 34018
rect 45894 33954 45946 33966
rect 34190 33906 34242 33918
rect 24266 33854 24278 33906
rect 24330 33854 24342 33906
rect 23326 33842 23378 33854
rect 34190 33842 34242 33854
rect 34862 33906 34914 33918
rect 34862 33842 34914 33854
rect 35422 33906 35474 33918
rect 35422 33842 35474 33854
rect 41134 33906 41186 33918
rect 41134 33842 41186 33854
rect 1344 33738 48608 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 48608 33738
rect 1344 33652 48608 33686
rect 27358 33570 27410 33582
rect 31166 33570 31218 33582
rect 12842 33518 12854 33570
rect 12906 33518 12918 33570
rect 15822 33514 15874 33526
rect 29642 33518 29654 33570
rect 29706 33518 29718 33570
rect 34190 33570 34242 33582
rect 27358 33506 27410 33518
rect 31166 33506 31218 33518
rect 32454 33514 32506 33526
rect 9986 33406 9998 33458
rect 10050 33406 10062 33458
rect 13570 33406 13582 33458
rect 13634 33406 13646 33458
rect 15822 33450 15874 33462
rect 16942 33458 16994 33470
rect 1598 33346 1650 33358
rect 5126 33346 5178 33358
rect 2370 33294 2382 33346
rect 2434 33294 2446 33346
rect 6190 33346 6242 33358
rect 9214 33346 9266 33358
rect 1598 33282 1650 33294
rect 5126 33282 5178 33294
rect 6078 33290 6130 33302
rect 4286 33234 4338 33246
rect 6962 33294 6974 33346
rect 7026 33294 7038 33346
rect 6190 33282 6242 33294
rect 9214 33282 9266 33294
rect 12462 33346 12514 33358
rect 12462 33282 12514 33294
rect 12574 33346 12626 33358
rect 16258 33350 16270 33402
rect 16322 33350 16334 33402
rect 16942 33394 16994 33406
rect 18510 33458 18562 33470
rect 18510 33394 18562 33406
rect 19742 33458 19794 33470
rect 25006 33458 25058 33470
rect 22530 33406 22542 33458
rect 22594 33406 22606 33458
rect 19742 33394 19794 33406
rect 25006 33394 25058 33406
rect 26966 33458 27018 33470
rect 34682 33518 34694 33570
rect 34746 33518 34758 33570
rect 42298 33518 42310 33570
rect 42362 33518 42374 33570
rect 34190 33506 34242 33518
rect 43486 33514 43538 33526
rect 32454 33450 32506 33462
rect 43922 33462 43934 33514
rect 43986 33462 43998 33514
rect 38882 33406 38894 33458
rect 38946 33406 38958 33458
rect 40786 33406 40798 33458
rect 40850 33406 40862 33458
rect 43486 33450 43538 33462
rect 48066 33406 48078 33458
rect 48130 33406 48142 33458
rect 26966 33394 27018 33406
rect 17390 33346 17442 33358
rect 12574 33282 12626 33294
rect 13638 33254 13650 33306
rect 13702 33254 13714 33306
rect 13794 33257 13806 33309
rect 13858 33257 13870 33309
rect 6078 33226 6130 33238
rect 8878 33234 8930 33246
rect 4286 33170 4338 33182
rect 8878 33170 8930 33182
rect 11902 33234 11954 33246
rect 14242 33238 14254 33290
rect 14306 33238 14318 33290
rect 14578 33261 14590 33313
rect 14642 33261 14654 33313
rect 15022 33256 15034 33308
rect 15086 33256 15098 33308
rect 15698 33294 15710 33346
rect 15762 33294 15774 33346
rect 17110 33290 17162 33302
rect 16482 33238 16494 33290
rect 16546 33238 16558 33290
rect 19406 33346 19458 33358
rect 21758 33346 21810 33358
rect 29262 33346 29314 33358
rect 17390 33282 17442 33294
rect 18254 33263 18266 33315
rect 18318 33263 18330 33315
rect 19406 33282 19458 33294
rect 19630 33307 19682 33319
rect 20066 33294 20078 33346
rect 20130 33294 20142 33346
rect 21522 33294 21534 33346
rect 21586 33294 21598 33346
rect 21758 33282 21810 33294
rect 24838 33290 24890 33302
rect 25218 33294 25230 33346
rect 25282 33294 25294 33346
rect 19630 33243 19682 33255
rect 17110 33226 17162 33238
rect 24446 33234 24498 33246
rect 11902 33170 11954 33182
rect 21366 33178 21418 33190
rect 5910 33122 5962 33134
rect 5910 33058 5962 33070
rect 20806 33122 20858 33134
rect 25442 33266 25454 33318
rect 25506 33266 25518 33318
rect 27638 33290 27690 33302
rect 24838 33226 24890 33238
rect 27906 33238 27918 33290
rect 27970 33238 27982 33290
rect 28130 33238 28142 33290
rect 28194 33238 28206 33290
rect 29262 33282 29314 33294
rect 29374 33346 29426 33358
rect 29374 33282 29426 33294
rect 30046 33346 30098 33358
rect 31502 33346 31554 33358
rect 30910 33294 30922 33346
rect 30974 33294 30986 33346
rect 30046 33282 30098 33294
rect 31502 33282 31554 33294
rect 31726 33346 31778 33358
rect 33070 33346 33122 33358
rect 34974 33346 35026 33358
rect 31726 33282 31778 33294
rect 32286 33290 32338 33302
rect 33934 33294 33946 33346
rect 33998 33294 34010 33346
rect 33070 33282 33122 33294
rect 34974 33282 35026 33294
rect 35198 33346 35250 33358
rect 36318 33346 36370 33358
rect 35198 33282 35250 33294
rect 35366 33290 35418 33302
rect 27638 33226 27690 33238
rect 31994 33182 32006 33234
rect 32058 33182 32070 33234
rect 32286 33226 32338 33238
rect 35522 33238 35534 33290
rect 35586 33238 35598 33290
rect 35858 33238 35870 33290
rect 35922 33238 35934 33290
rect 36318 33282 36370 33294
rect 36934 33346 36986 33358
rect 38110 33346 38162 33358
rect 37314 33294 37326 33346
rect 37378 33294 37390 33346
rect 36934 33282 36986 33294
rect 37662 33290 37714 33302
rect 35366 33226 35418 33238
rect 37102 33234 37154 33246
rect 38110 33282 38162 33294
rect 41806 33346 41858 33358
rect 41806 33282 41858 33294
rect 41918 33346 41970 33358
rect 41918 33282 41970 33294
rect 42590 33346 42642 33358
rect 42590 33282 42642 33294
rect 42702 33346 42754 33358
rect 44718 33346 44770 33358
rect 43138 33294 43150 33346
rect 43202 33294 43214 33346
rect 43362 33294 43374 33346
rect 43426 33294 43438 33346
rect 43922 33294 43934 33346
rect 43986 33294 43998 33346
rect 44146 33294 44158 33346
rect 44210 33294 44222 33346
rect 42702 33282 42754 33294
rect 44718 33282 44770 33294
rect 45390 33346 45442 33358
rect 46162 33294 46174 33346
rect 46226 33294 46238 33346
rect 45390 33282 45442 33294
rect 37662 33226 37714 33238
rect 41514 33182 41526 33234
rect 41578 33182 41590 33234
rect 24446 33170 24498 33182
rect 37102 33170 37154 33182
rect 21366 33114 21418 33126
rect 26294 33122 26346 33134
rect 20806 33058 20858 33070
rect 26294 33058 26346 33070
rect 45054 33122 45106 33134
rect 45054 33058 45106 33070
rect 1344 32954 48608 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 48608 32954
rect 1344 32868 48608 32902
rect 2270 32786 2322 32798
rect 2270 32722 2322 32734
rect 3222 32786 3274 32798
rect 3222 32722 3274 32734
rect 3670 32786 3722 32798
rect 3670 32722 3722 32734
rect 4118 32786 4170 32798
rect 4118 32722 4170 32734
rect 7198 32786 7250 32798
rect 7198 32722 7250 32734
rect 9774 32786 9826 32798
rect 7858 32678 7870 32730
rect 7922 32678 7934 32730
rect 9774 32722 9826 32734
rect 12798 32786 12850 32798
rect 10770 32678 10782 32730
rect 10834 32678 10846 32730
rect 12798 32722 12850 32734
rect 32566 32786 32618 32798
rect 32566 32722 32618 32734
rect 37438 32786 37490 32798
rect 37438 32722 37490 32734
rect 40126 32786 40178 32798
rect 40126 32722 40178 32734
rect 15150 32674 15202 32686
rect 2606 32562 2658 32574
rect 2606 32498 2658 32510
rect 4398 32562 4450 32574
rect 5966 32562 6018 32574
rect 6244 32562 6296 32574
rect 5262 32510 5274 32562
rect 5326 32510 5338 32562
rect 6066 32510 6078 32562
rect 6130 32510 6142 32562
rect 4398 32498 4450 32510
rect 5966 32498 6018 32510
rect 6244 32498 6296 32510
rect 7534 32562 7586 32574
rect 7858 32510 7870 32562
rect 7922 32510 7934 32562
rect 8082 32537 8094 32589
rect 8146 32537 8158 32589
rect 8430 32562 8482 32574
rect 7534 32498 7586 32510
rect 8430 32498 8482 32510
rect 9438 32562 9490 32574
rect 9438 32498 9490 32510
rect 10334 32562 10386 32574
rect 10882 32510 10894 32562
rect 10946 32510 10958 32562
rect 11666 32537 11678 32589
rect 11730 32537 11742 32589
rect 14354 32566 14366 32618
rect 14418 32566 14430 32618
rect 15150 32610 15202 32622
rect 17502 32674 17554 32686
rect 14578 32549 14590 32601
rect 14642 32549 14654 32601
rect 15941 32566 15953 32618
rect 16005 32566 16017 32618
rect 17502 32610 17554 32622
rect 21198 32674 21250 32686
rect 23550 32674 23602 32686
rect 22698 32622 22710 32674
rect 22762 32622 22774 32674
rect 16830 32562 16882 32574
rect 18050 32549 18062 32601
rect 18114 32549 18126 32601
rect 18274 32566 18286 32618
rect 18338 32566 18350 32618
rect 19394 32566 19406 32618
rect 19458 32566 19470 32618
rect 20178 32566 20190 32618
rect 20242 32566 20254 32618
rect 21198 32610 21250 32622
rect 21858 32566 21870 32618
rect 21922 32566 21934 32618
rect 23550 32610 23602 32622
rect 30382 32674 30434 32686
rect 22990 32562 23042 32574
rect 18610 32510 18622 32562
rect 18674 32510 18686 32562
rect 20738 32510 20750 32562
rect 20802 32510 20814 32562
rect 10334 32498 10386 32510
rect 14858 32454 14870 32506
rect 14922 32454 14934 32506
rect 16830 32498 16882 32510
rect 17770 32454 17782 32506
rect 17834 32454 17846 32506
rect 22990 32498 23042 32510
rect 23214 32562 23266 32574
rect 23781 32541 23793 32593
rect 23845 32541 23857 32593
rect 24670 32562 24722 32574
rect 23214 32498 23266 32510
rect 24670 32498 24722 32510
rect 25342 32562 25394 32574
rect 25342 32498 25394 32510
rect 28814 32562 28866 32574
rect 28814 32498 28866 32510
rect 29038 32562 29090 32574
rect 29038 32498 29090 32510
rect 29262 32562 29314 32574
rect 30126 32566 30138 32618
rect 30190 32566 30202 32618
rect 30382 32610 30434 32622
rect 33182 32674 33234 32686
rect 33182 32610 33234 32622
rect 47294 32618 47346 32630
rect 35870 32562 35922 32574
rect 30930 32510 30942 32562
rect 30994 32510 31006 32562
rect 31154 32510 31166 32562
rect 31218 32510 31230 32562
rect 35074 32510 35086 32562
rect 35138 32510 35150 32562
rect 36418 32537 36430 32589
rect 36482 32537 36494 32589
rect 38894 32562 38946 32574
rect 39174 32562 39226 32574
rect 29262 32498 29314 32510
rect 35870 32498 35922 32510
rect 38994 32510 39006 32562
rect 39058 32510 39070 32562
rect 38894 32498 38946 32510
rect 39174 32498 39226 32510
rect 40462 32562 40514 32574
rect 40842 32526 40854 32578
rect 40906 32526 40918 32578
rect 41010 32566 41022 32618
rect 41074 32566 41086 32618
rect 41234 32566 41246 32618
rect 41298 32566 41310 32618
rect 41458 32566 41470 32618
rect 41522 32566 41534 32618
rect 41750 32562 41802 32574
rect 44942 32562 44994 32574
rect 40462 32498 40514 32510
rect 44146 32510 44158 32562
rect 44210 32510 44222 32562
rect 41750 32498 41802 32510
rect 44942 32498 44994 32510
rect 45614 32562 45666 32574
rect 46478 32566 46490 32618
rect 46542 32566 46554 32618
rect 47294 32554 47346 32566
rect 48022 32618 48074 32630
rect 47618 32510 47630 32562
rect 47682 32510 47694 32562
rect 48022 32554 48074 32566
rect 45614 32498 45666 32510
rect 22374 32450 22426 32462
rect 32118 32450 32170 32462
rect 18790 32394 18842 32406
rect 5518 32338 5570 32350
rect 5518 32274 5570 32286
rect 6638 32338 6690 32350
rect 6638 32274 6690 32286
rect 15710 32338 15762 32350
rect 26114 32398 26126 32450
rect 26178 32398 26190 32450
rect 28018 32398 28030 32450
rect 28082 32398 28094 32450
rect 22374 32386 22426 32398
rect 30830 32394 30882 32406
rect 18790 32330 18842 32342
rect 32118 32386 32170 32398
rect 39566 32450 39618 32462
rect 45334 32450 45386 32462
rect 42242 32398 42254 32450
rect 42306 32398 42318 32450
rect 39566 32386 39618 32398
rect 45334 32386 45386 32398
rect 47854 32450 47906 32462
rect 47854 32386 47906 32398
rect 28522 32286 28534 32338
rect 28586 32286 28598 32338
rect 30830 32330 30882 32342
rect 46734 32338 46786 32350
rect 15710 32274 15762 32286
rect 46734 32274 46786 32286
rect 1344 32170 48608 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 48608 32170
rect 1344 32084 48608 32118
rect 4846 32002 4898 32014
rect 4846 31938 4898 31950
rect 7086 32002 7138 32014
rect 7086 31938 7138 31950
rect 13582 32002 13634 32014
rect 13582 31938 13634 31950
rect 22542 32002 22594 32014
rect 22542 31938 22594 31950
rect 26686 32002 26738 32014
rect 31166 32002 31218 32014
rect 29530 31950 29542 32002
rect 29594 31950 29606 32002
rect 26686 31938 26738 31950
rect 31166 31938 31218 31950
rect 38558 32002 38610 32014
rect 38558 31938 38610 31950
rect 43878 32002 43930 32014
rect 43878 31938 43930 31950
rect 21982 31890 22034 31902
rect 8082 31838 8094 31890
rect 8146 31838 8158 31890
rect 9258 31838 9270 31890
rect 9322 31838 9334 31890
rect 17782 31834 17834 31846
rect 2606 31778 2658 31790
rect 3614 31778 3666 31790
rect 2930 31726 2942 31778
rect 2994 31726 3006 31778
rect 2606 31714 2658 31726
rect 3266 31670 3278 31722
rect 3330 31670 3342 31722
rect 3614 31714 3666 31726
rect 4174 31778 4226 31790
rect 5630 31778 5682 31790
rect 7422 31778 7474 31790
rect 8318 31778 8370 31790
rect 4274 31726 4286 31778
rect 4338 31726 4350 31778
rect 6178 31726 6190 31778
rect 6242 31726 6254 31778
rect 7746 31726 7758 31778
rect 7810 31726 7822 31778
rect 4174 31714 4226 31726
rect 4442 31670 4454 31722
rect 4506 31670 4518 31722
rect 5630 31714 5682 31726
rect 7422 31714 7474 31726
rect 7970 31711 7982 31763
rect 8034 31711 8046 31763
rect 8318 31714 8370 31726
rect 8542 31778 8594 31790
rect 8542 31714 8594 31726
rect 9550 31778 9602 31790
rect 9550 31714 9602 31726
rect 9774 31778 9826 31790
rect 11342 31778 11394 31790
rect 14254 31778 14306 31790
rect 15878 31778 15930 31790
rect 9774 31714 9826 31726
rect 11062 31722 11114 31734
rect 10110 31666 10162 31678
rect 10490 31670 10502 31722
rect 10554 31670 10566 31722
rect 10770 31670 10782 31722
rect 10834 31670 10846 31722
rect 14130 31726 14142 31778
rect 14194 31726 14206 31778
rect 14466 31726 14478 31778
rect 14530 31726 14542 31778
rect 11342 31714 11394 31726
rect 12206 31670 12218 31722
rect 12270 31670 12282 31722
rect 8810 31614 8822 31666
rect 8874 31614 8886 31666
rect 11062 31658 11114 31670
rect 12462 31666 12514 31678
rect 13964 31670 13976 31722
rect 14028 31670 14040 31722
rect 14254 31714 14306 31726
rect 15878 31714 15930 31726
rect 16494 31778 16546 31790
rect 16494 31714 16546 31726
rect 16606 31778 16658 31790
rect 21982 31826 22034 31838
rect 26294 31890 26346 31902
rect 37158 31890 37210 31902
rect 33338 31838 33350 31890
rect 33402 31838 33414 31890
rect 41570 31838 41582 31890
rect 41634 31838 41646 31890
rect 48066 31838 48078 31890
rect 48130 31838 48142 31890
rect 26294 31826 26346 31838
rect 37158 31826 37210 31838
rect 17378 31726 17390 31778
rect 17442 31726 17454 31778
rect 17782 31770 17834 31782
rect 21310 31778 21362 31790
rect 22878 31778 22930 31790
rect 27022 31778 27074 31790
rect 16606 31714 16658 31726
rect 17154 31670 17166 31722
rect 17218 31670 17230 31722
rect 18610 31698 18622 31750
rect 18674 31698 18686 31750
rect 20514 31726 20526 31778
rect 20578 31726 20590 31778
rect 21410 31726 21422 31778
rect 21474 31726 21486 31778
rect 21310 31714 21362 31726
rect 17614 31666 17666 31678
rect 21576 31670 21588 31722
rect 21640 31670 21652 31722
rect 22878 31714 22930 31726
rect 24278 31722 24330 31734
rect 2270 31554 2322 31566
rect 3042 31558 3054 31610
rect 3106 31558 3118 31610
rect 6290 31558 6302 31610
rect 6354 31558 6366 31610
rect 10110 31602 10162 31614
rect 16202 31614 16214 31666
rect 16266 31614 16278 31666
rect 12462 31602 12514 31614
rect 17614 31602 17666 31614
rect 23998 31666 24050 31678
rect 24546 31687 24558 31739
rect 24610 31687 24622 31739
rect 25106 31726 25118 31778
rect 25170 31726 25182 31778
rect 24770 31670 24782 31722
rect 24834 31670 24846 31722
rect 27022 31714 27074 31726
rect 27246 31778 27298 31790
rect 28366 31778 28418 31790
rect 28110 31726 28122 31778
rect 28174 31726 28186 31778
rect 27246 31714 27298 31726
rect 28366 31714 28418 31726
rect 29038 31778 29090 31790
rect 29038 31714 29090 31726
rect 29262 31778 29314 31790
rect 31614 31778 31666 31790
rect 29262 31714 29314 31726
rect 30214 31722 30266 31734
rect 30426 31670 30438 31722
rect 30490 31670 30502 31722
rect 30594 31670 30606 31722
rect 30658 31670 30670 31722
rect 31614 31714 31666 31726
rect 31838 31778 31890 31790
rect 33630 31778 33682 31790
rect 33058 31726 33070 31778
rect 33122 31726 33134 31778
rect 31838 31714 31890 31726
rect 33630 31714 33682 31726
rect 33742 31778 33794 31790
rect 35198 31778 35250 31790
rect 42254 31778 42306 31790
rect 33954 31726 33966 31778
rect 34018 31726 34030 31778
rect 36062 31726 36074 31778
rect 36126 31726 36138 31778
rect 40910 31750 40962 31762
rect 33742 31714 33794 31726
rect 35198 31714 35250 31726
rect 37538 31698 37550 31750
rect 37602 31698 37614 31750
rect 24278 31658 24330 31670
rect 30214 31658 30266 31670
rect 36318 31666 36370 31678
rect 32106 31614 32118 31666
rect 32170 31614 32182 31666
rect 23998 31602 24050 31614
rect 32902 31610 32954 31622
rect 2270 31490 2322 31502
rect 23606 31554 23658 31566
rect 23606 31490 23658 31502
rect 25286 31554 25338 31566
rect 25286 31490 25338 31502
rect 25846 31554 25898 31566
rect 36318 31602 36370 31614
rect 40406 31666 40458 31678
rect 40674 31670 40686 31722
rect 40738 31670 40750 31722
rect 40910 31686 40962 31698
rect 41134 31750 41186 31762
rect 41134 31686 41186 31698
rect 41246 31743 41298 31755
rect 41246 31679 41298 31691
rect 41682 31682 41694 31734
rect 41746 31682 41758 31734
rect 42018 31726 42030 31778
rect 42082 31726 42094 31778
rect 44718 31778 44770 31790
rect 42254 31714 42306 31726
rect 43038 31743 43090 31755
rect 43038 31679 43090 31691
rect 43150 31750 43202 31762
rect 43150 31686 43202 31698
rect 43374 31750 43426 31762
rect 43374 31686 43426 31698
rect 43598 31750 43650 31762
rect 44718 31714 44770 31726
rect 45390 31778 45442 31790
rect 46162 31726 46174 31778
rect 46226 31726 46238 31778
rect 45390 31714 45442 31726
rect 43598 31686 43650 31698
rect 40406 31602 40458 31614
rect 32902 31546 32954 31558
rect 42590 31554 42642 31566
rect 25846 31490 25898 31502
rect 42590 31490 42642 31502
rect 45054 31554 45106 31566
rect 45054 31490 45106 31502
rect 1344 31386 48608 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 48608 31386
rect 1344 31300 48608 31334
rect 11062 31218 11114 31230
rect 11062 31154 11114 31166
rect 26294 31218 26346 31230
rect 26294 31154 26346 31166
rect 26742 31218 26794 31230
rect 26742 31154 26794 31166
rect 10446 31106 10498 31118
rect 27806 31106 27858 31118
rect 5114 31054 5126 31106
rect 5178 31054 5190 31106
rect 6582 31050 6634 31062
rect 7802 31054 7814 31106
rect 7866 31054 7878 31106
rect 1598 30994 1650 31006
rect 4286 30994 4338 31006
rect 2370 30942 2382 30994
rect 2434 30942 2446 30994
rect 1598 30930 1650 30942
rect 4286 30930 4338 30942
rect 4734 30994 4786 31006
rect 4734 30930 4786 30942
rect 4846 30994 4898 31006
rect 4846 30930 4898 30942
rect 6190 30994 6242 31006
rect 6190 30930 6242 30942
rect 6414 30994 6466 31006
rect 9494 31050 9546 31062
rect 7310 31032 7362 31044
rect 6582 30986 6634 30998
rect 6750 30994 6802 31006
rect 6414 30930 6466 30942
rect 6962 30942 6974 30994
rect 7026 30942 7038 30994
rect 7310 30968 7362 30980
rect 8094 30994 8146 31006
rect 6750 30930 6802 30942
rect 8094 30930 8146 30942
rect 8206 30994 8258 31006
rect 8206 30930 8258 30942
rect 8430 30994 8482 31006
rect 21242 31054 21254 31106
rect 21306 31054 21318 31106
rect 10446 31042 10498 31054
rect 27806 31042 27858 31054
rect 35758 31106 35810 31118
rect 9494 30986 9546 30998
rect 9650 30972 9662 31024
rect 9714 30972 9726 31024
rect 9874 30981 9886 31033
rect 9938 30981 9950 31033
rect 11442 30969 11454 31021
rect 11506 30969 11518 31021
rect 13358 30994 13410 31006
rect 8430 30930 8482 30942
rect 13358 30930 13410 30942
rect 14142 30994 14194 31006
rect 16158 30994 16210 31006
rect 15006 30942 15018 30994
rect 15070 30942 15082 30994
rect 14142 30930 14194 30942
rect 16158 30930 16210 30942
rect 16718 30994 16770 31006
rect 16718 30930 16770 30942
rect 16830 30994 16882 31006
rect 16830 30930 16882 30942
rect 17670 30994 17722 31006
rect 17938 30942 17950 30994
rect 18002 30942 18014 30994
rect 18274 30986 18286 31038
rect 18338 30986 18350 31038
rect 28366 31032 28418 31044
rect 20414 30994 20466 31006
rect 18610 30942 18622 30994
rect 18674 30942 18686 30994
rect 17670 30930 17722 30942
rect 20414 30930 20466 30942
rect 20526 30994 20578 31006
rect 20526 30930 20578 30942
rect 20750 30994 20802 31006
rect 20750 30930 20802 30942
rect 20974 30994 21026 31006
rect 23214 30994 23266 31006
rect 24558 30994 24610 31006
rect 21746 30942 21758 30994
rect 21810 30942 21822 30994
rect 21970 30942 21982 30994
rect 22034 30942 22046 30994
rect 22306 30942 22318 30994
rect 22370 30991 22382 30994
rect 22530 30991 22542 30994
rect 22370 30945 22542 30991
rect 22370 30942 22382 30945
rect 22530 30942 22542 30945
rect 22594 30942 22606 30994
rect 23538 30942 23550 30994
rect 23602 30942 23614 30994
rect 23874 30942 23886 30994
rect 23938 30942 23950 30994
rect 24266 30942 24278 30994
rect 24330 30942 24342 30994
rect 20974 30930 21026 30942
rect 23214 30930 23266 30942
rect 24558 30930 24610 30942
rect 24670 30994 24722 31006
rect 25566 30994 25618 31006
rect 25274 30942 25286 30994
rect 25338 30942 25350 30994
rect 24670 30930 24722 30942
rect 25566 30930 25618 30942
rect 25678 30994 25730 31006
rect 25678 30930 25730 30942
rect 26910 30994 26962 31006
rect 26910 30930 26962 30942
rect 27638 30938 27690 30950
rect 28018 30942 28030 30994
rect 28082 30942 28094 30994
rect 29598 30994 29650 31006
rect 30462 30998 30474 31050
rect 30526 30998 30538 31050
rect 28366 30968 28418 30980
rect 29362 30942 29374 30994
rect 29426 30942 29438 30994
rect 29598 30930 29650 30942
rect 30718 30994 30770 31006
rect 30718 30930 30770 30942
rect 31166 30994 31218 31006
rect 32286 30994 32338 31006
rect 32030 30942 32042 30994
rect 32094 30942 32106 30994
rect 31166 30930 31218 30942
rect 32286 30930 32338 30942
rect 33070 30994 33122 31006
rect 33934 30998 33946 31050
rect 33998 30998 34010 31050
rect 35758 31042 35810 31054
rect 40238 31106 40290 31118
rect 36840 31032 36892 31044
rect 40238 31042 40290 31054
rect 41022 31106 41074 31118
rect 41022 31042 41074 31054
rect 48078 31106 48130 31118
rect 48078 31042 48130 31054
rect 33070 30930 33122 30942
rect 34190 30994 34242 31006
rect 34190 30930 34242 30942
rect 34638 30994 34690 31006
rect 36542 30994 36594 31006
rect 35502 30942 35514 30994
rect 35566 30942 35578 30994
rect 36642 30942 36654 30994
rect 36706 30942 36718 30994
rect 36840 30968 36892 30980
rect 37550 30994 37602 31006
rect 43710 30994 43762 31006
rect 44718 30994 44770 31006
rect 42914 30942 42926 30994
rect 42978 30942 42990 30994
rect 44034 30942 44046 30994
rect 44098 30942 44110 30994
rect 34638 30930 34690 30942
rect 36542 30930 36594 30942
rect 37550 30930 37602 30942
rect 43710 30930 43762 30942
rect 44718 30930 44770 30942
rect 45222 30994 45274 31006
rect 45222 30930 45274 30942
rect 45390 30994 45442 31006
rect 45390 30930 45442 30942
rect 5898 30830 5910 30882
rect 5962 30830 5974 30882
rect 18386 30830 18398 30882
rect 18450 30830 18462 30882
rect 20122 30830 20134 30882
rect 20186 30830 20198 30882
rect 27638 30874 27690 30886
rect 37214 30882 37266 30894
rect 22094 30826 22146 30838
rect 29206 30826 29258 30838
rect 8766 30770 8818 30782
rect 8766 30706 8818 30718
rect 15262 30770 15314 30782
rect 15262 30706 15314 30718
rect 15822 30770 15874 30782
rect 16426 30718 16438 30770
rect 16490 30718 16502 30770
rect 22094 30762 22146 30774
rect 22878 30770 22930 30782
rect 23762 30774 23774 30826
rect 23826 30774 23838 30826
rect 15822 30706 15874 30718
rect 22878 30706 22930 30718
rect 27246 30770 27298 30782
rect 38322 30830 38334 30882
rect 38386 30830 38398 30882
rect 46162 30830 46174 30882
rect 46226 30830 46238 30882
rect 37214 30818 37266 30830
rect 43922 30774 43934 30826
rect 43986 30774 43998 30826
rect 29206 30762 29258 30774
rect 27246 30706 27298 30718
rect 1344 30602 48608 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 48608 30602
rect 1344 30516 48608 30550
rect 10110 30434 10162 30446
rect 11790 30434 11842 30446
rect 10110 30370 10162 30382
rect 10894 30378 10946 30390
rect 11790 30370 11842 30382
rect 14590 30434 14642 30446
rect 19114 30382 19126 30434
rect 19178 30382 19190 30434
rect 29530 30382 29542 30434
rect 29594 30382 29606 30434
rect 14590 30370 14642 30382
rect 30606 30378 30658 30390
rect 3154 30270 3166 30322
rect 3218 30270 3230 30322
rect 6290 30270 6302 30322
rect 6354 30270 6366 30322
rect 10894 30314 10946 30326
rect 18342 30322 18394 30334
rect 27906 30326 27918 30378
rect 27970 30326 27982 30378
rect 15810 30270 15822 30322
rect 15874 30270 15886 30322
rect 17714 30270 17726 30322
rect 17778 30270 17790 30322
rect 23314 30270 23326 30322
rect 23378 30270 23390 30322
rect 30606 30314 30658 30326
rect 30942 30378 30994 30390
rect 34526 30378 34578 30390
rect 45658 30382 45670 30434
rect 45722 30382 45734 30434
rect 33394 30326 33406 30378
rect 33458 30326 33470 30378
rect 30942 30314 30994 30326
rect 34526 30314 34578 30326
rect 41010 30270 41022 30322
rect 41074 30270 41086 30322
rect 44818 30270 44830 30322
rect 44882 30270 44894 30322
rect 46386 30270 46398 30322
rect 46450 30270 46462 30322
rect 47618 30270 47630 30322
rect 47682 30270 47694 30322
rect 18342 30258 18394 30270
rect 3502 30210 3554 30222
rect 5518 30210 5570 30222
rect 2818 30158 2830 30210
rect 2882 30158 2894 30210
rect 3042 30143 3054 30195
rect 3106 30143 3118 30195
rect 4366 30158 4378 30210
rect 4430 30158 4442 30210
rect 3502 30146 3554 30158
rect 5518 30146 5570 30158
rect 8206 30210 8258 30222
rect 12910 30210 12962 30222
rect 8978 30158 8990 30210
rect 9042 30158 9054 30210
rect 8206 30146 8258 30158
rect 9158 30154 9210 30166
rect 10994 30158 11006 30210
rect 11058 30158 11070 30210
rect 11330 30158 11342 30210
rect 11394 30158 11406 30210
rect 4622 30098 4674 30110
rect 9314 30102 9326 30154
rect 9378 30102 9390 30154
rect 9538 30102 9550 30154
rect 9602 30102 9614 30154
rect 12021 30102 12033 30154
rect 12085 30102 12097 30154
rect 12910 30146 12962 30158
rect 13470 30210 13522 30222
rect 15038 30210 15090 30222
rect 14334 30158 14346 30210
rect 14398 30158 14410 30210
rect 13470 30146 13522 30158
rect 15038 30146 15090 30158
rect 18734 30210 18786 30222
rect 18734 30146 18786 30158
rect 18846 30210 18898 30222
rect 21422 30210 21474 30222
rect 22542 30210 22594 30222
rect 18846 30146 18898 30158
rect 19506 30125 19518 30177
rect 19570 30125 19582 30177
rect 19786 30102 19798 30154
rect 19850 30102 19862 30154
rect 20402 30102 20414 30154
rect 20466 30102 20478 30154
rect 20558 30118 20570 30170
rect 20622 30118 20634 30170
rect 21254 30154 21306 30166
rect 9158 30090 9210 30102
rect 20750 30098 20802 30110
rect 4622 30034 4674 30046
rect 21634 30158 21646 30210
rect 21698 30158 21710 30210
rect 21422 30146 21474 30158
rect 21858 30102 21870 30154
rect 21922 30102 21934 30154
rect 22542 30146 22594 30158
rect 25678 30210 25730 30222
rect 25678 30146 25730 30158
rect 26798 30210 26850 30222
rect 29150 30210 29202 30222
rect 27906 30158 27918 30210
rect 27970 30158 27982 30210
rect 28242 30158 28254 30210
rect 28306 30158 28318 30210
rect 21254 30090 21306 30102
rect 25230 30098 25282 30110
rect 26542 30102 26554 30154
rect 26606 30102 26618 30154
rect 26798 30146 26850 30158
rect 29150 30146 29202 30158
rect 29262 30210 29314 30222
rect 34190 30210 34242 30222
rect 35814 30210 35866 30222
rect 30146 30158 30158 30210
rect 30210 30158 30222 30210
rect 30482 30158 30494 30210
rect 30546 30158 30558 30210
rect 31042 30158 31054 30210
rect 31106 30158 31118 30210
rect 31266 30158 31278 30210
rect 31330 30158 31342 30210
rect 29262 30146 29314 30158
rect 32006 30154 32058 30166
rect 32162 30128 32174 30180
rect 32226 30128 32238 30180
rect 32386 30119 32398 30171
rect 32450 30119 32462 30171
rect 33618 30158 33630 30210
rect 33682 30158 33694 30210
rect 34626 30158 34638 30210
rect 34690 30158 34702 30210
rect 34190 30146 34242 30158
rect 35302 30120 35314 30172
rect 35366 30120 35378 30172
rect 35814 30146 35866 30158
rect 36206 30210 36258 30222
rect 36206 30146 36258 30158
rect 36542 30210 36594 30222
rect 38502 30210 38554 30222
rect 36542 30146 36594 30158
rect 37382 30154 37434 30166
rect 20750 30034 20802 30046
rect 32006 30090 32058 30102
rect 32958 30098 33010 30110
rect 25230 30034 25282 30046
rect 32958 30034 33010 30046
rect 37102 30098 37154 30110
rect 37538 30102 37550 30154
rect 37602 30102 37614 30154
rect 37874 30102 37886 30154
rect 37938 30102 37950 30154
rect 38502 30146 38554 30158
rect 38950 30210 39002 30222
rect 38950 30146 39002 30158
rect 39230 30210 39282 30222
rect 39678 30210 39730 30222
rect 43710 30210 43762 30222
rect 45950 30210 46002 30222
rect 39330 30158 39342 30210
rect 39394 30158 39406 30210
rect 39230 30146 39282 30158
rect 39498 30102 39510 30154
rect 39562 30102 39574 30154
rect 39678 30146 39730 30158
rect 40226 30130 40238 30182
rect 40290 30130 40302 30182
rect 43026 30158 43038 30210
rect 43090 30158 43102 30210
rect 43486 30171 43538 30183
rect 43710 30146 43762 30158
rect 44930 30143 44942 30195
rect 44994 30143 45006 30195
rect 45154 30158 45166 30210
rect 45218 30158 45230 30210
rect 45950 30146 46002 30158
rect 46062 30210 46114 30222
rect 46062 30146 46114 30158
rect 46498 30143 46510 30195
rect 46562 30143 46574 30195
rect 46834 30158 46846 30210
rect 46898 30158 46910 30210
rect 47170 30158 47182 30210
rect 47234 30158 47246 30210
rect 47506 30143 47518 30195
rect 47570 30143 47582 30195
rect 43486 30107 43538 30119
rect 37382 30090 37434 30102
rect 37102 30034 37154 30046
rect 8822 29986 8874 29998
rect 8822 29922 8874 29934
rect 27414 29986 27466 29998
rect 43586 29990 43598 30042
rect 43650 29990 43662 30042
rect 27414 29922 27466 29934
rect 48134 29986 48186 29998
rect 48134 29922 48186 29934
rect 1344 29818 48608 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 48608 29818
rect 1344 29732 48608 29766
rect 2102 29650 2154 29662
rect 7478 29650 7530 29662
rect 2102 29586 2154 29598
rect 5350 29594 5402 29606
rect 2494 29538 2546 29550
rect 7478 29586 7530 29598
rect 23830 29650 23882 29662
rect 23830 29586 23882 29598
rect 30550 29650 30602 29662
rect 30550 29586 30602 29598
rect 32566 29650 32618 29662
rect 32566 29586 32618 29598
rect 35926 29650 35978 29662
rect 35926 29586 35978 29598
rect 42198 29650 42250 29662
rect 42198 29586 42250 29598
rect 5350 29530 5402 29542
rect 7870 29538 7922 29550
rect 2494 29474 2546 29486
rect 3042 29430 3054 29482
rect 3106 29430 3118 29482
rect 3266 29430 3278 29482
rect 3330 29430 3342 29482
rect 7870 29474 7922 29486
rect 10670 29538 10722 29550
rect 18958 29538 19010 29550
rect 15754 29486 15766 29538
rect 15818 29486 15830 29538
rect 16202 29486 16214 29538
rect 16266 29486 16278 29538
rect 3726 29426 3778 29438
rect 4590 29374 4602 29426
rect 4654 29374 4666 29426
rect 5506 29374 5518 29426
rect 5570 29374 5582 29426
rect 5842 29418 5854 29470
rect 5906 29418 5918 29470
rect 8101 29430 8113 29482
rect 8165 29430 8177 29482
rect 10670 29474 10722 29486
rect 8990 29426 9042 29438
rect 6178 29374 6190 29426
rect 6242 29374 6254 29426
rect 6626 29374 6638 29426
rect 6690 29374 6702 29426
rect 6850 29374 6862 29426
rect 6914 29374 6926 29426
rect 2762 29318 2774 29370
rect 2826 29318 2838 29370
rect 3726 29362 3778 29374
rect 8990 29362 9042 29374
rect 9550 29426 9602 29438
rect 11330 29430 11342 29482
rect 11394 29430 11406 29482
rect 12786 29430 12798 29482
rect 12850 29430 12862 29482
rect 13794 29430 13806 29482
rect 13858 29430 13870 29482
rect 18958 29474 19010 29486
rect 19350 29538 19402 29550
rect 25342 29538 25394 29550
rect 19350 29474 19402 29486
rect 25174 29482 25226 29494
rect 10414 29374 10426 29426
rect 10478 29374 10490 29426
rect 12226 29374 12238 29426
rect 12290 29374 12302 29426
rect 14740 29399 14752 29451
rect 14804 29399 14816 29451
rect 15038 29426 15090 29438
rect 14914 29374 14926 29426
rect 14978 29374 14990 29426
rect 9550 29362 9602 29374
rect 15038 29362 15090 29374
rect 15374 29426 15426 29438
rect 15374 29362 15426 29374
rect 15486 29426 15538 29438
rect 15486 29362 15538 29374
rect 16494 29426 16546 29438
rect 16494 29362 16546 29374
rect 16718 29426 16770 29438
rect 18622 29426 18674 29438
rect 17938 29374 17950 29426
rect 18002 29374 18014 29426
rect 18162 29374 18174 29426
rect 18226 29374 18238 29426
rect 19070 29426 19122 29438
rect 16718 29362 16770 29374
rect 18622 29362 18674 29374
rect 18790 29370 18842 29382
rect 12014 29314 12066 29326
rect 5730 29262 5742 29314
rect 5794 29262 5806 29314
rect 6526 29258 6578 29270
rect 4846 29202 4898 29214
rect 12014 29250 12066 29262
rect 14366 29314 14418 29326
rect 14366 29250 14418 29262
rect 17558 29314 17610 29326
rect 19070 29362 19122 29374
rect 19742 29426 19794 29438
rect 20022 29426 20074 29438
rect 21422 29426 21474 29438
rect 19842 29374 19854 29426
rect 19906 29374 19918 29426
rect 21074 29374 21086 29426
rect 21138 29374 21150 29426
rect 19742 29362 19794 29374
rect 20022 29362 20074 29374
rect 21422 29362 21474 29374
rect 21534 29426 21586 29438
rect 22206 29426 22258 29438
rect 22654 29426 22706 29438
rect 25342 29474 25394 29486
rect 29878 29538 29930 29550
rect 25722 29430 25734 29482
rect 25786 29430 25798 29482
rect 29878 29474 29930 29486
rect 34862 29538 34914 29550
rect 42702 29538 42754 29550
rect 39050 29486 39062 29538
rect 39114 29486 39126 29538
rect 29038 29461 29090 29473
rect 21802 29374 21814 29426
rect 21866 29374 21878 29426
rect 21534 29362 21586 29374
rect 22206 29362 22258 29374
rect 22374 29370 22426 29382
rect 22530 29374 22542 29426
rect 22594 29374 22606 29426
rect 24322 29374 24334 29426
rect 24386 29374 24398 29426
rect 24658 29374 24670 29426
rect 24722 29374 24734 29426
rect 25174 29418 25226 29430
rect 27190 29426 27242 29438
rect 27918 29426 27970 29438
rect 25554 29374 25566 29426
rect 25618 29374 25630 29426
rect 27570 29374 27582 29426
rect 27634 29374 27646 29426
rect 28242 29374 28254 29426
rect 28306 29374 28318 29426
rect 28578 29374 28590 29426
rect 28642 29374 28654 29426
rect 29038 29397 29090 29409
rect 29150 29454 29202 29466
rect 29150 29390 29202 29402
rect 29374 29454 29426 29466
rect 29374 29390 29426 29402
rect 29598 29454 29650 29466
rect 29598 29390 29650 29402
rect 30830 29426 30882 29438
rect 31694 29430 31706 29482
rect 31758 29430 31770 29482
rect 34862 29474 34914 29486
rect 18790 29306 18842 29318
rect 20414 29314 20466 29326
rect 17558 29250 17610 29262
rect 22654 29362 22706 29374
rect 27190 29362 27242 29374
rect 27918 29362 27970 29374
rect 30830 29362 30882 29374
rect 31950 29426 32002 29438
rect 31950 29362 32002 29374
rect 33742 29426 33794 29438
rect 36318 29426 36370 29438
rect 37182 29430 37194 29482
rect 37246 29430 37258 29482
rect 42702 29474 42754 29486
rect 34606 29374 34618 29426
rect 34670 29374 34682 29426
rect 36082 29374 36094 29426
rect 36146 29374 36158 29426
rect 33742 29362 33794 29374
rect 36318 29362 36370 29374
rect 37886 29426 37938 29438
rect 37886 29362 37938 29374
rect 37998 29426 38050 29438
rect 37998 29362 38050 29374
rect 38558 29426 38610 29438
rect 38558 29362 38610 29374
rect 38782 29426 38834 29438
rect 45390 29426 45442 29438
rect 39778 29374 39790 29426
rect 39842 29374 39854 29426
rect 40786 29374 40798 29426
rect 40850 29374 40862 29426
rect 44594 29374 44606 29426
rect 44658 29374 44670 29426
rect 38782 29362 38834 29374
rect 45390 29362 45442 29374
rect 45950 29426 46002 29438
rect 45950 29362 46002 29374
rect 46174 29426 46226 29438
rect 46734 29426 46786 29438
rect 46442 29374 46454 29426
rect 46506 29374 46518 29426
rect 46174 29362 46226 29374
rect 46734 29362 46786 29374
rect 48302 29426 48354 29438
rect 48302 29362 48354 29374
rect 22374 29306 22426 29318
rect 26742 29314 26794 29326
rect 18162 29206 18174 29258
rect 18226 29206 18238 29258
rect 20414 29250 20466 29262
rect 6526 29194 6578 29206
rect 20918 29202 20970 29214
rect 4846 29138 4898 29150
rect 20918 29138 20970 29150
rect 23214 29202 23266 29214
rect 24434 29206 24446 29258
rect 24498 29206 24510 29258
rect 26742 29250 26794 29262
rect 27358 29314 27410 29326
rect 27358 29250 27410 29262
rect 33462 29314 33514 29326
rect 33462 29250 33514 29262
rect 35478 29314 35530 29326
rect 35478 29250 35530 29262
rect 39622 29314 39674 29326
rect 39622 29250 39674 29262
rect 45782 29314 45834 29326
rect 45782 29250 45834 29262
rect 23214 29138 23266 29150
rect 37438 29202 37490 29214
rect 47070 29202 47122 29214
rect 38266 29150 38278 29202
rect 38330 29150 38342 29202
rect 37438 29138 37490 29150
rect 47070 29138 47122 29150
rect 47966 29202 48018 29214
rect 47966 29138 48018 29150
rect 1344 29034 48608 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 48608 29034
rect 1344 28948 48608 28982
rect 10110 28866 10162 28878
rect 10110 28802 10162 28814
rect 12686 28866 12738 28878
rect 15934 28866 15986 28878
rect 12686 28802 12738 28814
rect 14814 28810 14866 28822
rect 6302 28754 6354 28766
rect 1810 28702 1822 28754
rect 1874 28702 1886 28754
rect 3714 28702 3726 28754
rect 3778 28702 3790 28754
rect 15934 28802 15986 28814
rect 18902 28866 18954 28878
rect 23102 28866 23154 28878
rect 31054 28866 31106 28878
rect 21690 28814 21702 28866
rect 21754 28814 21766 28866
rect 28074 28814 28086 28866
rect 28138 28814 28150 28866
rect 14814 28746 14866 28758
rect 17446 28754 17498 28766
rect 18274 28758 18286 28810
rect 18338 28758 18350 28810
rect 18902 28802 18954 28814
rect 19506 28758 19518 28810
rect 19570 28758 19582 28810
rect 20402 28758 20414 28810
rect 20466 28758 20478 28810
rect 23102 28802 23154 28814
rect 29150 28810 29202 28822
rect 27750 28754 27802 28766
rect 6302 28690 6354 28702
rect 6470 28698 6522 28710
rect 4510 28642 4562 28654
rect 4510 28578 4562 28590
rect 4902 28642 4954 28654
rect 23650 28702 23662 28754
rect 23714 28702 23726 28754
rect 31054 28802 31106 28814
rect 36318 28866 36370 28878
rect 31826 28758 31838 28810
rect 31890 28758 31902 28810
rect 36318 28802 36370 28814
rect 43710 28866 43762 28878
rect 43710 28802 43762 28814
rect 44942 28866 44994 28878
rect 44942 28802 44994 28814
rect 29150 28746 29202 28758
rect 37158 28754 37210 28766
rect 44326 28754 44378 28766
rect 17446 28690 17498 28702
rect 27750 28690 27802 28702
rect 40562 28702 40574 28754
rect 40626 28702 40638 28754
rect 42466 28702 42478 28754
rect 42530 28702 42542 28754
rect 47506 28702 47518 28754
rect 47570 28702 47582 28754
rect 37158 28690 37210 28702
rect 44326 28690 44378 28702
rect 4902 28578 4954 28590
rect 5742 28604 5794 28616
rect 6066 28590 6078 28642
rect 6130 28590 6142 28642
rect 6470 28634 6522 28646
rect 7422 28642 7474 28654
rect 8990 28642 9042 28654
rect 10614 28642 10666 28654
rect 8286 28590 8298 28642
rect 8350 28590 8362 28642
rect 9854 28590 9866 28642
rect 9918 28590 9930 28642
rect 11678 28642 11730 28654
rect 7422 28578 7474 28590
rect 8990 28578 9042 28590
rect 10614 28578 10666 28590
rect 11342 28614 11394 28626
rect 5742 28540 5794 28552
rect 8542 28530 8594 28542
rect 10882 28534 10894 28586
rect 10946 28534 10958 28586
rect 11106 28534 11118 28586
rect 11170 28534 11182 28586
rect 11342 28550 11394 28562
rect 11454 28586 11506 28598
rect 11678 28578 11730 28590
rect 11902 28642 11954 28654
rect 13022 28642 13074 28654
rect 16270 28642 16322 28654
rect 21198 28642 21250 28654
rect 12170 28590 12182 28642
rect 12234 28590 12246 28642
rect 11902 28578 11954 28590
rect 13022 28578 13074 28590
rect 13638 28586 13690 28598
rect 14018 28590 14030 28642
rect 14082 28590 14094 28642
rect 14366 28604 14418 28616
rect 11454 28522 11506 28534
rect 14914 28590 14926 28642
rect 14978 28590 14990 28642
rect 15138 28590 15150 28642
rect 15202 28590 15214 28642
rect 16270 28578 16322 28590
rect 17710 28552 17722 28604
rect 17774 28552 17786 28604
rect 18386 28590 18398 28642
rect 18450 28590 18462 28642
rect 19058 28590 19070 28642
rect 19122 28590 19134 28642
rect 19394 28590 19406 28642
rect 19458 28590 19470 28642
rect 19730 28590 19742 28642
rect 19794 28590 19806 28642
rect 20290 28590 20302 28642
rect 20354 28590 20366 28642
rect 20514 28590 20526 28642
rect 20578 28590 20590 28642
rect 21198 28578 21250 28590
rect 21422 28642 21474 28654
rect 22262 28642 22314 28654
rect 22542 28642 22594 28654
rect 24222 28642 24274 28654
rect 21422 28578 21474 28590
rect 22094 28586 22146 28598
rect 13638 28522 13690 28534
rect 13806 28530 13858 28542
rect 14366 28540 14418 28552
rect 8542 28466 8594 28478
rect 22418 28590 22430 28642
rect 22482 28590 22494 28642
rect 23538 28590 23550 28642
rect 23602 28590 23614 28642
rect 22262 28578 22314 28590
rect 22542 28578 22594 28590
rect 23874 28563 23886 28615
rect 23938 28563 23950 28615
rect 24222 28578 24274 28590
rect 25454 28642 25506 28654
rect 25454 28578 25506 28590
rect 27302 28642 27354 28654
rect 26318 28534 26330 28586
rect 26382 28534 26394 28586
rect 27302 28578 27354 28590
rect 28366 28642 28418 28654
rect 28366 28578 28418 28590
rect 28478 28642 28530 28654
rect 29934 28642 29986 28654
rect 32566 28642 32618 28654
rect 29250 28590 29262 28642
rect 29314 28590 29326 28642
rect 29586 28590 29598 28642
rect 29650 28590 29662 28642
rect 31602 28590 31614 28642
rect 31666 28590 31678 28642
rect 31826 28590 31838 28642
rect 31890 28590 31902 28642
rect 28478 28578 28530 28590
rect 29934 28578 29986 28590
rect 22094 28522 22146 28534
rect 26574 28530 26626 28542
rect 30798 28534 30810 28586
rect 30862 28534 30874 28586
rect 32566 28578 32618 28590
rect 33014 28642 33066 28654
rect 33014 28578 33066 28590
rect 33630 28642 33682 28654
rect 34750 28642 34802 28654
rect 34494 28590 34506 28642
rect 34558 28590 34570 28642
rect 33630 28578 33682 28590
rect 34750 28578 34802 28590
rect 35198 28642 35250 28654
rect 37550 28642 37602 28654
rect 40238 28642 40290 28654
rect 36062 28590 36074 28642
rect 36126 28590 36138 28642
rect 39442 28590 39454 28642
rect 39506 28590 39518 28642
rect 35198 28578 35250 28590
rect 37550 28578 37602 28590
rect 40238 28578 40290 28590
rect 43262 28642 43314 28654
rect 43262 28578 43314 28590
rect 43374 28642 43426 28654
rect 43374 28578 43426 28590
rect 45278 28642 45330 28654
rect 45278 28578 45330 28590
rect 48302 28642 48354 28654
rect 48302 28578 48354 28590
rect 13806 28466 13858 28478
rect 26574 28466 26626 28478
rect 45614 28530 45666 28542
rect 45614 28466 45666 28478
rect 7142 28418 7194 28430
rect 7142 28354 7194 28366
rect 16998 28418 17050 28430
rect 16998 28354 17050 28366
rect 25174 28418 25226 28430
rect 25174 28354 25226 28366
rect 1344 28250 48608 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 48608 28250
rect 1344 28164 48608 28198
rect 7478 28082 7530 28094
rect 4902 28026 4954 28038
rect 16438 28082 16490 28094
rect 7478 28018 7530 28030
rect 8934 28026 8986 28038
rect 4902 27962 4954 27974
rect 16438 28018 16490 28030
rect 19518 28082 19570 28094
rect 19518 28018 19570 28030
rect 25398 28082 25450 28094
rect 25398 28018 25450 28030
rect 30774 28082 30826 28094
rect 30774 28018 30826 28030
rect 31278 28082 31330 28094
rect 31278 28018 31330 28030
rect 32566 28082 32618 28094
rect 32566 28018 32618 28030
rect 39342 28082 39394 28094
rect 39342 28018 39394 28030
rect 5450 27918 5462 27970
rect 5514 27918 5526 27970
rect 8934 27962 8986 27974
rect 9718 27970 9770 27982
rect 13470 27970 13522 27982
rect 1598 27858 1650 27870
rect 1598 27794 1650 27806
rect 4286 27858 4338 27870
rect 5742 27858 5794 27870
rect 4722 27806 4734 27858
rect 4786 27806 4798 27858
rect 4286 27794 4338 27806
rect 5742 27794 5794 27806
rect 5966 27858 6018 27870
rect 5966 27794 6018 27806
rect 6526 27858 6578 27870
rect 6794 27862 6806 27914
rect 6858 27862 6870 27914
rect 9718 27906 9770 27918
rect 10894 27914 10946 27926
rect 14590 27970 14642 27982
rect 9998 27886 10050 27898
rect 6974 27858 7026 27870
rect 6626 27806 6638 27858
rect 6690 27806 6702 27858
rect 6526 27794 6578 27806
rect 6974 27794 7026 27806
rect 7758 27858 7810 27870
rect 8038 27858 8090 27870
rect 7858 27806 7870 27858
rect 7922 27806 7934 27858
rect 9090 27806 9102 27858
rect 9154 27806 9166 27858
rect 10210 27862 10222 27914
rect 10274 27862 10286 27914
rect 10446 27886 10498 27898
rect 9998 27822 10050 27834
rect 10446 27822 10498 27834
rect 10558 27893 10610 27905
rect 10994 27862 11006 27914
rect 11058 27862 11070 27914
rect 11218 27862 11230 27914
rect 11282 27862 11294 27914
rect 11454 27886 11506 27898
rect 10894 27850 10946 27862
rect 10558 27829 10610 27841
rect 11454 27822 11506 27834
rect 12014 27897 12066 27909
rect 13470 27906 13522 27918
rect 13638 27914 13690 27926
rect 12014 27833 12066 27845
rect 13010 27834 13022 27886
rect 13074 27834 13086 27886
rect 13234 27806 13246 27858
rect 13298 27806 13310 27858
rect 13638 27850 13690 27862
rect 14030 27896 14082 27908
rect 14590 27906 14642 27918
rect 20638 27970 20690 27982
rect 14758 27858 14810 27870
rect 17950 27858 18002 27870
rect 14030 27832 14082 27844
rect 14354 27806 14366 27858
rect 14418 27806 14430 27858
rect 15138 27806 15150 27858
rect 15202 27806 15214 27858
rect 15362 27806 15374 27858
rect 15426 27806 15438 27858
rect 18274 27806 18286 27858
rect 18338 27806 18350 27858
rect 18950 27844 18962 27896
rect 19014 27844 19026 27896
rect 19182 27858 19234 27870
rect 20234 27862 20246 27914
rect 20298 27862 20310 27914
rect 20638 27906 20690 27918
rect 22766 27970 22818 27982
rect 32118 27970 32170 27982
rect 26842 27918 26854 27970
rect 26906 27918 26918 27970
rect 34190 27970 34242 27982
rect 41122 27974 41134 28026
rect 41186 27974 41198 28026
rect 21702 27887 21754 27899
rect 7758 27794 7810 27806
rect 8038 27794 8090 27806
rect 14758 27794 14810 27806
rect 17950 27794 18002 27806
rect 19182 27794 19234 27806
rect 20806 27802 20858 27814
rect 21298 27806 21310 27858
rect 21362 27806 21374 27858
rect 22530 27862 22542 27914
rect 22594 27862 22606 27914
rect 22766 27906 22818 27918
rect 23650 27862 23662 27914
rect 23714 27862 23726 27914
rect 24098 27862 24110 27914
rect 24162 27862 24174 27914
rect 29038 27897 29090 27909
rect 32118 27906 32170 27918
rect 33910 27914 33962 27926
rect 21702 27823 21754 27835
rect 23090 27806 23102 27858
rect 23154 27806 23166 27858
rect 25778 27806 25790 27858
rect 25842 27806 25854 27858
rect 26002 27821 26014 27873
rect 26066 27821 26078 27873
rect 26350 27858 26402 27870
rect 8430 27746 8482 27758
rect 2370 27694 2382 27746
rect 2434 27694 2446 27746
rect 8430 27682 8482 27694
rect 16886 27746 16938 27758
rect 19954 27750 19966 27802
rect 20018 27750 20030 27802
rect 26350 27794 26402 27806
rect 26574 27858 26626 27870
rect 26574 27794 26626 27806
rect 27470 27858 27522 27870
rect 27470 27794 27522 27806
rect 27638 27858 27690 27870
rect 27918 27858 27970 27870
rect 27794 27806 27806 27858
rect 27858 27806 27870 27858
rect 27638 27794 27690 27806
rect 27918 27794 27970 27806
rect 28814 27858 28866 27870
rect 30942 27858 30994 27870
rect 33394 27862 33406 27914
rect 33458 27862 33470 27914
rect 33730 27862 33742 27914
rect 33794 27862 33806 27914
rect 34190 27906 34242 27918
rect 46510 27970 46562 27982
rect 29038 27833 29090 27845
rect 29362 27806 29374 27858
rect 29426 27806 29438 27858
rect 29922 27806 29934 27858
rect 29986 27806 29998 27858
rect 30146 27806 30158 27858
rect 30210 27806 30222 27858
rect 33910 27850 33962 27862
rect 34526 27858 34578 27870
rect 28814 27794 28866 27806
rect 30942 27794 30994 27806
rect 34526 27794 34578 27806
rect 34750 27858 34802 27870
rect 34750 27794 34802 27806
rect 35870 27858 35922 27870
rect 37326 27858 37378 27870
rect 37706 27862 37718 27914
rect 37770 27862 37782 27914
rect 38334 27858 38386 27870
rect 35870 27794 35922 27806
rect 37158 27802 37210 27814
rect 20806 27738 20858 27750
rect 28198 27746 28250 27758
rect 36486 27746 36538 27758
rect 6246 27634 6298 27646
rect 15250 27638 15262 27690
rect 15314 27638 15326 27690
rect 16886 27682 16938 27694
rect 18174 27690 18226 27702
rect 21746 27694 21758 27746
rect 21810 27694 21822 27746
rect 26114 27694 26126 27746
rect 26178 27694 26190 27746
rect 29250 27694 29262 27746
rect 29314 27694 29326 27746
rect 6246 27570 6298 27582
rect 17614 27634 17666 27646
rect 28198 27682 28250 27694
rect 29822 27690 29874 27702
rect 18174 27626 18226 27638
rect 36486 27682 36538 27694
rect 36934 27746 36986 27758
rect 37538 27806 37550 27858
rect 37602 27806 37614 27858
rect 37326 27794 37378 27806
rect 38334 27794 38386 27806
rect 38446 27858 38498 27870
rect 39006 27858 39058 27870
rect 38714 27806 38726 27858
rect 38778 27806 38790 27858
rect 38446 27794 38498 27806
rect 39006 27794 39058 27806
rect 40238 27858 40290 27870
rect 40238 27794 40290 27806
rect 40462 27858 40514 27870
rect 40462 27794 40514 27806
rect 41134 27858 41186 27870
rect 41346 27862 41358 27914
rect 41410 27862 41422 27914
rect 46510 27906 46562 27918
rect 42030 27858 42082 27870
rect 45390 27858 45442 27870
rect 48302 27858 48354 27870
rect 41794 27806 41806 27858
rect 41858 27806 41870 27858
rect 42802 27806 42814 27858
rect 42866 27806 42878 27858
rect 46254 27806 46266 27858
rect 46318 27806 46330 27858
rect 47058 27806 47070 27858
rect 47122 27806 47134 27858
rect 47282 27806 47294 27858
rect 47346 27806 47358 27858
rect 41134 27794 41186 27806
rect 42030 27794 42082 27806
rect 45390 27794 45442 27806
rect 48302 27794 48354 27806
rect 37158 27738 37210 27750
rect 44706 27694 44718 27746
rect 44770 27694 44782 27746
rect 36934 27682 36986 27694
rect 46958 27690 47010 27702
rect 29822 27626 29874 27638
rect 35534 27634 35586 27646
rect 35018 27582 35030 27634
rect 35082 27582 35094 27634
rect 39946 27582 39958 27634
rect 40010 27582 40022 27634
rect 46958 27626 47010 27638
rect 47966 27634 48018 27646
rect 17614 27570 17666 27582
rect 35534 27570 35586 27582
rect 47966 27570 48018 27582
rect 1344 27466 48608 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 48608 27466
rect 1344 27380 48608 27414
rect 14982 27298 15034 27310
rect 5002 27246 5014 27298
rect 5066 27246 5078 27298
rect 12462 27242 12514 27254
rect 7522 27190 7534 27242
rect 7586 27190 7598 27242
rect 9326 27186 9378 27198
rect 2706 27134 2718 27186
rect 2770 27134 2782 27186
rect 9326 27122 9378 27134
rect 11118 27186 11170 27198
rect 14982 27234 15034 27246
rect 23382 27298 23434 27310
rect 28366 27298 28418 27310
rect 26506 27246 26518 27298
rect 26570 27246 26582 27298
rect 27514 27246 27526 27298
rect 27578 27246 27590 27298
rect 33518 27298 33570 27310
rect 41358 27298 41410 27310
rect 12462 27178 12514 27190
rect 18958 27186 19010 27198
rect 20290 27190 20302 27242
rect 20354 27190 20366 27242
rect 23382 27234 23434 27246
rect 28366 27234 28418 27246
rect 30382 27242 30434 27254
rect 24614 27186 24666 27198
rect 11118 27122 11170 27134
rect 14422 27130 14474 27142
rect 18162 27134 18174 27186
rect 18226 27134 18238 27186
rect 21690 27134 21702 27186
rect 21754 27134 21766 27186
rect 3726 27074 3778 27086
rect 2818 27007 2830 27059
rect 2882 27007 2894 27059
rect 3042 27022 3054 27074
rect 3106 27022 3118 27074
rect 3726 27010 3778 27022
rect 3950 27074 4002 27086
rect 4510 27074 4562 27086
rect 4218 27022 4230 27074
rect 4282 27022 4294 27074
rect 3950 27010 4002 27022
rect 4510 27010 4562 27022
rect 4734 27074 4786 27086
rect 4734 27010 4786 27022
rect 5630 27074 5682 27086
rect 8542 27074 8594 27086
rect 6178 27022 6190 27074
rect 6242 27022 6254 27074
rect 5630 27010 5682 27022
rect 7070 26984 7082 27036
rect 7134 26984 7146 27036
rect 7746 27022 7758 27074
rect 7810 27022 7822 27074
rect 8542 27010 8594 27022
rect 8654 27074 8706 27086
rect 13862 27074 13914 27086
rect 9538 27022 9550 27074
rect 9602 27022 9614 27074
rect 9762 27022 9774 27074
rect 9826 27022 9838 27074
rect 10322 27022 10334 27074
rect 10386 27022 10398 27074
rect 10658 27022 10670 27074
rect 10722 27022 10734 27074
rect 8654 27010 8706 27022
rect 10950 27018 11002 27030
rect 11330 27022 11342 27074
rect 11394 27022 11406 27074
rect 12562 27022 12574 27074
rect 12626 27022 12638 27074
rect 12898 27022 12910 27074
rect 12962 27022 12974 27074
rect 11498 26966 11510 27018
rect 11562 26966 11574 27018
rect 13862 27010 13914 27022
rect 14142 27074 14194 27086
rect 18958 27122 19010 27134
rect 24614 27122 24666 27134
rect 25566 27186 25618 27198
rect 36250 27246 36262 27298
rect 36314 27246 36326 27298
rect 45098 27246 45110 27298
rect 45162 27246 45174 27298
rect 33518 27234 33570 27246
rect 30382 27178 30434 27190
rect 35422 27186 35474 27198
rect 25566 27122 25618 27134
rect 35422 27122 35474 27134
rect 38390 27186 38442 27198
rect 38882 27190 38894 27242
rect 38946 27190 38958 27242
rect 41358 27234 41410 27246
rect 38390 27122 38442 27134
rect 48134 27186 48186 27198
rect 48134 27122 48186 27134
rect 14422 27066 14474 27078
rect 14590 27074 14642 27086
rect 15486 27074 15538 27086
rect 18622 27074 18674 27086
rect 21198 27074 21250 27086
rect 14142 27010 14194 27022
rect 14802 27022 14814 27074
rect 14866 27022 14878 27074
rect 16258 27022 16270 27074
rect 16322 27022 16334 27074
rect 14590 27010 14642 27022
rect 15486 27010 15538 27022
rect 18622 27010 18674 27022
rect 19550 26984 19562 27036
rect 19614 26984 19626 27036
rect 20290 27022 20302 27074
rect 20354 27022 20366 27074
rect 21198 27010 21250 27022
rect 21422 27074 21474 27086
rect 21422 27010 21474 27022
rect 22262 27074 22314 27086
rect 26798 27074 26850 27086
rect 22654 27046 22706 27058
rect 22262 27010 22314 27022
rect 22542 27018 22594 27030
rect 8250 26910 8262 26962
rect 8314 26910 8326 26962
rect 10950 26954 11002 26966
rect 14254 26962 14306 26974
rect 22654 26982 22706 26994
rect 22878 27046 22930 27058
rect 22878 26982 22930 26994
rect 23102 27046 23154 27058
rect 24882 27022 24894 27074
rect 24946 27022 24958 27074
rect 25330 27022 25342 27074
rect 25394 27022 25406 27074
rect 25778 27022 25790 27074
rect 25842 27022 25854 27074
rect 26114 27022 26126 27074
rect 26178 27022 26190 27074
rect 26798 27010 26850 27022
rect 27022 27074 27074 27086
rect 27022 27010 27074 27022
rect 27806 27074 27858 27086
rect 27806 27010 27858 27022
rect 27918 27074 27970 27086
rect 27918 27010 27970 27022
rect 28702 27074 28754 27086
rect 29990 27074 30042 27086
rect 31838 27074 31890 27086
rect 35758 27074 35810 27086
rect 28702 27010 28754 27022
rect 29150 27039 29202 27051
rect 23102 26982 23154 26994
rect 29150 26975 29202 26987
rect 29262 27046 29314 27058
rect 29710 27046 29762 27058
rect 29262 26982 29314 26994
rect 29474 26966 29486 27018
rect 29538 26966 29550 27018
rect 30482 27022 30494 27074
rect 30546 27022 30558 27074
rect 30706 27022 30718 27074
rect 30770 27022 30782 27074
rect 31602 27022 31614 27074
rect 31666 27022 31678 27074
rect 32702 27022 32714 27074
rect 32766 27022 32778 27074
rect 29990 27010 30042 27022
rect 31838 27010 31890 27022
rect 33798 27018 33850 27030
rect 29710 26982 29762 26994
rect 22542 26954 22594 26966
rect 32958 26962 33010 26974
rect 6066 26854 6078 26906
rect 6130 26854 6142 26906
rect 14254 26898 14306 26910
rect 31446 26906 31498 26918
rect 33954 26992 33966 27044
rect 34018 26992 34030 27044
rect 34862 27036 34914 27048
rect 34178 26983 34190 27035
rect 34242 26983 34254 27035
rect 35186 27022 35198 27074
rect 35250 27022 35262 27074
rect 34862 26972 34914 26984
rect 35590 27018 35642 27030
rect 33798 26954 33850 26966
rect 35758 27010 35810 27022
rect 35982 27074 36034 27086
rect 35982 27010 36034 27022
rect 37942 27074 37994 27086
rect 39342 27074 39394 27086
rect 38770 27022 38782 27074
rect 38834 27022 38846 27074
rect 39106 27022 39118 27074
rect 39170 27022 39182 27074
rect 37942 27010 37994 27022
rect 39342 27010 39394 27022
rect 39566 27074 39618 27086
rect 43822 27074 43874 27086
rect 39566 27010 39618 27022
rect 40338 26994 40350 27046
rect 40402 26994 40414 27046
rect 43138 27022 43150 27074
rect 43202 27022 43214 27074
rect 43474 26966 43486 27018
rect 43538 26966 43550 27018
rect 43822 27010 43874 27022
rect 45390 27074 45442 27086
rect 45390 27010 45442 27022
rect 45614 27074 45666 27086
rect 45614 27010 45666 27022
rect 46174 27074 46226 27086
rect 47070 27074 47122 27086
rect 46834 27022 46846 27074
rect 46898 27022 46910 27074
rect 46174 27010 46226 27022
rect 46386 26966 46398 27018
rect 46450 26966 46462 27018
rect 47070 27010 47122 27022
rect 47294 27074 47346 27086
rect 47294 27010 47346 27022
rect 35590 26954 35642 26966
rect 39834 26910 39846 26962
rect 39898 26910 39910 26962
rect 47562 26910 47574 26962
rect 47626 26910 47638 26962
rect 32958 26898 33010 26910
rect 31446 26842 31498 26854
rect 37494 26850 37546 26862
rect 43362 26854 43374 26906
rect 43426 26854 43438 26906
rect 46610 26854 46622 26906
rect 46674 26854 46686 26906
rect 37494 26786 37546 26798
rect 1344 26682 48608 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 48608 26682
rect 1344 26596 48608 26630
rect 10278 26514 10330 26526
rect 10278 26450 10330 26462
rect 10782 26514 10834 26526
rect 10782 26450 10834 26462
rect 15374 26514 15426 26526
rect 15374 26450 15426 26462
rect 16606 26514 16658 26526
rect 16606 26450 16658 26462
rect 20638 26514 20690 26526
rect 4080 26402 4132 26414
rect 4080 26338 4132 26350
rect 8318 26402 8370 26414
rect 19730 26406 19742 26458
rect 19794 26406 19806 26458
rect 20638 26450 20690 26462
rect 21310 26514 21362 26526
rect 21310 26450 21362 26462
rect 21982 26514 22034 26526
rect 21982 26450 22034 26462
rect 27470 26514 27522 26526
rect 27470 26450 27522 26462
rect 31670 26514 31722 26526
rect 26070 26402 26122 26414
rect 29138 26406 29150 26458
rect 29202 26406 29214 26458
rect 31670 26450 31722 26462
rect 32118 26514 32170 26526
rect 32118 26450 32170 26462
rect 32566 26514 32618 26526
rect 32566 26450 32618 26462
rect 34582 26514 34634 26526
rect 34582 26450 34634 26462
rect 40070 26514 40122 26526
rect 40070 26450 40122 26462
rect 41918 26514 41970 26526
rect 41918 26450 41970 26462
rect 33966 26402 34018 26414
rect 11722 26350 11734 26402
rect 11786 26350 11798 26402
rect 23482 26350 23494 26402
rect 23546 26350 23558 26402
rect 29978 26350 29990 26402
rect 30042 26350 30054 26402
rect 1598 26290 1650 26302
rect 1598 26226 1650 26238
rect 3166 26290 3218 26302
rect 3838 26290 3890 26302
rect 3166 26226 3218 26238
rect 3334 26234 3386 26246
rect 2550 26178 2602 26190
rect 4834 26238 4846 26290
rect 4898 26238 4910 26290
rect 5170 26238 5182 26290
rect 5234 26238 5246 26290
rect 5730 26238 5742 26290
rect 5794 26238 5806 26290
rect 5954 26253 5966 26305
rect 6018 26253 6030 26305
rect 6962 26294 6974 26346
rect 7026 26294 7038 26346
rect 7522 26294 7534 26346
rect 7586 26294 7598 26346
rect 8318 26338 8370 26350
rect 8530 26294 8542 26346
rect 8594 26294 8606 26346
rect 12294 26319 12346 26331
rect 11118 26290 11170 26302
rect 8082 26238 8094 26290
rect 8146 26238 8158 26290
rect 9426 26238 9438 26290
rect 9490 26238 9502 26290
rect 10434 26238 10446 26290
rect 10498 26238 10510 26290
rect 3838 26226 3890 26238
rect 11118 26226 11170 26238
rect 11230 26290 11282 26302
rect 11230 26226 11282 26238
rect 11454 26290 11506 26302
rect 12294 26255 12346 26267
rect 12450 26238 12462 26290
rect 12514 26238 12526 26290
rect 12830 26276 12842 26328
rect 12894 26276 12906 26328
rect 14288 26327 14340 26339
rect 14030 26290 14082 26302
rect 13570 26238 13582 26290
rect 13634 26238 13646 26290
rect 14130 26238 14142 26290
rect 14194 26238 14206 26290
rect 18324 26327 18376 26339
rect 14288 26263 14340 26275
rect 15038 26290 15090 26302
rect 11454 26226 11506 26238
rect 14030 26226 14082 26238
rect 15038 26226 15090 26238
rect 16942 26290 16994 26302
rect 25230 26325 25282 26337
rect 18622 26290 18674 26302
rect 18324 26263 18376 26275
rect 18498 26238 18510 26290
rect 18562 26238 18574 26290
rect 16942 26226 16994 26238
rect 18622 26226 18674 26238
rect 18958 26290 19010 26302
rect 20302 26290 20354 26302
rect 19618 26238 19630 26290
rect 19682 26238 19694 26290
rect 18958 26226 19010 26238
rect 20302 26226 20354 26238
rect 20974 26290 21026 26302
rect 20974 26226 21026 26238
rect 21646 26290 21698 26302
rect 21646 26226 21698 26238
rect 23774 26290 23826 26302
rect 23774 26226 23826 26238
rect 23998 26290 24050 26302
rect 24322 26238 24334 26290
rect 24386 26238 24398 26290
rect 24546 26238 24558 26290
rect 24610 26238 24622 26290
rect 25330 26294 25342 26346
rect 25394 26294 25406 26346
rect 25554 26294 25566 26346
rect 25618 26294 25630 26346
rect 25778 26294 25790 26346
rect 25842 26294 25854 26346
rect 26070 26338 26122 26350
rect 33014 26346 33066 26358
rect 27134 26290 27186 26302
rect 28970 26294 28982 26346
rect 29034 26294 29046 26346
rect 29486 26290 29538 26302
rect 25230 26261 25282 26273
rect 26562 26238 26574 26290
rect 26626 26238 26638 26290
rect 26898 26238 26910 26290
rect 26962 26238 26974 26290
rect 28018 26238 28030 26290
rect 28082 26238 28094 26290
rect 28354 26238 28366 26290
rect 28418 26238 28430 26290
rect 29250 26238 29262 26290
rect 29314 26238 29326 26290
rect 23998 26226 24050 26238
rect 27134 26226 27186 26238
rect 29486 26226 29538 26238
rect 29710 26290 29762 26302
rect 29710 26226 29762 26238
rect 30830 26290 30882 26302
rect 33966 26338 34018 26350
rect 35086 26402 35138 26414
rect 45166 26402 45218 26414
rect 40954 26350 40966 26402
rect 41018 26350 41030 26402
rect 45994 26350 46006 26402
rect 46058 26350 46070 26402
rect 35086 26338 35138 26350
rect 45166 26338 45218 26350
rect 47798 26346 47850 26358
rect 30930 26238 30942 26290
rect 30994 26238 31006 26290
rect 33014 26282 33066 26294
rect 33170 26268 33182 26320
rect 33234 26268 33246 26320
rect 33506 26268 33518 26320
rect 33570 26268 33582 26320
rect 47406 26318 47458 26330
rect 37774 26290 37826 26302
rect 30830 26226 30882 26238
rect 37774 26226 37826 26238
rect 38166 26290 38218 26302
rect 38166 26226 38218 26238
rect 38894 26290 38946 26302
rect 38894 26226 38946 26238
rect 39118 26290 39170 26302
rect 39118 26226 39170 26238
rect 39230 26290 39282 26302
rect 39230 26226 39282 26238
rect 41246 26290 41298 26302
rect 41246 26226 41298 26238
rect 41358 26290 41410 26302
rect 41358 26226 41410 26238
rect 41582 26290 41634 26302
rect 41582 26226 41634 26238
rect 42478 26290 42530 26302
rect 42478 26226 42530 26238
rect 45502 26290 45554 26302
rect 45502 26226 45554 26238
rect 45726 26290 45778 26302
rect 45726 26226 45778 26238
rect 46286 26290 46338 26302
rect 47406 26254 47458 26266
rect 47630 26318 47682 26330
rect 47798 26282 47850 26294
rect 47966 26325 48018 26337
rect 47630 26254 47682 26266
rect 47966 26261 48018 26273
rect 46286 26226 46338 26238
rect 3334 26170 3386 26182
rect 14702 26178 14754 26190
rect 2550 26114 2602 26126
rect 5294 26122 5346 26134
rect 6066 26126 6078 26178
rect 6130 26126 6142 26178
rect 12114 26126 12126 26178
rect 12178 26126 12190 26178
rect 1934 26066 1986 26078
rect 5294 26058 5346 26070
rect 9606 26066 9658 26078
rect 13458 26070 13470 26122
rect 13522 26070 13534 26122
rect 14702 26114 14754 26126
rect 16214 26178 16266 26190
rect 16214 26114 16266 26126
rect 17558 26178 17610 26190
rect 17558 26114 17610 26126
rect 17950 26178 18002 26190
rect 17950 26114 18002 26126
rect 22598 26178 22650 26190
rect 30494 26178 30546 26190
rect 22598 26114 22650 26126
rect 26462 26122 26514 26134
rect 24434 26070 24446 26122
rect 24498 26070 24510 26122
rect 1934 26002 1986 26014
rect 26462 26058 26514 26070
rect 28478 26122 28530 26134
rect 36978 26126 36990 26178
rect 37042 26126 37054 26178
rect 39498 26126 39510 26178
rect 39562 26126 39574 26178
rect 43250 26126 43262 26178
rect 43314 26126 43326 26178
rect 30494 26114 30546 26126
rect 28478 26058 28530 26070
rect 31110 26066 31162 26078
rect 9606 26002 9658 26014
rect 31110 26002 31162 26014
rect 38558 26066 38610 26078
rect 38558 26002 38610 26014
rect 46622 26066 46674 26078
rect 46622 26002 46674 26014
rect 47126 26066 47178 26078
rect 47126 26002 47178 26014
rect 1344 25898 48608 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 48608 25898
rect 1344 25812 48608 25846
rect 5854 25730 5906 25742
rect 2650 25678 2662 25730
rect 2714 25678 2726 25730
rect 3726 25618 3778 25630
rect 4834 25622 4846 25674
rect 4898 25622 4910 25674
rect 5854 25666 5906 25678
rect 8822 25730 8874 25742
rect 8822 25666 8874 25678
rect 10334 25730 10386 25742
rect 10334 25666 10386 25678
rect 13564 25730 13616 25742
rect 26798 25730 26850 25742
rect 34190 25730 34242 25742
rect 13564 25666 13616 25678
rect 14814 25674 14866 25686
rect 3726 25554 3778 25566
rect 6862 25618 6914 25630
rect 29530 25678 29542 25730
rect 29594 25678 29606 25730
rect 26798 25666 26850 25678
rect 14814 25610 14866 25622
rect 19518 25618 19570 25630
rect 28018 25622 28030 25674
rect 28082 25622 28094 25674
rect 34190 25666 34242 25678
rect 44046 25730 44098 25742
rect 45210 25678 45222 25730
rect 45274 25678 45286 25730
rect 46778 25678 46790 25730
rect 46842 25678 46854 25730
rect 47674 25678 47686 25730
rect 47738 25678 47750 25730
rect 44046 25666 44098 25678
rect 18386 25566 18398 25618
rect 18450 25566 18462 25618
rect 6862 25554 6914 25566
rect 19518 25554 19570 25566
rect 30830 25618 30882 25630
rect 48246 25618 48298 25630
rect 30830 25554 30882 25566
rect 35478 25562 35530 25574
rect 38434 25566 38446 25618
rect 38498 25566 38510 25618
rect 40338 25566 40350 25618
rect 40402 25566 40414 25618
rect 41458 25566 41470 25618
rect 41522 25566 41534 25618
rect 45602 25566 45614 25618
rect 45666 25566 45678 25618
rect 2270 25506 2322 25518
rect 2270 25442 2322 25454
rect 2382 25506 2434 25518
rect 5518 25506 5570 25518
rect 8094 25506 8146 25518
rect 2382 25442 2434 25454
rect 3166 25450 3218 25462
rect 3490 25454 3502 25506
rect 3554 25454 3566 25506
rect 3166 25386 3218 25398
rect 3894 25450 3946 25462
rect 4094 25416 4106 25468
rect 4158 25416 4170 25468
rect 4834 25454 4846 25506
rect 4898 25454 4910 25506
rect 6290 25454 6302 25506
rect 6354 25454 6366 25506
rect 6626 25454 6638 25506
rect 6690 25454 6702 25506
rect 7074 25454 7086 25506
rect 7138 25454 7150 25506
rect 7522 25454 7534 25506
rect 7586 25454 7598 25506
rect 5518 25442 5570 25454
rect 8094 25442 8146 25454
rect 8542 25506 8594 25518
rect 8250 25398 8262 25450
rect 8314 25398 8326 25450
rect 8542 25442 8594 25454
rect 9214 25506 9266 25518
rect 9214 25442 9266 25454
rect 13806 25506 13858 25518
rect 3894 25386 3946 25398
rect 8430 25394 8482 25406
rect 10078 25398 10090 25450
rect 10142 25398 10154 25450
rect 11442 25398 11454 25450
rect 11506 25398 11518 25450
rect 12114 25398 12126 25450
rect 12178 25398 12190 25450
rect 12674 25398 12686 25450
rect 12738 25398 12750 25450
rect 13806 25442 13858 25454
rect 14310 25506 14362 25518
rect 15710 25506 15762 25518
rect 18846 25506 18898 25518
rect 19854 25506 19906 25518
rect 14914 25454 14926 25506
rect 14978 25454 14990 25506
rect 15138 25454 15150 25506
rect 15202 25454 15214 25506
rect 16482 25454 16494 25506
rect 16546 25454 16558 25506
rect 18946 25454 18958 25506
rect 19010 25454 19022 25506
rect 14310 25442 14362 25454
rect 15710 25442 15762 25454
rect 18846 25442 18898 25454
rect 8430 25330 8482 25342
rect 14478 25394 14530 25406
rect 19112 25398 19124 25450
rect 19176 25398 19188 25450
rect 19854 25442 19906 25454
rect 21534 25506 21586 25518
rect 29038 25506 29090 25518
rect 22306 25454 22318 25506
rect 22370 25454 22382 25506
rect 21534 25442 21586 25454
rect 25106 25426 25118 25478
rect 25170 25426 25182 25478
rect 27906 25454 27918 25506
rect 27970 25454 27982 25506
rect 28242 25454 28254 25506
rect 28306 25454 28318 25506
rect 29038 25442 29090 25454
rect 29262 25506 29314 25518
rect 33070 25506 33122 25518
rect 34626 25510 34638 25562
rect 34690 25510 34702 25562
rect 48246 25554 48298 25566
rect 31042 25454 31054 25506
rect 31106 25454 31118 25506
rect 35478 25498 35530 25510
rect 35646 25506 35698 25518
rect 29262 25442 29314 25454
rect 11890 25286 11902 25338
rect 11954 25286 11966 25338
rect 14478 25330 14530 25342
rect 20806 25394 20858 25406
rect 20806 25330 20858 25342
rect 24222 25394 24274 25406
rect 30482 25398 30494 25450
rect 30546 25398 30558 25450
rect 31602 25398 31614 25450
rect 31666 25398 31678 25450
rect 32162 25398 32174 25450
rect 32226 25398 32238 25450
rect 33070 25442 33122 25454
rect 34750 25468 34802 25480
rect 33934 25398 33946 25450
rect 33998 25398 34010 25450
rect 35646 25442 35698 25454
rect 35870 25506 35922 25518
rect 36878 25506 36930 25518
rect 36138 25454 36150 25506
rect 36202 25454 36214 25506
rect 35870 25442 35922 25454
rect 36878 25442 36930 25454
rect 37662 25506 37714 25518
rect 37662 25442 37714 25454
rect 40686 25506 40738 25518
rect 40686 25442 40738 25454
rect 43710 25506 43762 25518
rect 43710 25442 43762 25454
rect 44718 25506 44770 25518
rect 44718 25442 44770 25454
rect 44942 25506 44994 25518
rect 46398 25506 46450 25518
rect 46050 25454 46062 25506
rect 46114 25454 46126 25506
rect 44942 25442 44994 25454
rect 34750 25404 34802 25416
rect 24222 25330 24274 25342
rect 35310 25394 35362 25406
rect 35310 25330 35362 25342
rect 43374 25394 43426 25406
rect 45770 25398 45782 25450
rect 45834 25398 45846 25450
rect 46398 25442 46450 25454
rect 46510 25506 46562 25518
rect 46510 25442 46562 25454
rect 47182 25506 47234 25518
rect 47182 25442 47234 25454
rect 47406 25506 47458 25518
rect 47406 25442 47458 25454
rect 43374 25330 43426 25342
rect 20190 25282 20242 25294
rect 20190 25218 20242 25230
rect 24838 25282 24890 25294
rect 24838 25218 24890 25230
rect 37214 25282 37266 25294
rect 37214 25218 37266 25230
rect 1344 25114 48608 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 48608 25114
rect 1344 25028 48608 25062
rect 2158 24946 2210 24958
rect 2158 24882 2210 24894
rect 15486 24946 15538 24958
rect 15486 24882 15538 24894
rect 17502 24946 17554 24958
rect 17502 24882 17554 24894
rect 22654 24946 22706 24958
rect 22654 24882 22706 24894
rect 35254 24946 35306 24958
rect 35254 24882 35306 24894
rect 38894 24946 38946 24958
rect 38894 24882 38946 24894
rect 44326 24946 44378 24958
rect 5406 24834 5458 24846
rect 8542 24834 8594 24846
rect 12126 24834 12178 24846
rect 2494 24722 2546 24734
rect 2494 24658 2546 24670
rect 3166 24722 3218 24734
rect 3166 24658 3218 24670
rect 3390 24722 3442 24734
rect 3390 24658 3442 24670
rect 3558 24722 3610 24734
rect 3558 24658 3610 24670
rect 4062 24722 4114 24734
rect 4834 24726 4846 24778
rect 4898 24726 4910 24778
rect 5406 24770 5458 24782
rect 7982 24778 8034 24790
rect 6514 24726 6526 24778
rect 6578 24726 6590 24778
rect 6962 24726 6974 24778
rect 7026 24726 7038 24778
rect 9930 24782 9942 24834
rect 9994 24782 10006 24834
rect 8542 24770 8594 24782
rect 12126 24770 12178 24782
rect 21982 24834 22034 24846
rect 5618 24670 5630 24722
rect 5682 24670 5694 24722
rect 7982 24714 8034 24726
rect 8710 24722 8762 24734
rect 8306 24670 8318 24722
rect 8370 24670 8382 24722
rect 4062 24658 4114 24670
rect 8710 24658 8762 24670
rect 9438 24722 9490 24734
rect 9438 24658 9490 24670
rect 9662 24722 9714 24734
rect 12238 24722 12290 24734
rect 10770 24670 10782 24722
rect 10834 24670 10846 24722
rect 10994 24670 11006 24722
rect 11058 24670 11070 24722
rect 11442 24670 11454 24722
rect 11506 24670 11518 24722
rect 11778 24670 11790 24722
rect 11842 24670 11854 24722
rect 12562 24670 12574 24722
rect 12626 24670 12638 24722
rect 13682 24670 13694 24722
rect 13746 24670 13758 24722
rect 14358 24708 14370 24760
rect 14422 24708 14434 24760
rect 18548 24759 18600 24771
rect 21982 24770 22034 24782
rect 24558 24834 24610 24846
rect 26350 24834 26402 24846
rect 24558 24770 24610 24782
rect 25790 24778 25842 24790
rect 15150 24722 15202 24734
rect 9662 24658 9714 24670
rect 12238 24658 12290 24670
rect 15150 24658 15202 24670
rect 16046 24722 16098 24734
rect 16046 24658 16098 24670
rect 17838 24722 17890 24734
rect 18846 24722 18898 24734
rect 18548 24695 18600 24707
rect 18722 24670 18734 24722
rect 18786 24670 18798 24722
rect 17838 24658 17890 24670
rect 18846 24658 18898 24670
rect 19294 24722 19346 24734
rect 22318 24722 22370 24734
rect 20066 24670 20078 24722
rect 20130 24670 20142 24722
rect 19294 24658 19346 24670
rect 22318 24658 22370 24670
rect 23662 24722 23714 24734
rect 24098 24698 24110 24750
rect 24162 24698 24174 24750
rect 24726 24722 24778 24734
rect 31334 24834 31386 24846
rect 35646 24834 35698 24846
rect 41570 24838 41582 24890
rect 41634 24838 41646 24890
rect 44326 24882 44378 24894
rect 26350 24770 26402 24782
rect 30419 24778 30471 24790
rect 31110 24778 31162 24790
rect 24322 24670 24334 24722
rect 24386 24670 24398 24722
rect 25442 24670 25454 24722
rect 25506 24670 25518 24722
rect 25790 24714 25842 24726
rect 26518 24722 26570 24734
rect 27806 24722 27858 24734
rect 30594 24726 30606 24778
rect 30658 24726 30670 24778
rect 30886 24757 30938 24769
rect 27010 24670 27022 24722
rect 27074 24670 27086 24722
rect 27458 24670 27470 24722
rect 27522 24670 27534 24722
rect 28242 24670 28254 24722
rect 28306 24670 28318 24722
rect 29138 24670 29150 24722
rect 29202 24670 29214 24722
rect 29474 24670 29486 24722
rect 29538 24670 29550 24722
rect 30419 24714 30471 24726
rect 34682 24782 34694 24834
rect 34746 24782 34758 24834
rect 31334 24770 31386 24782
rect 35646 24770 35698 24782
rect 48078 24834 48130 24846
rect 41358 24761 41410 24773
rect 48078 24770 48130 24782
rect 31110 24714 31162 24726
rect 34302 24722 34354 24734
rect 30886 24693 30938 24705
rect 31826 24670 31838 24722
rect 31890 24670 31902 24722
rect 32050 24670 32062 24722
rect 32114 24670 32126 24722
rect 33170 24670 33182 24722
rect 33234 24670 33246 24722
rect 33394 24670 33406 24722
rect 33458 24670 33470 24722
rect 23662 24658 23714 24670
rect 24726 24658 24778 24670
rect 4304 24610 4356 24622
rect 18174 24610 18226 24622
rect 25666 24614 25678 24666
rect 25730 24614 25742 24666
rect 26518 24658 26570 24670
rect 27806 24658 27858 24670
rect 34302 24658 34354 24670
rect 34414 24722 34466 24734
rect 38334 24722 38386 24734
rect 37538 24670 37550 24722
rect 37602 24670 37614 24722
rect 34414 24658 34466 24670
rect 38334 24658 38386 24670
rect 38558 24722 38610 24734
rect 38558 24658 38610 24670
rect 40126 24722 40178 24734
rect 40898 24670 40910 24722
rect 40962 24670 40974 24722
rect 41358 24697 41410 24709
rect 41582 24722 41634 24734
rect 42242 24714 42254 24766
rect 42306 24714 42318 24766
rect 43262 24722 43314 24734
rect 42466 24670 42478 24722
rect 42530 24670 42542 24722
rect 40126 24658 40178 24670
rect 41582 24658 41634 24670
rect 43262 24658 43314 24670
rect 43374 24722 43426 24734
rect 43374 24658 43426 24670
rect 43878 24722 43930 24734
rect 44818 24670 44830 24722
rect 44882 24670 44894 24722
rect 45042 24685 45054 24737
rect 45106 24685 45118 24737
rect 45390 24722 45442 24734
rect 46162 24670 46174 24722
rect 46226 24670 46238 24722
rect 43878 24658 43930 24670
rect 45390 24658 45442 24670
rect 28870 24610 28922 24622
rect 4304 24546 4356 24558
rect 13582 24554 13634 24566
rect 2830 24498 2882 24510
rect 10882 24502 10894 24554
rect 10946 24502 10958 24554
rect 18174 24546 18226 24558
rect 25286 24554 25338 24566
rect 28018 24558 28030 24610
rect 28082 24558 28094 24610
rect 13582 24490 13634 24502
rect 16382 24498 16434 24510
rect 2830 24434 2882 24446
rect 16382 24434 16434 24446
rect 23326 24498 23378 24510
rect 28870 24546 28922 24558
rect 30214 24610 30266 24622
rect 34022 24610 34074 24622
rect 29250 24502 29262 24554
rect 29314 24502 29326 24554
rect 30214 24546 30266 24558
rect 33070 24554 33122 24566
rect 31938 24502 31950 24554
rect 32002 24502 32014 24554
rect 42130 24558 42142 24610
rect 42194 24558 42206 24610
rect 45154 24558 45166 24610
rect 45218 24558 45230 24610
rect 34022 24546 34074 24558
rect 25286 24490 25338 24502
rect 33070 24490 33122 24502
rect 39790 24498 39842 24510
rect 23326 24434 23378 24446
rect 42970 24446 42982 24498
rect 43034 24446 43046 24498
rect 39790 24434 39842 24446
rect 1344 24330 48608 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 48608 24330
rect 1344 24244 48608 24278
rect 8430 24162 8482 24174
rect 3390 24106 3442 24118
rect 8430 24098 8482 24110
rect 11454 24162 11506 24174
rect 3390 24042 3442 24054
rect 4398 24050 4450 24062
rect 9202 24054 9214 24106
rect 9266 24054 9278 24106
rect 11454 24098 11506 24110
rect 11996 24162 12048 24174
rect 11996 24098 12048 24110
rect 38222 24162 38274 24174
rect 14242 24054 14254 24106
rect 14306 24054 14318 24106
rect 22374 24050 22426 24062
rect 26562 24054 26574 24106
rect 26626 24054 26638 24106
rect 28466 24054 28478 24106
rect 28530 24054 28542 24106
rect 29474 24054 29486 24106
rect 29538 24054 29550 24106
rect 38222 24098 38274 24110
rect 38894 24162 38946 24174
rect 38894 24098 38946 24110
rect 42086 24050 42138 24062
rect 15138 23998 15150 24050
rect 15202 23998 15214 24050
rect 17042 23998 17054 24050
rect 17106 23998 17118 24050
rect 20626 23998 20638 24050
rect 20690 23998 20702 24050
rect 36978 23998 36990 24050
rect 37042 23998 37054 24050
rect 41122 23998 41134 24050
rect 41186 23998 41198 24050
rect 4398 23986 4450 23998
rect 22374 23986 22426 23998
rect 42086 23986 42138 23998
rect 42534 24050 42586 24062
rect 42914 23998 42926 24050
rect 42978 23998 42990 24050
rect 42534 23986 42586 23998
rect 2382 23938 2434 23950
rect 7758 23938 7810 23950
rect 8036 23938 8088 23950
rect 10110 23938 10162 23950
rect 2382 23874 2434 23886
rect 2590 23848 2602 23900
rect 2654 23848 2666 23900
rect 3266 23886 3278 23938
rect 3330 23886 3342 23938
rect 3938 23858 3950 23910
rect 4002 23858 4014 23910
rect 4162 23886 4174 23938
rect 4226 23886 4238 23938
rect 4566 23882 4618 23894
rect 7858 23886 7870 23938
rect 7922 23886 7934 23938
rect 8866 23886 8878 23938
rect 8930 23886 8942 23938
rect 9202 23886 9214 23938
rect 9266 23886 9278 23938
rect 6626 23830 6638 23882
rect 6690 23830 6702 23882
rect 6850 23830 6862 23882
rect 6914 23830 6926 23882
rect 7298 23830 7310 23882
rect 7362 23830 7374 23882
rect 7758 23874 7810 23886
rect 8036 23874 8088 23886
rect 10110 23874 10162 23886
rect 11118 23938 11170 23950
rect 11118 23874 11170 23886
rect 12238 23938 12290 23950
rect 12238 23874 12290 23886
rect 12742 23938 12794 23950
rect 12742 23874 12794 23886
rect 12910 23938 12962 23950
rect 12910 23874 12962 23886
rect 13470 23938 13522 23950
rect 17838 23938 17890 23950
rect 14130 23886 14142 23938
rect 14194 23886 14206 23938
rect 13470 23874 13522 23886
rect 17838 23874 17890 23886
rect 17950 23938 18002 23950
rect 21926 23938 21978 23950
rect 18722 23886 18734 23938
rect 18786 23886 18798 23938
rect 21522 23886 21534 23938
rect 21586 23886 21598 23938
rect 17950 23874 18002 23886
rect 21926 23874 21978 23886
rect 22878 23938 22930 23950
rect 27694 23938 27746 23950
rect 34302 23938 34354 23950
rect 23650 23886 23662 23938
rect 23714 23886 23726 23938
rect 22878 23874 22930 23886
rect 26110 23848 26122 23900
rect 26174 23848 26186 23900
rect 26786 23886 26798 23938
rect 26850 23886 26862 23938
rect 28354 23886 28366 23938
rect 28418 23886 28430 23938
rect 29250 23886 29262 23938
rect 29314 23886 29326 23938
rect 27694 23874 27746 23886
rect 29990 23848 30002 23900
rect 30054 23848 30066 23900
rect 30594 23858 30606 23910
rect 30658 23858 30670 23910
rect 30818 23886 30830 23938
rect 30882 23886 30894 23938
rect 31222 23882 31274 23894
rect 33506 23886 33518 23938
rect 33570 23886 33582 23938
rect 4566 23818 4618 23830
rect 25566 23826 25618 23838
rect 2046 23714 2098 23726
rect 6514 23718 6526 23770
rect 6578 23718 6590 23770
rect 25566 23762 25618 23774
rect 31054 23826 31106 23838
rect 34302 23874 34354 23886
rect 35310 23938 35362 23950
rect 35310 23874 35362 23886
rect 35758 23938 35810 23950
rect 37886 23938 37938 23950
rect 35758 23874 35810 23886
rect 36082 23859 36094 23911
rect 36146 23859 36158 23911
rect 36418 23886 36430 23938
rect 36482 23886 36494 23938
rect 37090 23871 37102 23923
rect 37154 23871 37166 23923
rect 37314 23886 37326 23938
rect 37378 23886 37390 23938
rect 37886 23874 37938 23886
rect 38558 23938 38610 23950
rect 38558 23874 38610 23886
rect 40126 23938 40178 23950
rect 43598 23938 43650 23950
rect 40674 23886 40686 23938
rect 40738 23886 40750 23938
rect 40126 23874 40178 23886
rect 31222 23818 31274 23830
rect 31614 23826 31666 23838
rect 40506 23830 40518 23882
rect 40570 23830 40582 23882
rect 41234 23871 41246 23923
rect 41298 23871 41310 23923
rect 41458 23886 41470 23938
rect 41522 23886 41534 23938
rect 43026 23842 43038 23894
rect 43090 23842 43102 23894
rect 43250 23886 43262 23938
rect 43314 23886 43326 23938
rect 43598 23874 43650 23886
rect 45278 23938 45330 23950
rect 46174 23938 46226 23950
rect 45490 23886 45502 23938
rect 45554 23886 45566 23938
rect 45278 23874 45330 23886
rect 45826 23859 45838 23911
rect 45890 23859 45902 23911
rect 46174 23874 46226 23886
rect 47182 23938 47234 23950
rect 47730 23886 47742 23938
rect 47794 23886 47806 23938
rect 47182 23874 47234 23886
rect 47562 23830 47574 23882
rect 47626 23830 47638 23882
rect 31054 23762 31106 23774
rect 31614 23762 31666 23774
rect 2046 23650 2098 23662
rect 9774 23714 9826 23726
rect 9774 23650 9826 23662
rect 21366 23714 21418 23726
rect 21366 23650 21418 23662
rect 34974 23714 35026 23726
rect 35634 23718 35646 23770
rect 35698 23718 35710 23770
rect 40226 23718 40238 23770
rect 40290 23718 40302 23770
rect 34974 23650 35026 23662
rect 43934 23714 43986 23726
rect 43934 23650 43986 23662
rect 44942 23714 44994 23726
rect 46274 23718 46286 23770
rect 46338 23718 46350 23770
rect 47282 23718 47294 23770
rect 47346 23718 47358 23770
rect 44942 23650 44994 23662
rect 1344 23546 48608 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 48608 23546
rect 1344 23460 48608 23494
rect 17558 23378 17610 23390
rect 4286 23266 4338 23278
rect 5954 23270 5966 23322
rect 6018 23270 6030 23322
rect 4286 23202 4338 23214
rect 8486 23266 8538 23278
rect 12674 23270 12686 23322
rect 12738 23270 12750 23322
rect 17558 23314 17610 23326
rect 17950 23378 18002 23390
rect 17950 23314 18002 23326
rect 24446 23378 24498 23390
rect 24446 23314 24498 23326
rect 26462 23378 26514 23390
rect 26462 23314 26514 23326
rect 34638 23378 34690 23390
rect 34638 23314 34690 23326
rect 39006 23378 39058 23390
rect 39006 23314 39058 23326
rect 39678 23378 39730 23390
rect 39678 23314 39730 23326
rect 40294 23378 40346 23390
rect 40294 23314 40346 23326
rect 1598 23154 1650 23166
rect 5518 23154 5570 23166
rect 5730 23158 5742 23210
rect 5794 23158 5806 23210
rect 8486 23202 8538 23214
rect 25790 23266 25842 23278
rect 31614 23266 31666 23278
rect 30314 23214 30326 23266
rect 30378 23214 30390 23266
rect 33966 23266 34018 23278
rect 45714 23270 45726 23322
rect 45778 23270 45790 23322
rect 19036 23191 19088 23203
rect 4610 23102 4622 23154
rect 4674 23102 4686 23154
rect 6066 23102 6078 23154
rect 6130 23102 6142 23154
rect 6514 23102 6526 23154
rect 6578 23102 6590 23154
rect 6850 23129 6862 23181
rect 6914 23129 6926 23181
rect 7198 23154 7250 23166
rect 1598 23090 1650 23102
rect 5518 23090 5570 23102
rect 7198 23090 7250 23102
rect 7758 23154 7810 23166
rect 8206 23154 8258 23166
rect 7758 23090 7810 23102
rect 7926 23098 7978 23110
rect 8082 23102 8094 23154
rect 8146 23102 8158 23154
rect 8206 23090 8258 23102
rect 9438 23154 9490 23166
rect 13358 23154 13410 23166
rect 10210 23102 10222 23154
rect 10274 23102 10286 23154
rect 12674 23102 12686 23154
rect 12738 23102 12750 23154
rect 9438 23090 9490 23102
rect 13358 23090 13410 23102
rect 13918 23154 13970 23166
rect 14198 23154 14250 23166
rect 14018 23102 14030 23154
rect 14082 23102 14094 23154
rect 13918 23090 13970 23102
rect 14198 23090 14250 23102
rect 16440 23154 16492 23166
rect 16718 23154 16770 23166
rect 16594 23102 16606 23154
rect 16658 23102 16670 23154
rect 16440 23090 16492 23102
rect 16718 23090 16770 23102
rect 18286 23154 18338 23166
rect 22468 23191 22520 23203
rect 19294 23154 19346 23166
rect 19036 23127 19088 23139
rect 19170 23102 19182 23154
rect 19234 23102 19246 23154
rect 18286 23090 18338 23102
rect 19294 23090 19346 23102
rect 20414 23154 20466 23166
rect 20414 23090 20466 23102
rect 21086 23154 21138 23166
rect 21086 23090 21138 23102
rect 21198 23154 21250 23166
rect 21198 23090 21250 23102
rect 21534 23154 21586 23166
rect 23628 23191 23680 23203
rect 25790 23202 25842 23214
rect 31614 23202 31666 23214
rect 33014 23210 33066 23222
rect 40954 23214 40966 23266
rect 41018 23214 41030 23266
rect 46890 23214 46902 23266
rect 46954 23214 46966 23266
rect 48010 23214 48022 23266
rect 48074 23214 48086 23266
rect 22766 23154 22818 23166
rect 22468 23127 22520 23139
rect 22642 23102 22654 23154
rect 22706 23102 22718 23154
rect 23886 23154 23938 23166
rect 23628 23127 23680 23139
rect 23762 23102 23774 23154
rect 23826 23102 23838 23154
rect 21534 23090 21586 23102
rect 22766 23090 22818 23102
rect 23886 23090 23938 23102
rect 24110 23154 24162 23166
rect 24110 23090 24162 23102
rect 26126 23154 26178 23166
rect 26126 23090 26178 23102
rect 26798 23154 26850 23166
rect 26798 23090 26850 23102
rect 26910 23154 26962 23166
rect 27950 23140 27962 23192
rect 28014 23140 28026 23192
rect 29934 23154 29986 23166
rect 28690 23102 28702 23154
rect 28754 23102 28766 23154
rect 29250 23102 29262 23154
rect 29314 23102 29326 23154
rect 29474 23102 29486 23154
rect 29538 23102 29550 23154
rect 26910 23090 26962 23102
rect 29934 23090 29986 23102
rect 30046 23154 30098 23166
rect 30046 23090 30098 23102
rect 30998 23154 31050 23166
rect 30998 23090 31050 23102
rect 31278 23154 31330 23166
rect 31726 23154 31778 23166
rect 31278 23090 31330 23102
rect 31446 23098 31498 23110
rect 2370 22990 2382 23042
rect 2434 22990 2446 23042
rect 6738 22990 6750 23042
rect 6802 22990 6814 23042
rect 7926 23034 7978 23046
rect 16046 23042 16098 23054
rect 12114 22990 12126 23042
rect 12178 22990 12190 23042
rect 16046 22978 16098 22990
rect 18622 23042 18674 23054
rect 18622 22978 18674 22990
rect 22094 23042 22146 23054
rect 33170 23158 33182 23210
rect 33234 23158 33246 23210
rect 33966 23202 34018 23214
rect 46062 23193 46114 23205
rect 33014 23146 33066 23158
rect 33394 23141 33406 23193
rect 33458 23141 33470 23193
rect 34302 23154 34354 23166
rect 31726 23090 31778 23102
rect 34302 23090 34354 23102
rect 34974 23154 35026 23166
rect 37998 23154 38050 23166
rect 35746 23102 35758 23154
rect 35810 23102 35822 23154
rect 34974 23090 35026 23102
rect 37998 23090 38050 23102
rect 38670 23154 38722 23166
rect 38670 23090 38722 23102
rect 39342 23154 39394 23166
rect 39342 23090 39394 23102
rect 41246 23154 41298 23166
rect 41246 23090 41298 23102
rect 41470 23154 41522 23166
rect 41470 23090 41522 23102
rect 42142 23154 42194 23166
rect 44830 23154 44882 23166
rect 44034 23102 44046 23154
rect 44098 23102 44110 23154
rect 45602 23102 45614 23154
rect 45666 23102 45678 23154
rect 46062 23129 46114 23141
rect 46286 23154 46338 23166
rect 42142 23090 42194 23102
rect 44830 23090 44882 23102
rect 46286 23090 46338 23102
rect 47182 23154 47234 23166
rect 47182 23090 47234 23102
rect 47406 23154 47458 23166
rect 47406 23090 47458 23102
rect 47630 23154 47682 23166
rect 47630 23090 47682 23102
rect 47742 23154 47794 23166
rect 47742 23090 47794 23102
rect 31446 23034 31498 23046
rect 32566 23042 32618 23054
rect 45222 23042 45274 23054
rect 22094 22978 22146 22990
rect 28814 22986 28866 22998
rect 37650 22990 37662 23042
rect 37714 22990 37726 23042
rect 4790 22930 4842 22942
rect 4790 22866 4842 22878
rect 14590 22930 14642 22942
rect 14590 22866 14642 22878
rect 20078 22930 20130 22942
rect 20078 22866 20130 22878
rect 20750 22930 20802 22942
rect 20750 22866 20802 22878
rect 23214 22930 23266 22942
rect 23214 22866 23266 22878
rect 27246 22930 27298 22942
rect 29474 22934 29486 22986
rect 29538 22934 29550 22986
rect 32566 22978 32618 22990
rect 45222 22978 45274 22990
rect 28814 22922 28866 22934
rect 32006 22930 32058 22942
rect 27246 22866 27298 22878
rect 32006 22866 32058 22878
rect 38334 22930 38386 22942
rect 38334 22866 38386 22878
rect 1344 22762 48608 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 48608 22762
rect 1344 22676 48608 22710
rect 3894 22594 3946 22606
rect 3894 22530 3946 22542
rect 5854 22594 5906 22606
rect 5854 22530 5906 22542
rect 6974 22594 7026 22606
rect 6974 22530 7026 22542
rect 7646 22594 7698 22606
rect 7646 22530 7698 22542
rect 11230 22594 11282 22606
rect 14702 22594 14754 22606
rect 11230 22530 11282 22542
rect 12574 22538 12626 22550
rect 4958 22482 5010 22494
rect 14702 22530 14754 22542
rect 16382 22594 16434 22606
rect 16382 22530 16434 22542
rect 18342 22594 18394 22606
rect 18342 22530 18394 22542
rect 20414 22594 20466 22606
rect 3334 22426 3386 22438
rect 2830 22370 2882 22382
rect 2146 22318 2158 22370
rect 2210 22318 2222 22370
rect 2830 22306 2882 22318
rect 3166 22370 3218 22382
rect 4958 22418 5010 22430
rect 5126 22426 5178 22438
rect 9090 22430 9102 22482
rect 9154 22430 9166 22482
rect 12574 22474 12626 22486
rect 14142 22482 14194 22494
rect 19058 22486 19070 22538
rect 19122 22486 19134 22538
rect 20414 22530 20466 22542
rect 21534 22594 21586 22606
rect 21534 22530 21586 22542
rect 22094 22594 22146 22606
rect 22094 22530 22146 22542
rect 23774 22594 23826 22606
rect 31054 22594 31106 22606
rect 33966 22594 34018 22606
rect 23774 22530 23826 22542
rect 30494 22538 30546 22550
rect 19910 22482 19962 22494
rect 3334 22362 3386 22374
rect 3614 22370 3666 22382
rect 14142 22418 14194 22430
rect 17782 22426 17834 22438
rect 3166 22306 3218 22318
rect 4722 22318 4734 22370
rect 4786 22318 4798 22370
rect 5126 22362 5178 22374
rect 5518 22370 5570 22382
rect 3614 22306 3666 22318
rect 3502 22258 3554 22270
rect 4498 22262 4510 22314
rect 4562 22262 4574 22314
rect 5518 22306 5570 22318
rect 6302 22370 6354 22382
rect 6582 22370 6634 22382
rect 6402 22318 6414 22370
rect 6466 22318 6478 22370
rect 6302 22306 6354 22318
rect 6582 22306 6634 22318
rect 7310 22370 7362 22382
rect 10894 22370 10946 22382
rect 7310 22306 7362 22318
rect 9202 22303 9214 22355
rect 9266 22303 9278 22355
rect 9426 22318 9438 22370
rect 9490 22318 9502 22370
rect 10894 22306 10946 22318
rect 11566 22370 11618 22382
rect 13470 22370 13522 22382
rect 13750 22370 13802 22382
rect 11566 22306 11618 22318
rect 11774 22280 11786 22332
rect 11838 22280 11850 22332
rect 12450 22318 12462 22370
rect 12514 22318 12526 22370
rect 13570 22318 13582 22370
rect 13634 22318 13646 22370
rect 13470 22306 13522 22318
rect 13750 22306 13802 22318
rect 15094 22370 15146 22382
rect 15374 22370 15426 22382
rect 15250 22318 15262 22370
rect 15314 22318 15326 22370
rect 15094 22306 15146 22318
rect 15374 22306 15426 22318
rect 15710 22370 15762 22382
rect 15990 22370 16042 22382
rect 15810 22318 15822 22370
rect 15874 22318 15886 22370
rect 15710 22306 15762 22318
rect 15990 22306 16042 22318
rect 16998 22370 17050 22382
rect 16998 22306 17050 22318
rect 17614 22370 17666 22382
rect 19910 22418 19962 22430
rect 25454 22482 25506 22494
rect 31546 22542 31558 22594
rect 31610 22542 31622 22594
rect 33450 22542 33462 22594
rect 33514 22542 33526 22594
rect 31054 22530 31106 22542
rect 33966 22530 34018 22542
rect 26562 22430 26574 22482
rect 26626 22430 26638 22482
rect 28466 22430 28478 22482
rect 28530 22430 28542 22482
rect 30494 22474 30546 22486
rect 36262 22482 36314 22494
rect 32722 22430 32734 22482
rect 32786 22430 32798 22482
rect 39218 22430 39230 22482
rect 39282 22430 39294 22482
rect 41122 22430 41134 22482
rect 41186 22430 41198 22482
rect 43642 22430 43654 22482
rect 43706 22430 43718 22482
rect 45826 22430 45838 22482
rect 45890 22430 45902 22482
rect 25454 22418 25506 22430
rect 36262 22418 36314 22430
rect 17782 22362 17834 22374
rect 18062 22370 18114 22382
rect 20078 22370 20130 22382
rect 17614 22306 17666 22318
rect 18834 22318 18846 22370
rect 18898 22318 18910 22370
rect 19058 22318 19070 22370
rect 19122 22318 19134 22370
rect 18062 22306 18114 22318
rect 20078 22306 20130 22318
rect 21198 22370 21250 22382
rect 21198 22306 21250 22318
rect 22488 22370 22540 22382
rect 22766 22370 22818 22382
rect 22642 22318 22654 22370
rect 22706 22318 22718 22370
rect 22488 22306 22540 22318
rect 22766 22306 22818 22318
rect 23102 22370 23154 22382
rect 23380 22370 23432 22382
rect 23202 22318 23214 22370
rect 23266 22318 23278 22370
rect 23102 22306 23154 22318
rect 23380 22306 23432 22318
rect 24782 22370 24834 22382
rect 25790 22370 25842 22382
rect 30718 22370 30770 22382
rect 24882 22318 24894 22370
rect 24946 22318 24958 22370
rect 24782 22306 24834 22318
rect 2258 22150 2270 22202
rect 2322 22150 2334 22202
rect 3502 22194 3554 22206
rect 17950 22258 18002 22270
rect 25050 22262 25062 22314
rect 25114 22262 25126 22314
rect 25790 22306 25842 22318
rect 29630 22280 29642 22332
rect 29694 22280 29706 22332
rect 30370 22318 30382 22370
rect 30434 22318 30446 22370
rect 30718 22306 30770 22318
rect 31838 22370 31890 22382
rect 31838 22306 31890 22318
rect 32062 22370 32114 22382
rect 32958 22370 33010 22382
rect 32274 22318 32286 22370
rect 32338 22318 32350 22370
rect 32566 22340 32618 22352
rect 32062 22306 32114 22318
rect 32958 22306 33010 22318
rect 33182 22370 33234 22382
rect 33182 22306 33234 22318
rect 34302 22370 34354 22382
rect 34302 22306 34354 22318
rect 34414 22370 34466 22382
rect 34414 22306 34466 22318
rect 34638 22370 34690 22382
rect 35646 22370 35698 22382
rect 34906 22318 34918 22370
rect 34970 22318 34982 22370
rect 34638 22306 34690 22318
rect 35646 22306 35698 22318
rect 35870 22370 35922 22382
rect 35870 22306 35922 22318
rect 37326 22370 37378 22382
rect 37326 22306 37378 22318
rect 37438 22370 37490 22382
rect 37438 22306 37490 22318
rect 37942 22370 37994 22382
rect 37942 22306 37994 22318
rect 38446 22370 38498 22382
rect 38446 22306 38498 22318
rect 42030 22370 42082 22382
rect 43038 22370 43090 22382
rect 42354 22318 42366 22370
rect 42418 22318 42430 22370
rect 42814 22331 42866 22343
rect 42030 22306 42082 22318
rect 32566 22276 32618 22288
rect 43038 22306 43090 22318
rect 43934 22370 43986 22382
rect 43934 22306 43986 22318
rect 44046 22370 44098 22382
rect 44046 22306 44098 22318
rect 45054 22370 45106 22382
rect 45054 22306 45106 22318
rect 42814 22267 42866 22279
rect 47742 22258 47794 22270
rect 35354 22206 35366 22258
rect 35418 22206 35430 22258
rect 37034 22206 37046 22258
rect 37098 22206 37110 22258
rect 17950 22194 18002 22206
rect 10558 22146 10610 22158
rect 10558 22082 10610 22094
rect 24502 22146 24554 22158
rect 24502 22082 24554 22094
rect 41694 22146 41746 22158
rect 42914 22150 42926 22202
rect 42978 22150 42990 22202
rect 47742 22194 47794 22206
rect 41694 22082 41746 22094
rect 1344 21978 48608 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 48608 21978
rect 1344 21892 48608 21926
rect 2270 21810 2322 21822
rect 2270 21746 2322 21758
rect 13022 21810 13074 21822
rect 3614 21698 3666 21710
rect 6962 21702 6974 21754
rect 7026 21702 7038 21754
rect 13022 21746 13074 21758
rect 19182 21810 19234 21822
rect 19182 21746 19234 21758
rect 20246 21810 20298 21822
rect 20246 21746 20298 21758
rect 20694 21810 20746 21822
rect 20694 21746 20746 21758
rect 23046 21810 23098 21822
rect 23046 21746 23098 21758
rect 27974 21810 28026 21822
rect 27974 21746 28026 21758
rect 38166 21810 38218 21822
rect 3614 21634 3666 21646
rect 12350 21698 12402 21710
rect 12350 21634 12402 21646
rect 18286 21698 18338 21710
rect 2606 21586 2658 21598
rect 2606 21522 2658 21534
rect 3278 21586 3330 21598
rect 4046 21572 4058 21624
rect 4110 21572 4122 21624
rect 4722 21534 4734 21586
rect 4786 21534 4798 21586
rect 5394 21534 5406 21586
rect 5458 21534 5470 21586
rect 6629 21573 6641 21625
rect 6693 21573 6705 21625
rect 13840 21624 13892 21636
rect 7758 21586 7810 21598
rect 7186 21534 7198 21586
rect 7250 21534 7262 21586
rect 3278 21522 3330 21534
rect 7758 21522 7810 21534
rect 8766 21586 8818 21598
rect 8766 21522 8818 21534
rect 9662 21586 9714 21598
rect 12686 21586 12738 21598
rect 10434 21534 10446 21586
rect 10498 21534 10510 21586
rect 9662 21522 9714 21534
rect 12686 21522 12738 21534
rect 13582 21586 13634 21598
rect 13682 21534 13694 21586
rect 13746 21534 13758 21586
rect 13840 21560 13892 21572
rect 15188 21624 15240 21636
rect 18286 21634 18338 21646
rect 18678 21698 18730 21710
rect 18678 21634 18730 21646
rect 21702 21698 21754 21710
rect 21702 21634 21754 21646
rect 24278 21698 24330 21710
rect 28578 21702 28590 21754
rect 28642 21702 28654 21754
rect 38166 21746 38218 21758
rect 24278 21634 24330 21646
rect 32398 21698 32450 21710
rect 21982 21614 22034 21626
rect 15486 21586 15538 21598
rect 15188 21560 15240 21572
rect 15362 21534 15374 21586
rect 15426 21534 15438 21586
rect 13582 21522 13634 21534
rect 15486 21522 15538 21534
rect 16886 21586 16938 21598
rect 16886 21522 16938 21534
rect 17950 21586 18002 21598
rect 18398 21586 18450 21598
rect 17950 21522 18002 21534
rect 18118 21530 18170 21542
rect 14814 21474 14866 21486
rect 5618 21422 5630 21474
rect 5682 21422 5694 21474
rect 4498 21366 4510 21418
rect 4562 21366 4574 21418
rect 14814 21410 14866 21422
rect 15990 21474 16042 21486
rect 15990 21410 16042 21422
rect 16438 21474 16490 21486
rect 16438 21410 16490 21422
rect 17670 21474 17722 21486
rect 18398 21522 18450 21534
rect 19518 21586 19570 21598
rect 19518 21522 19570 21534
rect 21422 21586 21474 21598
rect 21982 21550 22034 21562
rect 22150 21621 22202 21633
rect 22150 21557 22202 21569
rect 22430 21614 22482 21626
rect 22430 21550 22482 21562
rect 22542 21621 22594 21633
rect 25824 21624 25876 21636
rect 22542 21557 22594 21569
rect 24726 21586 24778 21598
rect 21422 21522 21474 21534
rect 24726 21522 24778 21534
rect 25566 21586 25618 21598
rect 25666 21534 25678 21586
rect 25730 21534 25742 21586
rect 27188 21584 27200 21636
rect 27252 21584 27264 21636
rect 32398 21634 32450 21646
rect 36094 21698 36146 21710
rect 36094 21634 36146 21646
rect 40294 21698 40346 21710
rect 46106 21646 46118 21698
rect 46170 21646 46182 21698
rect 40294 21634 40346 21646
rect 47350 21615 47402 21627
rect 27470 21586 27522 21598
rect 29374 21586 29426 21598
rect 25824 21560 25876 21572
rect 27346 21534 27358 21586
rect 27410 21534 27422 21586
rect 28690 21534 28702 21586
rect 28754 21534 28766 21586
rect 25566 21522 25618 21534
rect 27470 21522 27522 21534
rect 29374 21522 29426 21534
rect 29710 21586 29762 21598
rect 29710 21522 29762 21534
rect 33238 21586 33290 21598
rect 33238 21522 33290 21534
rect 33406 21586 33458 21598
rect 37214 21586 37266 21598
rect 36530 21534 36542 21586
rect 36594 21534 36606 21586
rect 36866 21534 36878 21586
rect 36930 21534 36942 21586
rect 33406 21522 33458 21534
rect 37214 21522 37266 21534
rect 38894 21586 38946 21598
rect 38894 21522 38946 21534
rect 39342 21586 39394 21598
rect 39342 21522 39394 21534
rect 39678 21586 39730 21598
rect 39678 21522 39730 21534
rect 40798 21586 40850 21598
rect 43486 21586 43538 21598
rect 41570 21534 41582 21586
rect 41634 21534 41646 21586
rect 44034 21549 44046 21601
rect 44098 21549 44110 21601
rect 44606 21586 44658 21598
rect 44258 21534 44270 21586
rect 44322 21534 44334 21586
rect 40798 21522 40850 21534
rect 43486 21522 43538 21534
rect 44606 21522 44658 21534
rect 45614 21586 45666 21598
rect 45614 21522 45666 21534
rect 45838 21586 45890 21598
rect 46610 21549 46622 21601
rect 46674 21549 46686 21601
rect 46946 21534 46958 21586
rect 47010 21534 47022 21586
rect 47350 21551 47402 21563
rect 47730 21534 47742 21586
rect 47794 21534 47806 21586
rect 45838 21522 45890 21534
rect 18118 21466 18170 21478
rect 26238 21474 26290 21486
rect 48246 21474 48298 21486
rect 17670 21410 17722 21422
rect 30482 21422 30494 21474
rect 30546 21422 30558 21474
rect 34178 21422 34190 21474
rect 34242 21422 34254 21474
rect 43922 21422 43934 21474
rect 43986 21422 43998 21474
rect 46498 21422 46510 21474
rect 46562 21422 46574 21474
rect 47282 21422 47294 21474
rect 47346 21422 47358 21474
rect 26238 21410 26290 21422
rect 8430 21362 8482 21374
rect 8430 21298 8482 21310
rect 14254 21362 14306 21374
rect 14254 21298 14306 21310
rect 21086 21362 21138 21374
rect 21086 21298 21138 21310
rect 26798 21362 26850 21374
rect 36642 21366 36654 21418
rect 36706 21366 36718 21418
rect 48246 21410 48298 21422
rect 26798 21298 26850 21310
rect 37550 21362 37602 21374
rect 37550 21298 37602 21310
rect 38558 21362 38610 21374
rect 38558 21298 38610 21310
rect 44942 21362 44994 21374
rect 44942 21298 44994 21310
rect 1344 21194 48608 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 48608 21194
rect 1344 21108 48608 21142
rect 4846 21026 4898 21038
rect 4846 20962 4898 20974
rect 5854 21026 5906 21038
rect 5854 20962 5906 20974
rect 10558 21026 10610 21038
rect 10558 20962 10610 20974
rect 11230 21026 11282 21038
rect 11230 20962 11282 20974
rect 18342 21026 18394 21038
rect 11778 20918 11790 20970
rect 11842 20918 11854 20970
rect 18342 20962 18394 20974
rect 19462 21026 19514 21038
rect 19462 20962 19514 20974
rect 19910 21026 19962 21038
rect 19910 20962 19962 20974
rect 29374 21026 29426 21038
rect 29374 20962 29426 20974
rect 34526 21026 34578 21038
rect 14366 20914 14418 20926
rect 4274 20862 4286 20914
rect 4338 20862 4350 20914
rect 6962 20862 6974 20914
rect 7026 20862 7038 20914
rect 8866 20862 8878 20914
rect 8930 20862 8942 20914
rect 14366 20850 14418 20862
rect 15542 20914 15594 20926
rect 15542 20850 15594 20862
rect 15990 20914 16042 20926
rect 24894 20914 24946 20926
rect 33282 20918 33294 20970
rect 33346 20918 33358 20970
rect 34526 20962 34578 20974
rect 40910 21026 40962 21038
rect 43082 20974 43094 21026
rect 43146 20974 43158 21026
rect 40910 20962 40962 20974
rect 41526 20914 41578 20926
rect 15990 20850 16042 20862
rect 18902 20858 18954 20870
rect 1598 20802 1650 20814
rect 5182 20802 5234 20814
rect 6526 20802 6578 20814
rect 2370 20750 2382 20802
rect 2434 20750 2446 20802
rect 6402 20750 6414 20802
rect 6466 20750 6478 20802
rect 1598 20738 1650 20750
rect 5182 20738 5234 20750
rect 6236 20694 6248 20746
rect 6300 20694 6312 20746
rect 6526 20738 6578 20750
rect 9662 20802 9714 20814
rect 9662 20738 9714 20750
rect 9886 20802 9938 20814
rect 11566 20802 11618 20814
rect 12574 20802 12626 20814
rect 9986 20750 9998 20802
rect 10050 20750 10062 20802
rect 12002 20750 12014 20802
rect 12066 20750 12078 20802
rect 9886 20738 9938 20750
rect 10152 20694 10164 20746
rect 10216 20694 10228 20746
rect 11566 20738 11618 20750
rect 12574 20738 12626 20750
rect 13358 20802 13410 20814
rect 13358 20738 13410 20750
rect 14758 20802 14810 20814
rect 15038 20802 15090 20814
rect 14914 20750 14926 20802
rect 14978 20750 14990 20802
rect 14758 20738 14810 20750
rect 15038 20738 15090 20750
rect 16158 20802 16210 20814
rect 16158 20738 16210 20750
rect 16830 20802 16882 20814
rect 16830 20738 16882 20750
rect 17166 20802 17218 20814
rect 17166 20738 17218 20750
rect 17614 20802 17666 20814
rect 18062 20802 18114 20814
rect 17938 20750 17950 20802
rect 18002 20750 18014 20802
rect 17614 20738 17666 20750
rect 17770 20694 17782 20746
rect 17834 20694 17846 20746
rect 18062 20738 18114 20750
rect 18734 20802 18786 20814
rect 28466 20862 28478 20914
rect 28530 20862 28542 20914
rect 32386 20862 32398 20914
rect 32450 20862 32462 20914
rect 37090 20862 37102 20914
rect 37154 20862 37166 20914
rect 43810 20862 43822 20914
rect 43874 20862 43886 20914
rect 45490 20862 45502 20914
rect 45554 20862 45566 20914
rect 24894 20850 24946 20862
rect 41526 20850 41578 20862
rect 18902 20794 18954 20806
rect 19182 20802 19234 20814
rect 23326 20802 23378 20814
rect 18734 20738 18786 20750
rect 19182 20738 19234 20750
rect 20190 20774 20242 20786
rect 20750 20767 20802 20779
rect 20190 20710 20242 20722
rect 19070 20690 19122 20702
rect 20402 20694 20414 20746
rect 20466 20694 20478 20746
rect 20626 20694 20638 20746
rect 20690 20694 20702 20746
rect 22094 20746 22146 20758
rect 23090 20750 23102 20802
rect 23154 20750 23166 20802
rect 20750 20703 20802 20715
rect 21746 20694 21758 20746
rect 21810 20694 21822 20746
rect 23326 20738 23378 20750
rect 24558 20802 24610 20814
rect 25790 20802 25842 20814
rect 29038 20802 29090 20814
rect 25106 20750 25118 20802
rect 25170 20750 25182 20802
rect 26562 20750 26574 20802
rect 26626 20750 26638 20802
rect 23538 20694 23550 20746
rect 23602 20694 23614 20746
rect 24558 20738 24610 20750
rect 24938 20694 24950 20746
rect 25002 20694 25014 20746
rect 25790 20738 25842 20750
rect 29038 20738 29090 20750
rect 30942 20802 30994 20814
rect 30942 20738 30994 20750
rect 31390 20802 31442 20814
rect 34862 20802 34914 20814
rect 35422 20802 35474 20814
rect 31390 20738 31442 20750
rect 31714 20723 31726 20775
rect 31778 20723 31790 20775
rect 32050 20750 32062 20802
rect 32114 20750 32126 20802
rect 32722 20750 32734 20802
rect 32786 20750 32798 20802
rect 33170 20750 33182 20802
rect 33234 20750 33246 20802
rect 33506 20750 33518 20802
rect 33570 20750 33582 20802
rect 35130 20750 35142 20802
rect 35194 20750 35206 20802
rect 32554 20694 32566 20746
rect 32618 20694 32630 20746
rect 34862 20738 34914 20750
rect 35422 20738 35474 20750
rect 35646 20802 35698 20814
rect 35646 20738 35698 20750
rect 36318 20802 36370 20814
rect 39790 20802 39842 20814
rect 38994 20750 39006 20802
rect 39058 20750 39070 20802
rect 36318 20738 36370 20750
rect 39790 20738 39842 20750
rect 39902 20802 39954 20814
rect 39902 20738 39954 20750
rect 40574 20802 40626 20814
rect 42478 20802 42530 20814
rect 41794 20750 41806 20802
rect 41858 20750 41870 20802
rect 42254 20763 42306 20775
rect 40574 20738 40626 20750
rect 42478 20738 42530 20750
rect 43374 20802 43426 20814
rect 43374 20738 43426 20750
rect 43486 20802 43538 20814
rect 44718 20802 44770 20814
rect 43486 20738 43538 20750
rect 42254 20699 42306 20711
rect 43922 20706 43934 20758
rect 43986 20706 43998 20758
rect 44258 20750 44270 20802
rect 44322 20750 44334 20802
rect 44718 20738 44770 20750
rect 48302 20802 48354 20814
rect 48302 20738 48354 20750
rect 22094 20682 22146 20694
rect 47406 20690 47458 20702
rect 19070 20626 19122 20638
rect 13694 20578 13746 20590
rect 13694 20514 13746 20526
rect 16494 20578 16546 20590
rect 16494 20514 16546 20526
rect 30606 20578 30658 20590
rect 31266 20582 31278 20634
rect 31330 20582 31342 20634
rect 30606 20514 30658 20526
rect 34134 20578 34186 20590
rect 34134 20514 34186 20526
rect 35982 20578 36034 20590
rect 35982 20514 36034 20526
rect 40238 20578 40290 20590
rect 42018 20582 42030 20634
rect 42082 20582 42094 20634
rect 47406 20626 47458 20638
rect 40238 20514 40290 20526
rect 47966 20578 48018 20590
rect 47966 20514 48018 20526
rect 1344 20410 48608 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 48608 20410
rect 1344 20324 48608 20358
rect 1822 20242 1874 20254
rect 1822 20178 1874 20190
rect 18510 20242 18562 20254
rect 18510 20178 18562 20190
rect 28422 20242 28474 20254
rect 28422 20178 28474 20190
rect 28870 20242 28922 20254
rect 28870 20178 28922 20190
rect 12350 20130 12402 20142
rect 6492 20055 6544 20067
rect 12350 20066 12402 20078
rect 13414 20130 13466 20142
rect 13414 20066 13466 20078
rect 16718 20130 16770 20142
rect 21870 20130 21922 20142
rect 19562 20078 19574 20130
rect 19626 20078 19638 20130
rect 2158 20018 2210 20030
rect 2158 19954 2210 19966
rect 2270 20018 2322 20030
rect 6750 20018 6802 20030
rect 6492 19991 6544 20003
rect 6626 19966 6638 20018
rect 6690 19966 6702 20018
rect 2270 19954 2322 19966
rect 6750 19954 6802 19966
rect 7534 20018 7586 20030
rect 7534 19954 7586 19966
rect 7758 20018 7810 20030
rect 8038 20018 8090 20030
rect 7858 19966 7870 20018
rect 7922 19966 7934 20018
rect 7758 19954 7810 19966
rect 8038 19954 8090 19966
rect 9662 20018 9714 20030
rect 13694 20018 13746 20030
rect 13962 20022 13974 20074
rect 14026 20022 14038 20074
rect 16718 20066 16770 20078
rect 20638 20074 20690 20086
rect 14142 20018 14194 20030
rect 13010 19966 13022 20018
rect 13074 19966 13086 20018
rect 13794 19966 13806 20018
rect 13858 19966 13870 20018
rect 9662 19954 9714 19966
rect 13694 19954 13746 19966
rect 14142 19954 14194 19966
rect 14814 20018 14866 20030
rect 15094 20018 15146 20030
rect 14914 19966 14926 20018
rect 14978 19966 14990 20018
rect 14814 19954 14866 19966
rect 15094 19954 15146 19966
rect 15262 20018 15314 20030
rect 16382 20018 16434 20030
rect 15698 19966 15710 20018
rect 15762 19966 15774 20018
rect 15922 19966 15934 20018
rect 15986 19966 15998 20018
rect 15262 19954 15314 19966
rect 16382 19954 16434 19966
rect 17502 20018 17554 20030
rect 17502 19954 17554 19966
rect 17838 20018 17890 20030
rect 17838 19954 17890 19966
rect 18846 20018 18898 20030
rect 18846 19954 18898 19966
rect 19070 20018 19122 20030
rect 19070 19954 19122 19966
rect 19294 20018 19346 20030
rect 20178 20022 20190 20074
rect 20242 20022 20254 20074
rect 21870 20066 21922 20078
rect 27134 20130 27186 20142
rect 22530 20022 22542 20074
rect 22594 20022 22606 20074
rect 20638 20010 20690 20022
rect 22766 20018 22818 20030
rect 21634 19966 21646 20018
rect 21698 19966 21710 20018
rect 19294 19954 19346 19966
rect 22766 19954 22818 19966
rect 23774 20018 23826 20030
rect 24098 20022 24110 20074
rect 24162 20022 24174 20074
rect 26088 20056 26140 20068
rect 27134 20066 27186 20078
rect 31222 20130 31274 20142
rect 36878 20130 36930 20142
rect 31222 20066 31274 20078
rect 33742 20074 33794 20086
rect 36026 20078 36038 20130
rect 36090 20078 36102 20130
rect 25790 20018 25842 20030
rect 24434 19966 24446 20018
rect 24498 19966 24510 20018
rect 25442 19966 25454 20018
rect 25506 19966 25518 20018
rect 25890 19966 25902 20018
rect 25954 19966 25966 20018
rect 26088 19992 26140 20004
rect 26798 20018 26850 20030
rect 23774 19954 23826 19966
rect 25790 19954 25842 19966
rect 26798 19954 26850 19966
rect 28030 20018 28082 20030
rect 33014 20018 33066 20030
rect 30258 19966 30270 20018
rect 30322 19966 30334 20018
rect 30594 19966 30606 20018
rect 30658 19966 30670 20018
rect 31714 19966 31726 20018
rect 31778 19966 31790 20018
rect 32050 19966 32062 20018
rect 32114 19966 32126 20018
rect 32274 19966 32286 20018
rect 32338 19966 32350 20018
rect 33394 19966 33406 20018
rect 33458 19966 33470 20018
rect 33742 20010 33794 20022
rect 34414 20018 34466 20030
rect 35278 20022 35290 20074
rect 35342 20022 35354 20074
rect 36878 20066 36930 20078
rect 38110 20130 38162 20142
rect 28030 19954 28082 19966
rect 33014 19954 33066 19966
rect 34414 19954 34466 19966
rect 35534 20018 35586 20030
rect 35534 19954 35586 19966
rect 36318 20018 36370 20030
rect 36318 19954 36370 19966
rect 36542 20018 36594 20030
rect 36542 19954 36594 19966
rect 37214 20018 37266 20030
rect 37706 20022 37718 20074
rect 37770 20022 37782 20074
rect 38110 20066 38162 20078
rect 38782 20018 38834 20030
rect 43822 20018 43874 20030
rect 44718 20018 44770 20030
rect 37874 19966 37886 20018
rect 37938 19966 37950 20018
rect 37214 19954 37266 19966
rect 38278 19962 38330 19974
rect 5686 19906 5738 19918
rect 3042 19854 3054 19906
rect 3106 19854 3118 19906
rect 4946 19854 4958 19906
rect 5010 19854 5022 19906
rect 5686 19842 5738 19854
rect 7198 19906 7250 19918
rect 7198 19842 7250 19854
rect 8430 19906 8482 19918
rect 8430 19842 8482 19854
rect 9046 19906 9098 19918
rect 14534 19906 14586 19918
rect 10434 19854 10446 19906
rect 10498 19854 10510 19906
rect 24110 19906 24162 19918
rect 9046 19842 9098 19854
rect 14534 19842 14586 19854
rect 15598 19850 15650 19862
rect 6078 19794 6130 19806
rect 6078 19730 6130 19742
rect 12854 19794 12906 19806
rect 26462 19906 26514 19918
rect 24110 19842 24162 19854
rect 25286 19850 25338 19862
rect 15598 19786 15650 19798
rect 23102 19794 23154 19806
rect 12854 19730 12906 19742
rect 33182 19906 33234 19918
rect 26462 19842 26514 19854
rect 30718 19850 30770 19862
rect 25286 19786 25338 19798
rect 27694 19794 27746 19806
rect 23102 19730 23154 19742
rect 32398 19850 32450 19862
rect 30718 19786 30770 19798
rect 31558 19794 31610 19806
rect 27694 19730 27746 19742
rect 40002 19966 40014 20018
rect 40066 19966 40078 20018
rect 40338 19966 40350 20018
rect 40402 19966 40414 20018
rect 44146 19966 44158 20018
rect 44210 19966 44222 20018
rect 44482 19966 44494 20018
rect 44546 19966 44558 20018
rect 38782 19954 38834 19966
rect 43822 19954 43874 19966
rect 44718 19954 44770 19966
rect 45390 20018 45442 20030
rect 48078 20018 48130 20030
rect 46162 19966 46174 20018
rect 46226 19966 46238 20018
rect 45390 19954 45442 19966
rect 48078 19954 48130 19966
rect 38278 19898 38330 19910
rect 33182 19842 33234 19854
rect 39902 19850 39954 19862
rect 41122 19854 41134 19906
rect 41186 19854 41198 19906
rect 43026 19854 43038 19906
rect 43090 19854 43102 19906
rect 32398 19786 32450 19798
rect 39118 19794 39170 19806
rect 31558 19730 31610 19742
rect 39902 19786 39954 19798
rect 44046 19850 44098 19862
rect 44046 19786 44098 19798
rect 45054 19794 45106 19806
rect 39118 19730 39170 19742
rect 45054 19730 45106 19742
rect 1344 19626 48608 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 48608 19626
rect 1344 19540 48608 19574
rect 6974 19458 7026 19470
rect 5058 19350 5070 19402
rect 5122 19350 5134 19402
rect 6178 19350 6190 19402
rect 6242 19350 6254 19402
rect 6974 19394 7026 19406
rect 8990 19458 9042 19470
rect 8990 19394 9042 19406
rect 12798 19458 12850 19470
rect 12798 19394 12850 19406
rect 13694 19458 13746 19470
rect 13694 19394 13746 19406
rect 15430 19458 15482 19470
rect 15430 19394 15482 19406
rect 20526 19458 20578 19470
rect 20526 19394 20578 19406
rect 21366 19458 21418 19470
rect 21366 19394 21418 19406
rect 23494 19458 23546 19470
rect 23494 19394 23546 19406
rect 27134 19458 27186 19470
rect 40238 19458 40290 19470
rect 38042 19406 38054 19458
rect 38106 19406 38118 19458
rect 43978 19406 43990 19458
rect 44042 19406 44054 19458
rect 27134 19394 27186 19406
rect 40238 19394 40290 19406
rect 45614 19402 45666 19414
rect 16774 19346 16826 19358
rect 14870 19290 14922 19302
rect 4286 19234 4338 19246
rect 6638 19234 6690 19246
rect 4946 19182 4958 19234
rect 5010 19182 5022 19234
rect 6066 19182 6078 19234
rect 6130 19182 6142 19234
rect 6402 19182 6414 19234
rect 6466 19182 6478 19234
rect 4286 19170 4338 19182
rect 6638 19170 6690 19182
rect 7870 19234 7922 19246
rect 7870 19170 7922 19182
rect 9326 19234 9378 19246
rect 9326 19170 9378 19182
rect 9438 19234 9490 19246
rect 12126 19234 12178 19246
rect 10210 19182 10222 19234
rect 10274 19182 10286 19234
rect 9438 19170 9490 19182
rect 12126 19170 12178 19182
rect 12462 19234 12514 19246
rect 12462 19170 12514 19182
rect 14030 19234 14082 19246
rect 14030 19170 14082 19182
rect 14590 19234 14642 19246
rect 15990 19290 16042 19302
rect 14690 19182 14702 19234
rect 14754 19182 14766 19234
rect 14870 19226 14922 19238
rect 15038 19234 15090 19246
rect 14590 19170 14642 19182
rect 15038 19170 15090 19182
rect 15710 19234 15762 19246
rect 16774 19282 16826 19294
rect 17166 19346 17218 19358
rect 22262 19346 22314 19358
rect 17166 19282 17218 19294
rect 18342 19290 18394 19302
rect 15990 19226 16042 19238
rect 16158 19234 16210 19246
rect 15710 19170 15762 19182
rect 16158 19170 16210 19182
rect 17502 19234 17554 19246
rect 17502 19170 17554 19182
rect 18062 19234 18114 19246
rect 22262 19282 22314 19294
rect 22710 19346 22762 19358
rect 22710 19282 22762 19294
rect 23158 19346 23210 19358
rect 38614 19346 38666 19358
rect 23158 19282 23210 19294
rect 24054 19290 24106 19302
rect 18342 19226 18394 19238
rect 18510 19234 18562 19246
rect 18062 19170 18114 19182
rect 18510 19170 18562 19182
rect 19070 19234 19122 19246
rect 20190 19234 20242 19246
rect 23774 19234 23826 19246
rect 24726 19290 24778 19302
rect 31714 19294 31726 19346
rect 31778 19294 31790 19346
rect 33842 19294 33854 19346
rect 33906 19294 33918 19346
rect 35746 19294 35758 19346
rect 35810 19294 35822 19346
rect 45614 19338 45666 19350
rect 47182 19402 47234 19414
rect 47898 19406 47910 19458
rect 47962 19406 47974 19458
rect 47182 19338 47234 19350
rect 19070 19170 19122 19182
rect 19294 19195 19346 19207
rect 19618 19182 19630 19234
rect 19682 19182 19694 19234
rect 21522 19182 21534 19234
rect 21586 19182 21598 19234
rect 23874 19182 23886 19234
rect 23938 19182 23950 19234
rect 24054 19226 24106 19238
rect 24222 19234 24274 19246
rect 20190 19170 20242 19182
rect 23774 19170 23826 19182
rect 24222 19170 24274 19182
rect 24558 19234 24610 19246
rect 38614 19282 38666 19294
rect 24726 19226 24778 19238
rect 25006 19234 25058 19246
rect 26126 19234 26178 19246
rect 24882 19182 24894 19234
rect 24946 19182 24958 19234
rect 25666 19182 25678 19234
rect 25730 19182 25742 19234
rect 24558 19170 24610 19182
rect 25006 19170 25058 19182
rect 26126 19170 26178 19182
rect 26350 19234 26402 19246
rect 26350 19170 26402 19182
rect 27470 19234 27522 19246
rect 27470 19170 27522 19182
rect 29038 19234 29090 19246
rect 36542 19234 36594 19246
rect 29810 19182 29822 19234
rect 29874 19182 29886 19234
rect 32622 19206 32674 19218
rect 29038 19170 29090 19182
rect 14310 19122 14362 19134
rect 14310 19058 14362 19070
rect 15822 19122 15874 19134
rect 15822 19058 15874 19070
rect 17782 19122 17834 19134
rect 17782 19058 17834 19070
rect 18174 19122 18226 19134
rect 19294 19131 19346 19143
rect 32622 19142 32674 19154
rect 32846 19206 32898 19218
rect 33182 19199 33234 19211
rect 32846 19142 32898 19154
rect 25286 19122 25338 19134
rect 32342 19122 32394 19134
rect 33058 19126 33070 19178
rect 33122 19126 33134 19178
rect 36542 19170 36594 19182
rect 37438 19234 37490 19246
rect 37438 19170 37490 19182
rect 37550 19234 37602 19246
rect 37550 19170 37602 19182
rect 37774 19234 37826 19246
rect 43486 19234 43538 19246
rect 37774 19170 37826 19182
rect 39218 19154 39230 19206
rect 39282 19154 39294 19206
rect 33182 19135 33234 19147
rect 41794 19126 41806 19178
rect 41858 19126 41870 19178
rect 42130 19126 42142 19178
rect 42194 19126 42206 19178
rect 42578 19126 42590 19178
rect 42642 19126 42654 19178
rect 42776 19149 42788 19201
rect 42840 19149 42852 19201
rect 43486 19170 43538 19182
rect 43710 19234 43762 19246
rect 43710 19170 43762 19182
rect 44830 19234 44882 19246
rect 44830 19170 44882 19182
rect 44942 19234 44994 19246
rect 47406 19234 47458 19246
rect 45210 19182 45222 19234
rect 45274 19182 45286 19234
rect 45714 19182 45726 19234
rect 45778 19182 45790 19234
rect 45938 19182 45950 19234
rect 46002 19182 46014 19234
rect 46834 19182 46846 19234
rect 46898 19182 46910 19234
rect 47058 19182 47070 19234
rect 47122 19182 47134 19234
rect 44942 19170 44994 19182
rect 47406 19170 47458 19182
rect 47630 19234 47682 19246
rect 47630 19170 47682 19182
rect 18174 19058 18226 19070
rect 19406 19066 19458 19078
rect 4006 19010 4058 19022
rect 4006 18946 4058 18958
rect 7534 19010 7586 19022
rect 7534 18946 7586 18958
rect 8598 19010 8650 19022
rect 26618 19070 26630 19122
rect 26682 19070 26694 19122
rect 25286 19058 25338 19070
rect 32342 19058 32394 19070
rect 42926 19122 42978 19134
rect 42926 19058 42978 19070
rect 19406 19002 19458 19014
rect 25846 19010 25898 19022
rect 8598 18946 8650 18958
rect 25846 18946 25898 18958
rect 27862 19010 27914 19022
rect 27862 18946 27914 18958
rect 28310 19010 28362 19022
rect 28310 18946 28362 18958
rect 37102 19010 37154 19022
rect 37102 18946 37154 18958
rect 1344 18842 48608 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 48608 18842
rect 1344 18756 48608 18790
rect 14814 18674 14866 18686
rect 14814 18610 14866 18622
rect 15486 18674 15538 18686
rect 15486 18610 15538 18622
rect 21030 18674 21082 18686
rect 21030 18610 21082 18622
rect 23718 18674 23770 18686
rect 23718 18610 23770 18622
rect 31726 18562 31778 18574
rect 6134 18506 6186 18518
rect 33182 18562 33234 18574
rect 3054 18450 3106 18462
rect 3054 18386 3106 18398
rect 5742 18450 5794 18462
rect 6134 18442 6186 18454
rect 6862 18488 6914 18500
rect 6514 18398 6526 18450
rect 6578 18398 6590 18450
rect 14310 18479 14362 18491
rect 6862 18424 6914 18436
rect 7926 18450 7978 18462
rect 8306 18413 8318 18465
rect 8370 18413 8382 18465
rect 8530 18398 8542 18450
rect 8594 18398 8606 18450
rect 9762 18398 9774 18450
rect 9826 18398 9838 18450
rect 13122 18425 13134 18477
rect 13186 18425 13198 18477
rect 13906 18398 13918 18450
rect 13970 18398 13982 18450
rect 14310 18415 14362 18427
rect 15150 18450 15202 18462
rect 5742 18386 5794 18398
rect 7926 18386 7978 18398
rect 15150 18386 15202 18398
rect 15822 18450 15874 18462
rect 15922 18398 15934 18450
rect 15986 18398 15998 18450
rect 17378 18425 17390 18477
rect 17442 18425 17454 18477
rect 18734 18450 18786 18462
rect 15822 18386 15874 18398
rect 18734 18386 18786 18398
rect 20078 18450 20130 18462
rect 20078 18386 20130 18398
rect 20414 18450 20466 18462
rect 21578 18454 21590 18506
rect 21642 18454 21654 18506
rect 22654 18488 22706 18500
rect 31726 18498 31778 18510
rect 33014 18506 33066 18518
rect 21982 18450 22034 18462
rect 21298 18398 21310 18450
rect 21362 18398 21374 18450
rect 24110 18450 24162 18462
rect 22654 18424 22706 18436
rect 22978 18398 22990 18450
rect 23042 18398 23054 18450
rect 20414 18386 20466 18398
rect 21982 18386 22034 18398
rect 23382 18394 23434 18406
rect 23538 18398 23550 18450
rect 23602 18398 23614 18450
rect 6302 18338 6354 18350
rect 3826 18286 3838 18338
rect 3890 18286 3902 18338
rect 6302 18274 6354 18286
rect 7478 18338 7530 18350
rect 23214 18338 23266 18350
rect 8194 18286 8206 18338
rect 8258 18286 8270 18338
rect 14354 18286 14366 18338
rect 14418 18286 14430 18338
rect 21410 18286 21422 18338
rect 21474 18286 21486 18338
rect 24110 18386 24162 18398
rect 24222 18450 24274 18462
rect 25330 18442 25342 18494
rect 25394 18442 25406 18494
rect 26350 18450 26402 18462
rect 26798 18450 26850 18462
rect 25554 18398 25566 18450
rect 25618 18398 25630 18450
rect 26450 18398 26462 18450
rect 26514 18398 26526 18450
rect 24222 18386 24274 18398
rect 26350 18386 26402 18398
rect 26630 18394 26682 18406
rect 23382 18330 23434 18342
rect 26798 18386 26850 18398
rect 27022 18450 27074 18462
rect 28142 18450 28194 18462
rect 27022 18386 27074 18398
rect 27974 18394 28026 18406
rect 25218 18286 25230 18338
rect 25282 18286 25294 18338
rect 26630 18330 26682 18342
rect 28578 18426 28590 18478
rect 28642 18426 28654 18478
rect 29038 18450 29090 18462
rect 33182 18498 33234 18510
rect 33742 18506 33794 18518
rect 28142 18386 28194 18398
rect 32386 18398 32398 18450
rect 32450 18398 32462 18450
rect 33014 18442 33066 18454
rect 38390 18506 38442 18518
rect 33394 18398 33406 18450
rect 33458 18398 33470 18450
rect 33742 18442 33794 18454
rect 34470 18450 34522 18462
rect 28802 18342 28814 18394
rect 28866 18342 28878 18394
rect 29038 18386 29090 18398
rect 34470 18386 34522 18398
rect 35198 18450 35250 18462
rect 35198 18386 35250 18398
rect 35310 18450 35362 18462
rect 39118 18488 39170 18500
rect 38390 18442 38442 18454
rect 38558 18450 38610 18462
rect 35310 18386 35362 18398
rect 38770 18398 38782 18450
rect 38834 18398 38846 18450
rect 39118 18424 39170 18436
rect 39566 18450 39618 18462
rect 39846 18450 39898 18462
rect 39666 18398 39678 18450
rect 39730 18398 39742 18450
rect 38558 18386 38610 18398
rect 39566 18386 39618 18398
rect 39846 18386 39898 18398
rect 40798 18450 40850 18462
rect 40798 18386 40850 18398
rect 41022 18450 41074 18462
rect 42366 18450 42418 18462
rect 41290 18398 41302 18450
rect 41354 18398 41366 18450
rect 41682 18398 41694 18450
rect 41746 18398 41758 18450
rect 42018 18398 42030 18450
rect 42082 18398 42094 18450
rect 41022 18386 41074 18398
rect 42366 18386 42418 18398
rect 42590 18450 42642 18462
rect 43698 18454 43710 18506
rect 43762 18454 43774 18506
rect 43922 18431 43934 18483
rect 43986 18431 43998 18483
rect 44482 18434 44494 18486
rect 44546 18434 44558 18486
rect 44680 18438 44692 18490
rect 44744 18438 44756 18490
rect 45054 18450 45106 18462
rect 42590 18386 42642 18398
rect 45054 18386 45106 18398
rect 27974 18330 28026 18342
rect 34862 18338 34914 18350
rect 40238 18338 40290 18350
rect 29810 18286 29822 18338
rect 29874 18286 29886 18338
rect 36082 18286 36094 18338
rect 36146 18286 36158 18338
rect 37986 18286 37998 18338
rect 38050 18286 38062 18338
rect 7478 18274 7530 18286
rect 23214 18274 23266 18286
rect 34862 18274 34914 18286
rect 40238 18274 40290 18286
rect 42142 18282 42194 18294
rect 42858 18286 42870 18338
rect 42922 18286 42934 18338
rect 44706 18286 44718 18338
rect 44770 18286 44782 18338
rect 45826 18286 45838 18338
rect 45890 18286 45902 18338
rect 47730 18286 47742 18338
rect 47794 18286 47806 18338
rect 12126 18226 12178 18238
rect 26070 18226 26122 18238
rect 24490 18174 24502 18226
rect 24554 18174 24566 18226
rect 12126 18162 12178 18174
rect 26070 18162 26122 18174
rect 27358 18226 27410 18238
rect 27358 18162 27410 18174
rect 32230 18226 32282 18238
rect 42142 18218 42194 18230
rect 32230 18162 32282 18174
rect 1344 18058 48608 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 48608 18058
rect 1344 17972 48608 18006
rect 9662 17890 9714 17902
rect 6010 17838 6022 17890
rect 6074 17838 6086 17890
rect 9662 17826 9714 17838
rect 18454 17890 18506 17902
rect 24782 17890 24834 17902
rect 18454 17826 18506 17838
rect 23326 17834 23378 17846
rect 5126 17778 5178 17790
rect 13806 17778 13858 17790
rect 35422 17890 35474 17902
rect 24782 17826 24834 17838
rect 28030 17834 28082 17846
rect 7186 17726 7198 17778
rect 7250 17726 7262 17778
rect 16034 17726 16046 17778
rect 16098 17726 16110 17778
rect 20514 17726 20526 17778
rect 20578 17726 20590 17778
rect 21970 17726 21982 17778
rect 22034 17726 22046 17778
rect 23326 17770 23378 17782
rect 24390 17778 24442 17790
rect 35422 17826 35474 17838
rect 42030 17890 42082 17902
rect 42030 17826 42082 17838
rect 28030 17770 28082 17782
rect 29262 17778 29314 17790
rect 5126 17714 5178 17726
rect 13806 17714 13858 17726
rect 24390 17714 24442 17726
rect 29262 17714 29314 17726
rect 30550 17778 30602 17790
rect 43150 17778 43202 17790
rect 43922 17782 43934 17834
rect 43986 17782 43998 17834
rect 38994 17726 39006 17778
rect 39058 17726 39070 17778
rect 40898 17726 40910 17778
rect 40962 17726 40974 17778
rect 30550 17714 30602 17726
rect 43150 17714 43202 17726
rect 5518 17666 5570 17678
rect 5518 17602 5570 17614
rect 5742 17666 5794 17678
rect 5742 17602 5794 17614
rect 6414 17666 6466 17678
rect 6414 17602 6466 17614
rect 9998 17666 10050 17678
rect 9998 17602 10050 17614
rect 10110 17666 10162 17678
rect 12798 17666 12850 17678
rect 10882 17614 10894 17666
rect 10946 17614 10958 17666
rect 10110 17602 10162 17614
rect 12798 17602 12850 17614
rect 14200 17666 14252 17678
rect 14478 17666 14530 17678
rect 14354 17614 14366 17666
rect 14418 17614 14430 17666
rect 14200 17602 14252 17614
rect 14478 17602 14530 17614
rect 15262 17666 15314 17678
rect 15262 17602 15314 17614
rect 17950 17666 18002 17678
rect 17950 17602 18002 17614
rect 18734 17666 18786 17678
rect 19014 17666 19066 17678
rect 18834 17614 18846 17666
rect 18898 17614 18910 17666
rect 18734 17602 18786 17614
rect 19014 17602 19066 17614
rect 19182 17666 19234 17678
rect 19182 17602 19234 17614
rect 20078 17666 20130 17678
rect 22430 17666 22482 17678
rect 20078 17602 20130 17614
rect 20302 17627 20354 17639
rect 20738 17614 20750 17666
rect 20802 17614 20814 17666
rect 21186 17614 21198 17666
rect 21250 17614 21262 17666
rect 21746 17614 21758 17666
rect 21810 17614 21822 17666
rect 4230 17554 4282 17566
rect 4230 17490 4282 17502
rect 4678 17554 4730 17566
rect 4678 17490 4730 17502
rect 9102 17554 9154 17566
rect 20302 17563 20354 17575
rect 22082 17558 22094 17610
rect 22146 17558 22158 17610
rect 22430 17602 22482 17614
rect 22766 17666 22818 17678
rect 25118 17666 25170 17678
rect 23426 17614 23438 17666
rect 23490 17614 23502 17666
rect 23650 17614 23662 17666
rect 23714 17614 23726 17666
rect 22766 17602 22818 17614
rect 25118 17602 25170 17614
rect 25230 17666 25282 17678
rect 25230 17602 25282 17614
rect 25454 17666 25506 17678
rect 25454 17602 25506 17614
rect 26462 17666 26514 17678
rect 26910 17666 26962 17678
rect 26786 17614 26798 17666
rect 26850 17614 26862 17666
rect 26462 17602 26514 17614
rect 26618 17558 26630 17610
rect 26682 17558 26694 17610
rect 26910 17602 26962 17614
rect 27190 17666 27242 17678
rect 32174 17666 32226 17678
rect 35814 17666 35866 17678
rect 36094 17666 36146 17678
rect 28130 17614 28142 17666
rect 28194 17614 28206 17666
rect 28466 17614 28478 17666
rect 28530 17614 28542 17666
rect 27190 17602 27242 17614
rect 29094 17610 29146 17622
rect 29474 17614 29486 17666
rect 29538 17614 29550 17666
rect 29698 17586 29710 17638
rect 29762 17586 29774 17638
rect 30706 17614 30718 17666
rect 30770 17614 30782 17666
rect 32946 17614 32958 17666
rect 33010 17614 33022 17666
rect 35970 17614 35982 17666
rect 36034 17614 36046 17666
rect 32174 17602 32226 17614
rect 35814 17602 35866 17614
rect 36094 17602 36146 17614
rect 38110 17666 38162 17678
rect 38110 17602 38162 17614
rect 38222 17666 38274 17678
rect 38222 17602 38274 17614
rect 41358 17666 41410 17678
rect 41636 17666 41688 17678
rect 41458 17614 41470 17666
rect 41522 17614 41534 17666
rect 41358 17602 41410 17614
rect 41636 17602 41688 17614
rect 42478 17666 42530 17678
rect 42756 17666 42808 17678
rect 45278 17666 45330 17678
rect 42578 17614 42590 17666
rect 42642 17614 42654 17666
rect 43698 17614 43710 17666
rect 43762 17614 43774 17666
rect 43922 17614 43934 17666
rect 43986 17614 43998 17666
rect 42478 17602 42530 17614
rect 42756 17602 42808 17614
rect 45278 17602 45330 17614
rect 45390 17666 45442 17678
rect 46162 17614 46174 17666
rect 46226 17614 46238 17666
rect 45390 17602 45442 17614
rect 9102 17490 9154 17502
rect 21366 17498 21418 17510
rect 25722 17502 25734 17554
rect 25786 17502 25798 17554
rect 29094 17546 29146 17558
rect 34862 17554 34914 17566
rect 15094 17442 15146 17454
rect 34862 17490 34914 17502
rect 48078 17554 48130 17566
rect 48078 17490 48130 17502
rect 21366 17434 21418 17446
rect 27750 17442 27802 17454
rect 15094 17378 15146 17390
rect 27750 17378 27802 17390
rect 44942 17442 44994 17454
rect 44942 17378 44994 17390
rect 1344 17274 48608 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 48608 17274
rect 1344 17188 48608 17222
rect 4342 17106 4394 17118
rect 4342 17042 4394 17054
rect 16606 17106 16658 17118
rect 16606 17042 16658 17054
rect 21198 17106 21250 17118
rect 21198 17042 21250 17054
rect 23382 17106 23434 17118
rect 12126 16994 12178 17006
rect 22530 16998 22542 17050
rect 22594 16998 22606 17050
rect 23382 17042 23434 17054
rect 23718 17106 23770 17118
rect 23718 17042 23770 17054
rect 24334 17106 24386 17118
rect 24334 17042 24386 17054
rect 25342 17106 25394 17118
rect 25342 17042 25394 17054
rect 26686 17106 26738 17118
rect 26686 17042 26738 17054
rect 27246 17106 27298 17118
rect 27246 17042 27298 17054
rect 29430 17106 29482 17118
rect 40182 17106 40234 17118
rect 29430 17042 29482 17054
rect 34246 17050 34298 17062
rect 12126 16930 12178 16942
rect 28478 16994 28530 17006
rect 5070 16882 5122 16894
rect 5070 16818 5122 16830
rect 5182 16882 5234 16894
rect 5182 16818 5234 16830
rect 8766 16882 8818 16894
rect 8766 16818 8818 16830
rect 8990 16882 9042 16894
rect 8990 16818 9042 16830
rect 9438 16882 9490 16894
rect 9438 16818 9490 16830
rect 12910 16882 12962 16894
rect 12910 16818 12962 16830
rect 13022 16882 13074 16894
rect 13022 16818 13074 16830
rect 13358 16882 13410 16894
rect 13358 16818 13410 16830
rect 16942 16882 16994 16894
rect 17602 16830 17614 16882
rect 17666 16830 17678 16882
rect 17938 16874 17950 16926
rect 18002 16874 18014 16926
rect 18924 16919 18976 16931
rect 19182 16882 19234 16894
rect 18924 16855 18976 16867
rect 19058 16830 19070 16882
rect 19122 16830 19134 16882
rect 16942 16818 16994 16830
rect 19182 16818 19234 16830
rect 19686 16882 19738 16894
rect 20178 16886 20190 16938
rect 20242 16886 20254 16938
rect 21534 16882 21586 16894
rect 22194 16886 22206 16938
rect 22258 16886 22270 16938
rect 22430 16882 22482 16894
rect 23998 16882 24050 16894
rect 20402 16830 20414 16882
rect 20466 16830 20478 16882
rect 19686 16818 19738 16830
rect 20806 16826 20858 16838
rect 3894 16770 3946 16782
rect 3894 16706 3946 16718
rect 4734 16770 4786 16782
rect 20638 16770 20690 16782
rect 5954 16718 5966 16770
rect 6018 16718 6030 16770
rect 7858 16718 7870 16770
rect 7922 16718 7934 16770
rect 10210 16718 10222 16770
rect 10274 16718 10286 16770
rect 14130 16718 14142 16770
rect 14194 16718 14206 16770
rect 16034 16718 16046 16770
rect 16098 16718 16110 16770
rect 18050 16718 18062 16770
rect 18114 16718 18126 16770
rect 21746 16830 21758 16882
rect 21810 16830 21822 16882
rect 23874 16830 23886 16882
rect 23938 16830 23950 16882
rect 21534 16818 21586 16830
rect 22430 16818 22482 16830
rect 23998 16818 24050 16830
rect 25678 16882 25730 16894
rect 26350 16882 26402 16894
rect 26114 16830 26126 16882
rect 26178 16830 26190 16882
rect 25678 16818 25730 16830
rect 26350 16818 26402 16830
rect 27582 16882 27634 16894
rect 27582 16818 27634 16830
rect 28142 16882 28194 16894
rect 28298 16886 28310 16938
rect 28362 16886 28374 16938
rect 28478 16930 28530 16942
rect 28870 16994 28922 17006
rect 28870 16930 28922 16942
rect 33182 16994 33234 17006
rect 34246 16986 34298 16998
rect 34694 17050 34746 17062
rect 40182 17042 40234 17054
rect 34694 16986 34746 16998
rect 37662 16994 37714 17006
rect 33182 16930 33234 16942
rect 33854 16938 33906 16950
rect 28142 16818 28194 16830
rect 28590 16882 28642 16894
rect 28590 16818 28642 16830
rect 32622 16882 32674 16894
rect 32622 16818 32674 16830
rect 33014 16882 33066 16894
rect 33618 16886 33630 16938
rect 33682 16886 33694 16938
rect 37662 16930 37714 16942
rect 46510 16994 46562 17006
rect 46510 16930 46562 16942
rect 33854 16874 33906 16886
rect 34862 16902 34914 16914
rect 34402 16830 34414 16882
rect 34466 16830 34478 16882
rect 34862 16838 34914 16850
rect 34974 16882 35026 16894
rect 33014 16818 33066 16830
rect 34974 16818 35026 16830
rect 38446 16882 38498 16894
rect 38446 16818 38498 16830
rect 38558 16882 38610 16894
rect 38770 16830 38782 16882
rect 38834 16830 38846 16882
rect 40898 16857 40910 16909
rect 40962 16857 40974 16909
rect 43138 16830 43150 16882
rect 43202 16830 43214 16882
rect 43810 16874 43822 16926
rect 43874 16874 43886 16926
rect 44382 16882 44434 16894
rect 44034 16830 44046 16882
rect 44098 16830 44110 16882
rect 38558 16818 38610 16830
rect 44382 16818 44434 16830
rect 44606 16882 44658 16894
rect 44874 16830 44886 16882
rect 44938 16830 44950 16882
rect 45378 16863 45390 16915
rect 45442 16863 45454 16915
rect 45602 16863 45614 16915
rect 45666 16863 45678 16915
rect 46050 16863 46062 16915
rect 46114 16863 46126 16915
rect 46360 16863 46372 16915
rect 46424 16863 46436 16915
rect 47966 16882 48018 16894
rect 46946 16830 46958 16882
rect 47010 16830 47022 16882
rect 47282 16830 47294 16882
rect 47346 16830 47358 16882
rect 47674 16830 47686 16882
rect 47738 16830 47750 16882
rect 44606 16818 44658 16830
rect 47966 16818 48018 16830
rect 48078 16882 48130 16894
rect 48078 16818 48130 16830
rect 20806 16762 20858 16774
rect 29922 16718 29934 16770
rect 29986 16718 29998 16770
rect 31826 16718 31838 16770
rect 31890 16718 31902 16770
rect 35746 16718 35758 16770
rect 35810 16718 35822 16770
rect 43698 16718 43710 16770
rect 43762 16718 43774 16770
rect 4734 16706 4786 16718
rect 20638 16706 20690 16718
rect 46846 16714 46898 16726
rect 18510 16658 18562 16670
rect 2258 16606 2270 16658
rect 2322 16655 2334 16658
rect 3042 16655 3054 16658
rect 2322 16609 3054 16655
rect 2322 16606 2334 16609
rect 3042 16606 3054 16609
rect 3106 16606 3118 16658
rect 8474 16606 8486 16658
rect 8538 16606 8550 16658
rect 12618 16606 12630 16658
rect 12682 16606 12694 16658
rect 18510 16594 18562 16606
rect 25958 16658 26010 16670
rect 38154 16606 38166 16658
rect 38218 16606 38230 16658
rect 46846 16650 46898 16662
rect 25958 16594 26010 16606
rect 1344 16490 48608 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 48608 16490
rect 1344 16404 48608 16438
rect 22990 16322 23042 16334
rect 22990 16258 23042 16270
rect 25342 16322 25394 16334
rect 25342 16258 25394 16270
rect 32510 16322 32562 16334
rect 32510 16258 32562 16270
rect 44998 16322 45050 16334
rect 44998 16258 45050 16270
rect 14982 16210 15034 16222
rect 22038 16210 22090 16222
rect 7186 16158 7198 16210
rect 7250 16158 7262 16210
rect 8306 16158 8318 16210
rect 8370 16158 8382 16210
rect 12450 16158 12462 16210
rect 12514 16158 12526 16210
rect 16034 16158 16046 16210
rect 16098 16158 16110 16210
rect 16818 16158 16830 16210
rect 16882 16158 16894 16210
rect 33742 16210 33794 16222
rect 14982 16146 15034 16158
rect 22038 16146 22090 16158
rect 29654 16154 29706 16166
rect 2270 16098 2322 16110
rect 6638 16098 6690 16110
rect 9326 16098 9378 16110
rect 13582 16098 13634 16110
rect 15598 16098 15650 16110
rect 3042 16046 3054 16098
rect 3106 16046 3118 16098
rect 5954 16046 5966 16098
rect 6018 16046 6030 16098
rect 6414 16059 6466 16071
rect 2270 16034 2322 16046
rect 6638 16034 6690 16046
rect 4958 15986 5010 15998
rect 6414 15995 6466 16007
rect 7298 16002 7310 16054
rect 7362 16002 7374 16054
rect 7634 16046 7646 16098
rect 7698 16046 7710 16098
rect 8418 16031 8430 16083
rect 8482 16031 8494 16083
rect 8754 16046 8766 16098
rect 8818 16046 8830 16098
rect 10098 16046 10110 16098
rect 10162 16046 10174 16098
rect 9326 16034 9378 16046
rect 12562 16002 12574 16054
rect 12626 16002 12638 16054
rect 12898 16046 12910 16098
rect 12962 16046 12974 16098
rect 13414 16042 13466 16054
rect 4958 15922 5010 15934
rect 12014 15986 12066 15998
rect 13794 16046 13806 16098
rect 13858 16046 13870 16098
rect 13582 16034 13634 16046
rect 14142 16042 14194 16054
rect 13414 15978 13466 15990
rect 15598 16034 15650 16046
rect 15822 16098 15874 16110
rect 22318 16098 22370 16110
rect 23326 16098 23378 16110
rect 15822 16034 15874 16046
rect 16146 16031 16158 16083
rect 16210 16031 16222 16083
rect 16482 16046 16494 16098
rect 16546 16046 16558 16098
rect 16930 16031 16942 16083
rect 16994 16031 17006 16083
rect 17266 16046 17278 16098
rect 17330 16046 17342 16098
rect 17826 16046 17838 16098
rect 17890 16046 17902 16098
rect 19730 16018 19742 16070
rect 19794 16018 19806 16070
rect 20290 16046 20302 16098
rect 20354 16046 20366 16098
rect 21186 16046 21198 16098
rect 21250 16046 21262 16098
rect 22418 16046 22430 16098
rect 22482 16046 22494 16098
rect 22318 16034 22370 16046
rect 22586 15990 22598 16042
rect 22650 15990 22662 16042
rect 23326 16034 23378 16046
rect 24894 16098 24946 16110
rect 24894 16034 24946 16046
rect 25006 16098 25058 16110
rect 25006 16034 25058 16046
rect 26238 16098 26290 16110
rect 26238 16034 26290 16046
rect 26910 16098 26962 16110
rect 26910 16034 26962 16046
rect 27582 16098 27634 16110
rect 29486 16098 29538 16110
rect 28690 16046 28702 16098
rect 28754 16046 28766 16098
rect 36486 16210 36538 16222
rect 33742 16146 33794 16158
rect 34694 16154 34746 16166
rect 29654 16090 29706 16102
rect 29934 16098 29986 16110
rect 29810 16046 29822 16098
rect 29874 16046 29886 16098
rect 27582 16034 27634 16046
rect 29486 16034 29538 16046
rect 29934 16034 29986 16046
rect 30214 16098 30266 16110
rect 33574 16098 33626 16110
rect 36486 16146 36538 16158
rect 42926 16210 42978 16222
rect 48134 16210 48186 16222
rect 43362 16158 43374 16210
rect 43426 16158 43438 16210
rect 42926 16146 42978 16158
rect 48134 16146 48186 16158
rect 30214 16034 30266 16046
rect 31154 16018 31166 16070
rect 31218 16018 31230 16070
rect 33954 16046 33966 16098
rect 34018 16046 34030 16098
rect 34694 16090 34746 16102
rect 37662 16098 37714 16110
rect 42254 16098 42306 16110
rect 42534 16098 42586 16110
rect 47070 16098 47122 16110
rect 33574 16034 33626 16046
rect 34178 16018 34190 16070
rect 34242 16018 34254 16070
rect 35074 16046 35086 16098
rect 35138 16046 35150 16098
rect 35422 16042 35474 16054
rect 37202 16046 37214 16098
rect 37266 16046 37278 16098
rect 38434 16046 38446 16098
rect 38498 16046 38510 16098
rect 41570 16046 41582 16098
rect 41634 16046 41646 16098
rect 14142 15978 14194 15990
rect 34862 15986 34914 15998
rect 15306 15934 15318 15986
rect 15370 15934 15382 15986
rect 6066 15878 6078 15930
rect 6130 15878 6142 15930
rect 12014 15922 12066 15934
rect 28534 15930 28586 15942
rect 20470 15874 20522 15886
rect 20470 15810 20522 15822
rect 21366 15874 21418 15886
rect 21366 15810 21418 15822
rect 23662 15874 23714 15886
rect 23662 15810 23714 15822
rect 24558 15874 24610 15886
rect 24558 15810 24610 15822
rect 26070 15874 26122 15886
rect 26070 15810 26122 15822
rect 26574 15874 26626 15886
rect 26574 15810 26626 15822
rect 27246 15874 27298 15886
rect 27246 15810 27298 15822
rect 27918 15874 27970 15886
rect 37662 16034 37714 16046
rect 41974 16042 42026 16054
rect 35422 15978 35474 15990
rect 40350 15986 40402 15998
rect 41346 15990 41358 16042
rect 41410 15990 41422 16042
rect 34862 15922 34914 15934
rect 40350 15922 40402 15934
rect 41806 15986 41858 15998
rect 42354 16046 42366 16098
rect 42418 16046 42430 16098
rect 42254 16034 42306 16046
rect 42534 16034 42586 16046
rect 43474 16031 43486 16083
rect 43538 16031 43550 16083
rect 43698 16046 43710 16098
rect 43762 16046 43774 16098
rect 44034 16046 44046 16098
rect 44098 16046 44110 16098
rect 44818 16046 44830 16098
rect 44882 16046 44894 16098
rect 45378 15990 45390 16042
rect 45442 15990 45454 16042
rect 45714 15990 45726 16042
rect 45778 15990 45790 16042
rect 46162 15990 46174 16042
rect 46226 15990 46238 16042
rect 46430 16006 46442 16058
rect 46494 16006 46506 16058
rect 47070 16034 47122 16046
rect 47294 16098 47346 16110
rect 47294 16034 47346 16046
rect 41974 15978 42026 15990
rect 46622 15986 46674 15998
rect 41806 15922 41858 15934
rect 47562 15934 47574 15986
rect 47626 15934 47638 15986
rect 46622 15922 46674 15934
rect 28534 15866 28586 15878
rect 36038 15874 36090 15886
rect 27918 15810 27970 15822
rect 36038 15810 36090 15822
rect 37046 15874 37098 15886
rect 37046 15810 37098 15822
rect 44214 15874 44266 15886
rect 44214 15810 44266 15822
rect 1344 15706 48608 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 48608 15706
rect 1344 15620 48608 15654
rect 3502 15538 3554 15550
rect 3502 15474 3554 15486
rect 7142 15538 7194 15550
rect 5058 15430 5070 15482
rect 5122 15430 5134 15482
rect 7142 15474 7194 15486
rect 11790 15538 11842 15550
rect 11790 15474 11842 15486
rect 13582 15538 13634 15550
rect 13582 15474 13634 15486
rect 15766 15538 15818 15550
rect 15766 15474 15818 15486
rect 16606 15538 16658 15550
rect 16606 15474 16658 15486
rect 9662 15426 9714 15438
rect 9662 15362 9714 15374
rect 16214 15426 16266 15438
rect 3838 15314 3890 15326
rect 4274 15262 4286 15314
rect 4338 15262 4350 15314
rect 4498 15306 4510 15358
rect 4562 15306 4574 15358
rect 4946 15262 4958 15314
rect 5010 15262 5022 15314
rect 5282 15289 5294 15341
rect 5346 15289 5358 15341
rect 5630 15314 5682 15326
rect 6178 15262 6190 15314
rect 6242 15262 6254 15314
rect 6514 15277 6526 15329
rect 6578 15277 6590 15329
rect 7422 15314 7474 15326
rect 7298 15262 7310 15314
rect 7362 15262 7374 15314
rect 3838 15250 3890 15262
rect 5630 15250 5682 15262
rect 7422 15250 7474 15262
rect 7758 15314 7810 15326
rect 7758 15250 7810 15262
rect 8206 15314 8258 15326
rect 8486 15314 8538 15326
rect 8306 15262 8318 15314
rect 8370 15262 8382 15314
rect 8206 15250 8258 15262
rect 8486 15250 8538 15262
rect 9494 15314 9546 15326
rect 10098 15290 10110 15342
rect 10162 15290 10174 15342
rect 13122 15289 13134 15341
rect 13186 15289 13198 15341
rect 13918 15314 13970 15326
rect 9494 15250 9546 15262
rect 8878 15202 8930 15214
rect 10322 15206 10334 15258
rect 10386 15206 10398 15258
rect 13918 15250 13970 15262
rect 14198 15314 14250 15326
rect 14198 15250 14250 15262
rect 14478 15314 14530 15326
rect 14746 15318 14758 15370
rect 14810 15318 14822 15370
rect 16214 15362 16266 15374
rect 21422 15426 21474 15438
rect 21422 15362 21474 15374
rect 26182 15426 26234 15438
rect 22168 15352 22220 15364
rect 26182 15362 26234 15374
rect 27974 15426 28026 15438
rect 27974 15362 28026 15374
rect 35646 15426 35698 15438
rect 35646 15362 35698 15374
rect 36206 15426 36258 15438
rect 37382 15426 37434 15438
rect 36206 15362 36258 15374
rect 36766 15370 36818 15382
rect 14926 15314 14978 15326
rect 14578 15262 14590 15314
rect 14642 15262 14654 15314
rect 14478 15250 14530 15262
rect 14926 15250 14978 15262
rect 16942 15314 16994 15326
rect 18734 15314 18786 15326
rect 21870 15314 21922 15326
rect 17490 15262 17502 15314
rect 17554 15262 17566 15314
rect 19506 15262 19518 15314
rect 19570 15262 19582 15314
rect 21970 15262 21982 15314
rect 22034 15262 22046 15314
rect 22168 15288 22220 15300
rect 23774 15314 23826 15326
rect 16942 15250 16994 15262
rect 18734 15250 18786 15262
rect 21870 15250 21922 15262
rect 23774 15250 23826 15262
rect 23886 15314 23938 15326
rect 23886 15250 23938 15262
rect 27246 15314 27298 15326
rect 27694 15314 27746 15326
rect 27246 15250 27298 15262
rect 27414 15258 27466 15270
rect 27570 15262 27582 15314
rect 27634 15262 27646 15314
rect 4610 15150 4622 15202
rect 4674 15150 4686 15202
rect 6626 15150 6638 15202
rect 6690 15150 6702 15202
rect 8878 15138 8930 15150
rect 22542 15202 22594 15214
rect 22542 15138 22594 15150
rect 23438 15202 23490 15214
rect 23438 15138 23490 15150
rect 25734 15202 25786 15214
rect 25734 15138 25786 15150
rect 26630 15202 26682 15214
rect 27694 15250 27746 15262
rect 28534 15314 28586 15326
rect 28534 15250 28586 15262
rect 28926 15314 28978 15326
rect 29374 15314 29426 15326
rect 28926 15250 28978 15262
rect 29094 15258 29146 15270
rect 29250 15262 29262 15314
rect 29314 15262 29326 15314
rect 30370 15289 30382 15341
rect 30434 15289 30446 15341
rect 32958 15314 33010 15326
rect 27414 15194 27466 15206
rect 29374 15250 29426 15262
rect 33730 15262 33742 15314
rect 33794 15262 33806 15314
rect 36766 15306 36818 15318
rect 36878 15370 36930 15382
rect 37382 15362 37434 15374
rect 45614 15426 45666 15438
rect 36878 15306 36930 15318
rect 37550 15314 37602 15326
rect 32958 15250 33010 15262
rect 36038 15258 36090 15270
rect 29094 15194 29146 15206
rect 29654 15202 29706 15214
rect 26630 15138 26682 15150
rect 37550 15250 37602 15262
rect 40910 15314 40962 15326
rect 40910 15250 40962 15262
rect 41918 15314 41970 15326
rect 41918 15250 41970 15262
rect 42254 15314 42306 15326
rect 42634 15318 42646 15370
rect 42698 15318 42710 15370
rect 43520 15351 43572 15363
rect 45614 15362 45666 15374
rect 43262 15314 43314 15326
rect 42914 15262 42926 15314
rect 42978 15262 42990 15314
rect 43362 15262 43374 15314
rect 43426 15262 43438 15314
rect 43520 15287 43572 15299
rect 44482 15262 44494 15314
rect 44546 15262 44558 15314
rect 44706 15306 44718 15358
rect 44770 15306 44782 15358
rect 48302 15314 48354 15326
rect 47506 15262 47518 15314
rect 47570 15262 47582 15314
rect 42254 15250 42306 15262
rect 43262 15250 43314 15262
rect 48302 15250 48354 15262
rect 36038 15194 36090 15206
rect 41246 15202 41298 15214
rect 38322 15150 38334 15202
rect 38386 15150 38398 15202
rect 40226 15150 40238 15202
rect 40290 15150 40302 15202
rect 29654 15138 29706 15150
rect 41246 15138 41298 15150
rect 42590 15202 42642 15214
rect 42590 15138 42642 15150
rect 43934 15202 43986 15214
rect 44818 15150 44830 15202
rect 44882 15150 44894 15202
rect 43934 15138 43986 15150
rect 24222 15090 24274 15102
rect 24222 15026 24274 15038
rect 1344 14922 48608 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 48608 14922
rect 1344 14836 48608 14870
rect 11342 14754 11394 14766
rect 11342 14690 11394 14702
rect 12854 14754 12906 14766
rect 12854 14690 12906 14702
rect 23326 14754 23378 14766
rect 23326 14690 23378 14702
rect 23998 14754 24050 14766
rect 23998 14690 24050 14702
rect 28534 14754 28586 14766
rect 28534 14690 28586 14702
rect 30494 14754 30546 14766
rect 30494 14690 30546 14702
rect 43150 14754 43202 14766
rect 43150 14690 43202 14702
rect 46846 14698 46898 14710
rect 9662 14642 9714 14654
rect 5730 14590 5742 14642
rect 5794 14590 5806 14642
rect 9662 14578 9714 14590
rect 10222 14642 10274 14654
rect 22150 14642 22202 14654
rect 38110 14642 38162 14654
rect 16034 14590 16046 14642
rect 16098 14590 16110 14642
rect 17938 14590 17950 14642
rect 18002 14590 18014 14642
rect 18386 14590 18398 14642
rect 18450 14590 18462 14642
rect 10222 14578 10274 14590
rect 22150 14578 22202 14590
rect 29318 14586 29370 14598
rect 36306 14590 36318 14642
rect 36370 14590 36382 14642
rect 2046 14530 2098 14542
rect 4734 14530 4786 14542
rect 8094 14530 8146 14542
rect 2818 14478 2830 14530
rect 2882 14478 2894 14530
rect 2046 14466 2098 14478
rect 4734 14466 4786 14478
rect 5842 14463 5854 14515
rect 5906 14463 5918 14515
rect 6066 14478 6078 14530
rect 6130 14478 6142 14530
rect 6514 14478 6526 14530
rect 6578 14478 6590 14530
rect 6794 14422 6806 14474
rect 6858 14422 6870 14474
rect 8094 14466 8146 14478
rect 8766 14530 8818 14542
rect 10616 14530 10668 14542
rect 10894 14530 10946 14542
rect 12462 14530 12514 14542
rect 15262 14530 15314 14542
rect 19518 14530 19570 14542
rect 8766 14466 8818 14478
rect 9102 14474 9154 14486
rect 9426 14478 9438 14530
rect 9490 14478 9502 14530
rect 9102 14410 9154 14422
rect 9830 14474 9882 14486
rect 10770 14478 10782 14530
rect 10834 14478 10846 14530
rect 11573 14478 11585 14530
rect 11637 14478 11649 14530
rect 12674 14478 12686 14530
rect 12738 14478 12750 14530
rect 14018 14478 14030 14530
rect 14082 14478 14094 14530
rect 10616 14466 10668 14478
rect 10894 14466 10946 14478
rect 12462 14466 12514 14478
rect 14254 14474 14306 14486
rect 9830 14410 9882 14422
rect 14254 14410 14306 14422
rect 14366 14474 14418 14486
rect 15094 14474 15146 14486
rect 14366 14410 14418 14422
rect 14926 14418 14978 14430
rect 15262 14466 15314 14478
rect 18498 14463 18510 14515
rect 18562 14463 18574 14515
rect 18722 14478 18734 14530
rect 18786 14478 18798 14530
rect 19518 14466 19570 14478
rect 20190 14530 20242 14542
rect 20190 14466 20242 14478
rect 21758 14530 21810 14542
rect 21758 14466 21810 14478
rect 22318 14530 22370 14542
rect 22318 14466 22370 14478
rect 22990 14530 23042 14542
rect 22990 14466 23042 14478
rect 23662 14530 23714 14542
rect 23662 14466 23714 14478
rect 24334 14530 24386 14542
rect 24334 14466 24386 14478
rect 24670 14530 24722 14542
rect 24670 14466 24722 14478
rect 25902 14530 25954 14542
rect 25902 14466 25954 14478
rect 26686 14530 26738 14542
rect 26686 14466 26738 14478
rect 26854 14530 26906 14542
rect 26854 14466 26906 14478
rect 27134 14530 27186 14542
rect 27134 14466 27186 14478
rect 27806 14530 27858 14542
rect 27806 14466 27858 14478
rect 28254 14530 28306 14542
rect 15094 14410 15146 14422
rect 26238 14418 26290 14430
rect 6626 14310 6638 14362
rect 6690 14310 6702 14362
rect 14926 14354 14978 14366
rect 26238 14354 26290 14366
rect 27022 14418 27074 14430
rect 27022 14354 27074 14366
rect 27414 14418 27466 14430
rect 27962 14422 27974 14474
rect 28026 14422 28038 14474
rect 28254 14466 28306 14478
rect 29150 14530 29202 14542
rect 38110 14578 38162 14590
rect 39230 14642 39282 14654
rect 44146 14646 44158 14698
rect 44210 14646 44222 14698
rect 39230 14578 39282 14590
rect 45166 14642 45218 14654
rect 45166 14578 45218 14590
rect 46566 14642 46618 14654
rect 46846 14634 46898 14646
rect 47798 14642 47850 14654
rect 46566 14578 46618 14590
rect 47798 14578 47850 14590
rect 29318 14522 29370 14534
rect 29598 14530 29650 14542
rect 29150 14466 29202 14478
rect 29598 14466 29650 14478
rect 30158 14530 30210 14542
rect 33630 14530 33682 14542
rect 42366 14530 42418 14542
rect 30158 14466 30210 14478
rect 30930 14450 30942 14502
rect 30994 14450 31006 14502
rect 33170 14478 33182 14530
rect 33234 14478 33246 14530
rect 34402 14478 34414 14530
rect 34466 14478 34478 14530
rect 37202 14478 37214 14530
rect 37266 14478 37278 14530
rect 33630 14466 33682 14478
rect 37942 14474 37994 14486
rect 38322 14478 38334 14530
rect 38386 14478 38398 14530
rect 39062 14474 39114 14486
rect 39442 14478 39454 14530
rect 39506 14478 39518 14530
rect 40450 14478 40462 14530
rect 40514 14478 40526 14530
rect 41122 14478 41134 14530
rect 41186 14478 41198 14530
rect 41682 14478 41694 14530
rect 41746 14478 41758 14530
rect 27414 14354 27466 14366
rect 28142 14418 28194 14430
rect 28142 14354 28194 14366
rect 29486 14418 29538 14430
rect 29486 14354 29538 14366
rect 29878 14418 29930 14430
rect 38546 14422 38558 14474
rect 38610 14422 38622 14474
rect 39666 14422 39678 14474
rect 39730 14422 39742 14474
rect 42018 14422 42030 14474
rect 42082 14422 42094 14474
rect 42366 14466 42418 14478
rect 42814 14530 42866 14542
rect 45502 14530 45554 14542
rect 43922 14478 43934 14530
rect 43986 14478 43998 14530
rect 44258 14478 44270 14530
rect 44322 14478 44334 14530
rect 44818 14478 44830 14530
rect 44882 14478 44894 14530
rect 42814 14466 42866 14478
rect 45154 14422 45166 14474
rect 45218 14422 45230 14474
rect 45502 14466 45554 14478
rect 45838 14530 45890 14542
rect 46946 14478 46958 14530
rect 47010 14478 47022 14530
rect 47282 14478 47294 14530
rect 47346 14478 47358 14530
rect 45838 14466 45890 14478
rect 37942 14410 37994 14422
rect 39062 14410 39114 14422
rect 29878 14354 29930 14366
rect 40294 14362 40346 14374
rect 7758 14306 7810 14318
rect 7758 14242 7810 14254
rect 8430 14306 8482 14318
rect 8430 14242 8482 14254
rect 13862 14306 13914 14318
rect 13862 14242 13914 14254
rect 19350 14306 19402 14318
rect 19350 14242 19402 14254
rect 19854 14306 19906 14318
rect 19854 14242 19906 14254
rect 20526 14306 20578 14318
rect 20526 14242 20578 14254
rect 21422 14306 21474 14318
rect 21422 14242 21474 14254
rect 22654 14306 22706 14318
rect 22654 14242 22706 14254
rect 25734 14306 25786 14318
rect 25734 14242 25786 14254
rect 37046 14306 37098 14318
rect 37046 14242 37098 14254
rect 37718 14306 37770 14318
rect 40294 14298 40346 14310
rect 40966 14362 41018 14374
rect 42466 14310 42478 14362
rect 42530 14310 42542 14362
rect 40966 14298 41018 14310
rect 48246 14306 48298 14318
rect 37718 14242 37770 14254
rect 48246 14242 48298 14254
rect 1344 14138 48608 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 48608 14138
rect 1344 14052 48608 14086
rect 3166 13970 3218 13982
rect 3166 13906 3218 13918
rect 4902 13970 4954 13982
rect 4902 13906 4954 13918
rect 5406 13970 5458 13982
rect 5406 13906 5458 13918
rect 22934 13970 22986 13982
rect 5954 13862 5966 13914
rect 6018 13862 6030 13914
rect 22934 13906 22986 13918
rect 28870 13970 28922 13982
rect 28870 13906 28922 13918
rect 29318 13970 29370 13982
rect 29318 13906 29370 13918
rect 39958 13970 40010 13982
rect 39958 13906 40010 13918
rect 41414 13970 41466 13982
rect 41414 13906 41466 13918
rect 48134 13970 48186 13982
rect 48134 13906 48186 13918
rect 16718 13858 16770 13870
rect 6302 13785 6354 13797
rect 3502 13746 3554 13758
rect 3502 13682 3554 13694
rect 5070 13746 5122 13758
rect 5842 13694 5854 13746
rect 5906 13694 5918 13746
rect 10076 13784 10128 13796
rect 6302 13721 6354 13733
rect 6526 13746 6578 13758
rect 5070 13682 5122 13694
rect 6526 13682 6578 13694
rect 7758 13746 7810 13758
rect 7758 13682 7810 13694
rect 8430 13746 8482 13758
rect 8430 13682 8482 13694
rect 8542 13746 8594 13758
rect 16158 13784 16210 13796
rect 16718 13794 16770 13806
rect 30606 13858 30658 13870
rect 10334 13746 10386 13758
rect 10076 13720 10128 13732
rect 10210 13694 10222 13746
rect 10274 13694 10286 13746
rect 8542 13682 8594 13694
rect 10334 13682 10386 13694
rect 10558 13746 10610 13758
rect 10558 13682 10610 13694
rect 11566 13746 11618 13758
rect 14254 13746 14306 13758
rect 12338 13694 12350 13746
rect 12402 13694 12414 13746
rect 15138 13722 15150 13774
rect 15202 13722 15214 13774
rect 15766 13746 15818 13758
rect 15362 13694 15374 13746
rect 15426 13694 15438 13746
rect 17614 13746 17666 13758
rect 16158 13720 16210 13732
rect 16482 13694 16494 13746
rect 16546 13694 16558 13746
rect 11566 13682 11618 13694
rect 14254 13682 14306 13694
rect 15766 13682 15818 13694
rect 16886 13690 16938 13702
rect 8878 13634 8930 13646
rect 8878 13570 8930 13582
rect 9662 13634 9714 13646
rect 9662 13570 9714 13582
rect 15598 13634 15650 13646
rect 17614 13682 17666 13694
rect 17838 13746 17890 13758
rect 20862 13746 20914 13758
rect 21130 13750 21142 13802
rect 21194 13750 21206 13802
rect 21310 13746 21362 13758
rect 18106 13694 18118 13746
rect 18170 13694 18182 13746
rect 18610 13694 18622 13746
rect 18674 13694 18686 13746
rect 18946 13694 18958 13746
rect 19010 13694 19022 13746
rect 19506 13694 19518 13746
rect 19570 13694 19582 13746
rect 19842 13694 19854 13746
rect 19906 13694 19918 13746
rect 20962 13694 20974 13746
rect 21026 13694 21038 13746
rect 17838 13682 17890 13694
rect 20862 13682 20914 13694
rect 21310 13682 21362 13694
rect 21982 13746 22034 13758
rect 22430 13746 22482 13758
rect 22082 13694 22094 13746
rect 22146 13694 22158 13746
rect 21982 13682 22034 13694
rect 22262 13690 22314 13702
rect 16886 13626 16938 13638
rect 22430 13682 22482 13694
rect 24222 13746 24274 13758
rect 24222 13682 24274 13694
rect 25230 13746 25282 13758
rect 25678 13746 25730 13758
rect 27022 13746 27074 13758
rect 25230 13682 25282 13694
rect 25398 13690 25450 13702
rect 25554 13694 25566 13746
rect 25618 13694 25630 13746
rect 26338 13694 26350 13746
rect 26402 13694 26414 13746
rect 26674 13694 26686 13746
rect 26738 13694 26750 13746
rect 22262 13626 22314 13638
rect 25678 13682 25730 13694
rect 27022 13682 27074 13694
rect 29486 13746 29538 13758
rect 29486 13682 29538 13694
rect 30270 13746 30322 13758
rect 30426 13750 30438 13802
rect 30490 13750 30502 13802
rect 30606 13794 30658 13806
rect 32118 13858 32170 13870
rect 36206 13858 36258 13870
rect 43038 13858 43090 13870
rect 32118 13794 32170 13806
rect 36038 13802 36090 13814
rect 30270 13682 30322 13694
rect 30718 13746 30770 13758
rect 30718 13682 30770 13694
rect 31390 13746 31442 13758
rect 31838 13746 31890 13758
rect 31390 13682 31442 13694
rect 31558 13690 31610 13702
rect 31714 13694 31726 13746
rect 31778 13694 31790 13746
rect 25398 13626 25450 13638
rect 27358 13634 27410 13646
rect 15598 13570 15650 13582
rect 18510 13578 18562 13590
rect 7422 13522 7474 13534
rect 7422 13458 7474 13470
rect 8094 13522 8146 13534
rect 8094 13458 8146 13470
rect 10894 13522 10946 13534
rect 18510 13514 18562 13526
rect 19406 13578 19458 13590
rect 26798 13578 26850 13590
rect 19406 13514 19458 13526
rect 20582 13522 20634 13534
rect 10894 13458 10946 13470
rect 20582 13458 20634 13470
rect 21702 13522 21754 13534
rect 21702 13458 21754 13470
rect 23886 13522 23938 13534
rect 23886 13458 23938 13470
rect 25958 13522 26010 13534
rect 31838 13682 31890 13694
rect 32958 13746 33010 13758
rect 36206 13794 36258 13806
rect 36878 13802 36930 13814
rect 38714 13806 38726 13858
rect 38778 13806 38790 13858
rect 45222 13858 45274 13870
rect 36038 13738 36090 13750
rect 36642 13722 36654 13774
rect 36706 13722 36718 13774
rect 42478 13784 42530 13796
rect 43038 13794 43090 13806
rect 43206 13802 43258 13814
rect 36878 13738 36930 13750
rect 37426 13722 37438 13774
rect 37490 13722 37502 13774
rect 38222 13746 38274 13758
rect 32958 13682 33010 13694
rect 38054 13690 38106 13702
rect 37202 13638 37214 13690
rect 37266 13638 37278 13690
rect 31558 13626 31610 13638
rect 37886 13634 37938 13646
rect 33730 13582 33742 13634
rect 33794 13582 33806 13634
rect 35634 13582 35646 13634
rect 35698 13582 35710 13634
rect 38222 13682 38274 13694
rect 38446 13746 38498 13758
rect 38446 13682 38498 13694
rect 42142 13746 42194 13758
rect 45222 13794 45274 13806
rect 42478 13720 42530 13732
rect 42802 13694 42814 13746
rect 42866 13694 42878 13746
rect 43206 13738 43258 13750
rect 43586 13738 43598 13790
rect 43650 13738 43662 13790
rect 44494 13746 44546 13758
rect 44942 13746 44994 13758
rect 46286 13746 46338 13758
rect 43810 13694 43822 13746
rect 43874 13694 43886 13746
rect 42142 13682 42194 13694
rect 44494 13682 44546 13694
rect 44662 13690 44714 13702
rect 44818 13694 44830 13746
rect 44882 13694 44894 13746
rect 45714 13694 45726 13746
rect 45778 13694 45790 13746
rect 45938 13694 45950 13746
rect 46002 13694 46014 13746
rect 38054 13626 38106 13638
rect 39286 13634 39338 13646
rect 27358 13570 27410 13582
rect 37886 13570 37938 13582
rect 39286 13570 39338 13582
rect 40406 13634 40458 13646
rect 44942 13682 44994 13694
rect 46286 13682 46338 13694
rect 46510 13746 46562 13758
rect 47282 13694 47294 13746
rect 47346 13694 47358 13746
rect 47506 13694 47518 13746
rect 47570 13694 47582 13746
rect 46510 13682 46562 13694
rect 43474 13582 43486 13634
rect 43538 13582 43550 13634
rect 44662 13626 44714 13638
rect 40406 13570 40458 13582
rect 26798 13514 26850 13526
rect 29822 13522 29874 13534
rect 25958 13458 26010 13470
rect 29822 13458 29874 13470
rect 30998 13522 31050 13534
rect 30998 13458 31050 13470
rect 41806 13522 41858 13534
rect 45714 13526 45726 13578
rect 45778 13526 45790 13578
rect 47282 13526 47294 13578
rect 47346 13526 47358 13578
rect 46778 13470 46790 13522
rect 46842 13470 46854 13522
rect 41806 13458 41858 13470
rect 1344 13354 48608 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 48608 13354
rect 1344 13268 48608 13302
rect 15150 13186 15202 13198
rect 15150 13122 15202 13134
rect 19854 13186 19906 13198
rect 19854 13122 19906 13134
rect 27078 13186 27130 13198
rect 27078 13122 27130 13134
rect 33070 13186 33122 13198
rect 36206 13186 36258 13198
rect 34682 13134 34694 13186
rect 34746 13134 34758 13186
rect 33070 13122 33122 13134
rect 36206 13122 36258 13134
rect 12966 13074 13018 13086
rect 18790 13074 18842 13086
rect 6850 13022 6862 13074
rect 6914 13022 6926 13074
rect 8082 13022 8094 13074
rect 8146 13022 8158 13074
rect 11330 13022 11342 13074
rect 11394 13022 11406 13074
rect 16258 13022 16270 13074
rect 16322 13022 16334 13074
rect 18162 13022 18174 13074
rect 18226 13022 18238 13074
rect 12966 13010 13018 13022
rect 18790 13010 18842 13022
rect 19462 13074 19514 13086
rect 31838 13074 31890 13086
rect 19462 13010 19514 13022
rect 21478 13018 21530 13030
rect 5182 12962 5234 12974
rect 6302 12962 6354 12974
rect 8430 12962 8482 12974
rect 5618 12910 5630 12962
rect 5682 12910 5694 12962
rect 5182 12898 5234 12910
rect 6066 12854 6078 12906
rect 6130 12854 6142 12906
rect 6302 12898 6354 12910
rect 6962 12866 6974 12918
rect 7026 12866 7038 12918
rect 7186 12910 7198 12962
rect 7250 12910 7262 12962
rect 7634 12910 7646 12962
rect 7698 12910 7710 12962
rect 7970 12895 7982 12947
rect 8034 12895 8046 12947
rect 8430 12898 8482 12910
rect 12126 12962 12178 12974
rect 14030 12962 14082 12974
rect 15486 12962 15538 12974
rect 13458 12910 13470 12962
rect 13522 12910 13534 12962
rect 14894 12910 14906 12962
rect 14958 12910 14970 12962
rect 12126 12898 12178 12910
rect 14030 12898 14082 12910
rect 15486 12898 15538 12910
rect 20190 12962 20242 12974
rect 20190 12898 20242 12910
rect 20302 12962 20354 12974
rect 20302 12898 20354 12910
rect 20638 12962 20690 12974
rect 20638 12898 20690 12910
rect 21310 12962 21362 12974
rect 30550 13018 30602 13030
rect 21478 12954 21530 12966
rect 21758 12962 21810 12974
rect 21310 12898 21362 12910
rect 21758 12898 21810 12910
rect 22766 12962 22818 12974
rect 23214 12962 23266 12974
rect 22866 12910 22878 12962
rect 22930 12910 22942 12962
rect 22766 12898 22818 12910
rect 9438 12850 9490 12862
rect 21646 12850 21698 12862
rect 4846 12738 4898 12750
rect 5730 12742 5742 12794
rect 5794 12742 5806 12794
rect 9438 12786 9490 12798
rect 13638 12794 13690 12806
rect 4846 12674 4898 12686
rect 8766 12738 8818 12750
rect 8766 12674 8818 12686
rect 12518 12738 12570 12750
rect 21646 12786 21698 12798
rect 22038 12850 22090 12862
rect 22038 12786 22090 12798
rect 22486 12850 22538 12862
rect 23034 12854 23046 12906
rect 23098 12854 23110 12906
rect 23214 12898 23266 12910
rect 23438 12962 23490 12974
rect 23438 12898 23490 12910
rect 24446 12962 24498 12974
rect 24894 12962 24946 12974
rect 24770 12910 24782 12962
rect 24834 12910 24846 12962
rect 24446 12898 24498 12910
rect 24602 12854 24614 12906
rect 24666 12854 24678 12906
rect 24894 12898 24946 12910
rect 25174 12962 25226 12974
rect 31838 13010 31890 13022
rect 34134 13074 34186 13086
rect 41694 13074 41746 13086
rect 37650 13022 37662 13074
rect 37714 13022 37726 13074
rect 38658 13022 38670 13074
rect 38722 13022 38734 13074
rect 42578 13022 42590 13074
rect 42642 13022 42654 13074
rect 48066 13022 48078 13074
rect 48130 13022 48142 13074
rect 34134 13010 34186 13022
rect 41694 13010 41746 13022
rect 26898 12910 26910 12962
rect 26962 12910 26974 12962
rect 29586 12910 29598 12962
rect 29650 12910 29662 12962
rect 30550 12954 30602 12966
rect 31670 12962 31722 12974
rect 32734 12962 32786 12974
rect 34974 12962 35026 12974
rect 25174 12898 25226 12910
rect 29990 12906 30042 12918
rect 30930 12910 30942 12962
rect 30994 12910 31006 12962
rect 29418 12854 29430 12906
rect 29482 12854 29494 12906
rect 22486 12786 22538 12798
rect 29822 12850 29874 12862
rect 31154 12882 31166 12934
rect 31218 12882 31230 12934
rect 32050 12910 32062 12962
rect 32114 12910 32126 12962
rect 32398 12924 32450 12936
rect 31670 12898 31722 12910
rect 33730 12910 33742 12962
rect 33794 12910 33806 12962
rect 32734 12898 32786 12910
rect 34974 12898 35026 12910
rect 35198 12962 35250 12974
rect 35198 12898 35250 12910
rect 36542 12962 36594 12974
rect 37886 12962 37938 12974
rect 37314 12910 37326 12962
rect 37378 12910 37390 12962
rect 36542 12898 36594 12910
rect 29990 12842 30042 12854
rect 30718 12850 30770 12862
rect 32398 12860 32450 12872
rect 37538 12866 37550 12918
rect 37602 12866 37614 12918
rect 37886 12898 37938 12910
rect 41022 12962 41074 12974
rect 44270 12962 44322 12974
rect 41122 12910 41134 12962
rect 41186 12910 41198 12962
rect 42130 12910 42142 12962
rect 42194 12910 42206 12962
rect 41022 12898 41074 12910
rect 29822 12786 29874 12798
rect 40574 12850 40626 12862
rect 41288 12854 41300 12906
rect 41352 12854 41364 12906
rect 42466 12866 42478 12918
rect 42530 12866 42542 12918
rect 43381 12910 43393 12962
rect 43445 12910 43457 12962
rect 44270 12898 44322 12910
rect 44718 12962 44770 12974
rect 44718 12898 44770 12910
rect 45390 12962 45442 12974
rect 46162 12910 46174 12962
rect 46226 12910 46238 12962
rect 45390 12898 45442 12910
rect 30718 12786 30770 12798
rect 33574 12794 33626 12806
rect 13638 12730 13690 12742
rect 23774 12738 23826 12750
rect 12518 12674 12570 12686
rect 23774 12674 23826 12686
rect 27638 12738 27690 12750
rect 40574 12786 40626 12798
rect 43150 12850 43202 12862
rect 43150 12786 43202 12798
rect 33574 12730 33626 12742
rect 35814 12738 35866 12750
rect 27638 12674 27690 12686
rect 35814 12674 35866 12686
rect 45054 12738 45106 12750
rect 45054 12674 45106 12686
rect 1344 12570 48608 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 48608 12570
rect 1344 12484 48608 12518
rect 15318 12402 15370 12414
rect 15318 12338 15370 12350
rect 16886 12402 16938 12414
rect 16886 12338 16938 12350
rect 18566 12402 18618 12414
rect 18566 12338 18618 12350
rect 23998 12402 24050 12414
rect 23998 12338 24050 12350
rect 26014 12402 26066 12414
rect 26014 12338 26066 12350
rect 32342 12402 32394 12414
rect 32342 12338 32394 12350
rect 33462 12402 33514 12414
rect 33462 12338 33514 12350
rect 35758 12402 35810 12414
rect 35758 12338 35810 12350
rect 36486 12402 36538 12414
rect 36486 12338 36538 12350
rect 43878 12402 43930 12414
rect 43878 12338 43930 12350
rect 6638 12290 6690 12302
rect 22094 12290 22146 12302
rect 6638 12226 6690 12238
rect 13918 12234 13970 12246
rect 9848 12216 9900 12228
rect 3950 12178 4002 12190
rect 8094 12178 8146 12190
rect 4722 12126 4734 12178
rect 4786 12126 4798 12178
rect 8642 12141 8654 12193
rect 8706 12141 8718 12193
rect 9550 12178 9602 12190
rect 8978 12126 8990 12178
rect 9042 12126 9054 12178
rect 9650 12126 9662 12178
rect 9714 12126 9726 12178
rect 9848 12152 9900 12164
rect 10782 12178 10834 12190
rect 13918 12170 13970 12182
rect 14030 12234 14082 12246
rect 14030 12170 14082 12182
rect 14758 12234 14810 12246
rect 19686 12234 19738 12246
rect 14758 12170 14810 12182
rect 15698 12126 15710 12178
rect 15762 12126 15774 12178
rect 16034 12126 16046 12178
rect 16098 12126 16110 12178
rect 17490 12126 17502 12178
rect 17554 12126 17566 12178
rect 17714 12126 17726 12178
rect 17778 12126 17790 12178
rect 19058 12154 19070 12206
rect 19122 12154 19134 12206
rect 22094 12226 22146 12238
rect 23214 12290 23266 12302
rect 19282 12126 19294 12178
rect 19346 12126 19358 12178
rect 19686 12170 19738 12182
rect 19854 12178 19906 12190
rect 3950 12114 4002 12126
rect 8094 12114 8146 12126
rect 9550 12114 9602 12126
rect 10782 12114 10834 12126
rect 19854 12114 19906 12126
rect 21982 12178 22034 12190
rect 22250 12182 22262 12234
rect 22314 12182 22326 12234
rect 23214 12226 23266 12238
rect 34862 12290 34914 12302
rect 21982 12114 22034 12126
rect 22430 12178 22482 12190
rect 22430 12114 22482 12126
rect 23102 12178 23154 12190
rect 23370 12182 23382 12234
rect 23434 12182 23446 12234
rect 34862 12226 34914 12238
rect 38558 12290 38610 12302
rect 48122 12238 48134 12290
rect 48186 12238 48198 12290
rect 23102 12114 23154 12126
rect 23550 12178 23602 12190
rect 23550 12114 23602 12126
rect 24334 12178 24386 12190
rect 24334 12114 24386 12126
rect 25678 12178 25730 12190
rect 25678 12114 25730 12126
rect 26350 12178 26402 12190
rect 26350 12114 26402 12126
rect 27694 12178 27746 12190
rect 30830 12178 30882 12190
rect 31108 12178 31160 12190
rect 28466 12126 28478 12178
rect 28530 12126 28542 12178
rect 30930 12126 30942 12178
rect 30994 12126 31006 12178
rect 32498 12126 32510 12178
rect 32562 12126 32574 12178
rect 33842 12141 33854 12193
rect 33906 12141 33918 12193
rect 34526 12178 34578 12190
rect 34178 12126 34190 12178
rect 34242 12126 34254 12178
rect 34974 12178 35026 12190
rect 27694 12114 27746 12126
rect 30830 12114 30882 12126
rect 31108 12114 31160 12126
rect 34526 12114 34578 12126
rect 34694 12122 34746 12134
rect 7254 12066 7306 12078
rect 10222 12066 10274 12078
rect 14590 12066 14642 12078
rect 8530 12014 8542 12066
rect 8594 12014 8606 12066
rect 11554 12014 11566 12066
rect 11618 12014 11630 12066
rect 13458 12014 13470 12066
rect 13522 12014 13534 12066
rect 19518 12066 19570 12078
rect 7254 12002 7306 12014
rect 10222 12002 10274 12014
rect 14590 12002 14642 12014
rect 15598 12010 15650 12022
rect 7758 11954 7810 11966
rect 15598 11946 15650 11958
rect 17390 12010 17442 12022
rect 19518 12002 19570 12014
rect 20806 12066 20858 12078
rect 20806 12002 20858 12014
rect 21254 12066 21306 12078
rect 21254 12002 21306 12014
rect 27302 12066 27354 12078
rect 31502 12066 31554 12078
rect 34974 12114 35026 12126
rect 36094 12178 36146 12190
rect 36094 12114 36146 12126
rect 36990 12178 37042 12190
rect 37146 12182 37158 12234
rect 37210 12182 37222 12234
rect 38558 12226 38610 12238
rect 37438 12178 37490 12190
rect 37314 12126 37326 12178
rect 37378 12126 37390 12178
rect 36990 12114 37042 12126
rect 37438 12114 37490 12126
rect 37718 12178 37770 12190
rect 37718 12114 37770 12126
rect 38446 12178 38498 12190
rect 38894 12178 38946 12190
rect 40238 12178 40290 12190
rect 38446 12114 38498 12126
rect 38726 12122 38778 12134
rect 30370 12014 30382 12066
rect 30434 12014 30446 12066
rect 33730 12014 33742 12066
rect 33794 12014 33806 12066
rect 34694 12058 34746 12070
rect 39946 12126 39958 12178
rect 40010 12126 40022 12178
rect 38894 12114 38946 12126
rect 40238 12114 40290 12126
rect 40350 12178 40402 12190
rect 41010 12126 41022 12178
rect 41074 12126 41086 12178
rect 41234 12170 41246 12222
rect 41298 12170 41310 12222
rect 42888 12216 42940 12228
rect 41794 12141 41806 12193
rect 41858 12141 41870 12193
rect 42590 12178 42642 12190
rect 42018 12126 42030 12178
rect 42082 12126 42094 12178
rect 42690 12126 42702 12178
rect 42754 12126 42766 12178
rect 42888 12152 42940 12164
rect 44942 12178 44994 12190
rect 40350 12114 40402 12126
rect 42590 12114 42642 12126
rect 44942 12114 44994 12126
rect 45166 12178 45218 12190
rect 45378 12182 45390 12234
rect 45442 12182 45454 12234
rect 45826 12182 45838 12234
rect 45890 12182 45902 12234
rect 46162 12182 46174 12234
rect 46226 12182 46238 12234
rect 46472 12166 46484 12218
rect 46536 12166 46548 12218
rect 47630 12178 47682 12190
rect 47058 12126 47070 12178
rect 47122 12126 47134 12178
rect 47282 12126 47294 12178
rect 47346 12126 47358 12178
rect 45166 12114 45218 12126
rect 47630 12114 47682 12126
rect 47854 12178 47906 12190
rect 47854 12114 47906 12126
rect 38726 12058 38778 12070
rect 39398 12066 39450 12078
rect 43262 12066 43314 12078
rect 41346 12014 41358 12066
rect 41410 12014 41422 12066
rect 41682 12014 41694 12066
rect 41746 12014 41758 12066
rect 27302 12002 27354 12014
rect 31502 12002 31554 12014
rect 39398 12002 39450 12014
rect 43262 12002 43314 12014
rect 44326 12066 44378 12078
rect 46498 12014 46510 12066
rect 46562 12014 46574 12066
rect 44326 12002 44378 12014
rect 46958 12010 47010 12022
rect 17390 11946 17442 11958
rect 20190 11954 20242 11966
rect 7758 11890 7810 11902
rect 20190 11890 20242 11902
rect 21702 11954 21754 11966
rect 21702 11890 21754 11902
rect 22822 11954 22874 11966
rect 22822 11890 22874 11902
rect 26686 11954 26738 11966
rect 26686 11890 26738 11902
rect 35254 11954 35306 11966
rect 35254 11890 35306 11902
rect 38166 11954 38218 11966
rect 44650 11902 44662 11954
rect 44714 11902 44726 11954
rect 46958 11946 47010 11958
rect 38166 11890 38218 11902
rect 1344 11786 48608 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 48608 11786
rect 1344 11700 48608 11734
rect 22598 11618 22650 11630
rect 15978 11566 15990 11618
rect 16042 11566 16054 11618
rect 20694 11562 20746 11574
rect 5126 11506 5178 11518
rect 9718 11506 9770 11518
rect 6066 11454 6078 11506
rect 6130 11454 6142 11506
rect 6850 11454 6862 11506
rect 6914 11454 6926 11506
rect 5126 11442 5178 11454
rect 9718 11442 9770 11454
rect 13750 11506 13802 11518
rect 22598 11554 22650 11566
rect 26126 11618 26178 11630
rect 26126 11554 26178 11566
rect 30438 11618 30490 11630
rect 17154 11454 17166 11506
rect 17218 11454 17230 11506
rect 19506 11454 19518 11506
rect 19570 11454 19582 11506
rect 20694 11498 20746 11510
rect 23158 11506 23210 11518
rect 13750 11442 13802 11454
rect 22150 11450 22202 11462
rect 1822 11394 1874 11406
rect 4510 11394 4562 11406
rect 7534 11394 7586 11406
rect 2594 11342 2606 11394
rect 2658 11342 2670 11394
rect 5618 11342 5630 11394
rect 5682 11342 5694 11394
rect 1822 11330 1874 11342
rect 4510 11330 4562 11342
rect 5954 11298 5966 11350
rect 6018 11298 6030 11350
rect 6402 11342 6414 11394
rect 6466 11342 6478 11394
rect 6738 11327 6750 11379
rect 6802 11327 6814 11379
rect 7534 11330 7586 11342
rect 7870 11394 7922 11406
rect 7870 11330 7922 11342
rect 8542 11394 8594 11406
rect 10110 11394 10162 11406
rect 16270 11394 16322 11406
rect 9090 11342 9102 11394
rect 9154 11342 9166 11394
rect 10882 11342 10894 11394
rect 10946 11342 10958 11394
rect 8542 11330 8594 11342
rect 8922 11286 8934 11338
rect 8986 11286 8998 11338
rect 10110 11330 10162 11342
rect 14018 11309 14030 11361
rect 14082 11309 14094 11361
rect 12798 11282 12850 11294
rect 14354 11286 14366 11338
rect 14418 11286 14430 11338
rect 14802 11309 14814 11361
rect 14866 11309 14878 11361
rect 15112 11309 15124 11361
rect 15176 11309 15188 11361
rect 16270 11330 16322 11342
rect 16382 11394 16434 11406
rect 20302 11394 20354 11406
rect 21298 11398 21310 11450
rect 21362 11398 21374 11450
rect 25622 11506 25674 11518
rect 26898 11510 26910 11562
rect 26962 11510 26974 11562
rect 30438 11554 30490 11566
rect 35478 11618 35530 11630
rect 47182 11618 47234 11630
rect 35478 11554 35530 11566
rect 42926 11562 42978 11574
rect 34022 11506 34074 11518
rect 23158 11442 23210 11454
rect 24502 11450 24554 11462
rect 16706 11342 16718 11394
rect 16770 11342 16782 11394
rect 16382 11330 16434 11342
rect 17042 11327 17054 11379
rect 17106 11327 17118 11379
rect 20514 11342 20526 11394
rect 20578 11342 20590 11394
rect 22150 11386 22202 11398
rect 24054 11394 24106 11406
rect 21422 11356 21474 11368
rect 20302 11330 20354 11342
rect 22418 11342 22430 11394
rect 22482 11342 22494 11394
rect 24054 11330 24106 11342
rect 24334 11394 24386 11406
rect 31490 11454 31502 11506
rect 31554 11454 31566 11506
rect 33394 11454 33406 11506
rect 33458 11454 33470 11506
rect 40070 11506 40122 11518
rect 25622 11442 25674 11454
rect 34022 11442 34074 11454
rect 35142 11450 35194 11462
rect 24502 11386 24554 11398
rect 24782 11394 24834 11406
rect 24334 11330 24386 11342
rect 24782 11330 24834 11342
rect 26462 11394 26514 11406
rect 30718 11394 30770 11406
rect 34290 11398 34302 11450
rect 34354 11398 34366 11450
rect 26674 11342 26686 11394
rect 26738 11342 26750 11394
rect 27010 11342 27022 11394
rect 27074 11342 27086 11394
rect 30606 11373 30658 11385
rect 26462 11330 26514 11342
rect 30718 11330 30770 11342
rect 34974 11394 35026 11406
rect 36038 11450 36090 11462
rect 35142 11386 35194 11398
rect 35758 11394 35810 11406
rect 30606 11309 30658 11321
rect 8530 11174 8542 11226
rect 8594 11174 8606 11226
rect 12798 11218 12850 11230
rect 15262 11282 15314 11294
rect 15262 11218 15314 11230
rect 17614 11282 17666 11294
rect 21422 11292 21474 11304
rect 17614 11218 17666 11230
rect 21982 11282 22034 11294
rect 21982 11218 22034 11230
rect 24670 11282 24722 11294
rect 24670 11218 24722 11230
rect 25062 11282 25114 11294
rect 25062 11218 25114 11230
rect 30102 11282 30154 11294
rect 34514 11286 34526 11338
rect 34578 11286 34590 11338
rect 34974 11330 35026 11342
rect 47182 11554 47234 11566
rect 42926 11498 42978 11510
rect 47966 11506 48018 11518
rect 40070 11442 40122 11454
rect 41190 11450 41242 11462
rect 36038 11386 36090 11398
rect 36206 11394 36258 11406
rect 35758 11330 35810 11342
rect 36206 11330 36258 11342
rect 37438 11394 37490 11406
rect 37438 11330 37490 11342
rect 37550 11394 37602 11406
rect 37550 11330 37602 11342
rect 38222 11394 38274 11406
rect 38222 11330 38274 11342
rect 38894 11394 38946 11406
rect 43206 11450 43258 11462
rect 46498 11454 46510 11506
rect 46562 11454 46574 11506
rect 40786 11342 40798 11394
rect 40850 11342 40862 11394
rect 41190 11386 41242 11398
rect 41694 11394 41746 11406
rect 38894 11330 38946 11342
rect 30102 11218 30154 11230
rect 35870 11282 35922 11294
rect 40562 11286 40574 11338
rect 40626 11286 40638 11338
rect 41694 11330 41746 11342
rect 41806 11394 41858 11406
rect 47966 11442 48018 11454
rect 42578 11342 42590 11394
rect 42642 11342 42654 11394
rect 42802 11342 42814 11394
rect 42866 11342 42878 11394
rect 43206 11386 43258 11398
rect 46846 11394 46898 11406
rect 43586 11342 43598 11394
rect 43650 11342 43662 11394
rect 41806 11330 41858 11342
rect 43810 11314 43822 11366
rect 43874 11314 43886 11366
rect 45378 11309 45390 11361
rect 45442 11309 45454 11361
rect 45826 11305 45838 11357
rect 45890 11305 45902 11357
rect 46162 11309 46174 11361
rect 46226 11309 46238 11361
rect 46472 11302 46484 11354
rect 46536 11302 46548 11354
rect 46846 11330 46898 11342
rect 48302 11394 48354 11406
rect 48302 11330 48354 11342
rect 35870 11218 35922 11230
rect 41022 11282 41074 11294
rect 43374 11282 43426 11294
rect 42074 11230 42086 11282
rect 42138 11230 42150 11282
rect 41022 11218 41074 11230
rect 43374 11218 43426 11230
rect 27638 11170 27690 11182
rect 27638 11106 27690 11118
rect 28646 11170 28698 11182
rect 28646 11106 28698 11118
rect 29654 11170 29706 11182
rect 29654 11106 29706 11118
rect 37102 11170 37154 11182
rect 37102 11106 37154 11118
rect 37886 11170 37938 11182
rect 37886 11106 37938 11118
rect 38558 11170 38610 11182
rect 38558 11106 38610 11118
rect 39230 11170 39282 11182
rect 39230 11106 39282 11118
rect 44998 11170 45050 11182
rect 44998 11106 45050 11118
rect 1344 11002 48608 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 48608 11002
rect 1344 10916 48608 10950
rect 2942 10834 2994 10846
rect 2942 10770 2994 10782
rect 10838 10834 10890 10846
rect 5058 10726 5070 10778
rect 5122 10726 5134 10778
rect 9650 10726 9662 10778
rect 9714 10726 9726 10778
rect 10838 10770 10890 10782
rect 11286 10834 11338 10846
rect 11286 10770 11338 10782
rect 11734 10834 11786 10846
rect 11734 10770 11786 10782
rect 12182 10834 12234 10846
rect 12182 10770 12234 10782
rect 12630 10834 12682 10846
rect 12630 10770 12682 10782
rect 15766 10834 15818 10846
rect 15766 10770 15818 10782
rect 17558 10834 17610 10846
rect 17558 10770 17610 10782
rect 19014 10834 19066 10846
rect 19014 10770 19066 10782
rect 23102 10834 23154 10846
rect 23102 10770 23154 10782
rect 25454 10834 25506 10846
rect 25454 10770 25506 10782
rect 26070 10834 26122 10846
rect 36990 10834 37042 10846
rect 26070 10770 26122 10782
rect 32342 10778 32394 10790
rect 26686 10722 26738 10734
rect 15194 10670 15206 10722
rect 15258 10670 15270 10722
rect 16886 10666 16938 10678
rect 17882 10670 17894 10722
rect 17946 10670 17958 10722
rect 36990 10770 37042 10782
rect 39006 10834 39058 10846
rect 39006 10770 39058 10782
rect 39622 10834 39674 10846
rect 39622 10770 39674 10782
rect 32342 10714 32394 10726
rect 35646 10722 35698 10734
rect 2606 10610 2658 10622
rect 2606 10546 2658 10558
rect 3278 10610 3330 10622
rect 4162 10558 4174 10610
rect 4226 10558 4238 10610
rect 4386 10602 4398 10654
rect 4450 10602 4462 10654
rect 9942 10639 9994 10651
rect 4834 10558 4846 10610
rect 4898 10558 4910 10610
rect 5170 10585 5182 10637
rect 5234 10585 5246 10637
rect 5518 10610 5570 10622
rect 3278 10546 3330 10558
rect 5518 10546 5570 10558
rect 6190 10610 6242 10622
rect 6190 10546 6242 10558
rect 8878 10610 8930 10622
rect 9538 10558 9550 10610
rect 9602 10558 9614 10610
rect 13694 10610 13746 10622
rect 9942 10575 9994 10587
rect 13010 10558 13022 10610
rect 13074 10558 13086 10610
rect 13234 10558 13246 10610
rect 13298 10558 13310 10610
rect 13794 10558 13806 10610
rect 13858 10558 13870 10610
rect 13952 10608 13964 10660
rect 14016 10608 14028 10660
rect 16158 10648 16210 10660
rect 14702 10610 14754 10622
rect 8878 10546 8930 10558
rect 13694 10546 13746 10558
rect 14702 10546 14754 10558
rect 14926 10610 14978 10622
rect 16158 10584 16210 10596
rect 16482 10558 16494 10610
rect 16546 10558 16558 10610
rect 16886 10602 16938 10614
rect 18174 10610 18226 10622
rect 14926 10546 14978 10558
rect 18174 10546 18226 10558
rect 18286 10610 18338 10622
rect 22542 10610 22594 10622
rect 18834 10558 18846 10610
rect 18898 10558 18910 10610
rect 21746 10558 21758 10610
rect 21810 10558 21822 10610
rect 18286 10546 18338 10558
rect 22542 10546 22594 10558
rect 23438 10610 23490 10622
rect 23438 10546 23490 10558
rect 24782 10610 24834 10622
rect 24782 10546 24834 10558
rect 25118 10610 25170 10622
rect 25118 10546 25170 10558
rect 26350 10610 26402 10622
rect 26506 10614 26518 10666
rect 26570 10614 26582 10666
rect 26686 10658 26738 10670
rect 31652 10648 31704 10660
rect 35646 10658 35698 10670
rect 43486 10722 43538 10734
rect 43486 10658 43538 10670
rect 44046 10722 44098 10734
rect 44046 10658 44098 10670
rect 26350 10546 26402 10558
rect 26798 10610 26850 10622
rect 26798 10546 26850 10558
rect 27638 10610 27690 10622
rect 27638 10546 27690 10558
rect 28030 10610 28082 10622
rect 31950 10610 32002 10622
rect 32958 10610 33010 10622
rect 35982 10610 36034 10622
rect 31652 10584 31704 10596
rect 31826 10558 31838 10610
rect 31890 10558 31902 10610
rect 32498 10558 32510 10610
rect 32562 10558 32574 10610
rect 33730 10558 33742 10610
rect 33794 10558 33806 10610
rect 28030 10546 28082 10558
rect 31950 10546 32002 10558
rect 32958 10546 33010 10558
rect 35982 10546 36034 10558
rect 36654 10610 36706 10622
rect 36654 10546 36706 10558
rect 37326 10610 37378 10622
rect 37326 10546 37378 10558
rect 37998 10610 38050 10622
rect 37998 10546 38050 10558
rect 38670 10610 38722 10622
rect 38670 10546 38722 10558
rect 40238 10610 40290 10622
rect 40238 10546 40290 10558
rect 40350 10610 40402 10622
rect 40350 10546 40402 10558
rect 40798 10610 40850 10622
rect 46734 10610 46786 10622
rect 47742 10610 47794 10622
rect 41570 10558 41582 10610
rect 41634 10558 41646 10610
rect 45938 10558 45950 10610
rect 46002 10558 46014 10610
rect 47058 10558 47070 10610
rect 47122 10558 47134 10610
rect 47282 10558 47294 10610
rect 47346 10558 47358 10610
rect 40798 10546 40850 10558
rect 46734 10546 46786 10558
rect 47742 10546 47794 10558
rect 47854 10610 47906 10622
rect 48122 10558 48134 10610
rect 48186 10558 48198 10610
rect 47854 10546 47906 10558
rect 14366 10498 14418 10510
rect 4498 10446 4510 10498
rect 4562 10446 4574 10498
rect 6962 10446 6974 10498
rect 7026 10446 7038 10498
rect 13358 10442 13410 10454
rect 2270 10386 2322 10398
rect 14366 10434 14418 10446
rect 16718 10498 16770 10510
rect 19842 10446 19854 10498
rect 19906 10446 19918 10498
rect 28802 10446 28814 10498
rect 28866 10446 28878 10498
rect 30706 10446 30718 10498
rect 30770 10446 30782 10498
rect 16718 10434 16770 10446
rect 46958 10442 47010 10454
rect 13358 10378 13410 10390
rect 24446 10386 24498 10398
rect 2270 10322 2322 10334
rect 24446 10322 24498 10334
rect 27078 10386 27130 10398
rect 27078 10322 27130 10334
rect 31278 10386 31330 10398
rect 31278 10322 31330 10334
rect 36318 10386 36370 10398
rect 36318 10322 36370 10334
rect 37662 10386 37714 10398
rect 37662 10322 37714 10334
rect 38334 10386 38386 10398
rect 39946 10334 39958 10386
rect 40010 10334 40022 10386
rect 46958 10378 47010 10390
rect 38334 10322 38386 10334
rect 1344 10218 48608 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 48608 10218
rect 1344 10132 48608 10166
rect 8206 10050 8258 10062
rect 14366 10050 14418 10062
rect 43374 10050 43426 10062
rect 13514 9998 13526 10050
rect 13578 9998 13590 10050
rect 8206 9986 8258 9998
rect 14366 9986 14418 9998
rect 38558 9994 38610 10006
rect 39722 9998 39734 10050
rect 39786 9998 39798 10050
rect 10502 9938 10554 9950
rect 2370 9886 2382 9938
rect 2434 9886 2446 9938
rect 7298 9886 7310 9938
rect 7362 9886 7374 9938
rect 8866 9886 8878 9938
rect 8930 9886 8942 9938
rect 10502 9874 10554 9886
rect 11398 9938 11450 9950
rect 27918 9938 27970 9950
rect 16370 9886 16382 9938
rect 16434 9886 16446 9938
rect 11398 9874 11450 9886
rect 19574 9882 19626 9894
rect 1598 9826 1650 9838
rect 1598 9762 1650 9774
rect 4286 9826 4338 9838
rect 4286 9762 4338 9774
rect 5182 9826 5234 9838
rect 6302 9826 6354 9838
rect 8542 9826 8594 9838
rect 10110 9826 10162 9838
rect 5618 9774 5630 9826
rect 5682 9774 5694 9826
rect 6850 9774 6862 9826
rect 6914 9774 6926 9826
rect 5182 9762 5234 9774
rect 5954 9718 5966 9770
rect 6018 9718 6030 9770
rect 6302 9762 6354 9774
rect 7186 9730 7198 9782
rect 7250 9730 7262 9782
rect 8542 9762 8594 9774
rect 8978 9730 8990 9782
rect 9042 9730 9054 9782
rect 9202 9774 9214 9826
rect 9266 9774 9278 9826
rect 13806 9826 13858 9838
rect 10110 9762 10162 9774
rect 11678 9714 11730 9726
rect 11834 9718 11846 9770
rect 11898 9718 11910 9770
rect 12114 9741 12126 9793
rect 12178 9741 12190 9793
rect 12562 9718 12574 9770
rect 12626 9718 12638 9770
rect 12898 9718 12910 9770
rect 12962 9718 12974 9770
rect 13806 9762 13858 9774
rect 14030 9826 14082 9838
rect 15038 9826 15090 9838
rect 14914 9774 14926 9826
rect 14978 9774 14990 9826
rect 14030 9762 14082 9774
rect 14746 9718 14758 9770
rect 14810 9718 14822 9770
rect 15038 9762 15090 9774
rect 15598 9826 15650 9838
rect 19574 9818 19626 9830
rect 20806 9882 20858 9894
rect 22710 9882 22762 9894
rect 18846 9788 18898 9800
rect 15598 9762 15650 9774
rect 18734 9770 18786 9782
rect 4846 9602 4898 9614
rect 5730 9606 5742 9658
rect 5794 9606 5806 9658
rect 11678 9650 11730 9662
rect 18286 9714 18338 9726
rect 18846 9724 18898 9736
rect 20078 9788 20130 9800
rect 20402 9774 20414 9826
rect 20466 9774 20478 9826
rect 20806 9818 20858 9830
rect 22430 9826 22482 9838
rect 23382 9882 23434 9894
rect 22530 9774 22542 9826
rect 22594 9774 22606 9826
rect 22710 9818 22762 9830
rect 22878 9826 22930 9838
rect 22430 9762 22482 9774
rect 22878 9762 22930 9774
rect 23214 9826 23266 9838
rect 27918 9874 27970 9886
rect 29822 9938 29874 9950
rect 30550 9938 30602 9950
rect 23382 9818 23434 9830
rect 23662 9826 23714 9838
rect 23214 9762 23266 9774
rect 23662 9762 23714 9774
rect 24222 9826 24274 9838
rect 24222 9762 24274 9774
rect 25454 9826 25506 9838
rect 25454 9762 25506 9774
rect 27246 9826 27298 9838
rect 29138 9830 29150 9882
rect 29202 9830 29214 9882
rect 29822 9874 29874 9886
rect 29990 9882 30042 9894
rect 30550 9874 30602 9886
rect 32790 9938 32842 9950
rect 32790 9874 32842 9886
rect 33238 9938 33290 9950
rect 33238 9874 33290 9886
rect 34134 9938 34186 9950
rect 34134 9874 34186 9886
rect 35086 9938 35138 9950
rect 37606 9938 37658 9950
rect 36082 9886 36094 9938
rect 36146 9886 36158 9938
rect 35086 9874 35138 9886
rect 37606 9874 37658 9886
rect 38110 9938 38162 9950
rect 38558 9930 38610 9942
rect 40910 9994 40962 10006
rect 41906 9942 41918 9994
rect 41970 9942 41982 9994
rect 43374 9986 43426 9998
rect 45054 10050 45106 10062
rect 45054 9986 45106 9998
rect 40910 9930 40962 9942
rect 42646 9938 42698 9950
rect 38110 9874 38162 9886
rect 42646 9874 42698 9886
rect 44102 9938 44154 9950
rect 46162 9886 46174 9938
rect 46226 9886 46238 9938
rect 48066 9886 48078 9938
rect 48130 9886 48142 9938
rect 44102 9874 44154 9886
rect 27346 9774 27358 9826
rect 27410 9774 27422 9826
rect 29990 9818 30042 9830
rect 31838 9826 31890 9838
rect 27246 9762 27298 9774
rect 30942 9770 30994 9782
rect 31266 9774 31278 9826
rect 31330 9774 31342 9826
rect 18734 9706 18786 9718
rect 19406 9714 19458 9726
rect 20078 9724 20130 9736
rect 18286 9650 18338 9662
rect 19406 9650 19458 9662
rect 20638 9714 20690 9726
rect 20638 9650 20690 9662
rect 22150 9714 22202 9726
rect 22150 9650 22202 9662
rect 23550 9714 23602 9726
rect 23550 9650 23602 9662
rect 23942 9714 23994 9726
rect 27512 9718 27524 9770
rect 27576 9718 27588 9770
rect 29418 9718 29430 9770
rect 29482 9718 29494 9770
rect 31670 9770 31722 9782
rect 30942 9706 30994 9718
rect 31502 9714 31554 9726
rect 23942 9650 23994 9662
rect 31838 9762 31890 9774
rect 34414 9826 34466 9838
rect 34694 9826 34746 9838
rect 37774 9826 37826 9838
rect 39230 9826 39282 9838
rect 34514 9774 34526 9826
rect 34578 9774 34590 9826
rect 35634 9774 35646 9826
rect 35698 9774 35710 9826
rect 34414 9762 34466 9774
rect 34694 9762 34746 9774
rect 35970 9759 35982 9811
rect 36034 9759 36046 9811
rect 38658 9774 38670 9826
rect 38722 9774 38734 9826
rect 38994 9774 39006 9826
rect 39058 9774 39070 9826
rect 37774 9762 37826 9774
rect 39230 9762 39282 9774
rect 39454 9826 39506 9838
rect 39454 9762 39506 9774
rect 40686 9826 40738 9838
rect 43710 9826 43762 9838
rect 41010 9774 41022 9826
rect 41074 9774 41086 9826
rect 41346 9774 41358 9826
rect 41410 9774 41422 9826
rect 41682 9774 41694 9826
rect 41746 9774 41758 9826
rect 42018 9774 42030 9826
rect 42082 9774 42094 9826
rect 40686 9762 40738 9774
rect 43710 9762 43762 9774
rect 44718 9826 44770 9838
rect 44718 9762 44770 9774
rect 45390 9826 45442 9838
rect 45390 9762 45442 9774
rect 31670 9706 31722 9718
rect 31502 9650 31554 9662
rect 4846 9538 4898 9550
rect 9774 9602 9826 9614
rect 9774 9538 9826 9550
rect 21478 9602 21530 9614
rect 21478 9538 21530 9550
rect 24558 9602 24610 9614
rect 24558 9538 24610 9550
rect 25790 9602 25842 9614
rect 25790 9538 25842 9550
rect 26518 9602 26570 9614
rect 26518 9538 26570 9550
rect 26966 9602 27018 9614
rect 26966 9538 27018 9550
rect 28646 9602 28698 9614
rect 28646 9538 28698 9550
rect 32174 9602 32226 9614
rect 32174 9538 32226 9550
rect 33686 9602 33738 9614
rect 33686 9538 33738 9550
rect 37158 9602 37210 9614
rect 37158 9538 37210 9550
rect 40350 9602 40402 9614
rect 40350 9538 40402 9550
rect 1344 9434 48608 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 48608 9434
rect 1344 9348 48608 9382
rect 10502 9266 10554 9278
rect 5730 9158 5742 9210
rect 5794 9158 5806 9210
rect 8866 9158 8878 9210
rect 8930 9158 8942 9210
rect 10502 9202 10554 9214
rect 15038 9266 15090 9278
rect 15038 9202 15090 9214
rect 15598 9266 15650 9278
rect 15598 9202 15650 9214
rect 17670 9266 17722 9278
rect 17670 9202 17722 9214
rect 18118 9266 18170 9278
rect 18118 9202 18170 9214
rect 18678 9266 18730 9278
rect 18678 9202 18730 9214
rect 22990 9266 23042 9278
rect 22990 9202 23042 9214
rect 33686 9266 33738 9278
rect 33686 9202 33738 9214
rect 34134 9266 34186 9278
rect 34134 9202 34186 9214
rect 44550 9266 44602 9278
rect 44550 9202 44602 9214
rect 47126 9266 47178 9278
rect 47126 9202 47178 9214
rect 47574 9266 47626 9278
rect 47574 9202 47626 9214
rect 48246 9266 48298 9278
rect 48246 9202 48298 9214
rect 13358 9154 13410 9166
rect 1598 9042 1650 9054
rect 1598 8978 1650 8990
rect 4286 9042 4338 9054
rect 5450 9046 5462 9098
rect 5514 9046 5526 9098
rect 13358 9090 13410 9102
rect 16774 9154 16826 9166
rect 16774 9090 16826 9102
rect 24334 9154 24386 9166
rect 24334 9090 24386 9102
rect 36486 9154 36538 9166
rect 5854 9042 5906 9054
rect 5282 8990 5294 9042
rect 5346 8990 5358 9042
rect 6402 8990 6414 9042
rect 6466 8990 6478 9042
rect 6738 9034 6750 9086
rect 6802 9034 6814 9086
rect 7410 9005 7422 9057
rect 7474 9005 7486 9057
rect 7746 8990 7758 9042
rect 7810 8990 7822 9042
rect 8194 8990 8206 9042
rect 8258 8990 8270 9042
rect 8418 9017 8430 9069
rect 8482 9017 8494 9069
rect 8766 9042 8818 9054
rect 4286 8978 4338 8990
rect 5854 8978 5906 8990
rect 8766 8978 8818 8990
rect 9438 9042 9490 9054
rect 9438 8978 9490 8990
rect 10670 9042 10722 9054
rect 14702 9042 14754 9054
rect 11442 8990 11454 9042
rect 11506 8990 11518 9042
rect 13906 8990 13918 9042
rect 13970 8990 13982 9042
rect 14242 8990 14254 9042
rect 14306 8990 14318 9042
rect 10670 8978 10722 8990
rect 14702 8978 14754 8990
rect 15934 9042 15986 9054
rect 21982 9042 22034 9054
rect 18498 8990 18510 9042
rect 18562 8990 18574 9042
rect 21186 8990 21198 9042
rect 21250 8990 21262 9042
rect 15934 8978 15986 8990
rect 21982 8978 22034 8990
rect 22374 9042 22426 9054
rect 22374 8978 22426 8990
rect 22654 9042 22706 9054
rect 22654 8978 22706 8990
rect 24222 9042 24274 9054
rect 24490 9046 24502 9098
rect 24554 9046 24566 9098
rect 36486 9090 36538 9102
rect 39342 9154 39394 9166
rect 41134 9154 41186 9166
rect 40282 9102 40294 9154
rect 40346 9102 40358 9154
rect 39342 9090 39394 9102
rect 41134 9090 41186 9102
rect 24222 8978 24274 8990
rect 24670 9042 24722 9054
rect 26462 9042 26514 9054
rect 25778 8990 25790 9042
rect 25842 8990 25854 9042
rect 26002 8990 26014 9042
rect 26066 8990 26078 9042
rect 24670 8978 24722 8990
rect 26462 8978 26514 8990
rect 26630 9042 26682 9054
rect 26910 9042 26962 9054
rect 26786 8990 26798 9042
rect 26850 8990 26862 9042
rect 26630 8978 26682 8990
rect 26910 8978 26962 8990
rect 27806 9042 27858 9054
rect 27806 8978 27858 8990
rect 30830 9042 30882 9054
rect 30830 8978 30882 8990
rect 32232 9042 32284 9054
rect 32510 9042 32562 9054
rect 32386 8990 32398 9042
rect 32450 8990 32462 9042
rect 33282 8990 33294 9042
rect 33346 8990 33358 9042
rect 34626 8990 34638 9042
rect 34690 8990 34702 9042
rect 34962 9034 34974 9086
rect 35026 9034 35038 9086
rect 35310 9042 35362 9054
rect 32232 8978 32284 8990
rect 32510 8978 32562 8990
rect 35310 8978 35362 8990
rect 35534 9042 35586 9054
rect 35534 8978 35586 8990
rect 36654 9042 36706 9054
rect 36654 8978 36706 8990
rect 39902 9042 39954 9054
rect 39902 8978 39954 8990
rect 40014 9042 40066 9054
rect 40014 8978 40066 8990
rect 43822 9042 43874 9054
rect 43822 8978 43874 8990
rect 45278 9042 45330 9054
rect 45278 8978 45330 8990
rect 45614 9042 45666 9054
rect 46274 8990 46286 9042
rect 46338 8990 46350 9042
rect 46610 8990 46622 9042
rect 46674 8990 46686 9042
rect 45614 8978 45666 8990
rect 4902 8930 4954 8942
rect 16326 8930 16378 8942
rect 25398 8930 25450 8942
rect 31838 8930 31890 8942
rect 45110 8930 45162 8942
rect 2370 8878 2382 8930
rect 2434 8878 2446 8930
rect 6850 8878 6862 8930
rect 6914 8878 6926 8930
rect 7298 8878 7310 8930
rect 7362 8878 7374 8930
rect 4902 8866 4954 8878
rect 13806 8874 13858 8886
rect 9774 8818 9826 8830
rect 19282 8878 19294 8930
rect 19346 8878 19358 8930
rect 16326 8866 16378 8878
rect 25398 8866 25450 8878
rect 25678 8874 25730 8886
rect 28578 8878 28590 8930
rect 28642 8878 28654 8930
rect 30482 8878 30494 8930
rect 30546 8878 30558 8930
rect 13806 8810 13858 8822
rect 23942 8818 23994 8830
rect 9774 8754 9826 8766
rect 31838 8866 31890 8878
rect 33126 8874 33178 8886
rect 35074 8878 35086 8930
rect 35138 8878 35150 8930
rect 37426 8878 37438 8930
rect 37490 8878 37502 8930
rect 43026 8878 43038 8930
rect 43090 8878 43102 8930
rect 25678 8810 25730 8822
rect 27190 8818 27242 8830
rect 23942 8754 23994 8766
rect 27190 8754 27242 8766
rect 31166 8818 31218 8830
rect 45110 8866 45162 8878
rect 46174 8874 46226 8886
rect 33126 8810 33178 8822
rect 35802 8766 35814 8818
rect 35866 8766 35878 8818
rect 46174 8810 46226 8822
rect 31166 8754 31218 8766
rect 1344 8650 48608 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 48608 8650
rect 1344 8564 48608 8598
rect 2718 8482 2770 8494
rect 20470 8482 20522 8494
rect 2718 8418 2770 8430
rect 13470 8426 13522 8438
rect 3558 8370 3610 8382
rect 12182 8370 12234 8382
rect 4274 8318 4286 8370
rect 4338 8318 4350 8370
rect 5058 8318 5070 8370
rect 5122 8318 5134 8370
rect 6850 8318 6862 8370
rect 6914 8318 6926 8370
rect 8642 8318 8654 8370
rect 8706 8318 8718 8370
rect 10994 8318 11006 8370
rect 11058 8318 11070 8370
rect 27570 8430 27582 8482
rect 27634 8479 27646 8482
rect 27794 8479 27806 8482
rect 27634 8433 27806 8479
rect 27634 8430 27646 8433
rect 27794 8430 27806 8433
rect 27858 8430 27870 8482
rect 20470 8418 20522 8430
rect 13470 8362 13522 8374
rect 15542 8370 15594 8382
rect 28478 8370 28530 8382
rect 14914 8318 14926 8370
rect 14978 8318 14990 8370
rect 18050 8318 18062 8370
rect 18114 8318 18126 8370
rect 3558 8306 3610 8318
rect 12182 8306 12234 8318
rect 15542 8306 15594 8318
rect 21254 8314 21306 8326
rect 3054 8258 3106 8270
rect 6302 8258 6354 8270
rect 9102 8258 9154 8270
rect 3826 8206 3838 8258
rect 3890 8206 3902 8258
rect 4610 8206 4622 8258
rect 4674 8206 4686 8258
rect 3054 8194 3106 8206
rect 4106 8150 4118 8202
rect 4170 8150 4182 8202
rect 4946 8191 4958 8243
rect 5010 8191 5022 8243
rect 5618 8206 5630 8258
rect 5682 8206 5694 8258
rect 6078 8219 6130 8231
rect 6302 8194 6354 8206
rect 6962 8191 6974 8243
rect 7026 8191 7038 8243
rect 7186 8206 7198 8258
rect 7250 8206 7262 8258
rect 8194 8206 8206 8258
rect 8258 8206 8270 8258
rect 6078 8155 6130 8167
rect 8530 8162 8542 8214
rect 8594 8162 8606 8214
rect 9102 8194 9154 8206
rect 11790 8258 11842 8270
rect 12798 8258 12850 8270
rect 12506 8206 12518 8258
rect 12570 8206 12582 8258
rect 11790 8194 11842 8206
rect 12798 8194 12850 8206
rect 13022 8258 13074 8270
rect 18846 8258 18898 8270
rect 13570 8206 13582 8258
rect 13634 8206 13646 8258
rect 13794 8206 13806 8258
rect 13858 8206 13870 8258
rect 14466 8206 14478 8258
rect 14530 8206 14542 8258
rect 13022 8194 13074 8206
rect 14802 8162 14814 8214
rect 14866 8162 14878 8214
rect 18846 8194 18898 8206
rect 19238 8258 19290 8270
rect 19238 8194 19290 8206
rect 19686 8258 19738 8270
rect 19686 8194 19738 8206
rect 20134 8258 20186 8270
rect 26742 8314 26794 8326
rect 20290 8206 20302 8258
rect 20354 8206 20366 8258
rect 21254 8250 21306 8262
rect 22318 8258 22370 8270
rect 25454 8258 25506 8270
rect 25902 8258 25954 8270
rect 20134 8194 20186 8206
rect 21858 8178 21870 8230
rect 21922 8178 21934 8230
rect 22094 8202 22146 8214
rect 16158 8146 16210 8158
rect 5730 8038 5742 8090
rect 5794 8038 5806 8090
rect 16158 8082 16210 8094
rect 21422 8146 21474 8158
rect 23090 8206 23102 8258
rect 23154 8206 23166 8258
rect 25778 8206 25790 8258
rect 25842 8206 25854 8258
rect 22318 8194 22370 8206
rect 25454 8194 25506 8206
rect 22094 8138 22146 8150
rect 25006 8146 25058 8158
rect 25610 8150 25622 8202
rect 25674 8150 25686 8202
rect 25902 8194 25954 8206
rect 26574 8258 26626 8270
rect 28478 8306 28530 8318
rect 30102 8370 30154 8382
rect 37158 8370 37210 8382
rect 31490 8318 31502 8370
rect 31554 8318 31566 8370
rect 35298 8318 35310 8370
rect 35362 8318 35374 8370
rect 30102 8306 30154 8318
rect 37158 8306 37210 8318
rect 38110 8370 38162 8382
rect 39566 8370 39618 8382
rect 41806 8370 41858 8382
rect 38110 8306 38162 8318
rect 38278 8314 38330 8326
rect 26742 8250 26794 8262
rect 27022 8258 27074 8270
rect 26898 8206 26910 8258
rect 26962 8206 26974 8258
rect 26574 8194 26626 8206
rect 27022 8194 27074 8206
rect 28142 8258 28194 8270
rect 28142 8194 28194 8206
rect 29150 8258 29202 8270
rect 29150 8194 29202 8206
rect 30718 8258 30770 8270
rect 30718 8194 30770 8206
rect 34190 8258 34242 8270
rect 34190 8194 34242 8206
rect 34414 8258 34466 8270
rect 35982 8258 36034 8270
rect 40002 8318 40014 8370
rect 40066 8318 40078 8370
rect 39566 8306 39618 8318
rect 41806 8306 41858 8318
rect 41974 8314 42026 8326
rect 34682 8206 34694 8258
rect 34746 8206 34758 8258
rect 34414 8194 34466 8206
rect 35410 8162 35422 8214
rect 35474 8162 35486 8214
rect 35634 8206 35646 8258
rect 35698 8206 35710 8258
rect 35982 8194 36034 8206
rect 37550 8220 37602 8232
rect 37874 8206 37886 8258
rect 37938 8206 37950 8258
rect 38278 8250 38330 8262
rect 38894 8258 38946 8270
rect 38994 8206 39006 8258
rect 39058 8206 39070 8258
rect 38894 8194 38946 8206
rect 21422 8082 21474 8094
rect 25006 8082 25058 8094
rect 26182 8146 26234 8158
rect 26182 8082 26234 8094
rect 27302 8146 27354 8158
rect 27302 8082 27354 8094
rect 30550 8146 30602 8158
rect 30550 8082 30602 8094
rect 33406 8146 33458 8158
rect 37550 8156 37602 8168
rect 39160 8150 39172 8202
rect 39224 8150 39236 8202
rect 40114 8162 40126 8214
rect 40178 8162 40190 8214
rect 40450 8206 40462 8258
rect 40514 8206 40526 8258
rect 41570 8206 41582 8258
rect 41634 8206 41646 8258
rect 41974 8250 42026 8262
rect 44718 8258 44770 8270
rect 48302 8258 48354 8270
rect 41402 8150 41414 8202
rect 41466 8150 41478 8202
rect 43026 8150 43038 8202
rect 43090 8150 43102 8202
rect 43306 8150 43318 8202
rect 43370 8150 43382 8202
rect 43754 8150 43766 8202
rect 43818 8150 43830 8202
rect 44120 8173 44132 8225
rect 44184 8173 44196 8225
rect 45490 8206 45502 8258
rect 45554 8206 45566 8258
rect 44718 8194 44770 8206
rect 48302 8194 48354 8206
rect 33406 8082 33458 8094
rect 44270 8146 44322 8158
rect 44270 8082 44322 8094
rect 47406 8146 47458 8158
rect 47406 8082 47458 8094
rect 27974 8034 28026 8046
rect 27974 7970 28026 7982
rect 29486 8034 29538 8046
rect 29486 7970 29538 7982
rect 34022 8034 34074 8046
rect 34022 7970 34074 7982
rect 36318 8034 36370 8046
rect 36318 7970 36370 7982
rect 42422 8034 42474 8046
rect 42422 7970 42474 7982
rect 47966 8034 48018 8046
rect 47966 7970 48018 7982
rect 1344 7866 48608 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 48608 7866
rect 1344 7780 48608 7814
rect 12070 7698 12122 7710
rect 5966 7586 6018 7598
rect 6962 7590 6974 7642
rect 7026 7590 7038 7642
rect 7522 7590 7534 7642
rect 7586 7590 7598 7642
rect 9762 7590 9774 7642
rect 9826 7590 9838 7642
rect 12070 7634 12122 7646
rect 17558 7698 17610 7710
rect 17558 7634 17610 7646
rect 22150 7698 22202 7710
rect 22150 7634 22202 7646
rect 23774 7698 23826 7710
rect 23774 7634 23826 7646
rect 26742 7698 26794 7710
rect 26742 7634 26794 7646
rect 30214 7698 30266 7710
rect 30214 7634 30266 7646
rect 16158 7586 16210 7598
rect 34750 7586 34802 7598
rect 5966 7522 6018 7534
rect 13862 7530 13914 7542
rect 3278 7474 3330 7486
rect 6738 7466 6750 7518
rect 6802 7466 6814 7518
rect 7646 7474 7698 7486
rect 7074 7422 7086 7474
rect 7138 7422 7150 7474
rect 7970 7449 7982 7501
rect 8034 7449 8046 7501
rect 9874 7478 9886 7530
rect 9938 7478 9950 7530
rect 10222 7474 10274 7486
rect 8306 7422 8318 7474
rect 8370 7422 8382 7474
rect 9538 7422 9550 7474
rect 9602 7422 9614 7474
rect 10882 7466 10894 7518
rect 10946 7466 10958 7518
rect 12686 7474 12738 7486
rect 11106 7422 11118 7474
rect 11170 7422 11182 7474
rect 3278 7410 3330 7422
rect 7646 7410 7698 7422
rect 10222 7410 10274 7422
rect 12686 7410 12738 7422
rect 12910 7474 12962 7486
rect 12910 7410 12962 7422
rect 13470 7474 13522 7486
rect 13470 7410 13522 7422
rect 13694 7474 13746 7486
rect 13862 7466 13914 7478
rect 14590 7530 14642 7542
rect 33674 7534 33686 7586
rect 33738 7534 33750 7586
rect 38110 7586 38162 7598
rect 16158 7522 16210 7534
rect 18324 7511 18376 7523
rect 14242 7422 14254 7474
rect 14306 7422 14318 7474
rect 14590 7466 14642 7478
rect 15038 7474 15090 7486
rect 15902 7422 15914 7474
rect 15966 7422 15978 7474
rect 16930 7422 16942 7474
rect 16994 7422 17006 7474
rect 25488 7512 25540 7524
rect 21982 7494 22034 7506
rect 18622 7474 18674 7486
rect 18324 7447 18376 7459
rect 18498 7422 18510 7474
rect 18562 7422 18574 7474
rect 13694 7410 13746 7422
rect 15038 7410 15090 7422
rect 18622 7410 18674 7422
rect 19182 7474 19234 7486
rect 21870 7474 21922 7486
rect 21074 7422 21086 7474
rect 21138 7422 21150 7474
rect 21982 7430 22034 7442
rect 24110 7474 24162 7486
rect 19182 7410 19234 7422
rect 21870 7410 21922 7422
rect 24110 7410 24162 7422
rect 25230 7474 25282 7486
rect 25330 7422 25342 7474
rect 25394 7422 25406 7474
rect 25488 7448 25540 7460
rect 26910 7474 26962 7486
rect 30762 7478 30774 7530
rect 30826 7478 30838 7530
rect 32140 7512 32192 7524
rect 31334 7474 31386 7486
rect 30930 7422 30942 7474
rect 30994 7422 31006 7474
rect 34190 7512 34242 7524
rect 34750 7522 34802 7534
rect 34918 7530 34970 7542
rect 32398 7474 32450 7486
rect 32140 7448 32192 7460
rect 32274 7422 32286 7474
rect 32338 7422 32350 7474
rect 25230 7410 25282 7422
rect 26910 7410 26962 7422
rect 31334 7410 31386 7422
rect 32398 7410 32450 7422
rect 33182 7474 33234 7486
rect 33182 7410 33234 7422
rect 33406 7474 33458 7486
rect 43418 7534 43430 7586
rect 43482 7534 43494 7586
rect 38110 7522 38162 7534
rect 34190 7448 34242 7460
rect 34514 7422 34526 7474
rect 34578 7422 34590 7474
rect 34918 7466 34970 7478
rect 35422 7474 35474 7486
rect 33406 7410 33458 7422
rect 35422 7410 35474 7422
rect 39342 7474 39394 7486
rect 39342 7410 39394 7422
rect 39678 7474 39730 7486
rect 40002 7478 40014 7530
rect 40066 7478 40078 7530
rect 41022 7474 41074 7486
rect 41302 7474 41354 7486
rect 42926 7474 42978 7486
rect 40338 7422 40350 7474
rect 40402 7422 40414 7474
rect 41122 7422 41134 7474
rect 41186 7422 41198 7474
rect 42242 7422 42254 7474
rect 42306 7422 42318 7474
rect 42578 7422 42590 7474
rect 42642 7422 42654 7474
rect 39678 7410 39730 7422
rect 41022 7410 41074 7422
rect 41302 7410 41354 7422
rect 42926 7410 42978 7422
rect 43150 7474 43202 7486
rect 43922 7455 43934 7507
rect 43986 7455 43998 7507
rect 44202 7478 44214 7530
rect 44266 7478 44278 7530
rect 44650 7478 44662 7530
rect 44714 7478 44726 7530
rect 44974 7462 44986 7514
rect 45038 7462 45050 7514
rect 48302 7474 48354 7486
rect 43150 7410 43202 7422
rect 48302 7410 48354 7422
rect 14030 7362 14082 7374
rect 4050 7310 4062 7362
rect 4114 7310 4126 7362
rect 10770 7310 10782 7362
rect 10834 7310 10846 7362
rect 14030 7298 14082 7310
rect 17950 7362 18002 7374
rect 17950 7298 18002 7310
rect 24726 7362 24778 7374
rect 24726 7298 24778 7310
rect 25902 7362 25954 7374
rect 31166 7362 31218 7374
rect 27682 7310 27694 7362
rect 27746 7310 27758 7362
rect 29586 7310 29598 7362
rect 29650 7310 29662 7362
rect 25902 7298 25954 7310
rect 31166 7298 31218 7310
rect 31726 7362 31778 7374
rect 38726 7362 38778 7374
rect 36194 7310 36206 7362
rect 36258 7310 36270 7362
rect 31726 7298 31778 7310
rect 38726 7298 38778 7310
rect 40014 7362 40066 7374
rect 40014 7298 40066 7310
rect 41694 7362 41746 7374
rect 41694 7298 41746 7310
rect 42702 7306 42754 7318
rect 45042 7310 45054 7362
rect 45106 7310 45118 7362
rect 45602 7310 45614 7362
rect 45666 7310 45678 7362
rect 47506 7310 47518 7362
rect 47570 7310 47582 7362
rect 16774 7250 16826 7262
rect 12394 7198 12406 7250
rect 12458 7198 12470 7250
rect 13178 7198 13190 7250
rect 13242 7198 13254 7250
rect 42702 7242 42754 7254
rect 16774 7186 16826 7198
rect 1344 7082 48608 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 48608 7082
rect 1344 6996 48608 7030
rect 4174 6914 4226 6926
rect 25454 6914 25506 6926
rect 4174 6850 4226 6862
rect 13918 6858 13970 6870
rect 25454 6850 25506 6862
rect 47070 6858 47122 6870
rect 6514 6750 6526 6802
rect 6578 6750 6590 6802
rect 10882 6750 10894 6802
rect 10946 6750 10958 6802
rect 13918 6794 13970 6806
rect 15150 6802 15202 6814
rect 15150 6738 15202 6750
rect 18510 6802 18562 6814
rect 18510 6738 18562 6750
rect 20022 6802 20074 6814
rect 27358 6802 27410 6814
rect 43038 6802 43090 6814
rect 44034 6806 44046 6858
rect 44098 6806 44110 6858
rect 20022 6738 20074 6750
rect 22374 6746 22426 6758
rect 4510 6690 4562 6702
rect 4510 6626 4562 6638
rect 5182 6690 5234 6702
rect 5182 6626 5234 6638
rect 5798 6690 5850 6702
rect 7086 6690 7138 6702
rect 10110 6690 10162 6702
rect 6066 6638 6078 6690
rect 6130 6638 6142 6690
rect 5798 6626 5850 6638
rect 6402 6594 6414 6646
rect 6466 6594 6478 6646
rect 7858 6638 7870 6690
rect 7922 6638 7934 6690
rect 7086 6626 7138 6638
rect 10110 6626 10162 6638
rect 12798 6690 12850 6702
rect 14478 6690 14530 6702
rect 13794 6638 13806 6690
rect 13858 6638 13870 6690
rect 12798 6626 12850 6638
rect 9774 6578 9826 6590
rect 13570 6582 13582 6634
rect 13634 6582 13646 6634
rect 14478 6626 14530 6638
rect 14814 6690 14866 6702
rect 17054 6690 17106 6702
rect 14814 6626 14866 6638
rect 15038 6651 15090 6663
rect 15474 6638 15486 6690
rect 15538 6638 15550 6690
rect 15038 6587 15090 6599
rect 15766 6634 15818 6646
rect 16146 6638 16158 6690
rect 16210 6638 16222 6690
rect 16370 6610 16382 6662
rect 16434 6610 16446 6662
rect 17054 6626 17106 6638
rect 17390 6690 17442 6702
rect 17390 6626 17442 6638
rect 17838 6690 17890 6702
rect 17838 6626 17890 6638
rect 18174 6690 18226 6702
rect 19630 6690 19682 6702
rect 18722 6638 18734 6690
rect 18786 6638 18798 6690
rect 18174 6626 18226 6638
rect 15766 6570 15818 6582
rect 15934 6578 15986 6590
rect 18498 6582 18510 6634
rect 18562 6582 18574 6634
rect 19630 6626 19682 6638
rect 20470 6690 20522 6702
rect 22374 6682 22426 6694
rect 23942 6746 23994 6758
rect 25890 6750 25902 6802
rect 25954 6750 25966 6802
rect 27190 6746 27242 6758
rect 20470 6626 20522 6638
rect 21534 6634 21586 6646
rect 21746 6610 21758 6662
rect 21810 6610 21822 6662
rect 23314 6610 23326 6662
rect 23378 6610 23390 6662
rect 23538 6638 23550 6690
rect 23602 6638 23614 6690
rect 23942 6682 23994 6694
rect 24782 6690 24834 6702
rect 31042 6750 31054 6802
rect 31106 6750 31118 6802
rect 35410 6750 35422 6802
rect 35474 6750 35486 6802
rect 27358 6738 27410 6750
rect 37270 6746 37322 6758
rect 41570 6750 41582 6802
rect 41634 6750 41646 6802
rect 47070 6794 47122 6806
rect 24434 6638 24446 6690
rect 24498 6638 24510 6690
rect 24882 6638 24894 6690
rect 24946 6638 24958 6690
rect 24782 6626 24834 6638
rect 9774 6514 9826 6526
rect 21534 6570 21586 6582
rect 22206 6578 22258 6590
rect 15934 6514 15986 6526
rect 22206 6514 22258 6526
rect 23774 6578 23826 6590
rect 25050 6582 25062 6634
rect 25114 6582 25126 6634
rect 26002 6594 26014 6646
rect 26066 6594 26078 6646
rect 26226 6638 26238 6690
rect 26290 6638 26302 6690
rect 27190 6682 27242 6694
rect 29766 6690 29818 6702
rect 27570 6638 27582 6690
rect 27634 6638 27646 6690
rect 27794 6610 27806 6662
rect 27858 6610 27870 6662
rect 28578 6638 28590 6690
rect 28642 6638 28654 6690
rect 29362 6638 29374 6690
rect 29426 6638 29438 6690
rect 29766 6626 29818 6638
rect 30270 6690 30322 6702
rect 30270 6626 30322 6638
rect 36206 6690 36258 6702
rect 43038 6738 43090 6750
rect 37270 6682 37322 6694
rect 38334 6690 38386 6702
rect 37650 6638 37662 6690
rect 37714 6638 37726 6690
rect 37998 6652 38050 6664
rect 36206 6626 36258 6638
rect 38334 6626 38386 6638
rect 38670 6690 38722 6702
rect 39790 6690 39842 6702
rect 39106 6638 39118 6690
rect 39170 6638 39182 6690
rect 38670 6626 38722 6638
rect 39442 6611 39454 6663
rect 39506 6611 39518 6663
rect 39790 6626 39842 6638
rect 40238 6690 40290 6702
rect 42366 6690 42418 6702
rect 45390 6690 45442 6702
rect 40238 6626 40290 6638
rect 32958 6578 33010 6590
rect 23774 6514 23826 6526
rect 24278 6522 24330 6534
rect 4846 6466 4898 6478
rect 4846 6402 4898 6414
rect 19294 6466 19346 6478
rect 19294 6402 19346 6414
rect 22822 6466 22874 6478
rect 29206 6522 29258 6534
rect 24278 6458 24330 6470
rect 26854 6466 26906 6478
rect 22822 6402 22874 6414
rect 26854 6402 26906 6414
rect 28422 6466 28474 6478
rect 32958 6514 33010 6526
rect 33518 6578 33570 6590
rect 33518 6514 33570 6526
rect 37438 6578 37490 6590
rect 37998 6588 38050 6600
rect 41682 6594 41694 6646
rect 41746 6594 41758 6646
rect 42018 6638 42030 6690
rect 42082 6638 42094 6690
rect 42466 6638 42478 6690
rect 42530 6638 42542 6690
rect 43698 6638 43710 6690
rect 43762 6638 43774 6690
rect 44034 6638 44046 6690
rect 44098 6638 44110 6690
rect 44818 6638 44830 6690
rect 44882 6638 44894 6690
rect 42366 6626 42418 6638
rect 42634 6582 42646 6634
rect 42698 6582 42710 6634
rect 45390 6626 45442 6638
rect 45614 6690 45666 6702
rect 45614 6626 45666 6638
rect 46286 6690 46338 6702
rect 46286 6626 46338 6638
rect 46398 6690 46450 6702
rect 48134 6690 48186 6702
rect 46666 6638 46678 6690
rect 46730 6638 46742 6690
rect 47170 6638 47182 6690
rect 47234 6638 47246 6690
rect 47506 6638 47518 6690
rect 47570 6638 47582 6690
rect 46398 6626 46450 6638
rect 48134 6626 48186 6638
rect 45882 6526 45894 6578
rect 45946 6526 45958 6578
rect 37438 6514 37490 6526
rect 39218 6470 39230 6522
rect 39282 6470 39294 6522
rect 29206 6458 29258 6470
rect 40574 6466 40626 6478
rect 28422 6402 28474 6414
rect 40574 6402 40626 6414
rect 41190 6466 41242 6478
rect 41190 6402 41242 6414
rect 44998 6466 45050 6478
rect 44998 6402 45050 6414
rect 1344 6298 48608 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 48608 6298
rect 1344 6212 48608 6246
rect 8150 6130 8202 6142
rect 8150 6066 8202 6078
rect 9662 6130 9714 6142
rect 9662 6066 9714 6078
rect 10390 6130 10442 6142
rect 10390 6066 10442 6078
rect 12070 6130 12122 6142
rect 12070 6066 12122 6078
rect 32342 6130 32394 6142
rect 7534 6018 7586 6030
rect 7534 5954 7586 5966
rect 12350 6018 12402 6030
rect 12350 5954 12402 5966
rect 14926 6018 14978 6030
rect 18386 6022 18398 6074
rect 18450 6022 18462 6074
rect 32342 6066 32394 6078
rect 8710 5935 8762 5947
rect 4846 5906 4898 5918
rect 5618 5854 5630 5906
rect 5682 5854 5694 5906
rect 9998 5906 10050 5918
rect 8710 5871 8762 5883
rect 8978 5854 8990 5906
rect 9042 5854 9054 5906
rect 12497 5887 12509 5939
rect 12561 5887 12573 5939
rect 12786 5910 12798 5962
rect 12850 5910 12862 5962
rect 13122 5910 13134 5962
rect 13186 5910 13198 5962
rect 13458 5910 13470 5962
rect 13522 5910 13534 5962
rect 14926 5954 14978 5966
rect 24558 6018 24610 6030
rect 14814 5906 14866 5918
rect 4846 5842 4898 5854
rect 9998 5842 10050 5854
rect 15262 5906 15314 5918
rect 14814 5842 14866 5854
rect 15094 5850 15146 5862
rect 14198 5794 14250 5806
rect 8530 5742 8542 5794
rect 8594 5742 8606 5794
rect 15698 5854 15710 5906
rect 15762 5854 15774 5906
rect 16034 5854 16046 5906
rect 16098 5854 16110 5906
rect 16482 5869 16494 5921
rect 16546 5869 16558 5921
rect 18050 5910 18062 5962
rect 18114 5910 18126 5962
rect 24558 5954 24610 5966
rect 29150 6018 29202 6030
rect 45950 6018 46002 6030
rect 25528 5943 25580 5955
rect 29150 5954 29202 5966
rect 29934 5962 29986 5974
rect 18286 5906 18338 5918
rect 21646 5906 21698 5918
rect 16818 5854 16830 5906
rect 16882 5854 16894 5906
rect 17602 5854 17614 5906
rect 17666 5854 17678 5906
rect 20850 5854 20862 5906
rect 20914 5854 20926 5906
rect 15262 5842 15314 5854
rect 18286 5842 18338 5854
rect 21646 5842 21698 5854
rect 21870 5906 21922 5918
rect 25230 5906 25282 5918
rect 22642 5854 22654 5906
rect 22706 5854 22718 5906
rect 25330 5854 25342 5906
rect 25394 5854 25406 5906
rect 25528 5879 25580 5891
rect 26462 5906 26514 5918
rect 29934 5898 29986 5910
rect 30046 5962 30098 5974
rect 31166 5962 31218 5974
rect 37258 5966 37270 6018
rect 37322 5966 37334 6018
rect 43978 5966 43990 6018
rect 44042 5966 44054 6018
rect 46890 5966 46902 6018
rect 46954 5966 46966 6018
rect 30046 5898 30098 5910
rect 30774 5906 30826 5918
rect 21870 5842 21922 5854
rect 25230 5842 25282 5854
rect 26462 5842 26514 5854
rect 31166 5898 31218 5910
rect 33070 5906 33122 5918
rect 31490 5854 31502 5906
rect 31554 5854 31566 5906
rect 30774 5842 30826 5854
rect 31894 5850 31946 5862
rect 32498 5854 32510 5906
rect 32562 5854 32574 5906
rect 33170 5854 33182 5906
rect 33234 5854 33246 5906
rect 33328 5904 33340 5956
rect 33392 5904 33404 5956
rect 39304 5944 39356 5956
rect 34526 5906 34578 5918
rect 15094 5786 15146 5798
rect 30606 5794 30658 5806
rect 14198 5730 14250 5742
rect 15598 5738 15650 5750
rect 16370 5742 16382 5794
rect 16434 5742 16446 5794
rect 18946 5742 18958 5794
rect 19010 5742 19022 5794
rect 27234 5742 27246 5794
rect 27298 5742 27310 5794
rect 14534 5682 14586 5694
rect 30606 5730 30658 5742
rect 31726 5794 31778 5806
rect 33070 5842 33122 5854
rect 34526 5842 34578 5854
rect 34750 5906 34802 5918
rect 34750 5842 34802 5854
rect 34974 5906 35026 5918
rect 34974 5842 35026 5854
rect 35086 5906 35138 5918
rect 35086 5842 35138 5854
rect 36206 5906 36258 5918
rect 36206 5842 36258 5854
rect 36990 5906 37042 5918
rect 36990 5842 37042 5854
rect 37550 5906 37602 5918
rect 37550 5842 37602 5854
rect 37774 5906 37826 5918
rect 38334 5906 38386 5918
rect 38042 5854 38054 5906
rect 38106 5854 38118 5906
rect 37774 5842 37826 5854
rect 38334 5842 38386 5854
rect 38446 5906 38498 5918
rect 38446 5842 38498 5854
rect 39006 5906 39058 5918
rect 39106 5854 39118 5906
rect 39170 5854 39182 5906
rect 39304 5880 39356 5892
rect 40002 5854 40014 5906
rect 40066 5854 40078 5906
rect 40898 5854 40910 5906
rect 40962 5854 40974 5906
rect 41234 5869 41246 5921
rect 41298 5869 41310 5921
rect 41806 5906 41858 5918
rect 39006 5842 39058 5854
rect 41806 5842 41858 5854
rect 42142 5906 42194 5918
rect 42142 5842 42194 5854
rect 43374 5906 43426 5918
rect 43374 5842 43426 5854
rect 43598 5906 43650 5918
rect 43598 5842 43650 5854
rect 43710 5906 43762 5918
rect 44706 5910 44718 5962
rect 44770 5910 44782 5962
rect 44986 5910 44998 5962
rect 45050 5910 45062 5962
rect 45490 5910 45502 5962
rect 45554 5910 45566 5962
rect 45950 5954 46002 5966
rect 45800 5887 45812 5939
rect 45864 5887 45876 5939
rect 46398 5906 46450 5918
rect 43710 5842 43762 5854
rect 46398 5842 46450 5854
rect 46622 5906 46674 5918
rect 47394 5854 47406 5906
rect 47458 5854 47470 5906
rect 47618 5854 47630 5906
rect 47682 5854 47694 5906
rect 46622 5842 46674 5854
rect 31894 5786 31946 5798
rect 33742 5794 33794 5806
rect 31726 5730 31778 5742
rect 33742 5730 33794 5742
rect 35870 5794 35922 5806
rect 35870 5730 35922 5742
rect 36654 5794 36706 5806
rect 36654 5730 36706 5742
rect 39678 5794 39730 5806
rect 42534 5794 42586 5806
rect 39678 5730 39730 5742
rect 40182 5738 40234 5750
rect 41346 5742 41358 5794
rect 41410 5742 41422 5794
rect 48246 5794 48298 5806
rect 15598 5674 15650 5686
rect 25902 5682 25954 5694
rect 42534 5730 42586 5742
rect 47294 5738 47346 5750
rect 14534 5618 14586 5630
rect 34234 5630 34246 5682
rect 34298 5630 34310 5682
rect 35354 5630 35366 5682
rect 35418 5630 35430 5682
rect 40182 5674 40234 5686
rect 43038 5682 43090 5694
rect 48246 5730 48298 5742
rect 47294 5674 47346 5686
rect 25902 5618 25954 5630
rect 43038 5618 43090 5630
rect 1344 5514 48608 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 48608 5514
rect 1344 5428 48608 5462
rect 21366 5346 21418 5358
rect 32678 5346 32730 5358
rect 12562 5238 12574 5290
rect 12626 5238 12638 5290
rect 21366 5282 21418 5294
rect 21758 5290 21810 5302
rect 18510 5234 18562 5246
rect 18510 5170 18562 5182
rect 19630 5234 19682 5246
rect 19630 5170 19682 5182
rect 20806 5234 20858 5246
rect 21758 5226 21810 5238
rect 23214 5290 23266 5302
rect 32678 5282 32730 5294
rect 34302 5346 34354 5358
rect 41246 5346 41298 5358
rect 34302 5282 34354 5294
rect 34750 5290 34802 5302
rect 23214 5226 23266 5238
rect 27022 5234 27074 5246
rect 20806 5170 20858 5182
rect 26854 5178 26906 5190
rect 15262 5122 15314 5134
rect 17950 5122 18002 5134
rect 12562 5070 12574 5122
rect 12626 5070 12638 5122
rect 12786 5070 12798 5122
rect 12850 5070 12862 5122
rect 13638 5030 13650 5082
rect 13702 5030 13714 5082
rect 16034 5070 16046 5122
rect 16098 5070 16110 5122
rect 13470 5010 13522 5022
rect 13962 5014 13974 5066
rect 14026 5014 14038 5066
rect 14410 5014 14422 5066
rect 14474 5014 14486 5066
rect 14578 5014 14590 5066
rect 14642 5014 14654 5066
rect 15262 5058 15314 5070
rect 17950 5058 18002 5070
rect 18902 5122 18954 5134
rect 19182 5122 19234 5134
rect 20302 5122 20354 5134
rect 23438 5122 23490 5134
rect 27022 5170 27074 5182
rect 29318 5234 29370 5246
rect 33350 5234 33402 5246
rect 32162 5182 32174 5234
rect 32226 5182 32238 5234
rect 34750 5226 34802 5238
rect 35534 5290 35586 5302
rect 41246 5282 41298 5294
rect 45054 5346 45106 5358
rect 45054 5282 45106 5294
rect 35534 5226 35586 5238
rect 37662 5234 37714 5246
rect 27682 5126 27694 5178
rect 27746 5126 27758 5178
rect 29318 5170 29370 5182
rect 33350 5170 33402 5182
rect 40462 5234 40514 5246
rect 37662 5170 37714 5182
rect 39286 5178 39338 5190
rect 19058 5070 19070 5122
rect 19122 5070 19134 5122
rect 20178 5070 20190 5122
rect 20242 5070 20254 5122
rect 21186 5070 21198 5122
rect 21250 5070 21262 5122
rect 21858 5070 21870 5122
rect 21922 5070 21934 5122
rect 22194 5070 22206 5122
rect 22258 5070 22270 5122
rect 22866 5070 22878 5122
rect 22930 5070 22942 5122
rect 23090 5070 23102 5122
rect 23154 5070 23166 5122
rect 24210 5070 24222 5122
rect 24274 5070 24286 5122
rect 26854 5114 26906 5126
rect 27918 5122 27970 5134
rect 18902 5058 18954 5070
rect 19182 5058 19234 5070
rect 20010 5014 20022 5066
rect 20074 5014 20086 5066
rect 20302 5058 20354 5070
rect 23438 5058 23490 5070
rect 27458 5042 27470 5094
rect 27522 5042 27534 5094
rect 27918 5058 27970 5070
rect 28254 5122 28306 5134
rect 28254 5058 28306 5070
rect 29486 5122 29538 5134
rect 33630 5122 33682 5134
rect 33910 5122 33962 5134
rect 36486 5122 36538 5134
rect 37830 5122 37882 5134
rect 39118 5122 39170 5134
rect 30258 5070 30270 5122
rect 30322 5070 30334 5122
rect 32498 5070 32510 5122
rect 32562 5070 32574 5122
rect 33730 5070 33742 5122
rect 33794 5070 33806 5122
rect 34850 5070 34862 5122
rect 34914 5070 34926 5122
rect 35186 5070 35198 5122
rect 35250 5070 35262 5122
rect 35634 5070 35646 5122
rect 35698 5070 35710 5122
rect 35970 5070 35982 5122
rect 36034 5070 36046 5122
rect 29486 5058 29538 5070
rect 33630 5058 33682 5070
rect 33910 5058 33962 5070
rect 36486 5058 36538 5070
rect 37102 5084 37154 5096
rect 37426 5070 37438 5122
rect 37490 5070 37502 5122
rect 37830 5058 37882 5070
rect 38558 5084 38610 5096
rect 13470 4946 13522 4958
rect 26126 5010 26178 5022
rect 37102 5020 37154 5032
rect 38882 5070 38894 5122
rect 38946 5070 38958 5122
rect 40462 5170 40514 5182
rect 43374 5234 43426 5246
rect 43810 5182 43822 5234
rect 43874 5182 43886 5234
rect 45602 5182 45614 5234
rect 45666 5182 45678 5234
rect 47506 5182 47518 5234
rect 47570 5182 47582 5234
rect 43374 5170 43426 5182
rect 39286 5114 39338 5126
rect 39790 5122 39842 5134
rect 39118 5058 39170 5070
rect 39790 5058 39842 5070
rect 40126 5122 40178 5134
rect 42366 5122 42418 5134
rect 40786 5070 40798 5122
rect 40850 5070 40862 5122
rect 40126 5058 40178 5070
rect 38558 5020 38610 5032
rect 40338 5014 40350 5066
rect 40402 5014 40414 5066
rect 41477 5039 41489 5091
rect 41541 5039 41553 5091
rect 42366 5058 42418 5070
rect 42702 5122 42754 5134
rect 42980 5122 43032 5134
rect 44718 5122 44770 5134
rect 42802 5070 42814 5122
rect 42866 5070 42878 5122
rect 42702 5058 42754 5070
rect 42980 5058 43032 5070
rect 43922 5055 43934 5107
rect 43986 5055 43998 5107
rect 44258 5070 44270 5122
rect 44322 5070 44334 5122
rect 44718 5058 44770 5070
rect 48302 5122 48354 5134
rect 48302 5058 48354 5070
rect 26126 4946 26178 4958
rect 1344 4730 48608 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 48608 4730
rect 1344 4644 48608 4678
rect 11734 4562 11786 4574
rect 30102 4562 30154 4574
rect 11734 4498 11786 4510
rect 17446 4506 17498 4518
rect 14590 4450 14642 4462
rect 30102 4498 30154 4510
rect 33238 4562 33290 4574
rect 33238 4498 33290 4510
rect 47910 4562 47962 4574
rect 47910 4498 47962 4510
rect 17446 4442 17498 4454
rect 25230 4450 25282 4462
rect 23146 4398 23158 4450
rect 23210 4398 23222 4450
rect 14590 4386 14642 4398
rect 11902 4338 11954 4350
rect 15362 4342 15374 4394
rect 15426 4342 15438 4394
rect 15586 4342 15598 4394
rect 15650 4342 15662 4394
rect 16034 4342 16046 4394
rect 16098 4342 16110 4394
rect 25230 4386 25282 4398
rect 29486 4450 29538 4462
rect 12674 4286 12686 4338
rect 12738 4286 12750 4338
rect 16344 4326 16356 4378
rect 16408 4326 16420 4378
rect 17266 4286 17278 4338
rect 17330 4286 17342 4338
rect 17938 4286 17950 4338
rect 18002 4286 18014 4338
rect 18274 4330 18286 4382
rect 18338 4330 18350 4382
rect 19630 4338 19682 4350
rect 19058 4286 19070 4338
rect 19122 4286 19134 4338
rect 19282 4286 19294 4338
rect 19346 4286 19358 4338
rect 11902 4274 11954 4286
rect 19630 4274 19682 4286
rect 22318 4338 22370 4350
rect 22318 4274 22370 4286
rect 22654 4338 22706 4350
rect 22654 4274 22706 4286
rect 22878 4338 22930 4350
rect 22878 4274 22930 4286
rect 23438 4338 23490 4350
rect 23438 4274 23490 4286
rect 24558 4338 24610 4350
rect 24558 4274 24610 4286
rect 24782 4338 24834 4350
rect 25398 4319 25410 4371
rect 25462 4319 25474 4371
rect 25554 4322 25566 4374
rect 25618 4322 25630 4374
rect 26002 4342 26014 4394
rect 26066 4342 26078 4394
rect 26338 4342 26350 4394
rect 26402 4342 26414 4394
rect 29486 4386 29538 4398
rect 36318 4450 36370 4462
rect 31580 4376 31632 4388
rect 36318 4386 36370 4398
rect 39342 4450 39394 4462
rect 39342 4386 39394 4398
rect 45390 4450 45442 4462
rect 26798 4338 26850 4350
rect 24782 4274 24834 4286
rect 31838 4338 31890 4350
rect 33630 4338 33682 4350
rect 31580 4312 31632 4324
rect 31714 4286 31726 4338
rect 31778 4286 31790 4338
rect 32386 4286 32398 4338
rect 32450 4286 32462 4338
rect 26798 4274 26850 4286
rect 31838 4274 31890 4286
rect 33630 4274 33682 4286
rect 36654 4338 36706 4350
rect 41402 4342 41414 4394
rect 41466 4342 41478 4394
rect 41682 4342 41694 4394
rect 41746 4342 41758 4394
rect 42186 4342 42198 4394
rect 42250 4342 42262 4394
rect 42466 4342 42478 4394
rect 42530 4342 42542 4394
rect 45390 4386 45442 4398
rect 42702 4338 42754 4350
rect 39890 4286 39902 4338
rect 39954 4286 39966 4338
rect 40226 4286 40238 4338
rect 40290 4286 40302 4338
rect 36654 4274 36706 4286
rect 42702 4274 42754 4286
rect 45726 4338 45778 4350
rect 45726 4274 45778 4286
rect 45950 4338 46002 4350
rect 45950 4274 46002 4286
rect 46734 4338 46786 4350
rect 46734 4274 46786 4286
rect 47070 4338 47122 4350
rect 47070 4274 47122 4286
rect 30774 4226 30826 4238
rect 16370 4174 16382 4226
rect 16434 4174 16446 4226
rect 18386 4174 18398 4226
rect 18450 4174 18462 4226
rect 20402 4174 20414 4226
rect 20466 4174 20478 4226
rect 24266 4174 24278 4226
rect 24330 4174 24342 4226
rect 27570 4174 27582 4226
rect 27634 4174 27646 4226
rect 19170 4118 19182 4170
rect 19234 4118 19246 4170
rect 30774 4162 30826 4174
rect 31166 4226 31218 4238
rect 47462 4226 47514 4238
rect 31166 4162 31218 4174
rect 32230 4170 32282 4182
rect 34402 4174 34414 4226
rect 34466 4174 34478 4226
rect 37426 4174 37438 4226
rect 37490 4174 37502 4226
rect 23774 4114 23826 4126
rect 32230 4106 32282 4118
rect 39790 4170 39842 4182
rect 41346 4174 41358 4226
rect 41410 4174 41422 4226
rect 43474 4174 43486 4226
rect 43538 4174 43550 4226
rect 47462 4162 47514 4174
rect 39790 4106 39842 4118
rect 46218 4062 46230 4114
rect 46282 4062 46294 4114
rect 23774 4050 23826 4062
rect 1344 3946 48608 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 48608 3946
rect 1344 3860 48608 3894
rect 15038 3778 15090 3790
rect 13806 3722 13858 3734
rect 22430 3778 22482 3790
rect 15038 3714 15090 3726
rect 16382 3722 16434 3734
rect 13806 3658 13858 3670
rect 22430 3714 22482 3726
rect 25902 3722 25954 3734
rect 38602 3726 38614 3778
rect 38666 3726 38678 3778
rect 42186 3726 42198 3778
rect 42250 3726 42262 3778
rect 44830 3722 44882 3734
rect 16382 3658 16434 3670
rect 17222 3666 17274 3678
rect 17222 3602 17274 3614
rect 18398 3666 18450 3678
rect 18398 3602 18450 3614
rect 23270 3666 23322 3678
rect 23270 3602 23322 3614
rect 24838 3666 24890 3678
rect 25902 3658 25954 3670
rect 27134 3666 27186 3678
rect 32342 3666 32394 3678
rect 24838 3602 24890 3614
rect 26966 3610 27018 3622
rect 14478 3554 14530 3566
rect 13346 3502 13358 3554
rect 13410 3502 13422 3554
rect 13682 3502 13694 3554
rect 13746 3502 13758 3554
rect 14186 3502 14198 3554
rect 14250 3502 14262 3554
rect 14478 3490 14530 3502
rect 14702 3554 14754 3566
rect 14702 3490 14754 3502
rect 15374 3554 15426 3566
rect 17838 3554 17890 3566
rect 16034 3502 16046 3554
rect 16098 3502 16110 3554
rect 16258 3502 16270 3554
rect 16322 3502 16334 3554
rect 17546 3502 17558 3554
rect 17610 3502 17622 3554
rect 15374 3490 15426 3502
rect 17838 3490 17890 3502
rect 17950 3554 18002 3566
rect 17950 3490 18002 3502
rect 18734 3554 18786 3566
rect 20078 3554 20130 3566
rect 19786 3502 19798 3554
rect 19850 3502 19862 3554
rect 18734 3490 18786 3502
rect 20078 3490 20130 3502
rect 20302 3554 20354 3566
rect 22766 3554 22818 3566
rect 25454 3554 25506 3566
rect 20302 3490 20354 3502
rect 20918 3469 20930 3521
rect 20982 3469 20994 3521
rect 12630 3442 12682 3454
rect 12630 3378 12682 3390
rect 20750 3442 20802 3454
rect 21074 3446 21086 3498
rect 21138 3446 21150 3498
rect 21522 3465 21534 3517
rect 21586 3465 21598 3517
rect 21970 3469 21982 3521
rect 22034 3469 22046 3521
rect 25162 3502 25174 3554
rect 25226 3502 25238 3554
rect 22766 3490 22818 3502
rect 25454 3490 25506 3502
rect 25678 3554 25730 3566
rect 29586 3614 29598 3666
rect 29650 3614 29662 3666
rect 31490 3614 31502 3666
rect 31554 3614 31566 3666
rect 27134 3602 27186 3614
rect 32342 3602 32394 3614
rect 32790 3666 32842 3678
rect 32790 3602 32842 3614
rect 33238 3666 33290 3678
rect 35478 3666 35530 3678
rect 34626 3614 34638 3666
rect 34690 3614 34702 3666
rect 33238 3602 33290 3614
rect 35478 3602 35530 3614
rect 36374 3666 36426 3678
rect 39174 3666 39226 3678
rect 37762 3614 37774 3666
rect 37826 3614 37838 3666
rect 36374 3602 36426 3614
rect 39174 3602 39226 3614
rect 39958 3666 40010 3678
rect 41682 3670 41694 3722
rect 41746 3670 41758 3722
rect 43094 3666 43146 3678
rect 43698 3670 43710 3722
rect 43762 3670 43774 3722
rect 39958 3602 40010 3614
rect 40854 3610 40906 3622
rect 26002 3502 26014 3554
rect 26066 3502 26078 3554
rect 26226 3502 26238 3554
rect 26290 3502 26302 3554
rect 26966 3546 27018 3558
rect 28814 3554 28866 3566
rect 27694 3516 27746 3528
rect 25678 3490 25730 3502
rect 20750 3378 20802 3390
rect 24054 3442 24106 3454
rect 27694 3452 27746 3464
rect 27806 3498 27858 3510
rect 28578 3502 28590 3554
rect 28642 3502 28654 3554
rect 38222 3554 38274 3566
rect 28814 3490 28866 3502
rect 33618 3469 33630 3521
rect 33682 3469 33694 3521
rect 33954 3465 33966 3517
rect 34018 3465 34030 3517
rect 34234 3446 34246 3498
rect 34298 3446 34310 3498
rect 34600 3462 34612 3514
rect 34664 3462 34676 3514
rect 36754 3469 36766 3521
rect 36818 3469 36830 3521
rect 37090 3465 37102 3517
rect 37154 3465 37166 3517
rect 37426 3469 37438 3521
rect 37490 3469 37502 3521
rect 37736 3462 37748 3514
rect 37800 3462 37812 3514
rect 38222 3490 38274 3502
rect 38334 3554 38386 3566
rect 38334 3490 38386 3502
rect 40294 3554 40346 3566
rect 40294 3490 40346 3502
rect 40574 3554 40626 3566
rect 44830 3658 44882 3670
rect 45334 3666 45386 3678
rect 43094 3602 43146 3614
rect 45334 3602 45386 3614
rect 45782 3666 45834 3678
rect 45782 3602 45834 3614
rect 46678 3666 46730 3678
rect 46678 3602 46730 3614
rect 47574 3666 47626 3678
rect 47574 3602 47626 3614
rect 48022 3666 48074 3678
rect 48022 3602 48074 3614
rect 40854 3546 40906 3558
rect 41022 3554 41074 3566
rect 42478 3554 42530 3566
rect 40574 3490 40626 3502
rect 41458 3502 41470 3554
rect 41522 3502 41534 3554
rect 41682 3502 41694 3554
rect 41746 3502 41758 3554
rect 41022 3490 41074 3502
rect 42478 3490 42530 3502
rect 42590 3554 42642 3566
rect 43698 3502 43710 3554
rect 43762 3502 43774 3554
rect 44034 3502 44046 3554
rect 44098 3502 44110 3554
rect 44482 3502 44494 3554
rect 44546 3502 44558 3554
rect 44706 3502 44718 3554
rect 44770 3502 44782 3554
rect 42590 3490 42642 3502
rect 27806 3434 27858 3446
rect 40686 3442 40738 3454
rect 24054 3378 24106 3390
rect 28422 3386 28474 3398
rect 19462 3330 19514 3342
rect 40686 3378 40738 3390
rect 28422 3322 28474 3334
rect 46230 3330 46282 3342
rect 19462 3266 19514 3278
rect 46230 3266 46282 3278
rect 1344 3162 48608 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 48608 3162
rect 1344 3076 48608 3110
<< via1 >>
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 19182 46062 19234 46114
rect 22542 46062 22594 46114
rect 25846 46062 25898 46114
rect 28814 46006 28866 46058
rect 33182 46062 33234 46114
rect 36990 46062 37042 46114
rect 40798 46062 40850 46114
rect 44606 45950 44658 46002
rect 7310 45838 7362 45890
rect 10558 45838 10610 45890
rect 12686 45838 12738 45890
rect 13134 45838 13186 45890
rect 13918 45810 13970 45862
rect 16158 45838 16210 45890
rect 17502 45838 17554 45890
rect 20078 45810 20130 45862
rect 20750 45838 20802 45890
rect 21534 45810 21586 45862
rect 24446 45838 24498 45890
rect 24782 45838 24834 45890
rect 26126 45838 26178 45890
rect 26238 45838 26290 45890
rect 26462 45838 26514 45890
rect 27918 45838 27970 45890
rect 28366 45838 28418 45890
rect 28702 45838 28754 45890
rect 29486 45838 29538 45890
rect 29710 45838 29762 45890
rect 30270 45838 30322 45890
rect 30494 45838 30546 45890
rect 30606 45838 30658 45890
rect 30942 45838 30994 45890
rect 32174 45810 32226 45862
rect 35030 45838 35082 45890
rect 35310 45838 35362 45890
rect 35534 45838 35586 45890
rect 35982 45810 36034 45862
rect 38670 45838 38722 45890
rect 38894 45838 38946 45890
rect 39790 45810 39842 45862
rect 42478 45838 42530 45890
rect 42702 45838 42754 45890
rect 43598 45810 43650 45862
rect 46286 45838 46338 45890
rect 46510 45838 46562 45890
rect 47350 45782 47402 45834
rect 48078 45800 48130 45852
rect 3110 45614 3162 45666
rect 3558 45614 3610 45666
rect 3894 45670 3946 45722
rect 4566 45614 4618 45666
rect 5014 45614 5066 45666
rect 5574 45670 5626 45722
rect 6246 45614 6298 45666
rect 6694 45614 6746 45666
rect 7030 45670 7082 45722
rect 7646 45614 7698 45666
rect 8262 45614 8314 45666
rect 8598 45670 8650 45722
rect 9830 45614 9882 45666
rect 10166 45670 10218 45722
rect 10894 45614 10946 45666
rect 11398 45670 11450 45722
rect 11846 45670 11898 45722
rect 21086 45726 21138 45778
rect 29206 45726 29258 45778
rect 29990 45726 30042 45778
rect 12350 45614 12402 45666
rect 13470 45614 13522 45666
rect 17166 45614 17218 45666
rect 25398 45670 25450 45722
rect 39174 45726 39226 45778
rect 42982 45726 43034 45778
rect 46790 45726 46842 45778
rect 47518 45726 47570 45778
rect 48190 45782 48242 45834
rect 26798 45614 26850 45666
rect 27582 45614 27634 45666
rect 31446 45670 31498 45722
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 2662 45166 2714 45218
rect 13022 45166 13074 45218
rect 24446 45166 24498 45218
rect 32398 45166 32450 45218
rect 5854 45054 5906 45106
rect 6190 45054 6242 45106
rect 6974 45054 7026 45106
rect 9550 45054 9602 45106
rect 9886 45069 9938 45121
rect 10334 45054 10386 45106
rect 11118 45054 11170 45106
rect 15486 45054 15538 45106
rect 16270 45054 16322 45106
rect 16942 45054 16994 45106
rect 20750 45054 20802 45106
rect 20974 45054 21026 45106
rect 21198 45054 21250 45106
rect 21758 45054 21810 45106
rect 25230 45054 25282 45106
rect 26014 45054 26066 45106
rect 28870 45054 28922 45106
rect 29038 45054 29090 45106
rect 29150 45054 29202 45106
rect 29710 45054 29762 45106
rect 33070 45054 33122 45106
rect 36262 45110 36314 45162
rect 36430 45110 36482 45162
rect 36654 45110 36706 45162
rect 37550 45054 37602 45106
rect 40854 45110 40906 45162
rect 41022 45084 41074 45136
rect 41246 45093 41298 45145
rect 42254 45054 42306 45106
rect 45390 45054 45442 45106
rect 46174 45054 46226 45106
rect 2214 44942 2266 44994
rect 3110 44942 3162 44994
rect 3558 44942 3610 44994
rect 4006 44942 4058 44994
rect 4454 44942 4506 44994
rect 4902 44942 4954 44994
rect 5350 44942 5402 44994
rect 8878 44942 8930 44994
rect 9998 44942 10050 44994
rect 13582 44942 13634 44994
rect 17670 44942 17722 44994
rect 18062 44942 18114 44994
rect 19966 44942 20018 44994
rect 22542 44942 22594 44994
rect 27918 44942 27970 44994
rect 30494 44942 30546 44994
rect 33854 44942 33906 44994
rect 35758 44942 35810 44994
rect 38334 44942 38386 44994
rect 40238 44942 40290 44994
rect 43038 44942 43090 44994
rect 44942 44942 44994 44994
rect 48078 44942 48130 44994
rect 5686 44830 5738 44882
rect 16606 44830 16658 44882
rect 21478 44830 21530 44882
rect 28478 44830 28530 44882
rect 37214 44830 37266 44882
rect 41806 44830 41858 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 6806 44494 6858 44546
rect 12686 44494 12738 44546
rect 22318 44494 22370 44546
rect 25006 44494 25058 44546
rect 26742 44494 26794 44546
rect 29542 44494 29594 44546
rect 37998 44494 38050 44546
rect 40910 44494 40962 44546
rect 45614 44494 45666 44546
rect 10670 44382 10722 44434
rect 14478 44382 14530 44434
rect 18510 44382 18562 44434
rect 25678 44382 25730 44434
rect 2270 44270 2322 44322
rect 3054 44270 3106 44322
rect 5966 44270 6018 44322
rect 6078 44270 6130 44322
rect 7086 44270 7138 44322
rect 7310 44270 7362 44322
rect 7590 44270 7642 44322
rect 7870 44270 7922 44322
rect 8094 44270 8146 44322
rect 8262 44326 8314 44378
rect 9102 44326 9154 44378
rect 8430 44270 8482 44322
rect 8990 44214 9042 44266
rect 9662 44270 9714 44322
rect 9998 44243 10050 44295
rect 10222 44270 10274 44322
rect 10782 44226 10834 44278
rect 11006 44270 11058 44322
rect 11790 44270 11842 44322
rect 13022 44270 13074 44322
rect 14142 44270 14194 44322
rect 14366 44226 14418 44278
rect 16830 44270 16882 44322
rect 17614 44270 17666 44322
rect 17726 44270 17778 44322
rect 21310 44242 21362 44294
rect 23998 44270 24050 44322
rect 24222 44270 24274 44322
rect 25342 44270 25394 44322
rect 25902 44270 25954 44322
rect 4958 44158 5010 44210
rect 6358 44158 6410 44210
rect 14926 44158 14978 44210
rect 9774 44102 9826 44154
rect 25510 44214 25562 44266
rect 20414 44158 20466 44210
rect 24502 44158 24554 44210
rect 26238 44214 26290 44266
rect 27022 44270 27074 44322
rect 27246 44270 27298 44322
rect 27918 44270 27970 44322
rect 28198 44270 28250 44322
rect 28478 44270 28530 44322
rect 28590 44270 28642 44322
rect 29150 44270 29202 44322
rect 29262 44270 29314 44322
rect 31614 44270 31666 44322
rect 32286 44270 32338 44322
rect 30737 44214 30789 44266
rect 34190 44242 34242 44294
rect 35553 44270 35605 44322
rect 36430 44270 36482 44322
rect 36990 44242 37042 44294
rect 39902 44242 39954 44294
rect 43262 44240 43314 44292
rect 43486 44231 43538 44283
rect 44270 44270 44322 44322
rect 2102 44046 2154 44098
rect 11622 44046 11674 44098
rect 12126 44046 12178 44098
rect 13526 44046 13578 44098
rect 27582 44046 27634 44098
rect 29990 44102 30042 44154
rect 30494 44158 30546 44210
rect 35310 44158 35362 44210
rect 42814 44158 42866 44210
rect 43766 44214 43818 44266
rect 47182 44242 47234 44294
rect 47518 44270 47570 44322
rect 47742 44270 47794 44322
rect 48022 44158 48074 44210
rect 44102 44046 44154 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 19294 43710 19346 43762
rect 4062 43598 4114 43650
rect 7086 43654 7138 43706
rect 6526 43598 6578 43650
rect 15598 43654 15650 43706
rect 8318 43598 8370 43650
rect 17670 43598 17722 43650
rect 4398 43486 4450 43538
rect 4734 43486 4786 43538
rect 4958 43501 5010 43553
rect 5406 43486 5458 43538
rect 6282 43486 6334 43538
rect 7198 43486 7250 43538
rect 7422 43525 7474 43577
rect 7758 43486 7810 43538
rect 8542 43486 8594 43538
rect 8766 43514 8818 43566
rect 9438 43486 9490 43538
rect 1878 43374 1930 43426
rect 2326 43374 2378 43426
rect 2774 43374 2826 43426
rect 3222 43374 3274 43426
rect 8150 43430 8202 43482
rect 9662 43486 9714 43538
rect 10222 43486 10274 43538
rect 11006 43486 11058 43538
rect 11882 43486 11934 43538
rect 12126 43486 12178 43538
rect 12574 43486 12626 43538
rect 13450 43486 13502 43538
rect 14254 43516 14306 43568
rect 14478 43525 14530 43577
rect 15038 43486 15090 43538
rect 14758 43430 14810 43482
rect 15934 43542 15986 43594
rect 38054 43654 38106 43706
rect 23102 43598 23154 43650
rect 23942 43598 23994 43650
rect 15710 43486 15762 43538
rect 16382 43486 16434 43538
rect 16886 43486 16938 43538
rect 17950 43513 18002 43565
rect 20862 43486 20914 43538
rect 21738 43486 21790 43538
rect 22654 43514 22706 43566
rect 22878 43486 22930 43538
rect 23270 43430 23322 43482
rect 23438 43486 23490 43538
rect 23662 43486 23714 43538
rect 24222 43486 24274 43538
rect 25454 43486 25506 43538
rect 25902 43486 25954 43538
rect 26778 43486 26830 43538
rect 27358 43486 27410 43538
rect 27694 43486 27746 43538
rect 28086 43542 28138 43594
rect 41022 43598 41074 43650
rect 28254 43516 28306 43568
rect 28478 43525 28530 43577
rect 45054 43598 45106 43650
rect 29934 43486 29986 43538
rect 30158 43486 30210 43538
rect 30494 43516 30546 43568
rect 30830 43516 30882 43568
rect 31278 43486 31330 43538
rect 30998 43430 31050 43482
rect 31726 43486 31778 43538
rect 31838 43486 31890 43538
rect 31984 43523 32036 43575
rect 33070 43486 33122 43538
rect 33742 43486 33794 43538
rect 34414 43486 34466 43538
rect 35534 43513 35586 43565
rect 37886 43486 37938 43538
rect 38558 43486 38610 43538
rect 38801 43486 38853 43538
rect 39678 43486 39730 43538
rect 41265 43542 41317 43594
rect 39902 43486 39954 43538
rect 42142 43486 42194 43538
rect 42702 43516 42754 43568
rect 43038 43516 43090 43568
rect 43486 43486 43538 43538
rect 3670 43374 3722 43426
rect 5070 43374 5122 43426
rect 9942 43374 9994 43426
rect 43206 43430 43258 43482
rect 43934 43486 43986 43538
rect 44810 43486 44862 43538
rect 45390 43486 45442 43538
rect 29654 43374 29706 43426
rect 34078 43374 34130 43426
rect 36206 43374 36258 43426
rect 46174 43374 46226 43426
rect 48078 43374 48130 43426
rect 10558 43262 10610 43314
rect 13694 43262 13746 43314
rect 21982 43262 22034 43314
rect 24558 43262 24610 43314
rect 25286 43262 25338 43314
rect 27022 43262 27074 43314
rect 29038 43262 29090 43314
rect 32398 43262 32450 43314
rect 34750 43262 34802 43314
rect 40238 43262 40290 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 5686 42926 5738 42978
rect 7086 42926 7138 42978
rect 14198 42926 14250 42978
rect 20638 42926 20690 42978
rect 26574 42926 26626 42978
rect 28478 42926 28530 42978
rect 32454 42926 32506 42978
rect 12462 42814 12514 42866
rect 15262 42814 15314 42866
rect 35870 42870 35922 42922
rect 43038 42926 43090 42978
rect 45838 42926 45890 42978
rect 21982 42814 22034 42866
rect 23550 42814 23602 42866
rect 25454 42814 25506 42866
rect 32062 42814 32114 42866
rect 35422 42814 35474 42866
rect 42254 42814 42306 42866
rect 1598 42702 1650 42754
rect 3614 42687 3666 42739
rect 3950 42702 4002 42754
rect 4286 42702 4338 42754
rect 4398 42702 4450 42754
rect 5966 42702 6018 42754
rect 6190 42702 6242 42754
rect 6414 42702 6466 42754
rect 6526 42702 6578 42754
rect 6692 42702 6744 42754
rect 7646 42702 7698 42754
rect 7870 42702 7922 42754
rect 9102 42702 9154 42754
rect 9886 42702 9938 42754
rect 12574 42687 12626 42739
rect 12910 42702 12962 42754
rect 13806 42702 13858 42754
rect 13918 42702 13970 42754
rect 15038 42702 15090 42754
rect 4678 42590 4730 42642
rect 8150 42590 8202 42642
rect 11790 42590 11842 42642
rect 14702 42646 14754 42698
rect 16158 42702 16210 42754
rect 16382 42702 16434 42754
rect 15430 42646 15482 42698
rect 15934 42646 15986 42698
rect 16550 42646 16602 42698
rect 17166 42702 17218 42754
rect 17390 42702 17442 42754
rect 17502 42702 17554 42754
rect 17726 42702 17778 42754
rect 18006 42702 18058 42754
rect 19182 42702 19234 42754
rect 19742 42702 19794 42754
rect 19966 42702 20018 42754
rect 20078 42702 20130 42754
rect 20246 42702 20298 42754
rect 21758 42702 21810 42754
rect 22150 42702 22202 42754
rect 22318 42702 22370 42754
rect 22766 42702 22818 42754
rect 21534 42646 21586 42698
rect 25902 42702 25954 42754
rect 26014 42702 26066 42754
rect 27358 42702 27410 42754
rect 28234 42702 28286 42754
rect 29710 42702 29762 42754
rect 26180 42646 26232 42698
rect 29934 42702 29986 42754
rect 31614 42702 31666 42754
rect 30810 42646 30862 42698
rect 31950 42687 32002 42739
rect 32286 42702 32338 42754
rect 32734 42702 32786 42754
rect 33518 42702 33570 42754
rect 35982 42702 36034 42754
rect 36206 42702 36258 42754
rect 36878 42702 36930 42754
rect 41582 42758 41634 42810
rect 42422 42758 42474 42810
rect 37102 42702 37154 42754
rect 40014 42702 40066 42754
rect 40798 42702 40850 42754
rect 41022 42702 41074 42754
rect 41694 42664 41746 42716
rect 43430 42646 43482 42698
rect 43710 42646 43762 42698
rect 43990 42646 44042 42698
rect 45054 42674 45106 42726
rect 47518 42702 47570 42754
rect 47742 42702 47794 42754
rect 16886 42590 16938 42642
rect 1934 42478 1986 42530
rect 2774 42478 2826 42530
rect 3222 42478 3274 42530
rect 3614 42534 3666 42586
rect 8934 42478 8986 42530
rect 18846 42478 18898 42530
rect 19574 42534 19626 42586
rect 31054 42590 31106 42642
rect 37382 42590 37434 42642
rect 38110 42590 38162 42642
rect 48022 42590 48074 42642
rect 22486 42478 22538 42530
rect 29374 42478 29426 42530
rect 41190 42478 41242 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 9662 42142 9714 42194
rect 34582 42142 34634 42194
rect 4846 42030 4898 42082
rect 10334 42086 10386 42138
rect 24558 42086 24610 42138
rect 40182 42142 40234 42194
rect 43990 42142 44042 42194
rect 7870 42030 7922 42082
rect 1598 41918 1650 41970
rect 4286 41918 4338 41970
rect 5089 41918 5141 41970
rect 5966 41918 6018 41970
rect 6302 41918 6354 41970
rect 6862 41918 6914 41970
rect 7702 41918 7754 41970
rect 8094 41918 8146 41970
rect 8318 41946 8370 41998
rect 8766 41918 8818 41970
rect 9998 41918 10050 41970
rect 10334 41918 10386 41970
rect 10670 41957 10722 42009
rect 10894 41918 10946 41970
rect 11790 41918 11842 41970
rect 12014 41918 12066 41970
rect 12462 41918 12514 41970
rect 13022 41918 13074 41970
rect 13898 41918 13950 41970
rect 14870 41918 14922 41970
rect 15150 41918 15202 41970
rect 15374 41918 15426 41970
rect 15598 41918 15650 41970
rect 15710 41918 15762 41970
rect 15896 41955 15948 42007
rect 17614 41918 17666 41970
rect 18398 41918 18450 41970
rect 20750 41918 20802 41970
rect 21626 41918 21678 41970
rect 21870 41918 21922 41970
rect 22430 41956 22482 42008
rect 22766 41918 22818 41970
rect 23774 41918 23826 41970
rect 24222 41957 24274 42009
rect 24446 41918 24498 41970
rect 2382 41806 2434 41858
rect 16270 41806 16322 41858
rect 7086 41750 7138 41802
rect 16886 41806 16938 41858
rect 20302 41806 20354 41858
rect 22990 41806 23042 41858
rect 23158 41862 23210 41914
rect 25230 41918 25282 41970
rect 26106 41918 26158 41970
rect 26686 41918 26738 41970
rect 27638 41974 27690 42026
rect 28590 42030 28642 42082
rect 37998 42030 38050 42082
rect 26910 41918 26962 41970
rect 27190 41918 27242 41970
rect 27806 41948 27858 42000
rect 28142 41948 28194 42000
rect 29150 41918 29202 41970
rect 29486 41918 29538 41970
rect 30158 41918 30210 41970
rect 31818 41974 31870 42026
rect 30942 41918 30994 41970
rect 32062 41918 32114 41970
rect 32958 41918 33010 41970
rect 33294 41918 33346 41970
rect 33966 41918 34018 41970
rect 36654 41974 36706 42026
rect 34302 41918 34354 41970
rect 34750 41918 34802 41970
rect 34974 41918 35026 41970
rect 35850 41918 35902 41970
rect 36990 41948 37042 42000
rect 38222 41918 38274 41970
rect 38446 41946 38498 41998
rect 39118 41974 39170 42026
rect 44326 41974 44378 42026
rect 44494 41974 44546 42026
rect 44830 41974 44882 42026
rect 39454 41918 39506 41970
rect 37158 41862 37210 41914
rect 8934 41694 8986 41746
rect 11510 41694 11562 41746
rect 12294 41694 12346 41746
rect 14142 41694 14194 41746
rect 26350 41694 26402 41746
rect 29598 41750 29650 41802
rect 36094 41806 36146 41858
rect 37438 41806 37490 41858
rect 37830 41862 37882 41914
rect 40350 41918 40402 41970
rect 40798 41918 40850 41970
rect 44158 41918 44210 41970
rect 45726 41945 45778 41997
rect 39678 41806 39730 41858
rect 39846 41862 39898 41914
rect 41582 41806 41634 41858
rect 43486 41806 43538 41858
rect 46734 41806 46786 41858
rect 30494 41694 30546 41746
rect 45278 41694 45330 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 2382 41358 2434 41410
rect 12014 41358 12066 41410
rect 14366 41358 14418 41410
rect 16046 41358 16098 41410
rect 19742 41358 19794 41410
rect 22206 41358 22258 41410
rect 22710 41358 22762 41410
rect 33070 41358 33122 41410
rect 35926 41358 35978 41410
rect 20414 41302 20466 41354
rect 1990 41246 2042 41298
rect 12462 41246 12514 41298
rect 24670 41246 24722 41298
rect 25454 41246 25506 41298
rect 28646 41246 28698 41298
rect 37662 41246 37714 41298
rect 41358 41246 41410 41298
rect 2718 41134 2770 41186
rect 3278 41134 3330 41186
rect 3614 41107 3666 41159
rect 3950 41134 4002 41186
rect 4510 41134 4562 41186
rect 4622 41134 4674 41186
rect 5518 41134 5570 41186
rect 6302 41134 6354 41186
rect 9886 41134 9938 41186
rect 4902 41022 4954 41074
rect 8206 41022 8258 41074
rect 3390 40966 3442 41018
rect 9009 41078 9061 41130
rect 10894 41134 10946 41186
rect 11770 41103 11822 41155
rect 12574 41090 12626 41142
rect 12798 41134 12850 41186
rect 8766 41022 8818 41074
rect 10614 41022 10666 41074
rect 13414 41078 13466 41130
rect 13582 41104 13634 41156
rect 14926 41134 14978 41186
rect 13918 41078 13970 41130
rect 16718 41134 16770 41186
rect 18622 41134 18674 41186
rect 19406 41134 19458 41186
rect 15802 41078 15854 41130
rect 20078 41134 20130 41186
rect 20414 41134 20466 41186
rect 20638 41134 20690 41186
rect 21254 41078 21306 41130
rect 21534 41095 21586 41147
rect 22990 41134 23042 41186
rect 21814 41078 21866 41130
rect 23214 41134 23266 41186
rect 23326 41134 23378 41186
rect 23550 41134 23602 41186
rect 23830 41134 23882 41186
rect 24782 41119 24834 41171
rect 25118 41134 25170 41186
rect 25566 41090 25618 41142
rect 25902 41134 25954 41186
rect 26574 41134 26626 41186
rect 29038 41134 29090 41186
rect 27450 41078 27502 41130
rect 29822 41134 29874 41186
rect 30698 41134 30750 41186
rect 30942 41134 30994 41186
rect 31390 41134 31442 41186
rect 32266 41134 32318 41186
rect 33406 41134 33458 41186
rect 34078 41134 34130 41186
rect 34750 41134 34802 41186
rect 35086 41134 35138 41186
rect 36206 41134 36258 41186
rect 37830 41190 37882 41242
rect 36318 41134 36370 41186
rect 37214 41106 37266 41158
rect 37438 41134 37490 41186
rect 38110 41134 38162 41186
rect 38894 41134 38946 41186
rect 41470 41119 41522 41171
rect 41806 41134 41858 41186
rect 42198 41134 42250 41186
rect 42478 41134 42530 41186
rect 42758 41190 42810 41242
rect 48078 41246 48130 41298
rect 42926 41134 42978 41186
rect 43206 41190 43258 41242
rect 43598 41134 43650 41186
rect 43934 41096 43986 41148
rect 45278 41134 45330 41186
rect 45390 41134 45442 41186
rect 46174 41134 46226 41186
rect 24278 40966 24330 41018
rect 27694 41022 27746 41074
rect 32510 41022 32562 41074
rect 40798 41022 40850 41074
rect 42590 41022 42642 41074
rect 43374 41022 43426 41074
rect 29374 40910 29426 40962
rect 33742 40910 33794 40962
rect 34414 40910 34466 40962
rect 35422 40910 35474 40962
rect 44942 40910 44994 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 2886 40574 2938 40626
rect 6638 40574 6690 40626
rect 9718 40574 9770 40626
rect 10166 40574 10218 40626
rect 15318 40574 15370 40626
rect 17614 40574 17666 40626
rect 1990 40462 2042 40514
rect 6246 40462 6298 40514
rect 7254 40462 7306 40514
rect 2438 40350 2490 40402
rect 3390 40406 3442 40458
rect 4174 40380 4226 40432
rect 4398 40406 4450 40458
rect 8878 40462 8930 40514
rect 4846 40350 4898 40402
rect 4006 40294 4058 40346
rect 5070 40350 5122 40402
rect 5350 40350 5402 40402
rect 6974 40350 7026 40402
rect 7534 40350 7586 40402
rect 7758 40350 7810 40402
rect 7926 40406 7978 40458
rect 8094 40406 8146 40458
rect 8318 40406 8370 40458
rect 16494 40518 16546 40570
rect 19798 40574 19850 40626
rect 24726 40574 24778 40626
rect 32286 40574 32338 40626
rect 14702 40462 14754 40514
rect 10614 40350 10666 40402
rect 10894 40350 10946 40402
rect 11230 40394 11282 40446
rect 11678 40350 11730 40402
rect 11790 40350 11842 40402
rect 11976 40388 12028 40440
rect 14458 40406 14510 40458
rect 18230 40462 18282 40514
rect 20918 40462 20970 40514
rect 28926 40462 28978 40514
rect 12798 40350 12850 40402
rect 13134 40350 13186 40402
rect 13582 40350 13634 40402
rect 15486 40350 15538 40402
rect 16046 40350 16098 40402
rect 16270 40389 16322 40441
rect 16606 40350 16658 40402
rect 17278 40350 17330 40402
rect 19294 40350 19346 40402
rect 20302 40350 20354 40402
rect 20414 40350 20466 40402
rect 20638 40350 20690 40402
rect 21310 40350 21362 40402
rect 21422 40350 21474 40402
rect 21590 40350 21642 40402
rect 22430 40350 22482 40402
rect 22542 40350 22594 40402
rect 22822 40350 22874 40402
rect 24222 40350 24274 40402
rect 25454 40350 25506 40402
rect 25566 40350 25618 40402
rect 25712 40387 25764 40439
rect 26462 40350 26514 40402
rect 26686 40350 26738 40402
rect 27526 40350 27578 40402
rect 28682 40406 28734 40458
rect 27806 40350 27858 40402
rect 30158 40406 30210 40458
rect 29766 40350 29818 40402
rect 30494 40380 30546 40432
rect 30662 40406 30714 40458
rect 30942 40462 30994 40514
rect 31278 40350 31330 40402
rect 31502 40350 31554 40402
rect 31782 40350 31834 40402
rect 32622 40350 32674 40402
rect 36206 40406 36258 40458
rect 32958 40350 33010 40402
rect 33742 40350 33794 40402
rect 35646 40350 35698 40402
rect 36430 40389 36482 40441
rect 36710 40406 36762 40458
rect 36990 40462 37042 40514
rect 42758 40462 42810 40514
rect 46398 40462 46450 40514
rect 37326 40350 37378 40402
rect 37550 40350 37602 40402
rect 37830 40350 37882 40402
rect 38334 40350 38386 40402
rect 38446 40350 38498 40402
rect 39454 40350 39506 40402
rect 39678 40350 39730 40402
rect 40238 40350 40290 40402
rect 40462 40350 40514 40402
rect 41246 40350 41298 40402
rect 41358 40350 41410 40402
rect 41526 40350 41578 40402
rect 42254 40350 42306 40402
rect 42478 40350 42530 40402
rect 43654 40406 43706 40458
rect 45370 40406 45422 40458
rect 43374 40350 43426 40402
rect 43486 40350 43538 40402
rect 44494 40350 44546 40402
rect 45614 40350 45666 40402
rect 46062 40350 46114 40402
rect 46230 40350 46282 40402
rect 46510 40350 46562 40402
rect 47742 40406 47794 40458
rect 47126 40350 47178 40402
rect 47518 40350 47570 40402
rect 11342 40238 11394 40290
rect 12350 40238 12402 40290
rect 3222 40126 3274 40178
rect 3726 40126 3778 40178
rect 13246 40182 13298 40234
rect 21982 40238 22034 40290
rect 23494 40238 23546 40290
rect 26126 40238 26178 40290
rect 26966 40238 27018 40290
rect 41918 40238 41970 40290
rect 47294 40238 47346 40290
rect 18958 40126 19010 40178
rect 20134 40126 20186 40178
rect 23886 40126 23938 40178
rect 38726 40126 38778 40178
rect 39174 40126 39226 40178
rect 39958 40126 40010 40178
rect 44046 40126 44098 40178
rect 46790 40126 46842 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 8094 39790 8146 39842
rect 10334 39790 10386 39842
rect 12854 39790 12906 39842
rect 16830 39790 16882 39842
rect 36206 39790 36258 39842
rect 32622 39734 32674 39786
rect 37718 39790 37770 39842
rect 4286 39678 4338 39730
rect 6302 39678 6354 39730
rect 16270 39678 16322 39730
rect 17558 39678 17610 39730
rect 18622 39678 18674 39730
rect 20526 39678 20578 39730
rect 23550 39678 23602 39730
rect 25454 39678 25506 39730
rect 28534 39678 28586 39730
rect 31390 39678 31442 39730
rect 1598 39566 1650 39618
rect 2382 39566 2434 39618
rect 5854 39538 5906 39590
rect 6078 39566 6130 39618
rect 6974 39566 7026 39618
rect 5126 39454 5178 39506
rect 6470 39510 6522 39562
rect 9998 39566 10050 39618
rect 7142 39510 7194 39562
rect 7422 39510 7474 39562
rect 7702 39510 7754 39562
rect 10782 39510 10834 39562
rect 11118 39510 11170 39562
rect 11286 39510 11338 39562
rect 12126 39566 12178 39618
rect 12294 39566 12346 39618
rect 12574 39566 12626 39618
rect 13526 39566 13578 39618
rect 13806 39566 13858 39618
rect 13918 39566 13970 39618
rect 14254 39566 14306 39618
rect 15934 39566 15986 39618
rect 17166 39566 17218 39618
rect 15130 39510 15182 39562
rect 12462 39454 12514 39506
rect 16102 39510 16154 39562
rect 17838 39566 17890 39618
rect 21310 39566 21362 39618
rect 22766 39566 22818 39618
rect 22186 39510 22238 39562
rect 26238 39566 26290 39618
rect 27358 39566 27410 39618
rect 15374 39454 15426 39506
rect 27114 39510 27166 39562
rect 28142 39566 28194 39618
rect 28254 39566 28306 39618
rect 29038 39566 29090 39618
rect 29710 39566 29762 39618
rect 30830 39566 30882 39618
rect 30586 39510 30638 39562
rect 31614 39566 31666 39618
rect 32398 39566 32450 39618
rect 32734 39566 32786 39618
rect 33070 39566 33122 39618
rect 31222 39510 31274 39562
rect 31782 39510 31834 39562
rect 33294 39566 33346 39618
rect 33574 39566 33626 39618
rect 34302 39566 34354 39618
rect 34526 39566 34578 39618
rect 35402 39566 35454 39618
rect 36542 39566 36594 39618
rect 36990 39566 37042 39618
rect 37158 39622 37210 39674
rect 37326 39566 37378 39618
rect 37438 39566 37490 39618
rect 38222 39566 38274 39618
rect 39006 39566 39058 39618
rect 41358 39566 41410 39618
rect 42142 39566 42194 39618
rect 45278 39566 45330 39618
rect 45390 39566 45442 39618
rect 46174 39566 46226 39618
rect 22430 39454 22482 39506
rect 6806 39342 6858 39394
rect 9046 39342 9098 39394
rect 9494 39342 9546 39394
rect 9830 39342 9882 39394
rect 11846 39342 11898 39394
rect 29206 39398 29258 39450
rect 35646 39454 35698 39506
rect 40910 39454 40962 39506
rect 44046 39454 44098 39506
rect 48078 39454 48130 39506
rect 34134 39342 34186 39394
rect 44942 39342 44994 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 2270 39006 2322 39058
rect 15598 39006 15650 39058
rect 16606 39006 16658 39058
rect 23494 39006 23546 39058
rect 4062 38894 4114 38946
rect 2606 38782 2658 38834
rect 3818 38838 3870 38890
rect 5182 38894 5234 38946
rect 22318 38950 22370 39002
rect 27750 39006 27802 39058
rect 24558 38950 24610 39002
rect 37606 39006 37658 39058
rect 2942 38782 2994 38834
rect 7086 38782 7138 38834
rect 7870 38782 7922 38834
rect 8094 38838 8146 38890
rect 14926 38894 14978 38946
rect 30718 38950 30770 39002
rect 39902 39006 39954 39058
rect 41134 39006 41186 39058
rect 26350 38894 26402 38946
rect 8206 38820 8258 38872
rect 8766 38782 8818 38834
rect 4678 38670 4730 38722
rect 8934 38726 8986 38778
rect 9438 38782 9490 38834
rect 12730 38820 12782 38872
rect 13470 38782 13522 38834
rect 14366 38820 14418 38872
rect 14702 38782 14754 38834
rect 15094 38726 15146 38778
rect 15934 38782 15986 38834
rect 16942 38782 16994 38834
rect 17502 38782 17554 38834
rect 20862 38782 20914 38834
rect 21086 38826 21138 38878
rect 21758 38782 21810 38834
rect 21982 38821 22034 38873
rect 24054 38838 24106 38890
rect 31390 38894 31442 38946
rect 22318 38782 22370 38834
rect 23774 38782 23826 38834
rect 24446 38782 24498 38834
rect 25230 38782 25282 38834
rect 26106 38813 26158 38865
rect 28906 38838 28958 38890
rect 26798 38782 26850 38834
rect 27134 38782 27186 38834
rect 28030 38782 28082 38834
rect 29150 38782 29202 38834
rect 31782 38838 31834 38890
rect 29934 38782 29986 38834
rect 30494 38782 30546 38834
rect 32174 38812 32226 38864
rect 32342 38838 32394 38890
rect 39230 38894 39282 38946
rect 33070 38782 33122 38834
rect 33946 38782 33998 38834
rect 34806 38782 34858 38834
rect 35086 38782 35138 38834
rect 35310 38782 35362 38834
rect 35534 38838 35586 38890
rect 35814 38838 35866 38890
rect 42422 38894 42474 38946
rect 36374 38782 36426 38834
rect 36542 38782 36594 38834
rect 36766 38782 36818 38834
rect 37886 38782 37938 38834
rect 37998 38782 38050 38834
rect 38144 38819 38196 38871
rect 38894 38782 38946 38834
rect 39566 38782 39618 38834
rect 40798 38782 40850 38834
rect 41507 38838 41559 38890
rect 41694 38838 41746 38890
rect 41918 38810 41970 38862
rect 42142 38838 42194 38890
rect 43150 38782 43202 38834
rect 43374 38782 43426 38834
rect 43878 38782 43930 38834
rect 44158 38810 44210 38862
rect 44382 38810 44434 38862
rect 44606 38838 44658 38890
rect 44718 38838 44770 38890
rect 45894 38894 45946 38946
rect 47462 38894 47514 38946
rect 45054 38838 45106 38890
rect 45166 38810 45218 38862
rect 45390 38810 45442 38862
rect 45614 38838 45666 38890
rect 46286 38782 46338 38834
rect 46398 38782 46450 38834
rect 46564 38782 46616 38834
rect 47742 38782 47794 38834
rect 47854 38782 47906 38834
rect 10222 38670 10274 38722
rect 12126 38670 12178 38722
rect 18286 38670 18338 38722
rect 20190 38670 20242 38722
rect 21198 38670 21250 38722
rect 22934 38670 22986 38722
rect 13582 38614 13634 38666
rect 27246 38614 27298 38666
rect 36206 38670 36258 38722
rect 38558 38670 38610 38722
rect 43486 38614 43538 38666
rect 46958 38670 47010 38722
rect 34190 38558 34242 38610
rect 37046 38558 37098 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 7870 38222 7922 38274
rect 2998 38110 3050 38162
rect 3446 38110 3498 38162
rect 8654 38166 8706 38218
rect 9774 38166 9826 38218
rect 6470 38110 6522 38162
rect 12126 38166 12178 38218
rect 12574 38166 12626 38218
rect 13862 38110 13914 38162
rect 14590 38166 14642 38218
rect 18622 38222 18674 38274
rect 22206 38222 22258 38274
rect 28478 38222 28530 38274
rect 31838 38222 31890 38274
rect 32342 38222 32394 38274
rect 34526 38222 34578 38274
rect 35310 38222 35362 38274
rect 35982 38222 36034 38274
rect 39342 38222 39394 38274
rect 39902 38222 39954 38274
rect 42086 38222 42138 38274
rect 22822 38110 22874 38162
rect 23214 38110 23266 38162
rect 24614 38110 24666 38162
rect 25174 38110 25226 38162
rect 43262 38166 43314 38218
rect 48078 38110 48130 38162
rect 2606 37998 2658 38050
rect 3782 37998 3834 38050
rect 4062 37998 4114 38050
rect 4286 37998 4338 38050
rect 4566 37998 4618 38050
rect 4846 37998 4898 38050
rect 4958 37998 5010 38050
rect 6750 37998 6802 38050
rect 7626 37967 7678 38019
rect 8430 37998 8482 38050
rect 8766 37998 8818 38050
rect 9438 37998 9490 38050
rect 9662 37998 9714 38050
rect 10110 37998 10162 38050
rect 11678 37998 11730 38050
rect 12014 37998 12066 38050
rect 12574 37998 12626 38050
rect 12798 37998 12850 38050
rect 14254 37998 14306 38050
rect 14478 37998 14530 38050
rect 14926 37998 14978 38050
rect 15802 37998 15854 38050
rect 16046 37998 16098 38050
rect 10986 37942 11038 37994
rect 16942 37998 16994 38050
rect 18958 37998 19010 38050
rect 23550 37998 23602 38050
rect 11230 37886 11282 37938
rect 19686 37886 19738 37938
rect 21254 37942 21306 37994
rect 21478 37942 21530 37994
rect 21646 37942 21698 37994
rect 23662 37998 23714 38050
rect 26238 37998 26290 38050
rect 26350 37998 26402 38050
rect 26574 37998 26626 38050
rect 26798 37998 26850 38050
rect 27526 37942 27578 37994
rect 27806 37942 27858 37994
rect 28030 37968 28082 38020
rect 29150 37998 29202 38050
rect 30026 37998 30078 38050
rect 30270 37998 30322 38050
rect 30718 37998 30770 38050
rect 32174 37998 32226 38050
rect 32622 37998 32674 38050
rect 34190 37998 34242 38050
rect 31594 37942 31646 37994
rect 34862 37998 34914 38050
rect 34974 37998 35026 38050
rect 35646 37998 35698 38050
rect 37438 37998 37490 38050
rect 37998 37998 38050 38050
rect 38110 37998 38162 38050
rect 38334 37942 38386 37994
rect 39006 37998 39058 38050
rect 40238 37998 40290 38050
rect 41134 37970 41186 38022
rect 25958 37886 26010 37938
rect 27078 37886 27130 37938
rect 37718 37886 37770 37938
rect 41358 37942 41410 37994
rect 41582 37942 41634 37994
rect 41694 37963 41746 38015
rect 42366 37970 42418 38022
rect 42590 37970 42642 38022
rect 42814 37970 42866 38022
rect 43374 37998 43426 38050
rect 43710 37998 43762 38050
rect 44214 37998 44266 38050
rect 42926 37942 42978 37994
rect 45278 37998 45330 38050
rect 45390 37998 45442 38050
rect 46174 37998 46226 38050
rect 40854 37886 40906 37938
rect 2270 37774 2322 37826
rect 5798 37774 5850 37826
rect 16606 37774 16658 37826
rect 17334 37774 17386 37826
rect 17782 37774 17834 37826
rect 18230 37774 18282 37826
rect 20134 37774 20186 37826
rect 20582 37774 20634 37826
rect 23998 37774 24050 37826
rect 25622 37774 25674 37826
rect 32790 37830 32842 37882
rect 33462 37774 33514 37826
rect 33854 37774 33906 37826
rect 37102 37774 37154 37826
rect 38670 37774 38722 37826
rect 44942 37774 44994 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 9046 37438 9098 37490
rect 14646 37438 14698 37490
rect 20246 37438 20298 37490
rect 30662 37438 30714 37490
rect 35646 37438 35698 37490
rect 41246 37438 41298 37490
rect 41918 37438 41970 37490
rect 43374 37438 43426 37490
rect 4846 37326 4898 37378
rect 1598 37214 1650 37266
rect 2382 37214 2434 37266
rect 4286 37214 4338 37266
rect 5089 37214 5141 37266
rect 5966 37214 6018 37266
rect 6246 37270 6298 37322
rect 7198 37326 7250 37378
rect 8038 37326 8090 37378
rect 6414 37244 6466 37296
rect 6750 37244 6802 37296
rect 7646 37214 7698 37266
rect 7758 37214 7810 37266
rect 9942 37270 9994 37322
rect 10110 37326 10162 37378
rect 12854 37326 12906 37378
rect 13358 37326 13410 37378
rect 10670 37270 10722 37322
rect 16382 37326 16434 37378
rect 10334 37214 10386 37266
rect 11678 37214 11730 37266
rect 12014 37229 12066 37281
rect 12350 37214 12402 37266
rect 12574 37214 12626 37266
rect 13582 37214 13634 37266
rect 13806 37242 13858 37294
rect 14478 37214 14530 37266
rect 16718 37214 16770 37266
rect 18286 37242 18338 37294
rect 18510 37214 18562 37266
rect 8598 37102 8650 37154
rect 9718 37102 9770 37154
rect 13190 37158 13242 37210
rect 11286 37102 11338 37154
rect 12126 37102 12178 37154
rect 15206 37102 15258 37154
rect 15990 37102 16042 37154
rect 17782 37102 17834 37154
rect 18734 37102 18786 37154
rect 18902 37158 18954 37210
rect 19070 37214 19122 37266
rect 21514 37270 21566 37322
rect 19294 37214 19346 37266
rect 20414 37214 20466 37266
rect 20638 37214 20690 37266
rect 21758 37214 21810 37266
rect 22318 37270 22370 37322
rect 25678 37326 25730 37378
rect 28366 37326 28418 37378
rect 35030 37326 35082 37378
rect 40238 37326 40290 37378
rect 22654 37214 22706 37266
rect 22878 37102 22930 37154
rect 23046 37158 23098 37210
rect 24222 37214 24274 37266
rect 26126 37244 26178 37296
rect 26462 37244 26514 37296
rect 27246 37214 27298 37266
rect 28122 37214 28174 37266
rect 30214 37214 30266 37266
rect 23494 37102 23546 37154
rect 23886 37102 23938 37154
rect 25958 37158 26010 37210
rect 31054 37214 31106 37266
rect 31930 37214 31982 37266
rect 32174 37214 32226 37266
rect 33070 37214 33122 37266
rect 33946 37214 33998 37266
rect 34190 37214 34242 37266
rect 34638 37214 34690 37266
rect 34750 37214 34802 37266
rect 35310 37214 35362 37266
rect 37048 37214 37100 37266
rect 37214 37214 37266 37266
rect 37326 37214 37378 37266
rect 37550 37214 37602 37266
rect 38334 37214 38386 37266
rect 41582 37214 41634 37266
rect 42254 37214 42306 37266
rect 42926 37214 42978 37266
rect 43710 37214 43762 37266
rect 44270 37229 44322 37281
rect 44606 37214 44658 37266
rect 45166 37214 45218 37266
rect 46230 37270 46282 37322
rect 45390 37214 45442 37266
rect 46398 37214 46450 37266
rect 46734 37214 46786 37266
rect 46958 37214 47010 37266
rect 47238 37214 47290 37266
rect 47518 37214 47570 37266
rect 47742 37214 47794 37266
rect 24726 37102 24778 37154
rect 28982 37102 29034 37154
rect 29766 37102 29818 37154
rect 36262 37102 36314 37154
rect 36654 37102 36706 37154
rect 44158 37102 44210 37154
rect 46062 37102 46114 37154
rect 19574 36990 19626 37042
rect 42590 36990 42642 37042
rect 45670 36990 45722 37042
rect 48022 36990 48074 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 10502 36654 10554 36706
rect 18846 36654 18898 36706
rect 4398 36542 4450 36594
rect 5798 36542 5850 36594
rect 6246 36542 6298 36594
rect 13582 36598 13634 36650
rect 22486 36654 22538 36706
rect 28478 36654 28530 36706
rect 20302 36598 20354 36650
rect 30382 36654 30434 36706
rect 32286 36654 32338 36706
rect 8150 36542 8202 36594
rect 12686 36542 12738 36594
rect 14422 36542 14474 36594
rect 16382 36542 16434 36594
rect 23662 36542 23714 36594
rect 25566 36542 25618 36594
rect 32846 36542 32898 36594
rect 34302 36598 34354 36650
rect 40294 36654 40346 36706
rect 41526 36654 41578 36706
rect 2606 36430 2658 36482
rect 3502 36430 3554 36482
rect 3614 36430 3666 36482
rect 3894 36430 3946 36482
rect 4230 36430 4282 36482
rect 4622 36430 4674 36482
rect 4958 36374 5010 36426
rect 6974 36430 7026 36482
rect 7254 36430 7306 36482
rect 7534 36430 7586 36482
rect 7758 36430 7810 36482
rect 8430 36430 8482 36482
rect 9550 36430 9602 36482
rect 9886 36430 9938 36482
rect 10782 36430 10834 36482
rect 9306 36374 9358 36426
rect 10894 36430 10946 36482
rect 11454 36430 11506 36482
rect 11790 36430 11842 36482
rect 12238 36430 12290 36482
rect 12574 36430 12626 36482
rect 13582 36430 13634 36482
rect 13806 36430 13858 36482
rect 15486 36430 15538 36482
rect 15598 36430 15650 36482
rect 19966 36430 20018 36482
rect 20414 36430 20466 36482
rect 20750 36430 20802 36482
rect 21366 36430 21418 36482
rect 21646 36430 21698 36482
rect 19089 36374 19141 36426
rect 21870 36430 21922 36482
rect 21982 36430 22034 36482
rect 22206 36430 22258 36482
rect 22878 36430 22930 36482
rect 32006 36486 32058 36538
rect 26014 36430 26066 36482
rect 26890 36430 26942 36482
rect 18286 36318 18338 36370
rect 27694 36374 27746 36426
rect 27918 36374 27970 36426
rect 28198 36374 28250 36426
rect 29262 36430 29314 36482
rect 30138 36430 30190 36482
rect 31502 36400 31554 36452
rect 33406 36430 33458 36482
rect 33518 36430 33570 36482
rect 33854 36430 33906 36482
rect 34190 36430 34242 36482
rect 35198 36430 35250 36482
rect 35366 36486 35418 36538
rect 42870 36542 42922 36594
rect 46174 36542 46226 36594
rect 31726 36374 31778 36426
rect 33240 36374 33292 36426
rect 35646 36430 35698 36482
rect 36878 36430 36930 36482
rect 37662 36430 37714 36482
rect 39566 36430 39618 36482
rect 40574 36402 40626 36454
rect 27134 36318 27186 36370
rect 34918 36318 34970 36370
rect 35534 36318 35586 36370
rect 40798 36374 40850 36426
rect 41022 36374 41074 36426
rect 41134 36395 41186 36447
rect 41806 36402 41858 36454
rect 42030 36402 42082 36454
rect 42254 36402 42306 36454
rect 42366 36374 42418 36426
rect 43486 36402 43538 36454
rect 35926 36318 35978 36370
rect 43710 36374 43762 36426
rect 43934 36374 43986 36426
rect 44046 36395 44098 36447
rect 44718 36430 44770 36482
rect 45390 36430 45442 36482
rect 43206 36318 43258 36370
rect 48078 36318 48130 36370
rect 2270 36206 2322 36258
rect 6638 36206 6690 36258
rect 10054 36206 10106 36258
rect 15150 36206 15202 36258
rect 31110 36206 31162 36258
rect 36486 36206 36538 36258
rect 45054 36206 45106 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 5910 35870 5962 35922
rect 21030 35870 21082 35922
rect 30438 35870 30490 35922
rect 32566 35870 32618 35922
rect 40294 35870 40346 35922
rect 5406 35758 5458 35810
rect 1598 35646 1650 35698
rect 2382 35646 2434 35698
rect 4846 35684 4898 35736
rect 5574 35702 5626 35754
rect 8878 35758 8930 35810
rect 5182 35646 5234 35698
rect 6078 35666 6130 35718
rect 6246 35672 6298 35724
rect 9494 35702 9546 35754
rect 10446 35758 10498 35810
rect 18454 35758 18506 35810
rect 19742 35758 19794 35810
rect 6974 35646 7026 35698
rect 9662 35676 9714 35728
rect 9886 35685 9938 35737
rect 11006 35646 11058 35698
rect 11882 35646 11934 35698
rect 12126 35646 12178 35698
rect 12574 35646 12626 35698
rect 13450 35646 13502 35698
rect 14030 35646 14082 35698
rect 14814 35646 14866 35698
rect 17838 35646 17890 35698
rect 17950 35646 18002 35698
rect 18174 35646 18226 35698
rect 18790 35702 18842 35754
rect 19014 35702 19066 35754
rect 26686 35758 26738 35810
rect 29038 35758 29090 35810
rect 33406 35814 33458 35866
rect 41806 35870 41858 35922
rect 42478 35870 42530 35922
rect 46286 35814 46338 35866
rect 31838 35758 31890 35810
rect 34582 35758 34634 35810
rect 35422 35758 35474 35810
rect 38614 35758 38666 35810
rect 44438 35758 44490 35810
rect 19182 35685 19234 35737
rect 20190 35646 20242 35698
rect 20470 35675 20522 35727
rect 20862 35646 20914 35698
rect 21758 35646 21810 35698
rect 25342 35676 25394 35728
rect 25678 35676 25730 35728
rect 26126 35646 26178 35698
rect 25846 35590 25898 35642
rect 26910 35646 26962 35698
rect 27134 35674 27186 35726
rect 27918 35646 27970 35698
rect 28794 35646 28846 35698
rect 30718 35646 30770 35698
rect 31594 35646 31646 35698
rect 33182 35646 33234 35698
rect 33854 35646 33906 35698
rect 26518 35590 26570 35642
rect 34078 35646 34130 35698
rect 34302 35646 34354 35698
rect 35870 35676 35922 35728
rect 36094 35684 36146 35736
rect 36374 35702 36426 35754
rect 36654 35646 36706 35698
rect 36766 35646 36818 35698
rect 37438 35646 37490 35698
rect 37550 35646 37602 35698
rect 37718 35646 37770 35698
rect 38894 35646 38946 35698
rect 39118 35646 39170 35698
rect 39342 35646 39394 35698
rect 39454 35646 39506 35698
rect 39734 35646 39786 35698
rect 40798 35646 40850 35698
rect 41470 35646 41522 35698
rect 42142 35646 42194 35698
rect 43374 35646 43426 35698
rect 44046 35646 44098 35698
rect 44718 35646 44770 35698
rect 44830 35646 44882 35698
rect 45390 35702 45442 35754
rect 45166 35646 45218 35698
rect 46286 35646 46338 35698
rect 46622 35685 46674 35737
rect 46846 35646 46898 35698
rect 47406 35646 47458 35698
rect 47742 35690 47794 35742
rect 4286 35534 4338 35586
rect 13694 35534 13746 35586
rect 16718 35534 16770 35586
rect 20638 35534 20690 35586
rect 21590 35534 21642 35586
rect 22542 35534 22594 35586
rect 24446 35534 24498 35586
rect 29990 35534 30042 35586
rect 38110 35534 38162 35586
rect 43710 35534 43762 35586
rect 47854 35534 47906 35586
rect 17502 35422 17554 35474
rect 37046 35422 37098 35474
rect 41134 35422 41186 35474
rect 43038 35422 43090 35474
rect 45670 35422 45722 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 2662 35086 2714 35138
rect 8150 35086 8202 35138
rect 12798 35086 12850 35138
rect 15150 35086 15202 35138
rect 19630 35086 19682 35138
rect 6694 34974 6746 35026
rect 7086 34974 7138 35026
rect 21646 35030 21698 35082
rect 23326 35086 23378 35138
rect 28478 35086 28530 35138
rect 30270 35086 30322 35138
rect 32734 35086 32786 35138
rect 42422 35086 42474 35138
rect 45726 35086 45778 35138
rect 46398 35086 46450 35138
rect 48134 35086 48186 35138
rect 37662 34974 37714 35026
rect 2942 34862 2994 34914
rect 3166 34862 3218 34914
rect 3390 34862 3442 34914
rect 4266 34862 4318 34914
rect 4510 34862 4562 34914
rect 5182 34862 5234 34914
rect 5966 34862 6018 34914
rect 6190 34862 6242 34914
rect 7310 34862 7362 34914
rect 8430 34862 8482 34914
rect 6918 34806 6970 34858
rect 7534 34806 7586 34858
rect 8654 34862 8706 34914
rect 9214 34862 9266 34914
rect 9457 34862 9509 34914
rect 10334 34862 10386 34914
rect 10782 34862 10834 34914
rect 12518 34918 12570 34970
rect 11006 34862 11058 34914
rect 14030 34862 14082 34914
rect 12014 34806 12066 34858
rect 12350 34806 12402 34858
rect 16046 34862 16098 34914
rect 14906 34806 14958 34858
rect 16270 34862 16322 34914
rect 16494 34862 16546 34914
rect 19070 34862 19122 34914
rect 17222 34806 17274 34858
rect 17502 34806 17554 34858
rect 17782 34806 17834 34858
rect 19294 34862 19346 34914
rect 20750 34862 20802 34914
rect 21758 34862 21810 34914
rect 21982 34862 22034 34914
rect 22878 34862 22930 34914
rect 5686 34750 5738 34802
rect 11286 34750 11338 34802
rect 16774 34750 16826 34802
rect 19873 34806 19925 34858
rect 26910 34918 26962 34970
rect 22990 34862 23042 34914
rect 24334 34862 24386 34914
rect 24558 34862 24610 34914
rect 37830 34918 37882 34970
rect 38278 34974 38330 35026
rect 39230 34974 39282 35026
rect 41134 34974 41186 35026
rect 44942 34974 44994 35026
rect 25434 34831 25486 34883
rect 18174 34750 18226 34802
rect 18790 34750 18842 34802
rect 25678 34750 25730 34802
rect 26070 34806 26122 34858
rect 26238 34750 26290 34802
rect 26798 34806 26850 34858
rect 27526 34806 27578 34858
rect 27806 34806 27858 34858
rect 28030 34832 28082 34884
rect 29150 34862 29202 34914
rect 30026 34862 30078 34914
rect 33070 34862 33122 34914
rect 33854 34862 33906 34914
rect 35758 34862 35810 34914
rect 36094 34862 36146 34914
rect 31558 34750 31610 34802
rect 31782 34806 31834 34858
rect 31950 34806 32002 34858
rect 32286 34806 32338 34858
rect 36990 34806 37042 34858
rect 37102 34806 37154 34858
rect 38446 34862 38498 34914
rect 41526 34846 41578 34898
rect 41694 34834 41746 34886
rect 41918 34834 41970 34886
rect 42142 34834 42194 34886
rect 42926 34862 42978 34914
rect 43150 34862 43202 34914
rect 43430 34862 43482 34914
rect 43710 34862 43762 34914
rect 45278 34862 45330 34914
rect 45390 34862 45442 34914
rect 46062 34862 46114 34914
rect 47294 34862 47346 34914
rect 47518 34862 47570 34914
rect 47630 34862 47682 34914
rect 47854 34862 47906 34914
rect 47014 34750 47066 34802
rect 5014 34638 5066 34690
rect 13750 34638 13802 34690
rect 15710 34638 15762 34690
rect 22542 34638 22594 34690
rect 24166 34638 24218 34690
rect 31110 34638 31162 34690
rect 36262 34638 36314 34690
rect 44046 34638 44098 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 8094 34302 8146 34354
rect 9662 34302 9714 34354
rect 36990 34302 37042 34354
rect 41806 34302 41858 34354
rect 4846 34190 4898 34242
rect 3894 34134 3946 34186
rect 4062 34134 4114 34186
rect 4286 34134 4338 34186
rect 5574 34134 5626 34186
rect 5742 34190 5794 34242
rect 7142 34190 7194 34242
rect 10894 34190 10946 34242
rect 12966 34190 13018 34242
rect 14646 34190 14698 34242
rect 6302 34134 6354 34186
rect 22598 34190 22650 34242
rect 5966 34078 6018 34130
rect 6638 34078 6690 34130
rect 6862 34078 6914 34130
rect 8430 34078 8482 34130
rect 9102 34078 9154 34130
rect 9998 34078 10050 34130
rect 10334 34116 10386 34168
rect 11342 34078 11394 34130
rect 12462 34078 12514 34130
rect 3670 33966 3722 34018
rect 10222 34022 10274 34074
rect 11062 34022 11114 34074
rect 12686 34078 12738 34130
rect 13918 34078 13970 34130
rect 14254 34078 14306 34130
rect 14366 34078 14418 34130
rect 7702 33966 7754 34018
rect 13638 33966 13690 34018
rect 14086 34022 14138 34074
rect 14926 34078 14978 34130
rect 15150 34078 15202 34130
rect 16942 34078 16994 34130
rect 17278 34078 17330 34130
rect 18062 34078 18114 34130
rect 19966 34105 20018 34157
rect 20582 34094 20634 34146
rect 20750 34134 20802 34186
rect 20974 34106 21026 34158
rect 21198 34134 21250 34186
rect 28366 34190 28418 34242
rect 30326 34190 30378 34242
rect 46398 34246 46450 34298
rect 45278 34190 45330 34242
rect 21478 34078 21530 34130
rect 21870 34078 21922 34130
rect 22206 34078 22258 34130
rect 22318 34078 22370 34130
rect 22038 34022 22090 34074
rect 23662 34078 23714 34130
rect 23774 34078 23826 34130
rect 23998 34078 24050 34130
rect 25678 34078 25730 34130
rect 26014 34078 26066 34130
rect 26518 34078 26570 34130
rect 26798 34078 26850 34130
rect 26910 34078 26962 34130
rect 27246 34078 27298 34130
rect 28122 34078 28174 34130
rect 29598 34078 29650 34130
rect 29766 34078 29818 34130
rect 29934 34078 29986 34130
rect 30046 34078 30098 34130
rect 30718 34078 30770 34130
rect 31594 34078 31646 34130
rect 31838 34078 31890 34130
rect 33946 34134 33998 34186
rect 33070 34078 33122 34130
rect 34526 34078 34578 34130
rect 35665 34078 35717 34130
rect 36542 34078 36594 34130
rect 37326 34078 37378 34130
rect 37438 34078 37490 34130
rect 38950 34078 39002 34130
rect 39230 34078 39282 34130
rect 39454 34078 39506 34130
rect 39678 34078 39730 34130
rect 39790 34078 39842 34130
rect 40070 34078 40122 34130
rect 40798 34078 40850 34130
rect 41470 34078 41522 34130
rect 42590 34078 42642 34130
rect 43374 34078 43426 34130
rect 46510 34078 46562 34130
rect 46846 34105 46898 34157
rect 47182 34078 47234 34130
rect 47630 34122 47682 34174
rect 47854 34078 47906 34130
rect 25398 33966 25450 34018
rect 28982 33966 29034 34018
rect 8766 33854 8818 33906
rect 15430 33854 15482 33906
rect 17446 33854 17498 33906
rect 25902 33910 25954 33962
rect 32566 33966 32618 34018
rect 42422 33966 42474 34018
rect 45894 33966 45946 34018
rect 47518 33966 47570 34018
rect 23326 33854 23378 33906
rect 24278 33854 24330 33906
rect 34190 33854 34242 33906
rect 34862 33854 34914 33906
rect 35422 33854 35474 33906
rect 41134 33854 41186 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 12854 33518 12906 33570
rect 15822 33462 15874 33514
rect 27358 33518 27410 33570
rect 29654 33518 29706 33570
rect 31166 33518 31218 33570
rect 9998 33406 10050 33458
rect 13582 33406 13634 33458
rect 16942 33406 16994 33458
rect 1598 33294 1650 33346
rect 2382 33294 2434 33346
rect 5126 33294 5178 33346
rect 4286 33182 4338 33234
rect 6078 33238 6130 33290
rect 6190 33294 6242 33346
rect 6974 33294 7026 33346
rect 9214 33294 9266 33346
rect 12462 33294 12514 33346
rect 16270 33350 16322 33402
rect 18510 33406 18562 33458
rect 19742 33406 19794 33458
rect 22542 33406 22594 33458
rect 25006 33406 25058 33458
rect 26966 33406 27018 33458
rect 32454 33462 32506 33514
rect 34190 33518 34242 33570
rect 34694 33518 34746 33570
rect 42310 33518 42362 33570
rect 43486 33462 43538 33514
rect 43934 33462 43986 33514
rect 38894 33406 38946 33458
rect 40798 33406 40850 33458
rect 48078 33406 48130 33458
rect 12574 33294 12626 33346
rect 13650 33254 13702 33306
rect 13806 33257 13858 33309
rect 8878 33182 8930 33234
rect 14254 33238 14306 33290
rect 14590 33261 14642 33313
rect 15034 33256 15086 33308
rect 15710 33294 15762 33346
rect 16494 33238 16546 33290
rect 17110 33238 17162 33290
rect 17390 33294 17442 33346
rect 18266 33263 18318 33315
rect 19406 33294 19458 33346
rect 19630 33255 19682 33307
rect 20078 33294 20130 33346
rect 21534 33294 21586 33346
rect 21758 33294 21810 33346
rect 25230 33294 25282 33346
rect 11902 33182 11954 33234
rect 5910 33070 5962 33122
rect 20806 33070 20858 33122
rect 21366 33126 21418 33178
rect 24446 33182 24498 33234
rect 24838 33238 24890 33290
rect 25454 33266 25506 33318
rect 29262 33294 29314 33346
rect 27638 33238 27690 33290
rect 27918 33238 27970 33290
rect 28142 33238 28194 33290
rect 29374 33294 29426 33346
rect 30046 33294 30098 33346
rect 30922 33294 30974 33346
rect 31502 33294 31554 33346
rect 31726 33294 31778 33346
rect 32286 33238 32338 33290
rect 33070 33294 33122 33346
rect 33946 33294 33998 33346
rect 34974 33294 35026 33346
rect 35198 33294 35250 33346
rect 36318 33294 36370 33346
rect 32006 33182 32058 33234
rect 35366 33238 35418 33290
rect 35534 33238 35586 33290
rect 35870 33238 35922 33290
rect 36934 33294 36986 33346
rect 37326 33294 37378 33346
rect 37102 33182 37154 33234
rect 37662 33238 37714 33290
rect 38110 33294 38162 33346
rect 41806 33294 41858 33346
rect 41918 33294 41970 33346
rect 42590 33294 42642 33346
rect 42702 33294 42754 33346
rect 43150 33294 43202 33346
rect 43374 33294 43426 33346
rect 43934 33294 43986 33346
rect 44158 33294 44210 33346
rect 44718 33294 44770 33346
rect 45390 33294 45442 33346
rect 46174 33294 46226 33346
rect 41526 33182 41578 33234
rect 26294 33070 26346 33122
rect 45054 33070 45106 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 2270 32734 2322 32786
rect 3222 32734 3274 32786
rect 3670 32734 3722 32786
rect 4118 32734 4170 32786
rect 7198 32734 7250 32786
rect 9774 32734 9826 32786
rect 7870 32678 7922 32730
rect 12798 32734 12850 32786
rect 10782 32678 10834 32730
rect 32566 32734 32618 32786
rect 37438 32734 37490 32786
rect 40126 32734 40178 32786
rect 15150 32622 15202 32674
rect 2606 32510 2658 32562
rect 4398 32510 4450 32562
rect 5274 32510 5326 32562
rect 5966 32510 6018 32562
rect 6078 32510 6130 32562
rect 6244 32510 6296 32562
rect 7534 32510 7586 32562
rect 7870 32510 7922 32562
rect 8094 32537 8146 32589
rect 8430 32510 8482 32562
rect 9438 32510 9490 32562
rect 10334 32510 10386 32562
rect 10894 32510 10946 32562
rect 11678 32537 11730 32589
rect 14366 32566 14418 32618
rect 17502 32622 17554 32674
rect 14590 32549 14642 32601
rect 15953 32566 16005 32618
rect 21198 32622 21250 32674
rect 22710 32622 22762 32674
rect 23550 32622 23602 32674
rect 16830 32510 16882 32562
rect 18062 32549 18114 32601
rect 18286 32566 18338 32618
rect 19406 32566 19458 32618
rect 20190 32566 20242 32618
rect 21870 32566 21922 32618
rect 30382 32622 30434 32674
rect 18622 32510 18674 32562
rect 20750 32510 20802 32562
rect 22990 32510 23042 32562
rect 14870 32454 14922 32506
rect 17782 32454 17834 32506
rect 23214 32510 23266 32562
rect 23793 32541 23845 32593
rect 24670 32510 24722 32562
rect 25342 32510 25394 32562
rect 28814 32510 28866 32562
rect 29038 32510 29090 32562
rect 30138 32566 30190 32618
rect 33182 32622 33234 32674
rect 29262 32510 29314 32562
rect 30942 32510 30994 32562
rect 31166 32510 31218 32562
rect 35086 32510 35138 32562
rect 35870 32510 35922 32562
rect 36430 32537 36482 32589
rect 38894 32510 38946 32562
rect 39006 32510 39058 32562
rect 39174 32510 39226 32562
rect 40462 32510 40514 32562
rect 40854 32526 40906 32578
rect 41022 32566 41074 32618
rect 41246 32566 41298 32618
rect 41470 32566 41522 32618
rect 41750 32510 41802 32562
rect 44158 32510 44210 32562
rect 44942 32510 44994 32562
rect 46490 32566 46542 32618
rect 47294 32566 47346 32618
rect 45614 32510 45666 32562
rect 48022 32566 48074 32618
rect 47630 32510 47682 32562
rect 5518 32286 5570 32338
rect 6638 32286 6690 32338
rect 15710 32286 15762 32338
rect 18790 32342 18842 32394
rect 22374 32398 22426 32450
rect 26126 32398 26178 32450
rect 28030 32398 28082 32450
rect 30830 32342 30882 32394
rect 32118 32398 32170 32450
rect 39566 32398 39618 32450
rect 42254 32398 42306 32450
rect 45334 32398 45386 32450
rect 47854 32398 47906 32450
rect 28534 32286 28586 32338
rect 46734 32286 46786 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 4846 31950 4898 32002
rect 7086 31950 7138 32002
rect 13582 31950 13634 32002
rect 22542 31950 22594 32002
rect 26686 31950 26738 32002
rect 29542 31950 29594 32002
rect 31166 31950 31218 32002
rect 38558 31950 38610 32002
rect 43878 31950 43930 32002
rect 8094 31838 8146 31890
rect 9270 31838 9322 31890
rect 2606 31726 2658 31778
rect 2942 31726 2994 31778
rect 3614 31726 3666 31778
rect 3278 31670 3330 31722
rect 4174 31726 4226 31778
rect 4286 31726 4338 31778
rect 5630 31726 5682 31778
rect 6190 31726 6242 31778
rect 7422 31726 7474 31778
rect 7758 31726 7810 31778
rect 4454 31670 4506 31722
rect 7982 31711 8034 31763
rect 8318 31726 8370 31778
rect 8542 31726 8594 31778
rect 9550 31726 9602 31778
rect 9774 31726 9826 31778
rect 10502 31670 10554 31722
rect 10782 31670 10834 31722
rect 11062 31670 11114 31722
rect 11342 31726 11394 31778
rect 14142 31726 14194 31778
rect 14254 31726 14306 31778
rect 14478 31726 14530 31778
rect 15878 31726 15930 31778
rect 12218 31670 12270 31722
rect 8822 31614 8874 31666
rect 10110 31614 10162 31666
rect 13976 31670 14028 31722
rect 16494 31726 16546 31778
rect 17782 31782 17834 31834
rect 21982 31838 22034 31890
rect 26294 31838 26346 31890
rect 33350 31838 33402 31890
rect 37158 31838 37210 31890
rect 41582 31838 41634 31890
rect 48078 31838 48130 31890
rect 16606 31726 16658 31778
rect 17390 31726 17442 31778
rect 17166 31670 17218 31722
rect 18622 31698 18674 31750
rect 20526 31726 20578 31778
rect 21310 31726 21362 31778
rect 21422 31726 21474 31778
rect 22878 31726 22930 31778
rect 21588 31670 21640 31722
rect 3054 31558 3106 31610
rect 6302 31558 6354 31610
rect 12462 31614 12514 31666
rect 16214 31614 16266 31666
rect 17614 31614 17666 31666
rect 23998 31614 24050 31666
rect 24278 31670 24330 31722
rect 24558 31687 24610 31739
rect 25118 31726 25170 31778
rect 27022 31726 27074 31778
rect 24782 31670 24834 31722
rect 27246 31726 27298 31778
rect 28122 31726 28174 31778
rect 28366 31726 28418 31778
rect 29038 31726 29090 31778
rect 29262 31726 29314 31778
rect 31614 31726 31666 31778
rect 30214 31670 30266 31722
rect 30438 31670 30490 31722
rect 30606 31670 30658 31722
rect 31838 31726 31890 31778
rect 33070 31726 33122 31778
rect 33630 31726 33682 31778
rect 33742 31726 33794 31778
rect 33966 31726 34018 31778
rect 35198 31726 35250 31778
rect 36074 31726 36126 31778
rect 37550 31698 37602 31750
rect 32118 31614 32170 31666
rect 2270 31502 2322 31554
rect 23606 31502 23658 31554
rect 25286 31502 25338 31554
rect 25846 31502 25898 31554
rect 32902 31558 32954 31610
rect 36318 31614 36370 31666
rect 40686 31670 40738 31722
rect 40910 31698 40962 31750
rect 41134 31698 41186 31750
rect 41246 31691 41298 31743
rect 41694 31682 41746 31734
rect 42030 31726 42082 31778
rect 42254 31726 42306 31778
rect 43038 31691 43090 31743
rect 43150 31698 43202 31750
rect 43374 31698 43426 31750
rect 43598 31698 43650 31750
rect 44718 31726 44770 31778
rect 45390 31726 45442 31778
rect 46174 31726 46226 31778
rect 40406 31614 40458 31666
rect 42590 31502 42642 31554
rect 45054 31502 45106 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 11062 31166 11114 31218
rect 26294 31166 26346 31218
rect 26742 31166 26794 31218
rect 5126 31054 5178 31106
rect 7814 31054 7866 31106
rect 1598 30942 1650 30994
rect 2382 30942 2434 30994
rect 4286 30942 4338 30994
rect 4734 30942 4786 30994
rect 4846 30942 4898 30994
rect 6190 30942 6242 30994
rect 6414 30942 6466 30994
rect 6582 30998 6634 31050
rect 6750 30942 6802 30994
rect 6974 30942 7026 30994
rect 7310 30980 7362 31032
rect 8094 30942 8146 30994
rect 8206 30942 8258 30994
rect 8430 30942 8482 30994
rect 9494 30998 9546 31050
rect 10446 31054 10498 31106
rect 21254 31054 21306 31106
rect 27806 31054 27858 31106
rect 35758 31054 35810 31106
rect 9662 30972 9714 31024
rect 9886 30981 9938 31033
rect 11454 30969 11506 31021
rect 13358 30942 13410 30994
rect 14142 30942 14194 30994
rect 15018 30942 15070 30994
rect 16158 30942 16210 30994
rect 16718 30942 16770 30994
rect 16830 30942 16882 30994
rect 17670 30942 17722 30994
rect 17950 30942 18002 30994
rect 18286 30986 18338 31038
rect 18622 30942 18674 30994
rect 20414 30942 20466 30994
rect 20526 30942 20578 30994
rect 20750 30942 20802 30994
rect 20974 30942 21026 30994
rect 21758 30942 21810 30994
rect 21982 30942 22034 30994
rect 22318 30942 22370 30994
rect 22542 30942 22594 30994
rect 23214 30942 23266 30994
rect 23550 30942 23602 30994
rect 23886 30942 23938 30994
rect 24278 30942 24330 30994
rect 24558 30942 24610 30994
rect 24670 30942 24722 30994
rect 25286 30942 25338 30994
rect 25566 30942 25618 30994
rect 25678 30942 25730 30994
rect 26910 30942 26962 30994
rect 28030 30942 28082 30994
rect 28366 30980 28418 31032
rect 30474 30998 30526 31050
rect 29374 30942 29426 30994
rect 29598 30942 29650 30994
rect 27638 30886 27690 30938
rect 30718 30942 30770 30994
rect 31166 30942 31218 30994
rect 32042 30942 32094 30994
rect 32286 30942 32338 30994
rect 33946 30998 33998 31050
rect 40238 31054 40290 31106
rect 41022 31054 41074 31106
rect 48078 31054 48130 31106
rect 33070 30942 33122 30994
rect 34190 30942 34242 30994
rect 34638 30942 34690 30994
rect 35514 30942 35566 30994
rect 36542 30942 36594 30994
rect 36654 30942 36706 30994
rect 36840 30980 36892 31032
rect 37550 30942 37602 30994
rect 42926 30942 42978 30994
rect 43710 30942 43762 30994
rect 44046 30942 44098 30994
rect 44718 30942 44770 30994
rect 45222 30942 45274 30994
rect 45390 30942 45442 30994
rect 5910 30830 5962 30882
rect 18398 30830 18450 30882
rect 20134 30830 20186 30882
rect 8766 30718 8818 30770
rect 15262 30718 15314 30770
rect 22094 30774 22146 30826
rect 15822 30718 15874 30770
rect 16438 30718 16490 30770
rect 23774 30774 23826 30826
rect 22878 30718 22930 30770
rect 27246 30718 27298 30770
rect 29206 30774 29258 30826
rect 37214 30830 37266 30882
rect 38334 30830 38386 30882
rect 46174 30830 46226 30882
rect 43934 30774 43986 30826
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 10110 30382 10162 30434
rect 10894 30326 10946 30378
rect 11790 30382 11842 30434
rect 14590 30382 14642 30434
rect 19126 30382 19178 30434
rect 29542 30382 29594 30434
rect 3166 30270 3218 30322
rect 6302 30270 6354 30322
rect 27918 30326 27970 30378
rect 30606 30326 30658 30378
rect 15822 30270 15874 30322
rect 17726 30270 17778 30322
rect 18342 30270 18394 30322
rect 23326 30270 23378 30322
rect 45670 30382 45722 30434
rect 30942 30326 30994 30378
rect 33406 30326 33458 30378
rect 34526 30326 34578 30378
rect 41022 30270 41074 30322
rect 44830 30270 44882 30322
rect 46398 30270 46450 30322
rect 47630 30270 47682 30322
rect 2830 30158 2882 30210
rect 3054 30143 3106 30195
rect 3502 30158 3554 30210
rect 4378 30158 4430 30210
rect 5518 30158 5570 30210
rect 8206 30158 8258 30210
rect 8990 30158 9042 30210
rect 11006 30158 11058 30210
rect 11342 30158 11394 30210
rect 12910 30158 12962 30210
rect 4622 30046 4674 30098
rect 9158 30102 9210 30154
rect 9326 30102 9378 30154
rect 9550 30102 9602 30154
rect 12033 30102 12085 30154
rect 13470 30158 13522 30210
rect 14346 30158 14398 30210
rect 15038 30158 15090 30210
rect 18734 30158 18786 30210
rect 18846 30158 18898 30210
rect 19518 30125 19570 30177
rect 19798 30102 19850 30154
rect 20414 30102 20466 30154
rect 20570 30118 20622 30170
rect 20750 30046 20802 30098
rect 21254 30102 21306 30154
rect 21422 30158 21474 30210
rect 21646 30158 21698 30210
rect 22542 30158 22594 30210
rect 21870 30102 21922 30154
rect 25678 30158 25730 30210
rect 26798 30158 26850 30210
rect 27918 30158 27970 30210
rect 28254 30158 28306 30210
rect 29150 30158 29202 30210
rect 26554 30102 26606 30154
rect 29262 30158 29314 30210
rect 30158 30158 30210 30210
rect 30494 30158 30546 30210
rect 31054 30158 31106 30210
rect 31278 30158 31330 30210
rect 32006 30102 32058 30154
rect 32174 30128 32226 30180
rect 32398 30119 32450 30171
rect 33630 30158 33682 30210
rect 34190 30158 34242 30210
rect 34638 30158 34690 30210
rect 35314 30120 35366 30172
rect 35814 30158 35866 30210
rect 36206 30158 36258 30210
rect 36542 30158 36594 30210
rect 38502 30158 38554 30210
rect 25230 30046 25282 30098
rect 32958 30046 33010 30098
rect 37102 30046 37154 30098
rect 37382 30102 37434 30154
rect 37550 30102 37602 30154
rect 37886 30102 37938 30154
rect 38950 30158 39002 30210
rect 39230 30158 39282 30210
rect 39342 30158 39394 30210
rect 39678 30158 39730 30210
rect 39510 30102 39562 30154
rect 40238 30130 40290 30182
rect 43038 30158 43090 30210
rect 43486 30119 43538 30171
rect 43710 30158 43762 30210
rect 44942 30143 44994 30195
rect 45166 30158 45218 30210
rect 45950 30158 46002 30210
rect 46062 30158 46114 30210
rect 46510 30143 46562 30195
rect 46846 30158 46898 30210
rect 47182 30158 47234 30210
rect 47518 30143 47570 30195
rect 8822 29934 8874 29986
rect 43598 29990 43650 30042
rect 27414 29934 27466 29986
rect 48134 29934 48186 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 2102 29598 2154 29650
rect 2494 29486 2546 29538
rect 5350 29542 5402 29594
rect 7478 29598 7530 29650
rect 23830 29598 23882 29650
rect 30550 29598 30602 29650
rect 32566 29598 32618 29650
rect 35926 29598 35978 29650
rect 42198 29598 42250 29650
rect 7870 29486 7922 29538
rect 3054 29430 3106 29482
rect 3278 29430 3330 29482
rect 10670 29486 10722 29538
rect 15766 29486 15818 29538
rect 16214 29486 16266 29538
rect 18958 29486 19010 29538
rect 3726 29374 3778 29426
rect 4602 29374 4654 29426
rect 5518 29374 5570 29426
rect 5854 29418 5906 29470
rect 8113 29430 8165 29482
rect 6190 29374 6242 29426
rect 6638 29374 6690 29426
rect 6862 29374 6914 29426
rect 8990 29374 9042 29426
rect 2774 29318 2826 29370
rect 11342 29430 11394 29482
rect 12798 29430 12850 29482
rect 13806 29430 13858 29482
rect 19350 29486 19402 29538
rect 9550 29374 9602 29426
rect 10426 29374 10478 29426
rect 12238 29374 12290 29426
rect 14752 29399 14804 29451
rect 14926 29374 14978 29426
rect 15038 29374 15090 29426
rect 15374 29374 15426 29426
rect 15486 29374 15538 29426
rect 16494 29374 16546 29426
rect 16718 29374 16770 29426
rect 17950 29374 18002 29426
rect 18174 29374 18226 29426
rect 18622 29374 18674 29426
rect 5742 29262 5794 29314
rect 4846 29150 4898 29202
rect 6526 29206 6578 29258
rect 12014 29262 12066 29314
rect 14366 29262 14418 29314
rect 17558 29262 17610 29314
rect 18790 29318 18842 29370
rect 19070 29374 19122 29426
rect 19742 29374 19794 29426
rect 19854 29374 19906 29426
rect 20022 29374 20074 29426
rect 21086 29374 21138 29426
rect 21422 29374 21474 29426
rect 25174 29430 25226 29482
rect 25342 29486 25394 29538
rect 29878 29486 29930 29538
rect 25734 29430 25786 29482
rect 34862 29486 34914 29538
rect 39062 29486 39114 29538
rect 42702 29486 42754 29538
rect 21534 29374 21586 29426
rect 21814 29374 21866 29426
rect 22206 29374 22258 29426
rect 22542 29374 22594 29426
rect 22654 29374 22706 29426
rect 24334 29374 24386 29426
rect 24670 29374 24722 29426
rect 25566 29374 25618 29426
rect 27190 29374 27242 29426
rect 27582 29374 27634 29426
rect 27918 29374 27970 29426
rect 28254 29374 28306 29426
rect 28590 29374 28642 29426
rect 29038 29409 29090 29461
rect 29150 29402 29202 29454
rect 29374 29402 29426 29454
rect 29598 29402 29650 29454
rect 31706 29430 31758 29482
rect 30830 29374 30882 29426
rect 20414 29262 20466 29314
rect 22374 29318 22426 29370
rect 31950 29374 32002 29426
rect 37194 29430 37246 29482
rect 33742 29374 33794 29426
rect 34618 29374 34670 29426
rect 36094 29374 36146 29426
rect 36318 29374 36370 29426
rect 37886 29374 37938 29426
rect 37998 29374 38050 29426
rect 38558 29374 38610 29426
rect 38782 29374 38834 29426
rect 39790 29374 39842 29426
rect 40798 29374 40850 29426
rect 44606 29374 44658 29426
rect 45390 29374 45442 29426
rect 45950 29374 46002 29426
rect 46174 29374 46226 29426
rect 46454 29374 46506 29426
rect 46734 29374 46786 29426
rect 48302 29374 48354 29426
rect 18174 29206 18226 29258
rect 26742 29262 26794 29314
rect 20918 29150 20970 29202
rect 24446 29206 24498 29258
rect 27358 29262 27410 29314
rect 33462 29262 33514 29314
rect 35478 29262 35530 29314
rect 39622 29262 39674 29314
rect 45782 29262 45834 29314
rect 23214 29150 23266 29202
rect 37438 29150 37490 29202
rect 38278 29150 38330 29202
rect 47070 29150 47122 29202
rect 47966 29150 48018 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 10110 28814 10162 28866
rect 12686 28814 12738 28866
rect 1822 28702 1874 28754
rect 3726 28702 3778 28754
rect 6302 28702 6354 28754
rect 14814 28758 14866 28810
rect 15934 28814 15986 28866
rect 18902 28814 18954 28866
rect 21702 28814 21754 28866
rect 23102 28814 23154 28866
rect 28086 28814 28138 28866
rect 18286 28758 18338 28810
rect 19518 28758 19570 28810
rect 20414 28758 20466 28810
rect 4510 28590 4562 28642
rect 6470 28646 6522 28698
rect 17446 28702 17498 28754
rect 23662 28702 23714 28754
rect 27750 28702 27802 28754
rect 29150 28758 29202 28810
rect 31054 28814 31106 28866
rect 36318 28814 36370 28866
rect 31838 28758 31890 28810
rect 43710 28814 43762 28866
rect 44942 28814 44994 28866
rect 37158 28702 37210 28754
rect 40574 28702 40626 28754
rect 42478 28702 42530 28754
rect 44326 28702 44378 28754
rect 47518 28702 47570 28754
rect 4902 28590 4954 28642
rect 5742 28552 5794 28604
rect 6078 28590 6130 28642
rect 7422 28590 7474 28642
rect 8298 28590 8350 28642
rect 8990 28590 9042 28642
rect 9866 28590 9918 28642
rect 10614 28590 10666 28642
rect 10894 28534 10946 28586
rect 11118 28534 11170 28586
rect 11342 28562 11394 28614
rect 11454 28534 11506 28586
rect 11678 28590 11730 28642
rect 11902 28590 11954 28642
rect 12182 28590 12234 28642
rect 13022 28590 13074 28642
rect 14030 28590 14082 28642
rect 8542 28478 8594 28530
rect 13638 28534 13690 28586
rect 14366 28552 14418 28604
rect 14926 28590 14978 28642
rect 15150 28590 15202 28642
rect 16270 28590 16322 28642
rect 17722 28552 17774 28604
rect 18398 28590 18450 28642
rect 19070 28590 19122 28642
rect 19406 28590 19458 28642
rect 19742 28590 19794 28642
rect 20302 28590 20354 28642
rect 20526 28590 20578 28642
rect 21198 28590 21250 28642
rect 21422 28590 21474 28642
rect 13806 28478 13858 28530
rect 22094 28534 22146 28586
rect 22262 28590 22314 28642
rect 22430 28590 22482 28642
rect 22542 28590 22594 28642
rect 23550 28590 23602 28642
rect 23886 28563 23938 28615
rect 24222 28590 24274 28642
rect 25454 28590 25506 28642
rect 27302 28590 27354 28642
rect 26330 28534 26382 28586
rect 28366 28590 28418 28642
rect 28478 28590 28530 28642
rect 29262 28590 29314 28642
rect 29598 28590 29650 28642
rect 29934 28590 29986 28642
rect 31614 28590 31666 28642
rect 31838 28590 31890 28642
rect 32566 28590 32618 28642
rect 30810 28534 30862 28586
rect 33014 28590 33066 28642
rect 33630 28590 33682 28642
rect 34506 28590 34558 28642
rect 34750 28590 34802 28642
rect 35198 28590 35250 28642
rect 36074 28590 36126 28642
rect 37550 28590 37602 28642
rect 39454 28590 39506 28642
rect 40238 28590 40290 28642
rect 43262 28590 43314 28642
rect 43374 28590 43426 28642
rect 45278 28590 45330 28642
rect 48302 28590 48354 28642
rect 26574 28478 26626 28530
rect 45614 28478 45666 28530
rect 7142 28366 7194 28418
rect 16998 28366 17050 28418
rect 25174 28366 25226 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 4902 27974 4954 28026
rect 7478 28030 7530 28082
rect 8934 27974 8986 28026
rect 16438 28030 16490 28082
rect 19518 28030 19570 28082
rect 25398 28030 25450 28082
rect 30774 28030 30826 28082
rect 31278 28030 31330 28082
rect 32566 28030 32618 28082
rect 39342 28030 39394 28082
rect 5462 27918 5514 27970
rect 9718 27918 9770 27970
rect 1598 27806 1650 27858
rect 4286 27806 4338 27858
rect 4734 27806 4786 27858
rect 5742 27806 5794 27858
rect 5966 27806 6018 27858
rect 6806 27862 6858 27914
rect 13470 27918 13522 27970
rect 6526 27806 6578 27858
rect 6638 27806 6690 27858
rect 6974 27806 7026 27858
rect 7758 27806 7810 27858
rect 7870 27806 7922 27858
rect 8038 27806 8090 27858
rect 9102 27806 9154 27858
rect 9998 27834 10050 27886
rect 10222 27862 10274 27914
rect 10446 27834 10498 27886
rect 10558 27841 10610 27893
rect 10894 27862 10946 27914
rect 11006 27862 11058 27914
rect 11230 27862 11282 27914
rect 11454 27834 11506 27886
rect 12014 27845 12066 27897
rect 13022 27834 13074 27886
rect 13638 27862 13690 27914
rect 14590 27918 14642 27970
rect 13246 27806 13298 27858
rect 20638 27918 20690 27970
rect 14030 27844 14082 27896
rect 14366 27806 14418 27858
rect 14758 27806 14810 27858
rect 15150 27806 15202 27858
rect 15374 27806 15426 27858
rect 17950 27806 18002 27858
rect 18286 27806 18338 27858
rect 18962 27844 19014 27896
rect 20246 27862 20298 27914
rect 22766 27918 22818 27970
rect 26854 27918 26906 27970
rect 32118 27918 32170 27970
rect 41134 27974 41186 28026
rect 19182 27806 19234 27858
rect 21310 27806 21362 27858
rect 21702 27835 21754 27887
rect 22542 27862 22594 27914
rect 23662 27862 23714 27914
rect 24110 27862 24162 27914
rect 23102 27806 23154 27858
rect 25790 27806 25842 27858
rect 26014 27821 26066 27873
rect 26350 27806 26402 27858
rect 2382 27694 2434 27746
rect 8430 27694 8482 27746
rect 19966 27750 20018 27802
rect 20806 27750 20858 27802
rect 26574 27806 26626 27858
rect 27470 27806 27522 27858
rect 27638 27806 27690 27858
rect 27806 27806 27858 27858
rect 27918 27806 27970 27858
rect 28814 27806 28866 27858
rect 29038 27845 29090 27897
rect 33406 27862 33458 27914
rect 33742 27862 33794 27914
rect 33910 27862 33962 27914
rect 34190 27918 34242 27970
rect 46510 27918 46562 27970
rect 29374 27806 29426 27858
rect 29934 27806 29986 27858
rect 30158 27806 30210 27858
rect 30942 27806 30994 27858
rect 34526 27806 34578 27858
rect 34750 27806 34802 27858
rect 35870 27806 35922 27858
rect 37718 27862 37770 27914
rect 16886 27694 16938 27746
rect 15262 27638 15314 27690
rect 21758 27694 21810 27746
rect 26126 27694 26178 27746
rect 28198 27694 28250 27746
rect 29262 27694 29314 27746
rect 6246 27582 6298 27634
rect 17614 27582 17666 27634
rect 18174 27638 18226 27690
rect 29822 27638 29874 27690
rect 36486 27694 36538 27746
rect 36934 27694 36986 27746
rect 37158 27750 37210 27802
rect 37326 27806 37378 27858
rect 37550 27806 37602 27858
rect 38334 27806 38386 27858
rect 38446 27806 38498 27858
rect 38726 27806 38778 27858
rect 39006 27806 39058 27858
rect 40238 27806 40290 27858
rect 40462 27806 40514 27858
rect 41358 27862 41410 27914
rect 41134 27806 41186 27858
rect 41806 27806 41858 27858
rect 42030 27806 42082 27858
rect 42814 27806 42866 27858
rect 45390 27806 45442 27858
rect 46266 27806 46318 27858
rect 47070 27806 47122 27858
rect 47294 27806 47346 27858
rect 48302 27806 48354 27858
rect 44718 27694 44770 27746
rect 46958 27638 47010 27690
rect 35030 27582 35082 27634
rect 35534 27582 35586 27634
rect 39958 27582 40010 27634
rect 47966 27582 48018 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 5014 27246 5066 27298
rect 7534 27190 7586 27242
rect 2718 27134 2770 27186
rect 9326 27134 9378 27186
rect 11118 27134 11170 27186
rect 12462 27190 12514 27242
rect 14982 27246 15034 27298
rect 23382 27246 23434 27298
rect 26518 27246 26570 27298
rect 27526 27246 27578 27298
rect 28366 27246 28418 27298
rect 20302 27190 20354 27242
rect 18174 27134 18226 27186
rect 18958 27134 19010 27186
rect 21702 27134 21754 27186
rect 24614 27134 24666 27186
rect 2830 27007 2882 27059
rect 3054 27022 3106 27074
rect 3726 27022 3778 27074
rect 3950 27022 4002 27074
rect 4230 27022 4282 27074
rect 4510 27022 4562 27074
rect 4734 27022 4786 27074
rect 5630 27022 5682 27074
rect 6190 27022 6242 27074
rect 7082 26984 7134 27036
rect 7758 27022 7810 27074
rect 8542 27022 8594 27074
rect 8654 27022 8706 27074
rect 9550 27022 9602 27074
rect 9774 27022 9826 27074
rect 10334 27022 10386 27074
rect 10670 27022 10722 27074
rect 11342 27022 11394 27074
rect 12574 27022 12626 27074
rect 12910 27022 12962 27074
rect 13862 27022 13914 27074
rect 10950 26966 11002 27018
rect 11510 26966 11562 27018
rect 14142 27022 14194 27074
rect 14422 27078 14474 27130
rect 25566 27134 25618 27186
rect 30382 27190 30434 27242
rect 33518 27246 33570 27298
rect 36262 27246 36314 27298
rect 41358 27246 41410 27298
rect 45110 27246 45162 27298
rect 35422 27134 35474 27186
rect 38894 27190 38946 27242
rect 38390 27134 38442 27186
rect 48134 27134 48186 27186
rect 14590 27022 14642 27074
rect 14814 27022 14866 27074
rect 15486 27022 15538 27074
rect 16270 27022 16322 27074
rect 18622 27022 18674 27074
rect 19562 26984 19614 27036
rect 20302 27022 20354 27074
rect 21198 27022 21250 27074
rect 21422 27022 21474 27074
rect 22262 27022 22314 27074
rect 8262 26910 8314 26962
rect 14254 26910 14306 26962
rect 22542 26966 22594 27018
rect 22654 26994 22706 27046
rect 22878 26994 22930 27046
rect 23102 26994 23154 27046
rect 24894 27022 24946 27074
rect 25342 27022 25394 27074
rect 25790 27022 25842 27074
rect 26126 27022 26178 27074
rect 26798 27022 26850 27074
rect 27022 27022 27074 27074
rect 27806 27022 27858 27074
rect 27918 27022 27970 27074
rect 28702 27022 28754 27074
rect 29150 26987 29202 27039
rect 29262 26994 29314 27046
rect 29486 26966 29538 27018
rect 29710 26994 29762 27046
rect 29990 27022 30042 27074
rect 30494 27022 30546 27074
rect 30718 27022 30770 27074
rect 31614 27022 31666 27074
rect 31838 27022 31890 27074
rect 32714 27022 32766 27074
rect 6078 26854 6130 26906
rect 31446 26854 31498 26906
rect 32958 26910 33010 26962
rect 33798 26966 33850 27018
rect 33966 26992 34018 27044
rect 34190 26983 34242 27035
rect 34862 26984 34914 27036
rect 35198 27022 35250 27074
rect 35590 26966 35642 27018
rect 35758 27022 35810 27074
rect 35982 27022 36034 27074
rect 37942 27022 37994 27074
rect 38782 27022 38834 27074
rect 39118 27022 39170 27074
rect 39342 27022 39394 27074
rect 39566 27022 39618 27074
rect 40350 26994 40402 27046
rect 43150 27022 43202 27074
rect 43822 27022 43874 27074
rect 43486 26966 43538 27018
rect 45390 27022 45442 27074
rect 45614 27022 45666 27074
rect 46174 27022 46226 27074
rect 46846 27022 46898 27074
rect 47070 27022 47122 27074
rect 46398 26966 46450 27018
rect 47294 27022 47346 27074
rect 39846 26910 39898 26962
rect 47574 26910 47626 26962
rect 43374 26854 43426 26906
rect 46622 26854 46674 26906
rect 37494 26798 37546 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 10278 26462 10330 26514
rect 10782 26462 10834 26514
rect 15374 26462 15426 26514
rect 16606 26462 16658 26514
rect 20638 26462 20690 26514
rect 4080 26350 4132 26402
rect 19742 26406 19794 26458
rect 21310 26462 21362 26514
rect 21982 26462 22034 26514
rect 27470 26462 27522 26514
rect 31670 26462 31722 26514
rect 29150 26406 29202 26458
rect 32118 26462 32170 26514
rect 32566 26462 32618 26514
rect 34582 26462 34634 26514
rect 40070 26462 40122 26514
rect 41918 26462 41970 26514
rect 8318 26350 8370 26402
rect 11734 26350 11786 26402
rect 23494 26350 23546 26402
rect 26070 26350 26122 26402
rect 29990 26350 30042 26402
rect 1598 26238 1650 26290
rect 3166 26238 3218 26290
rect 2550 26126 2602 26178
rect 3334 26182 3386 26234
rect 3838 26238 3890 26290
rect 4846 26238 4898 26290
rect 5182 26238 5234 26290
rect 5742 26238 5794 26290
rect 5966 26253 6018 26305
rect 6974 26294 7026 26346
rect 7534 26294 7586 26346
rect 8542 26294 8594 26346
rect 8094 26238 8146 26290
rect 9438 26238 9490 26290
rect 10446 26238 10498 26290
rect 11118 26238 11170 26290
rect 11230 26238 11282 26290
rect 11454 26238 11506 26290
rect 12294 26267 12346 26319
rect 12462 26238 12514 26290
rect 12842 26276 12894 26328
rect 13582 26238 13634 26290
rect 14030 26238 14082 26290
rect 14142 26238 14194 26290
rect 14288 26275 14340 26327
rect 15038 26238 15090 26290
rect 16942 26238 16994 26290
rect 18324 26275 18376 26327
rect 18510 26238 18562 26290
rect 18622 26238 18674 26290
rect 18958 26238 19010 26290
rect 19630 26238 19682 26290
rect 20302 26238 20354 26290
rect 20974 26238 21026 26290
rect 21646 26238 21698 26290
rect 23774 26238 23826 26290
rect 23998 26238 24050 26290
rect 24334 26238 24386 26290
rect 24558 26238 24610 26290
rect 25230 26273 25282 26325
rect 25342 26294 25394 26346
rect 25566 26294 25618 26346
rect 25790 26294 25842 26346
rect 28982 26294 29034 26346
rect 26574 26238 26626 26290
rect 26910 26238 26962 26290
rect 27134 26238 27186 26290
rect 28030 26238 28082 26290
rect 28366 26238 28418 26290
rect 29262 26238 29314 26290
rect 29486 26238 29538 26290
rect 29710 26238 29762 26290
rect 33014 26294 33066 26346
rect 33966 26350 34018 26402
rect 35086 26350 35138 26402
rect 40966 26350 41018 26402
rect 45166 26350 45218 26402
rect 46006 26350 46058 26402
rect 30830 26238 30882 26290
rect 30942 26238 30994 26290
rect 33182 26268 33234 26320
rect 33518 26268 33570 26320
rect 37774 26238 37826 26290
rect 38166 26238 38218 26290
rect 38894 26238 38946 26290
rect 39118 26238 39170 26290
rect 39230 26238 39282 26290
rect 41246 26238 41298 26290
rect 41358 26238 41410 26290
rect 41582 26238 41634 26290
rect 42478 26238 42530 26290
rect 45502 26238 45554 26290
rect 45726 26238 45778 26290
rect 46286 26238 46338 26290
rect 47406 26266 47458 26318
rect 47630 26266 47682 26318
rect 47798 26294 47850 26346
rect 47966 26273 48018 26325
rect 6078 26126 6130 26178
rect 12126 26126 12178 26178
rect 14702 26126 14754 26178
rect 1934 26014 1986 26066
rect 5294 26070 5346 26122
rect 13470 26070 13522 26122
rect 16214 26126 16266 26178
rect 17558 26126 17610 26178
rect 17950 26126 18002 26178
rect 22598 26126 22650 26178
rect 24446 26070 24498 26122
rect 26462 26070 26514 26122
rect 9606 26014 9658 26066
rect 28478 26070 28530 26122
rect 30494 26126 30546 26178
rect 36990 26126 37042 26178
rect 39510 26126 39562 26178
rect 43262 26126 43314 26178
rect 31110 26014 31162 26066
rect 38558 26014 38610 26066
rect 46622 26014 46674 26066
rect 47126 26014 47178 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 2662 25678 2714 25730
rect 5854 25678 5906 25730
rect 4846 25622 4898 25674
rect 8822 25678 8874 25730
rect 10334 25678 10386 25730
rect 13564 25678 13616 25730
rect 3726 25566 3778 25618
rect 6862 25566 6914 25618
rect 14814 25622 14866 25674
rect 26798 25678 26850 25730
rect 29542 25678 29594 25730
rect 34190 25678 34242 25730
rect 28030 25622 28082 25674
rect 44046 25678 44098 25730
rect 45222 25678 45274 25730
rect 46790 25678 46842 25730
rect 47686 25678 47738 25730
rect 18398 25566 18450 25618
rect 19518 25566 19570 25618
rect 30830 25566 30882 25618
rect 38446 25566 38498 25618
rect 40350 25566 40402 25618
rect 41470 25566 41522 25618
rect 45614 25566 45666 25618
rect 48246 25566 48298 25618
rect 2270 25454 2322 25506
rect 2382 25454 2434 25506
rect 3502 25454 3554 25506
rect 3166 25398 3218 25450
rect 3894 25398 3946 25450
rect 4106 25416 4158 25468
rect 4846 25454 4898 25506
rect 5518 25454 5570 25506
rect 6302 25454 6354 25506
rect 6638 25454 6690 25506
rect 7086 25454 7138 25506
rect 7534 25454 7586 25506
rect 8094 25454 8146 25506
rect 8542 25454 8594 25506
rect 8262 25398 8314 25450
rect 9214 25454 9266 25506
rect 13806 25454 13858 25506
rect 10090 25398 10142 25450
rect 11454 25398 11506 25450
rect 12126 25398 12178 25450
rect 12686 25398 12738 25450
rect 14310 25454 14362 25506
rect 14926 25454 14978 25506
rect 15150 25454 15202 25506
rect 15710 25454 15762 25506
rect 16494 25454 16546 25506
rect 18846 25454 18898 25506
rect 18958 25454 19010 25506
rect 19854 25454 19906 25506
rect 8430 25342 8482 25394
rect 19124 25398 19176 25450
rect 21534 25454 21586 25506
rect 22318 25454 22370 25506
rect 25118 25426 25170 25478
rect 27918 25454 27970 25506
rect 28254 25454 28306 25506
rect 29038 25454 29090 25506
rect 34638 25510 34690 25562
rect 35478 25510 35530 25562
rect 29262 25454 29314 25506
rect 31054 25454 31106 25506
rect 33070 25454 33122 25506
rect 14478 25342 14530 25394
rect 11902 25286 11954 25338
rect 20806 25342 20858 25394
rect 30494 25398 30546 25450
rect 31614 25398 31666 25450
rect 32174 25398 32226 25450
rect 33946 25398 33998 25450
rect 34750 25416 34802 25468
rect 35646 25454 35698 25506
rect 35870 25454 35922 25506
rect 36150 25454 36202 25506
rect 36878 25454 36930 25506
rect 37662 25454 37714 25506
rect 40686 25454 40738 25506
rect 43710 25454 43762 25506
rect 44718 25454 44770 25506
rect 44942 25454 44994 25506
rect 46062 25454 46114 25506
rect 46398 25454 46450 25506
rect 24222 25342 24274 25394
rect 35310 25342 35362 25394
rect 45782 25398 45834 25450
rect 46510 25454 46562 25506
rect 47182 25454 47234 25506
rect 47406 25454 47458 25506
rect 43374 25342 43426 25394
rect 20190 25230 20242 25282
rect 24838 25230 24890 25282
rect 37214 25230 37266 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 2158 24894 2210 24946
rect 15486 24894 15538 24946
rect 17502 24894 17554 24946
rect 22654 24894 22706 24946
rect 35254 24894 35306 24946
rect 38894 24894 38946 24946
rect 44326 24894 44378 24946
rect 5406 24782 5458 24834
rect 2494 24670 2546 24722
rect 3166 24670 3218 24722
rect 3390 24670 3442 24722
rect 3558 24670 3610 24722
rect 4846 24726 4898 24778
rect 6526 24726 6578 24778
rect 6974 24726 7026 24778
rect 7982 24726 8034 24778
rect 8542 24782 8594 24834
rect 9942 24782 9994 24834
rect 12126 24782 12178 24834
rect 21982 24782 22034 24834
rect 4062 24670 4114 24722
rect 5630 24670 5682 24722
rect 8318 24670 8370 24722
rect 8710 24670 8762 24722
rect 9438 24670 9490 24722
rect 9662 24670 9714 24722
rect 10782 24670 10834 24722
rect 11006 24670 11058 24722
rect 11454 24670 11506 24722
rect 11790 24670 11842 24722
rect 12238 24670 12290 24722
rect 12574 24670 12626 24722
rect 13694 24670 13746 24722
rect 14370 24708 14422 24760
rect 24558 24782 24610 24834
rect 15150 24670 15202 24722
rect 16046 24670 16098 24722
rect 17838 24670 17890 24722
rect 18548 24707 18600 24759
rect 18734 24670 18786 24722
rect 18846 24670 18898 24722
rect 19294 24670 19346 24722
rect 20078 24670 20130 24722
rect 22318 24670 22370 24722
rect 23662 24670 23714 24722
rect 24110 24698 24162 24750
rect 25790 24726 25842 24778
rect 26350 24782 26402 24834
rect 41582 24838 41634 24890
rect 24334 24670 24386 24722
rect 24726 24670 24778 24722
rect 25454 24670 25506 24722
rect 30419 24726 30471 24778
rect 30606 24726 30658 24778
rect 26518 24670 26570 24722
rect 27022 24670 27074 24722
rect 27470 24670 27522 24722
rect 27806 24670 27858 24722
rect 28254 24670 28306 24722
rect 29150 24670 29202 24722
rect 29486 24670 29538 24722
rect 30886 24705 30938 24757
rect 31110 24726 31162 24778
rect 31334 24782 31386 24834
rect 34694 24782 34746 24834
rect 35646 24782 35698 24834
rect 48078 24782 48130 24834
rect 31838 24670 31890 24722
rect 32062 24670 32114 24722
rect 33182 24670 33234 24722
rect 33406 24670 33458 24722
rect 34302 24670 34354 24722
rect 4304 24558 4356 24610
rect 25678 24614 25730 24666
rect 34414 24670 34466 24722
rect 37550 24670 37602 24722
rect 38334 24670 38386 24722
rect 38558 24670 38610 24722
rect 40126 24670 40178 24722
rect 40910 24670 40962 24722
rect 41358 24709 41410 24761
rect 41582 24670 41634 24722
rect 42254 24714 42306 24766
rect 42478 24670 42530 24722
rect 43262 24670 43314 24722
rect 43374 24670 43426 24722
rect 43878 24670 43930 24722
rect 44830 24670 44882 24722
rect 45054 24685 45106 24737
rect 45390 24670 45442 24722
rect 46174 24670 46226 24722
rect 10894 24502 10946 24554
rect 13582 24502 13634 24554
rect 18174 24558 18226 24610
rect 28030 24558 28082 24610
rect 28870 24558 28922 24610
rect 2830 24446 2882 24498
rect 16382 24446 16434 24498
rect 23326 24446 23378 24498
rect 25286 24502 25338 24554
rect 30214 24558 30266 24610
rect 29262 24502 29314 24554
rect 31950 24502 32002 24554
rect 33070 24502 33122 24554
rect 34022 24558 34074 24610
rect 42142 24558 42194 24610
rect 45166 24558 45218 24610
rect 39790 24446 39842 24498
rect 42982 24446 43034 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 3390 24054 3442 24106
rect 8430 24110 8482 24162
rect 11454 24110 11506 24162
rect 9214 24054 9266 24106
rect 11996 24110 12048 24162
rect 38222 24110 38274 24162
rect 14254 24054 14306 24106
rect 26574 24054 26626 24106
rect 28478 24054 28530 24106
rect 29486 24054 29538 24106
rect 38894 24110 38946 24162
rect 4398 23998 4450 24050
rect 15150 23998 15202 24050
rect 17054 23998 17106 24050
rect 20638 23998 20690 24050
rect 22374 23998 22426 24050
rect 36990 23998 37042 24050
rect 41134 23998 41186 24050
rect 42086 23998 42138 24050
rect 42534 23998 42586 24050
rect 42926 23998 42978 24050
rect 2382 23886 2434 23938
rect 2602 23848 2654 23900
rect 3278 23886 3330 23938
rect 3950 23858 4002 23910
rect 4174 23886 4226 23938
rect 7758 23886 7810 23938
rect 7870 23886 7922 23938
rect 8036 23886 8088 23938
rect 8878 23886 8930 23938
rect 9214 23886 9266 23938
rect 10110 23886 10162 23938
rect 4566 23830 4618 23882
rect 6638 23830 6690 23882
rect 6862 23830 6914 23882
rect 7310 23830 7362 23882
rect 11118 23886 11170 23938
rect 12238 23886 12290 23938
rect 12742 23886 12794 23938
rect 12910 23886 12962 23938
rect 13470 23886 13522 23938
rect 14142 23886 14194 23938
rect 17838 23886 17890 23938
rect 17950 23886 18002 23938
rect 18734 23886 18786 23938
rect 21534 23886 21586 23938
rect 21926 23886 21978 23938
rect 22878 23886 22930 23938
rect 23662 23886 23714 23938
rect 26122 23848 26174 23900
rect 26798 23886 26850 23938
rect 27694 23886 27746 23938
rect 28366 23886 28418 23938
rect 29262 23886 29314 23938
rect 30002 23848 30054 23900
rect 30606 23858 30658 23910
rect 30830 23886 30882 23938
rect 33518 23886 33570 23938
rect 34302 23886 34354 23938
rect 25566 23774 25618 23826
rect 6526 23718 6578 23770
rect 31054 23774 31106 23826
rect 31222 23830 31274 23882
rect 35310 23886 35362 23938
rect 35758 23886 35810 23938
rect 36094 23859 36146 23911
rect 36430 23886 36482 23938
rect 37102 23871 37154 23923
rect 37326 23886 37378 23938
rect 37886 23886 37938 23938
rect 38558 23886 38610 23938
rect 40126 23886 40178 23938
rect 40686 23886 40738 23938
rect 40518 23830 40570 23882
rect 41246 23871 41298 23923
rect 41470 23886 41522 23938
rect 43038 23842 43090 23894
rect 43262 23886 43314 23938
rect 43598 23886 43650 23938
rect 45278 23886 45330 23938
rect 45502 23886 45554 23938
rect 45838 23859 45890 23911
rect 46174 23886 46226 23938
rect 47182 23886 47234 23938
rect 47742 23886 47794 23938
rect 47574 23830 47626 23882
rect 31614 23774 31666 23826
rect 2046 23662 2098 23714
rect 9774 23662 9826 23714
rect 21366 23662 21418 23714
rect 35646 23718 35698 23770
rect 40238 23718 40290 23770
rect 34974 23662 35026 23714
rect 43934 23662 43986 23714
rect 46286 23718 46338 23770
rect 47294 23718 47346 23770
rect 44942 23662 44994 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 17558 23326 17610 23378
rect 5966 23270 6018 23322
rect 4286 23214 4338 23266
rect 12686 23270 12738 23322
rect 17950 23326 18002 23378
rect 24446 23326 24498 23378
rect 26462 23326 26514 23378
rect 34638 23326 34690 23378
rect 39006 23326 39058 23378
rect 39678 23326 39730 23378
rect 40294 23326 40346 23378
rect 8486 23214 8538 23266
rect 5742 23158 5794 23210
rect 25790 23214 25842 23266
rect 30326 23214 30378 23266
rect 31614 23214 31666 23266
rect 45726 23270 45778 23322
rect 1598 23102 1650 23154
rect 4622 23102 4674 23154
rect 5518 23102 5570 23154
rect 6078 23102 6130 23154
rect 6526 23102 6578 23154
rect 6862 23129 6914 23181
rect 7198 23102 7250 23154
rect 7758 23102 7810 23154
rect 8094 23102 8146 23154
rect 8206 23102 8258 23154
rect 7926 23046 7978 23098
rect 9438 23102 9490 23154
rect 10222 23102 10274 23154
rect 12686 23102 12738 23154
rect 13358 23102 13410 23154
rect 13918 23102 13970 23154
rect 14030 23102 14082 23154
rect 14198 23102 14250 23154
rect 16440 23102 16492 23154
rect 16606 23102 16658 23154
rect 16718 23102 16770 23154
rect 18286 23102 18338 23154
rect 19036 23139 19088 23191
rect 19182 23102 19234 23154
rect 19294 23102 19346 23154
rect 20414 23102 20466 23154
rect 21086 23102 21138 23154
rect 21198 23102 21250 23154
rect 21534 23102 21586 23154
rect 22468 23139 22520 23191
rect 33966 23214 34018 23266
rect 40966 23214 41018 23266
rect 46902 23214 46954 23266
rect 48022 23214 48074 23266
rect 22654 23102 22706 23154
rect 22766 23102 22818 23154
rect 23628 23139 23680 23191
rect 23774 23102 23826 23154
rect 23886 23102 23938 23154
rect 24110 23102 24162 23154
rect 26126 23102 26178 23154
rect 26798 23102 26850 23154
rect 26910 23102 26962 23154
rect 27962 23140 28014 23192
rect 28702 23102 28754 23154
rect 29262 23102 29314 23154
rect 29486 23102 29538 23154
rect 29934 23102 29986 23154
rect 30046 23102 30098 23154
rect 30998 23102 31050 23154
rect 31278 23102 31330 23154
rect 2382 22990 2434 23042
rect 6750 22990 6802 23042
rect 12126 22990 12178 23042
rect 16046 22990 16098 23042
rect 18622 22990 18674 23042
rect 22094 22990 22146 23042
rect 31446 23046 31498 23098
rect 31726 23102 31778 23154
rect 33014 23158 33066 23210
rect 33182 23158 33234 23210
rect 33406 23141 33458 23193
rect 34302 23102 34354 23154
rect 34974 23102 35026 23154
rect 35758 23102 35810 23154
rect 37998 23102 38050 23154
rect 38670 23102 38722 23154
rect 39342 23102 39394 23154
rect 41246 23102 41298 23154
rect 41470 23102 41522 23154
rect 42142 23102 42194 23154
rect 44046 23102 44098 23154
rect 44830 23102 44882 23154
rect 45614 23102 45666 23154
rect 46062 23141 46114 23193
rect 46286 23102 46338 23154
rect 47182 23102 47234 23154
rect 47406 23102 47458 23154
rect 47630 23102 47682 23154
rect 47742 23102 47794 23154
rect 32566 22990 32618 23042
rect 37662 22990 37714 23042
rect 45222 22990 45274 23042
rect 4790 22878 4842 22930
rect 14590 22878 14642 22930
rect 20078 22878 20130 22930
rect 20750 22878 20802 22930
rect 23214 22878 23266 22930
rect 27246 22878 27298 22930
rect 28814 22934 28866 22986
rect 29486 22934 29538 22986
rect 32006 22878 32058 22930
rect 38334 22878 38386 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 3894 22542 3946 22594
rect 5854 22542 5906 22594
rect 6974 22542 7026 22594
rect 7646 22542 7698 22594
rect 11230 22542 11282 22594
rect 12574 22486 12626 22538
rect 14702 22542 14754 22594
rect 16382 22542 16434 22594
rect 18342 22542 18394 22594
rect 20414 22542 20466 22594
rect 2158 22318 2210 22370
rect 2830 22318 2882 22370
rect 3166 22318 3218 22370
rect 3334 22374 3386 22426
rect 4958 22430 5010 22482
rect 9102 22430 9154 22482
rect 19070 22486 19122 22538
rect 21534 22542 21586 22594
rect 22094 22542 22146 22594
rect 23774 22542 23826 22594
rect 14142 22430 14194 22482
rect 5126 22374 5178 22426
rect 3614 22318 3666 22370
rect 4734 22318 4786 22370
rect 5518 22318 5570 22370
rect 4510 22262 4562 22314
rect 6302 22318 6354 22370
rect 6414 22318 6466 22370
rect 6582 22318 6634 22370
rect 7310 22318 7362 22370
rect 9214 22303 9266 22355
rect 9438 22318 9490 22370
rect 10894 22318 10946 22370
rect 11566 22318 11618 22370
rect 11786 22280 11838 22332
rect 12462 22318 12514 22370
rect 13470 22318 13522 22370
rect 13582 22318 13634 22370
rect 13750 22318 13802 22370
rect 15094 22318 15146 22370
rect 15262 22318 15314 22370
rect 15374 22318 15426 22370
rect 15710 22318 15762 22370
rect 15822 22318 15874 22370
rect 15990 22318 16042 22370
rect 16998 22318 17050 22370
rect 17614 22318 17666 22370
rect 17782 22374 17834 22426
rect 19910 22430 19962 22482
rect 30494 22486 30546 22538
rect 31054 22542 31106 22594
rect 31558 22542 31610 22594
rect 33462 22542 33514 22594
rect 33966 22542 34018 22594
rect 25454 22430 25506 22482
rect 26574 22430 26626 22482
rect 28478 22430 28530 22482
rect 32734 22430 32786 22482
rect 36262 22430 36314 22482
rect 39230 22430 39282 22482
rect 41134 22430 41186 22482
rect 43654 22430 43706 22482
rect 45838 22430 45890 22482
rect 18062 22318 18114 22370
rect 18846 22318 18898 22370
rect 19070 22318 19122 22370
rect 20078 22318 20130 22370
rect 21198 22318 21250 22370
rect 22488 22318 22540 22370
rect 22654 22318 22706 22370
rect 22766 22318 22818 22370
rect 23102 22318 23154 22370
rect 23214 22318 23266 22370
rect 23380 22318 23432 22370
rect 24782 22318 24834 22370
rect 24894 22318 24946 22370
rect 25790 22318 25842 22370
rect 3502 22206 3554 22258
rect 2270 22150 2322 22202
rect 25062 22262 25114 22314
rect 29642 22280 29694 22332
rect 30382 22318 30434 22370
rect 30718 22318 30770 22370
rect 31838 22318 31890 22370
rect 32062 22318 32114 22370
rect 32286 22318 32338 22370
rect 32566 22288 32618 22340
rect 32958 22318 33010 22370
rect 33182 22318 33234 22370
rect 34302 22318 34354 22370
rect 34414 22318 34466 22370
rect 34638 22318 34690 22370
rect 34918 22318 34970 22370
rect 35646 22318 35698 22370
rect 35870 22318 35922 22370
rect 37326 22318 37378 22370
rect 37438 22318 37490 22370
rect 37942 22318 37994 22370
rect 38446 22318 38498 22370
rect 42030 22318 42082 22370
rect 42366 22318 42418 22370
rect 42814 22279 42866 22331
rect 43038 22318 43090 22370
rect 43934 22318 43986 22370
rect 44046 22318 44098 22370
rect 45054 22318 45106 22370
rect 17950 22206 18002 22258
rect 35366 22206 35418 22258
rect 37046 22206 37098 22258
rect 47742 22206 47794 22258
rect 10558 22094 10610 22146
rect 24502 22094 24554 22146
rect 42926 22150 42978 22202
rect 41694 22094 41746 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 2270 21758 2322 21810
rect 13022 21758 13074 21810
rect 6974 21702 7026 21754
rect 19182 21758 19234 21810
rect 20246 21758 20298 21810
rect 20694 21758 20746 21810
rect 23046 21758 23098 21810
rect 27974 21758 28026 21810
rect 38166 21758 38218 21810
rect 3614 21646 3666 21698
rect 12350 21646 12402 21698
rect 18286 21646 18338 21698
rect 2606 21534 2658 21586
rect 3278 21534 3330 21586
rect 4058 21572 4110 21624
rect 4734 21534 4786 21586
rect 5406 21534 5458 21586
rect 6641 21573 6693 21625
rect 7198 21534 7250 21586
rect 7758 21534 7810 21586
rect 8766 21534 8818 21586
rect 9662 21534 9714 21586
rect 10446 21534 10498 21586
rect 12686 21534 12738 21586
rect 13582 21534 13634 21586
rect 13694 21534 13746 21586
rect 13840 21572 13892 21624
rect 18678 21646 18730 21698
rect 21702 21646 21754 21698
rect 28590 21702 28642 21754
rect 24278 21646 24330 21698
rect 32398 21646 32450 21698
rect 15188 21572 15240 21624
rect 15374 21534 15426 21586
rect 15486 21534 15538 21586
rect 16886 21534 16938 21586
rect 17950 21534 18002 21586
rect 5630 21422 5682 21474
rect 14814 21422 14866 21474
rect 4510 21366 4562 21418
rect 15990 21422 16042 21474
rect 16438 21422 16490 21474
rect 17670 21422 17722 21474
rect 18118 21478 18170 21530
rect 18398 21534 18450 21586
rect 19518 21534 19570 21586
rect 21422 21534 21474 21586
rect 21982 21562 22034 21614
rect 22150 21569 22202 21621
rect 22430 21562 22482 21614
rect 22542 21569 22594 21621
rect 24726 21534 24778 21586
rect 25566 21534 25618 21586
rect 25678 21534 25730 21586
rect 25824 21572 25876 21624
rect 27200 21584 27252 21636
rect 36094 21646 36146 21698
rect 40294 21646 40346 21698
rect 46118 21646 46170 21698
rect 27358 21534 27410 21586
rect 27470 21534 27522 21586
rect 28702 21534 28754 21586
rect 29374 21534 29426 21586
rect 29710 21534 29762 21586
rect 33238 21534 33290 21586
rect 33406 21534 33458 21586
rect 36542 21534 36594 21586
rect 36878 21534 36930 21586
rect 37214 21534 37266 21586
rect 38894 21534 38946 21586
rect 39342 21534 39394 21586
rect 39678 21534 39730 21586
rect 40798 21534 40850 21586
rect 41582 21534 41634 21586
rect 43486 21534 43538 21586
rect 44046 21549 44098 21601
rect 44270 21534 44322 21586
rect 44606 21534 44658 21586
rect 45614 21534 45666 21586
rect 45838 21534 45890 21586
rect 46622 21549 46674 21601
rect 46958 21534 47010 21586
rect 47350 21563 47402 21615
rect 47742 21534 47794 21586
rect 26238 21422 26290 21474
rect 30494 21422 30546 21474
rect 34190 21422 34242 21474
rect 43934 21422 43986 21474
rect 46510 21422 46562 21474
rect 47294 21422 47346 21474
rect 48246 21422 48298 21474
rect 8430 21310 8482 21362
rect 14254 21310 14306 21362
rect 21086 21310 21138 21362
rect 36654 21366 36706 21418
rect 26798 21310 26850 21362
rect 37550 21310 37602 21362
rect 38558 21310 38610 21362
rect 44942 21310 44994 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 4846 20974 4898 21026
rect 5854 20974 5906 21026
rect 10558 20974 10610 21026
rect 11230 20974 11282 21026
rect 18342 20974 18394 21026
rect 11790 20918 11842 20970
rect 19462 20974 19514 21026
rect 19910 20974 19962 21026
rect 29374 20974 29426 21026
rect 34526 20974 34578 21026
rect 4286 20862 4338 20914
rect 6974 20862 7026 20914
rect 8878 20862 8930 20914
rect 14366 20862 14418 20914
rect 15542 20862 15594 20914
rect 15990 20862 16042 20914
rect 33294 20918 33346 20970
rect 40910 20974 40962 21026
rect 43094 20974 43146 21026
rect 1598 20750 1650 20802
rect 2382 20750 2434 20802
rect 5182 20750 5234 20802
rect 6414 20750 6466 20802
rect 6526 20750 6578 20802
rect 6248 20694 6300 20746
rect 9662 20750 9714 20802
rect 9886 20750 9938 20802
rect 9998 20750 10050 20802
rect 11566 20750 11618 20802
rect 12014 20750 12066 20802
rect 12574 20750 12626 20802
rect 10164 20694 10216 20746
rect 13358 20750 13410 20802
rect 14758 20750 14810 20802
rect 14926 20750 14978 20802
rect 15038 20750 15090 20802
rect 16158 20750 16210 20802
rect 16830 20750 16882 20802
rect 17166 20750 17218 20802
rect 17614 20750 17666 20802
rect 17950 20750 18002 20802
rect 18062 20750 18114 20802
rect 17782 20694 17834 20746
rect 18734 20750 18786 20802
rect 18902 20806 18954 20858
rect 24894 20862 24946 20914
rect 28478 20862 28530 20914
rect 32398 20862 32450 20914
rect 37102 20862 37154 20914
rect 41526 20862 41578 20914
rect 43822 20862 43874 20914
rect 45502 20862 45554 20914
rect 19182 20750 19234 20802
rect 20190 20722 20242 20774
rect 20414 20694 20466 20746
rect 20638 20694 20690 20746
rect 20750 20715 20802 20767
rect 23102 20750 23154 20802
rect 23326 20750 23378 20802
rect 21758 20694 21810 20746
rect 22094 20694 22146 20746
rect 24558 20750 24610 20802
rect 25118 20750 25170 20802
rect 25790 20750 25842 20802
rect 26574 20750 26626 20802
rect 29038 20750 29090 20802
rect 23550 20694 23602 20746
rect 24950 20694 25002 20746
rect 30942 20750 30994 20802
rect 31390 20750 31442 20802
rect 31726 20723 31778 20775
rect 32062 20750 32114 20802
rect 32734 20750 32786 20802
rect 33182 20750 33234 20802
rect 33518 20750 33570 20802
rect 34862 20750 34914 20802
rect 35142 20750 35194 20802
rect 35422 20750 35474 20802
rect 32566 20694 32618 20746
rect 35646 20750 35698 20802
rect 36318 20750 36370 20802
rect 39006 20750 39058 20802
rect 39790 20750 39842 20802
rect 39902 20750 39954 20802
rect 40574 20750 40626 20802
rect 41806 20750 41858 20802
rect 42254 20711 42306 20763
rect 42478 20750 42530 20802
rect 43374 20750 43426 20802
rect 43486 20750 43538 20802
rect 43934 20706 43986 20758
rect 44270 20750 44322 20802
rect 44718 20750 44770 20802
rect 48302 20750 48354 20802
rect 19070 20638 19122 20690
rect 47406 20638 47458 20690
rect 13694 20526 13746 20578
rect 16494 20526 16546 20578
rect 31278 20582 31330 20634
rect 30606 20526 30658 20578
rect 34134 20526 34186 20578
rect 35982 20526 36034 20578
rect 42030 20582 42082 20634
rect 40238 20526 40290 20578
rect 47966 20526 48018 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 1822 20190 1874 20242
rect 18510 20190 18562 20242
rect 28422 20190 28474 20242
rect 28870 20190 28922 20242
rect 12350 20078 12402 20130
rect 13414 20078 13466 20130
rect 16718 20078 16770 20130
rect 19574 20078 19626 20130
rect 2158 19966 2210 20018
rect 2270 19966 2322 20018
rect 6492 20003 6544 20055
rect 6638 19966 6690 20018
rect 6750 19966 6802 20018
rect 7534 19966 7586 20018
rect 7758 19966 7810 20018
rect 7870 19966 7922 20018
rect 8038 19966 8090 20018
rect 13974 20022 14026 20074
rect 9662 19966 9714 20018
rect 13022 19966 13074 20018
rect 13694 19966 13746 20018
rect 13806 19966 13858 20018
rect 14142 19966 14194 20018
rect 14814 19966 14866 20018
rect 14926 19966 14978 20018
rect 15094 19966 15146 20018
rect 15262 19966 15314 20018
rect 15710 19966 15762 20018
rect 15934 19966 15986 20018
rect 16382 19966 16434 20018
rect 17502 19966 17554 20018
rect 17838 19966 17890 20018
rect 18846 19966 18898 20018
rect 19070 19966 19122 20018
rect 20190 20022 20242 20074
rect 20638 20022 20690 20074
rect 21870 20078 21922 20130
rect 27134 20078 27186 20130
rect 22542 20022 22594 20074
rect 19294 19966 19346 20018
rect 21646 19966 21698 20018
rect 22766 19966 22818 20018
rect 24110 20022 24162 20074
rect 31222 20078 31274 20130
rect 36038 20078 36090 20130
rect 36878 20078 36930 20130
rect 23774 19966 23826 20018
rect 24446 19966 24498 20018
rect 25454 19966 25506 20018
rect 25790 19966 25842 20018
rect 25902 19966 25954 20018
rect 26088 20004 26140 20056
rect 26798 19966 26850 20018
rect 33742 20022 33794 20074
rect 28030 19966 28082 20018
rect 30270 19966 30322 20018
rect 30606 19966 30658 20018
rect 31726 19966 31778 20018
rect 32062 19966 32114 20018
rect 32286 19966 32338 20018
rect 33014 19966 33066 20018
rect 33406 19966 33458 20018
rect 35290 20022 35342 20074
rect 38110 20078 38162 20130
rect 34414 19966 34466 20018
rect 35534 19966 35586 20018
rect 36318 19966 36370 20018
rect 36542 19966 36594 20018
rect 37718 20022 37770 20074
rect 37214 19966 37266 20018
rect 37886 19966 37938 20018
rect 3054 19854 3106 19906
rect 4958 19854 5010 19906
rect 5686 19854 5738 19906
rect 7198 19854 7250 19906
rect 8430 19854 8482 19906
rect 9046 19854 9098 19906
rect 10446 19854 10498 19906
rect 14534 19854 14586 19906
rect 6078 19742 6130 19794
rect 12854 19742 12906 19794
rect 15598 19798 15650 19850
rect 24110 19854 24162 19906
rect 23102 19742 23154 19794
rect 25286 19798 25338 19850
rect 26462 19854 26514 19906
rect 27694 19742 27746 19794
rect 30718 19798 30770 19850
rect 31558 19742 31610 19794
rect 32398 19798 32450 19850
rect 33182 19854 33234 19906
rect 38278 19910 38330 19962
rect 38782 19966 38834 20018
rect 40014 19966 40066 20018
rect 40350 19966 40402 20018
rect 43822 19966 43874 20018
rect 44158 19966 44210 20018
rect 44494 19966 44546 20018
rect 44718 19966 44770 20018
rect 45390 19966 45442 20018
rect 46174 19966 46226 20018
rect 48078 19966 48130 20018
rect 41134 19854 41186 19906
rect 43038 19854 43090 19906
rect 39118 19742 39170 19794
rect 39902 19798 39954 19850
rect 44046 19798 44098 19850
rect 45054 19742 45106 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 6974 19406 7026 19458
rect 5070 19350 5122 19402
rect 6190 19350 6242 19402
rect 8990 19406 9042 19458
rect 12798 19406 12850 19458
rect 13694 19406 13746 19458
rect 15430 19406 15482 19458
rect 20526 19406 20578 19458
rect 21366 19406 21418 19458
rect 23494 19406 23546 19458
rect 27134 19406 27186 19458
rect 38054 19406 38106 19458
rect 40238 19406 40290 19458
rect 43990 19406 44042 19458
rect 4286 19182 4338 19234
rect 4958 19182 5010 19234
rect 6078 19182 6130 19234
rect 6414 19182 6466 19234
rect 6638 19182 6690 19234
rect 7870 19182 7922 19234
rect 9326 19182 9378 19234
rect 9438 19182 9490 19234
rect 10222 19182 10274 19234
rect 12126 19182 12178 19234
rect 12462 19182 12514 19234
rect 14030 19182 14082 19234
rect 14870 19238 14922 19290
rect 14590 19182 14642 19234
rect 14702 19182 14754 19234
rect 15038 19182 15090 19234
rect 15710 19182 15762 19234
rect 15990 19238 16042 19290
rect 16774 19294 16826 19346
rect 17166 19294 17218 19346
rect 16158 19182 16210 19234
rect 17502 19182 17554 19234
rect 18062 19182 18114 19234
rect 18342 19238 18394 19290
rect 22262 19294 22314 19346
rect 22710 19294 22762 19346
rect 23158 19294 23210 19346
rect 18510 19182 18562 19234
rect 24054 19238 24106 19290
rect 31726 19294 31778 19346
rect 33854 19294 33906 19346
rect 35758 19294 35810 19346
rect 38614 19294 38666 19346
rect 45614 19350 45666 19402
rect 47910 19406 47962 19458
rect 47182 19350 47234 19402
rect 19070 19182 19122 19234
rect 19294 19143 19346 19195
rect 19630 19182 19682 19234
rect 20190 19182 20242 19234
rect 21534 19182 21586 19234
rect 23774 19182 23826 19234
rect 23886 19182 23938 19234
rect 24222 19182 24274 19234
rect 24558 19182 24610 19234
rect 24726 19238 24778 19290
rect 24894 19182 24946 19234
rect 25006 19182 25058 19234
rect 25678 19182 25730 19234
rect 26126 19182 26178 19234
rect 26350 19182 26402 19234
rect 27470 19182 27522 19234
rect 29038 19182 29090 19234
rect 29822 19182 29874 19234
rect 14310 19070 14362 19122
rect 15822 19070 15874 19122
rect 17782 19070 17834 19122
rect 32622 19154 32674 19206
rect 32846 19154 32898 19206
rect 18174 19070 18226 19122
rect 33070 19126 33122 19178
rect 33182 19147 33234 19199
rect 36542 19182 36594 19234
rect 37438 19182 37490 19234
rect 37550 19182 37602 19234
rect 37774 19182 37826 19234
rect 39230 19154 39282 19206
rect 41806 19126 41858 19178
rect 42142 19126 42194 19178
rect 42590 19126 42642 19178
rect 42788 19149 42840 19201
rect 43486 19182 43538 19234
rect 43710 19182 43762 19234
rect 44830 19182 44882 19234
rect 44942 19182 44994 19234
rect 45222 19182 45274 19234
rect 45726 19182 45778 19234
rect 45950 19182 46002 19234
rect 46846 19182 46898 19234
rect 47070 19182 47122 19234
rect 47406 19182 47458 19234
rect 47630 19182 47682 19234
rect 4006 18958 4058 19010
rect 7534 18958 7586 19010
rect 8598 18958 8650 19010
rect 19406 19014 19458 19066
rect 25286 19070 25338 19122
rect 26630 19070 26682 19122
rect 32342 19070 32394 19122
rect 42926 19070 42978 19122
rect 25846 18958 25898 19010
rect 27862 18958 27914 19010
rect 28310 18958 28362 19010
rect 37102 18958 37154 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 14814 18622 14866 18674
rect 15486 18622 15538 18674
rect 21030 18622 21082 18674
rect 23718 18622 23770 18674
rect 31726 18510 31778 18562
rect 3054 18398 3106 18450
rect 5742 18398 5794 18450
rect 6134 18454 6186 18506
rect 6526 18398 6578 18450
rect 6862 18436 6914 18488
rect 7926 18398 7978 18450
rect 8318 18413 8370 18465
rect 8542 18398 8594 18450
rect 9774 18398 9826 18450
rect 13134 18425 13186 18477
rect 13918 18398 13970 18450
rect 14310 18427 14362 18479
rect 15150 18398 15202 18450
rect 15822 18398 15874 18450
rect 15934 18398 15986 18450
rect 17390 18425 17442 18477
rect 18734 18398 18786 18450
rect 20078 18398 20130 18450
rect 21590 18454 21642 18506
rect 20414 18398 20466 18450
rect 21310 18398 21362 18450
rect 21982 18398 22034 18450
rect 22654 18436 22706 18488
rect 22990 18398 23042 18450
rect 23550 18398 23602 18450
rect 24110 18398 24162 18450
rect 3838 18286 3890 18338
rect 6302 18286 6354 18338
rect 7478 18286 7530 18338
rect 8206 18286 8258 18338
rect 14366 18286 14418 18338
rect 21422 18286 21474 18338
rect 23214 18286 23266 18338
rect 23382 18342 23434 18394
rect 24222 18398 24274 18450
rect 25342 18442 25394 18494
rect 25566 18398 25618 18450
rect 26350 18398 26402 18450
rect 26462 18398 26514 18450
rect 26630 18342 26682 18394
rect 26798 18398 26850 18450
rect 27022 18398 27074 18450
rect 25230 18286 25282 18338
rect 27974 18342 28026 18394
rect 28142 18398 28194 18450
rect 28590 18426 28642 18478
rect 33014 18454 33066 18506
rect 33182 18510 33234 18562
rect 29038 18398 29090 18450
rect 32398 18398 32450 18450
rect 33742 18454 33794 18506
rect 33406 18398 33458 18450
rect 34470 18398 34522 18450
rect 28814 18342 28866 18394
rect 35198 18398 35250 18450
rect 35310 18398 35362 18450
rect 38390 18454 38442 18506
rect 38558 18398 38610 18450
rect 38782 18398 38834 18450
rect 39118 18436 39170 18488
rect 39566 18398 39618 18450
rect 39678 18398 39730 18450
rect 39846 18398 39898 18450
rect 40798 18398 40850 18450
rect 41022 18398 41074 18450
rect 41302 18398 41354 18450
rect 41694 18398 41746 18450
rect 42030 18398 42082 18450
rect 42366 18398 42418 18450
rect 43710 18454 43762 18506
rect 42590 18398 42642 18450
rect 43934 18431 43986 18483
rect 44494 18434 44546 18486
rect 44692 18438 44744 18490
rect 45054 18398 45106 18450
rect 29822 18286 29874 18338
rect 34862 18286 34914 18338
rect 36094 18286 36146 18338
rect 37998 18286 38050 18338
rect 40238 18286 40290 18338
rect 42870 18286 42922 18338
rect 44718 18286 44770 18338
rect 45838 18286 45890 18338
rect 47742 18286 47794 18338
rect 12126 18174 12178 18226
rect 24502 18174 24554 18226
rect 26070 18174 26122 18226
rect 27358 18174 27410 18226
rect 32230 18174 32282 18226
rect 42142 18230 42194 18282
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 6022 17838 6074 17890
rect 9662 17838 9714 17890
rect 18454 17838 18506 17890
rect 23326 17782 23378 17834
rect 24782 17838 24834 17890
rect 5126 17726 5178 17778
rect 7198 17726 7250 17778
rect 13806 17726 13858 17778
rect 16046 17726 16098 17778
rect 20526 17726 20578 17778
rect 21982 17726 22034 17778
rect 24390 17726 24442 17778
rect 28030 17782 28082 17834
rect 35422 17838 35474 17890
rect 42030 17838 42082 17890
rect 29262 17726 29314 17778
rect 43934 17782 43986 17834
rect 30550 17726 30602 17778
rect 39006 17726 39058 17778
rect 40910 17726 40962 17778
rect 43150 17726 43202 17778
rect 5518 17614 5570 17666
rect 5742 17614 5794 17666
rect 6414 17614 6466 17666
rect 9998 17614 10050 17666
rect 10110 17614 10162 17666
rect 10894 17614 10946 17666
rect 12798 17614 12850 17666
rect 14200 17614 14252 17666
rect 14366 17614 14418 17666
rect 14478 17614 14530 17666
rect 15262 17614 15314 17666
rect 17950 17614 18002 17666
rect 18734 17614 18786 17666
rect 18846 17614 18898 17666
rect 19014 17614 19066 17666
rect 19182 17614 19234 17666
rect 20078 17614 20130 17666
rect 20302 17575 20354 17627
rect 20750 17614 20802 17666
rect 21198 17614 21250 17666
rect 21758 17614 21810 17666
rect 22430 17614 22482 17666
rect 4230 17502 4282 17554
rect 4678 17502 4730 17554
rect 22094 17558 22146 17610
rect 22766 17614 22818 17666
rect 23438 17614 23490 17666
rect 23662 17614 23714 17666
rect 25118 17614 25170 17666
rect 25230 17614 25282 17666
rect 25454 17614 25506 17666
rect 26462 17614 26514 17666
rect 26798 17614 26850 17666
rect 26910 17614 26962 17666
rect 26630 17558 26682 17610
rect 27190 17614 27242 17666
rect 28142 17614 28194 17666
rect 28478 17614 28530 17666
rect 29486 17614 29538 17666
rect 29094 17558 29146 17610
rect 29710 17586 29762 17638
rect 30718 17614 30770 17666
rect 32174 17614 32226 17666
rect 32958 17614 33010 17666
rect 35814 17614 35866 17666
rect 35982 17614 36034 17666
rect 36094 17614 36146 17666
rect 38110 17614 38162 17666
rect 38222 17614 38274 17666
rect 41358 17614 41410 17666
rect 41470 17614 41522 17666
rect 41636 17614 41688 17666
rect 42478 17614 42530 17666
rect 42590 17614 42642 17666
rect 42756 17614 42808 17666
rect 43710 17614 43762 17666
rect 43934 17614 43986 17666
rect 45278 17614 45330 17666
rect 45390 17614 45442 17666
rect 46174 17614 46226 17666
rect 9102 17502 9154 17554
rect 25734 17502 25786 17554
rect 34862 17502 34914 17554
rect 15094 17390 15146 17442
rect 21366 17446 21418 17498
rect 48078 17502 48130 17554
rect 27750 17390 27802 17442
rect 44942 17390 44994 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 4342 17054 4394 17106
rect 16606 17054 16658 17106
rect 21198 17054 21250 17106
rect 23382 17054 23434 17106
rect 22542 16998 22594 17050
rect 23718 17054 23770 17106
rect 24334 17054 24386 17106
rect 25342 17054 25394 17106
rect 26686 17054 26738 17106
rect 27246 17054 27298 17106
rect 29430 17054 29482 17106
rect 12126 16942 12178 16994
rect 28478 16942 28530 16994
rect 5070 16830 5122 16882
rect 5182 16830 5234 16882
rect 8766 16830 8818 16882
rect 8990 16830 9042 16882
rect 9438 16830 9490 16882
rect 12910 16830 12962 16882
rect 13022 16830 13074 16882
rect 13358 16830 13410 16882
rect 16942 16830 16994 16882
rect 17614 16830 17666 16882
rect 17950 16874 18002 16926
rect 18924 16867 18976 16919
rect 19070 16830 19122 16882
rect 19182 16830 19234 16882
rect 20190 16886 20242 16938
rect 22206 16886 22258 16938
rect 19686 16830 19738 16882
rect 20414 16830 20466 16882
rect 3894 16718 3946 16770
rect 4734 16718 4786 16770
rect 5966 16718 6018 16770
rect 7870 16718 7922 16770
rect 10222 16718 10274 16770
rect 14142 16718 14194 16770
rect 16046 16718 16098 16770
rect 18062 16718 18114 16770
rect 20638 16718 20690 16770
rect 20806 16774 20858 16826
rect 21534 16830 21586 16882
rect 21758 16830 21810 16882
rect 22430 16830 22482 16882
rect 23886 16830 23938 16882
rect 23998 16830 24050 16882
rect 25678 16830 25730 16882
rect 26126 16830 26178 16882
rect 26350 16830 26402 16882
rect 27582 16830 27634 16882
rect 28310 16886 28362 16938
rect 28870 16942 28922 16994
rect 33182 16942 33234 16994
rect 34246 16998 34298 17050
rect 34694 16998 34746 17050
rect 40182 17054 40234 17106
rect 28142 16830 28194 16882
rect 28590 16830 28642 16882
rect 32622 16830 32674 16882
rect 33630 16886 33682 16938
rect 33854 16886 33906 16938
rect 37662 16942 37714 16994
rect 46510 16942 46562 16994
rect 33014 16830 33066 16882
rect 34414 16830 34466 16882
rect 34862 16850 34914 16902
rect 34974 16830 35026 16882
rect 38446 16830 38498 16882
rect 38558 16830 38610 16882
rect 38782 16830 38834 16882
rect 40910 16857 40962 16909
rect 43150 16830 43202 16882
rect 43822 16874 43874 16926
rect 44046 16830 44098 16882
rect 44382 16830 44434 16882
rect 44606 16830 44658 16882
rect 44886 16830 44938 16882
rect 45390 16863 45442 16915
rect 45614 16863 45666 16915
rect 46062 16863 46114 16915
rect 46372 16863 46424 16915
rect 46958 16830 47010 16882
rect 47294 16830 47346 16882
rect 47686 16830 47738 16882
rect 47966 16830 48018 16882
rect 48078 16830 48130 16882
rect 29934 16718 29986 16770
rect 31838 16718 31890 16770
rect 35758 16718 35810 16770
rect 43710 16718 43762 16770
rect 2270 16606 2322 16658
rect 3054 16606 3106 16658
rect 8486 16606 8538 16658
rect 12630 16606 12682 16658
rect 18510 16606 18562 16658
rect 46846 16662 46898 16714
rect 25958 16606 26010 16658
rect 38166 16606 38218 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 22990 16270 23042 16322
rect 25342 16270 25394 16322
rect 32510 16270 32562 16322
rect 44998 16270 45050 16322
rect 7198 16158 7250 16210
rect 8318 16158 8370 16210
rect 12462 16158 12514 16210
rect 14982 16158 15034 16210
rect 16046 16158 16098 16210
rect 16830 16158 16882 16210
rect 22038 16158 22090 16210
rect 2270 16046 2322 16098
rect 3054 16046 3106 16098
rect 5966 16046 6018 16098
rect 6414 16007 6466 16059
rect 6638 16046 6690 16098
rect 7310 16002 7362 16054
rect 7646 16046 7698 16098
rect 8430 16031 8482 16083
rect 8766 16046 8818 16098
rect 9326 16046 9378 16098
rect 10110 16046 10162 16098
rect 12574 16002 12626 16054
rect 12910 16046 12962 16098
rect 4958 15934 5010 15986
rect 12014 15934 12066 15986
rect 13414 15990 13466 16042
rect 13582 16046 13634 16098
rect 13806 16046 13858 16098
rect 14142 15990 14194 16042
rect 15598 16046 15650 16098
rect 15822 16046 15874 16098
rect 16158 16031 16210 16083
rect 16494 16046 16546 16098
rect 16942 16031 16994 16083
rect 17278 16046 17330 16098
rect 17838 16046 17890 16098
rect 19742 16018 19794 16070
rect 20302 16046 20354 16098
rect 21198 16046 21250 16098
rect 22318 16046 22370 16098
rect 22430 16046 22482 16098
rect 23326 16046 23378 16098
rect 22598 15990 22650 16042
rect 24894 16046 24946 16098
rect 25006 16046 25058 16098
rect 26238 16046 26290 16098
rect 26910 16046 26962 16098
rect 27582 16046 27634 16098
rect 28702 16046 28754 16098
rect 29486 16046 29538 16098
rect 29654 16102 29706 16154
rect 33742 16158 33794 16210
rect 29822 16046 29874 16098
rect 29934 16046 29986 16098
rect 30214 16046 30266 16098
rect 34694 16102 34746 16154
rect 36486 16158 36538 16210
rect 42926 16158 42978 16210
rect 43374 16158 43426 16210
rect 48134 16158 48186 16210
rect 31166 16018 31218 16070
rect 33574 16046 33626 16098
rect 33966 16046 34018 16098
rect 34190 16018 34242 16070
rect 35086 16046 35138 16098
rect 37214 16046 37266 16098
rect 37662 16046 37714 16098
rect 38446 16046 38498 16098
rect 41582 16046 41634 16098
rect 15318 15934 15370 15986
rect 6078 15878 6130 15930
rect 20470 15822 20522 15874
rect 21366 15822 21418 15874
rect 23662 15822 23714 15874
rect 24558 15822 24610 15874
rect 26070 15822 26122 15874
rect 26574 15822 26626 15874
rect 27246 15822 27298 15874
rect 27918 15822 27970 15874
rect 28534 15878 28586 15930
rect 34862 15934 34914 15986
rect 35422 15990 35474 16042
rect 41358 15990 41410 16042
rect 40350 15934 40402 15986
rect 41806 15934 41858 15986
rect 41974 15990 42026 16042
rect 42254 16046 42306 16098
rect 42366 16046 42418 16098
rect 42534 16046 42586 16098
rect 43486 16031 43538 16083
rect 43710 16046 43762 16098
rect 44046 16046 44098 16098
rect 44830 16046 44882 16098
rect 45390 15990 45442 16042
rect 45726 15990 45778 16042
rect 46174 15990 46226 16042
rect 46442 16006 46494 16058
rect 47070 16046 47122 16098
rect 47294 16046 47346 16098
rect 46622 15934 46674 15986
rect 47574 15934 47626 15986
rect 36038 15822 36090 15874
rect 37046 15822 37098 15874
rect 44214 15822 44266 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 3502 15486 3554 15538
rect 7142 15486 7194 15538
rect 5070 15430 5122 15482
rect 11790 15486 11842 15538
rect 13582 15486 13634 15538
rect 15766 15486 15818 15538
rect 16606 15486 16658 15538
rect 9662 15374 9714 15426
rect 16214 15374 16266 15426
rect 3838 15262 3890 15314
rect 4286 15262 4338 15314
rect 4510 15306 4562 15358
rect 4958 15262 5010 15314
rect 5294 15289 5346 15341
rect 5630 15262 5682 15314
rect 6190 15262 6242 15314
rect 6526 15277 6578 15329
rect 7310 15262 7362 15314
rect 7422 15262 7474 15314
rect 7758 15262 7810 15314
rect 8206 15262 8258 15314
rect 8318 15262 8370 15314
rect 8486 15262 8538 15314
rect 9494 15262 9546 15314
rect 10110 15290 10162 15342
rect 13134 15289 13186 15341
rect 13918 15262 13970 15314
rect 10334 15206 10386 15258
rect 14198 15262 14250 15314
rect 14758 15318 14810 15370
rect 21422 15374 21474 15426
rect 26182 15374 26234 15426
rect 27974 15374 28026 15426
rect 35646 15374 35698 15426
rect 36206 15374 36258 15426
rect 14478 15262 14530 15314
rect 14590 15262 14642 15314
rect 14926 15262 14978 15314
rect 16942 15262 16994 15314
rect 17502 15262 17554 15314
rect 18734 15262 18786 15314
rect 19518 15262 19570 15314
rect 21870 15262 21922 15314
rect 21982 15262 22034 15314
rect 22168 15300 22220 15352
rect 23774 15262 23826 15314
rect 23886 15262 23938 15314
rect 27246 15262 27298 15314
rect 27582 15262 27634 15314
rect 27694 15262 27746 15314
rect 4622 15150 4674 15202
rect 6638 15150 6690 15202
rect 8878 15150 8930 15202
rect 22542 15150 22594 15202
rect 23438 15150 23490 15202
rect 25734 15150 25786 15202
rect 26630 15150 26682 15202
rect 27414 15206 27466 15258
rect 28534 15262 28586 15314
rect 28926 15262 28978 15314
rect 29262 15262 29314 15314
rect 29374 15262 29426 15314
rect 30382 15289 30434 15341
rect 36766 15318 36818 15370
rect 29094 15206 29146 15258
rect 32958 15262 33010 15314
rect 33742 15262 33794 15314
rect 36878 15318 36930 15370
rect 37382 15374 37434 15426
rect 45614 15374 45666 15426
rect 29654 15150 29706 15202
rect 36038 15206 36090 15258
rect 37550 15262 37602 15314
rect 40910 15262 40962 15314
rect 41918 15262 41970 15314
rect 42646 15318 42698 15370
rect 42254 15262 42306 15314
rect 42926 15262 42978 15314
rect 43262 15262 43314 15314
rect 43374 15262 43426 15314
rect 43520 15299 43572 15351
rect 44494 15262 44546 15314
rect 44718 15306 44770 15358
rect 47518 15262 47570 15314
rect 48302 15262 48354 15314
rect 38334 15150 38386 15202
rect 40238 15150 40290 15202
rect 41246 15150 41298 15202
rect 42590 15150 42642 15202
rect 43934 15150 43986 15202
rect 44830 15150 44882 15202
rect 24222 15038 24274 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 11342 14702 11394 14754
rect 12854 14702 12906 14754
rect 23326 14702 23378 14754
rect 23998 14702 24050 14754
rect 28534 14702 28586 14754
rect 30494 14702 30546 14754
rect 43150 14702 43202 14754
rect 5742 14590 5794 14642
rect 9662 14590 9714 14642
rect 10222 14590 10274 14642
rect 16046 14590 16098 14642
rect 17950 14590 18002 14642
rect 18398 14590 18450 14642
rect 22150 14590 22202 14642
rect 36318 14590 36370 14642
rect 38110 14590 38162 14642
rect 2046 14478 2098 14530
rect 2830 14478 2882 14530
rect 4734 14478 4786 14530
rect 5854 14463 5906 14515
rect 6078 14478 6130 14530
rect 6526 14478 6578 14530
rect 8094 14478 8146 14530
rect 6806 14422 6858 14474
rect 8766 14478 8818 14530
rect 9438 14478 9490 14530
rect 9102 14422 9154 14474
rect 9830 14422 9882 14474
rect 10616 14478 10668 14530
rect 10782 14478 10834 14530
rect 10894 14478 10946 14530
rect 11585 14478 11637 14530
rect 12462 14478 12514 14530
rect 12686 14478 12738 14530
rect 14030 14478 14082 14530
rect 14254 14422 14306 14474
rect 14366 14422 14418 14474
rect 14926 14366 14978 14418
rect 15094 14422 15146 14474
rect 15262 14478 15314 14530
rect 18510 14463 18562 14515
rect 18734 14478 18786 14530
rect 19518 14478 19570 14530
rect 20190 14478 20242 14530
rect 21758 14478 21810 14530
rect 22318 14478 22370 14530
rect 22990 14478 23042 14530
rect 23662 14478 23714 14530
rect 24334 14478 24386 14530
rect 24670 14478 24722 14530
rect 25902 14478 25954 14530
rect 26686 14478 26738 14530
rect 26854 14478 26906 14530
rect 27134 14478 27186 14530
rect 27806 14478 27858 14530
rect 28254 14478 28306 14530
rect 6638 14310 6690 14362
rect 26238 14366 26290 14418
rect 27022 14366 27074 14418
rect 27974 14422 28026 14474
rect 29150 14478 29202 14530
rect 29318 14534 29370 14586
rect 44158 14646 44210 14698
rect 39230 14590 39282 14642
rect 45166 14590 45218 14642
rect 46566 14590 46618 14642
rect 46846 14646 46898 14698
rect 47798 14590 47850 14642
rect 29598 14478 29650 14530
rect 30158 14478 30210 14530
rect 30942 14450 30994 14502
rect 33182 14478 33234 14530
rect 33630 14478 33682 14530
rect 34414 14478 34466 14530
rect 37214 14478 37266 14530
rect 38334 14478 38386 14530
rect 39454 14478 39506 14530
rect 40462 14478 40514 14530
rect 41134 14478 41186 14530
rect 41694 14478 41746 14530
rect 42366 14478 42418 14530
rect 27414 14366 27466 14418
rect 28142 14366 28194 14418
rect 29486 14366 29538 14418
rect 29878 14366 29930 14418
rect 37942 14422 37994 14474
rect 38558 14422 38610 14474
rect 39062 14422 39114 14474
rect 39678 14422 39730 14474
rect 42030 14422 42082 14474
rect 42814 14478 42866 14530
rect 43934 14478 43986 14530
rect 44270 14478 44322 14530
rect 44830 14478 44882 14530
rect 45502 14478 45554 14530
rect 45166 14422 45218 14474
rect 45838 14478 45890 14530
rect 46958 14478 47010 14530
rect 47294 14478 47346 14530
rect 7758 14254 7810 14306
rect 8430 14254 8482 14306
rect 13862 14254 13914 14306
rect 19350 14254 19402 14306
rect 19854 14254 19906 14306
rect 20526 14254 20578 14306
rect 21422 14254 21474 14306
rect 22654 14254 22706 14306
rect 25734 14254 25786 14306
rect 37046 14254 37098 14306
rect 37718 14254 37770 14306
rect 40294 14310 40346 14362
rect 40966 14310 41018 14362
rect 42478 14310 42530 14362
rect 48246 14254 48298 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 3166 13918 3218 13970
rect 4902 13918 4954 13970
rect 5406 13918 5458 13970
rect 22934 13918 22986 13970
rect 5966 13862 6018 13914
rect 28870 13918 28922 13970
rect 29318 13918 29370 13970
rect 39958 13918 40010 13970
rect 41414 13918 41466 13970
rect 48134 13918 48186 13970
rect 16718 13806 16770 13858
rect 3502 13694 3554 13746
rect 5070 13694 5122 13746
rect 5854 13694 5906 13746
rect 6302 13733 6354 13785
rect 6526 13694 6578 13746
rect 7758 13694 7810 13746
rect 8430 13694 8482 13746
rect 8542 13694 8594 13746
rect 10076 13732 10128 13784
rect 30606 13806 30658 13858
rect 10222 13694 10274 13746
rect 10334 13694 10386 13746
rect 10558 13694 10610 13746
rect 11566 13694 11618 13746
rect 12350 13694 12402 13746
rect 14254 13694 14306 13746
rect 15150 13722 15202 13774
rect 15374 13694 15426 13746
rect 15766 13694 15818 13746
rect 16158 13732 16210 13784
rect 16494 13694 16546 13746
rect 8878 13582 8930 13634
rect 9662 13582 9714 13634
rect 15598 13582 15650 13634
rect 16886 13638 16938 13690
rect 17614 13694 17666 13746
rect 21142 13750 21194 13802
rect 17838 13694 17890 13746
rect 18118 13694 18170 13746
rect 18622 13694 18674 13746
rect 18958 13694 19010 13746
rect 19518 13694 19570 13746
rect 19854 13694 19906 13746
rect 20862 13694 20914 13746
rect 20974 13694 21026 13746
rect 21310 13694 21362 13746
rect 21982 13694 22034 13746
rect 22094 13694 22146 13746
rect 22262 13638 22314 13690
rect 22430 13694 22482 13746
rect 24222 13694 24274 13746
rect 25230 13694 25282 13746
rect 25566 13694 25618 13746
rect 25678 13694 25730 13746
rect 26350 13694 26402 13746
rect 26686 13694 26738 13746
rect 27022 13694 27074 13746
rect 25398 13638 25450 13690
rect 29486 13694 29538 13746
rect 30438 13750 30490 13802
rect 32118 13806 32170 13858
rect 30270 13694 30322 13746
rect 30718 13694 30770 13746
rect 31390 13694 31442 13746
rect 31726 13694 31778 13746
rect 31838 13694 31890 13746
rect 7422 13470 7474 13522
rect 8094 13470 8146 13522
rect 10894 13470 10946 13522
rect 18510 13526 18562 13578
rect 19406 13526 19458 13578
rect 20582 13470 20634 13522
rect 21702 13470 21754 13522
rect 23886 13470 23938 13522
rect 25958 13470 26010 13522
rect 26798 13526 26850 13578
rect 27358 13582 27410 13634
rect 31558 13638 31610 13690
rect 32958 13694 33010 13746
rect 36038 13750 36090 13802
rect 36206 13806 36258 13858
rect 38726 13806 38778 13858
rect 43038 13806 43090 13858
rect 36654 13722 36706 13774
rect 36878 13750 36930 13802
rect 37438 13722 37490 13774
rect 37214 13638 37266 13690
rect 33742 13582 33794 13634
rect 35646 13582 35698 13634
rect 37886 13582 37938 13634
rect 38054 13638 38106 13690
rect 38222 13694 38274 13746
rect 38446 13694 38498 13746
rect 42142 13694 42194 13746
rect 42478 13732 42530 13784
rect 43206 13750 43258 13802
rect 45222 13806 45274 13858
rect 42814 13694 42866 13746
rect 43598 13738 43650 13790
rect 43822 13694 43874 13746
rect 44494 13694 44546 13746
rect 44830 13694 44882 13746
rect 44942 13694 44994 13746
rect 45726 13694 45778 13746
rect 45950 13694 46002 13746
rect 46286 13694 46338 13746
rect 39286 13582 39338 13634
rect 44662 13638 44714 13690
rect 46510 13694 46562 13746
rect 47294 13694 47346 13746
rect 47518 13694 47570 13746
rect 40406 13582 40458 13634
rect 43486 13582 43538 13634
rect 29822 13470 29874 13522
rect 30998 13470 31050 13522
rect 45726 13526 45778 13578
rect 47294 13526 47346 13578
rect 41806 13470 41858 13522
rect 46790 13470 46842 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 15150 13134 15202 13186
rect 19854 13134 19906 13186
rect 27078 13134 27130 13186
rect 33070 13134 33122 13186
rect 34694 13134 34746 13186
rect 36206 13134 36258 13186
rect 6862 13022 6914 13074
rect 8094 13022 8146 13074
rect 11342 13022 11394 13074
rect 12966 13022 13018 13074
rect 16270 13022 16322 13074
rect 18174 13022 18226 13074
rect 18790 13022 18842 13074
rect 19462 13022 19514 13074
rect 5182 12910 5234 12962
rect 5630 12910 5682 12962
rect 6302 12910 6354 12962
rect 6078 12854 6130 12906
rect 6974 12866 7026 12918
rect 7198 12910 7250 12962
rect 7646 12910 7698 12962
rect 7982 12895 8034 12947
rect 8430 12910 8482 12962
rect 12126 12910 12178 12962
rect 13470 12910 13522 12962
rect 14030 12910 14082 12962
rect 14906 12910 14958 12962
rect 15486 12910 15538 12962
rect 20190 12910 20242 12962
rect 20302 12910 20354 12962
rect 20638 12910 20690 12962
rect 21310 12910 21362 12962
rect 21478 12966 21530 13018
rect 21758 12910 21810 12962
rect 22766 12910 22818 12962
rect 22878 12910 22930 12962
rect 23214 12910 23266 12962
rect 9438 12798 9490 12850
rect 5742 12742 5794 12794
rect 4846 12686 4898 12738
rect 8766 12686 8818 12738
rect 12518 12686 12570 12738
rect 13638 12742 13690 12794
rect 21646 12798 21698 12850
rect 22038 12798 22090 12850
rect 23046 12854 23098 12906
rect 23438 12910 23490 12962
rect 24446 12910 24498 12962
rect 24782 12910 24834 12962
rect 24894 12910 24946 12962
rect 24614 12854 24666 12906
rect 30550 12966 30602 13018
rect 31838 13022 31890 13074
rect 34134 13022 34186 13074
rect 37662 13022 37714 13074
rect 38670 13022 38722 13074
rect 41694 13022 41746 13074
rect 42590 13022 42642 13074
rect 48078 13022 48130 13074
rect 25174 12910 25226 12962
rect 26910 12910 26962 12962
rect 29598 12910 29650 12962
rect 30942 12910 30994 12962
rect 29430 12854 29482 12906
rect 22486 12798 22538 12850
rect 29822 12798 29874 12850
rect 29990 12854 30042 12906
rect 31166 12882 31218 12934
rect 31670 12910 31722 12962
rect 32062 12910 32114 12962
rect 32398 12872 32450 12924
rect 32734 12910 32786 12962
rect 33742 12910 33794 12962
rect 34974 12910 35026 12962
rect 35198 12910 35250 12962
rect 36542 12910 36594 12962
rect 37326 12910 37378 12962
rect 37550 12866 37602 12918
rect 37886 12910 37938 12962
rect 41022 12910 41074 12962
rect 41134 12910 41186 12962
rect 42142 12910 42194 12962
rect 30718 12798 30770 12850
rect 41300 12854 41352 12906
rect 42478 12866 42530 12918
rect 43393 12910 43445 12962
rect 44270 12910 44322 12962
rect 44718 12910 44770 12962
rect 45390 12910 45442 12962
rect 46174 12910 46226 12962
rect 23774 12686 23826 12738
rect 27638 12686 27690 12738
rect 33574 12742 33626 12794
rect 40574 12798 40626 12850
rect 43150 12798 43202 12850
rect 35814 12686 35866 12738
rect 45054 12686 45106 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 15318 12350 15370 12402
rect 16886 12350 16938 12402
rect 18566 12350 18618 12402
rect 23998 12350 24050 12402
rect 26014 12350 26066 12402
rect 32342 12350 32394 12402
rect 33462 12350 33514 12402
rect 35758 12350 35810 12402
rect 36486 12350 36538 12402
rect 43878 12350 43930 12402
rect 6638 12238 6690 12290
rect 3950 12126 4002 12178
rect 4734 12126 4786 12178
rect 8094 12126 8146 12178
rect 8654 12141 8706 12193
rect 8990 12126 9042 12178
rect 9550 12126 9602 12178
rect 9662 12126 9714 12178
rect 9848 12164 9900 12216
rect 10782 12126 10834 12178
rect 13918 12182 13970 12234
rect 14030 12182 14082 12234
rect 14758 12182 14810 12234
rect 15710 12126 15762 12178
rect 16046 12126 16098 12178
rect 17502 12126 17554 12178
rect 17726 12126 17778 12178
rect 19070 12154 19122 12206
rect 19686 12182 19738 12234
rect 22094 12238 22146 12290
rect 23214 12238 23266 12290
rect 19294 12126 19346 12178
rect 19854 12126 19906 12178
rect 22262 12182 22314 12234
rect 34862 12238 34914 12290
rect 21982 12126 22034 12178
rect 22430 12126 22482 12178
rect 23382 12182 23434 12234
rect 38558 12238 38610 12290
rect 48134 12238 48186 12290
rect 23102 12126 23154 12178
rect 23550 12126 23602 12178
rect 24334 12126 24386 12178
rect 25678 12126 25730 12178
rect 26350 12126 26402 12178
rect 27694 12126 27746 12178
rect 28478 12126 28530 12178
rect 30830 12126 30882 12178
rect 30942 12126 30994 12178
rect 31108 12126 31160 12178
rect 32510 12126 32562 12178
rect 33854 12141 33906 12193
rect 34190 12126 34242 12178
rect 34526 12126 34578 12178
rect 7254 12014 7306 12066
rect 8542 12014 8594 12066
rect 10222 12014 10274 12066
rect 11566 12014 11618 12066
rect 13470 12014 13522 12066
rect 14590 12014 14642 12066
rect 7758 11902 7810 11954
rect 15598 11958 15650 12010
rect 17390 11958 17442 12010
rect 19518 12014 19570 12066
rect 20806 12014 20858 12066
rect 21254 12014 21306 12066
rect 34694 12070 34746 12122
rect 34974 12126 35026 12178
rect 36094 12126 36146 12178
rect 37158 12182 37210 12234
rect 36990 12126 37042 12178
rect 37326 12126 37378 12178
rect 37438 12126 37490 12178
rect 37718 12126 37770 12178
rect 38446 12126 38498 12178
rect 27302 12014 27354 12066
rect 30382 12014 30434 12066
rect 31502 12014 31554 12066
rect 33742 12014 33794 12066
rect 38726 12070 38778 12122
rect 38894 12126 38946 12178
rect 39958 12126 40010 12178
rect 40238 12126 40290 12178
rect 40350 12126 40402 12178
rect 41022 12126 41074 12178
rect 41246 12170 41298 12222
rect 41806 12141 41858 12193
rect 42030 12126 42082 12178
rect 42590 12126 42642 12178
rect 42702 12126 42754 12178
rect 42888 12164 42940 12216
rect 44942 12126 44994 12178
rect 45390 12182 45442 12234
rect 45838 12182 45890 12234
rect 46174 12182 46226 12234
rect 45166 12126 45218 12178
rect 46484 12166 46536 12218
rect 47070 12126 47122 12178
rect 47294 12126 47346 12178
rect 47630 12126 47682 12178
rect 47854 12126 47906 12178
rect 39398 12014 39450 12066
rect 41358 12014 41410 12066
rect 41694 12014 41746 12066
rect 43262 12014 43314 12066
rect 44326 12014 44378 12066
rect 46510 12014 46562 12066
rect 20190 11902 20242 11954
rect 21702 11902 21754 11954
rect 22822 11902 22874 11954
rect 26686 11902 26738 11954
rect 35254 11902 35306 11954
rect 46958 11958 47010 12010
rect 38166 11902 38218 11954
rect 44662 11902 44714 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 15990 11566 16042 11618
rect 5126 11454 5178 11506
rect 6078 11454 6130 11506
rect 6862 11454 6914 11506
rect 9718 11454 9770 11506
rect 20694 11510 20746 11562
rect 22598 11566 22650 11618
rect 26126 11566 26178 11618
rect 30438 11566 30490 11618
rect 13750 11454 13802 11506
rect 17166 11454 17218 11506
rect 19518 11454 19570 11506
rect 1822 11342 1874 11394
rect 2606 11342 2658 11394
rect 4510 11342 4562 11394
rect 5630 11342 5682 11394
rect 5966 11298 6018 11350
rect 6414 11342 6466 11394
rect 6750 11327 6802 11379
rect 7534 11342 7586 11394
rect 7870 11342 7922 11394
rect 8542 11342 8594 11394
rect 9102 11342 9154 11394
rect 10110 11342 10162 11394
rect 10894 11342 10946 11394
rect 8934 11286 8986 11338
rect 14030 11309 14082 11361
rect 14366 11286 14418 11338
rect 14814 11309 14866 11361
rect 15124 11309 15176 11361
rect 16270 11342 16322 11394
rect 21310 11398 21362 11450
rect 22150 11398 22202 11450
rect 23158 11454 23210 11506
rect 26910 11510 26962 11562
rect 35478 11566 35530 11618
rect 16382 11342 16434 11394
rect 16718 11342 16770 11394
rect 17054 11327 17106 11379
rect 20302 11342 20354 11394
rect 20526 11342 20578 11394
rect 21422 11304 21474 11356
rect 22430 11342 22482 11394
rect 24054 11342 24106 11394
rect 24334 11342 24386 11394
rect 24502 11398 24554 11450
rect 25622 11454 25674 11506
rect 31502 11454 31554 11506
rect 33406 11454 33458 11506
rect 34022 11454 34074 11506
rect 24782 11342 24834 11394
rect 34302 11398 34354 11450
rect 26462 11342 26514 11394
rect 26686 11342 26738 11394
rect 27022 11342 27074 11394
rect 30606 11321 30658 11373
rect 30718 11342 30770 11394
rect 34974 11342 35026 11394
rect 35142 11398 35194 11450
rect 12798 11230 12850 11282
rect 8542 11174 8594 11226
rect 15262 11230 15314 11282
rect 17614 11230 17666 11282
rect 21982 11230 22034 11282
rect 24670 11230 24722 11282
rect 25062 11230 25114 11282
rect 34526 11286 34578 11338
rect 35758 11342 35810 11394
rect 36038 11398 36090 11450
rect 40070 11454 40122 11506
rect 42926 11510 42978 11562
rect 47182 11566 47234 11618
rect 36206 11342 36258 11394
rect 37438 11342 37490 11394
rect 37550 11342 37602 11394
rect 38222 11342 38274 11394
rect 41190 11398 41242 11450
rect 46510 11454 46562 11506
rect 47966 11454 48018 11506
rect 38894 11342 38946 11394
rect 40798 11342 40850 11394
rect 41694 11342 41746 11394
rect 30102 11230 30154 11282
rect 40574 11286 40626 11338
rect 43206 11398 43258 11450
rect 41806 11342 41858 11394
rect 42590 11342 42642 11394
rect 42814 11342 42866 11394
rect 43598 11342 43650 11394
rect 43822 11314 43874 11366
rect 45390 11309 45442 11361
rect 45838 11305 45890 11357
rect 46174 11309 46226 11361
rect 46484 11302 46536 11354
rect 46846 11342 46898 11394
rect 48302 11342 48354 11394
rect 35870 11230 35922 11282
rect 41022 11230 41074 11282
rect 42086 11230 42138 11282
rect 43374 11230 43426 11282
rect 27638 11118 27690 11170
rect 28646 11118 28698 11170
rect 29654 11118 29706 11170
rect 37102 11118 37154 11170
rect 37886 11118 37938 11170
rect 38558 11118 38610 11170
rect 39230 11118 39282 11170
rect 44998 11118 45050 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 2942 10782 2994 10834
rect 10838 10782 10890 10834
rect 5070 10726 5122 10778
rect 9662 10726 9714 10778
rect 11286 10782 11338 10834
rect 11734 10782 11786 10834
rect 12182 10782 12234 10834
rect 12630 10782 12682 10834
rect 15766 10782 15818 10834
rect 17558 10782 17610 10834
rect 19014 10782 19066 10834
rect 23102 10782 23154 10834
rect 25454 10782 25506 10834
rect 26070 10782 26122 10834
rect 15206 10670 15258 10722
rect 17894 10670 17946 10722
rect 26686 10670 26738 10722
rect 32342 10726 32394 10778
rect 36990 10782 37042 10834
rect 39006 10782 39058 10834
rect 39622 10782 39674 10834
rect 2606 10558 2658 10610
rect 3278 10558 3330 10610
rect 4174 10558 4226 10610
rect 4398 10602 4450 10654
rect 4846 10558 4898 10610
rect 5182 10585 5234 10637
rect 5518 10558 5570 10610
rect 6190 10558 6242 10610
rect 8878 10558 8930 10610
rect 9550 10558 9602 10610
rect 9942 10587 9994 10639
rect 13022 10558 13074 10610
rect 13246 10558 13298 10610
rect 13694 10558 13746 10610
rect 13806 10558 13858 10610
rect 13964 10608 14016 10660
rect 14702 10558 14754 10610
rect 14926 10558 14978 10610
rect 16158 10596 16210 10648
rect 16886 10614 16938 10666
rect 16494 10558 16546 10610
rect 18174 10558 18226 10610
rect 18286 10558 18338 10610
rect 18846 10558 18898 10610
rect 21758 10558 21810 10610
rect 22542 10558 22594 10610
rect 23438 10558 23490 10610
rect 24782 10558 24834 10610
rect 25118 10558 25170 10610
rect 26518 10614 26570 10666
rect 35646 10670 35698 10722
rect 43486 10670 43538 10722
rect 44046 10670 44098 10722
rect 26350 10558 26402 10610
rect 26798 10558 26850 10610
rect 27638 10558 27690 10610
rect 28030 10558 28082 10610
rect 31652 10596 31704 10648
rect 31838 10558 31890 10610
rect 31950 10558 32002 10610
rect 32510 10558 32562 10610
rect 32958 10558 33010 10610
rect 33742 10558 33794 10610
rect 35982 10558 36034 10610
rect 36654 10558 36706 10610
rect 37326 10558 37378 10610
rect 37998 10558 38050 10610
rect 38670 10558 38722 10610
rect 40238 10558 40290 10610
rect 40350 10558 40402 10610
rect 40798 10558 40850 10610
rect 41582 10558 41634 10610
rect 45950 10558 46002 10610
rect 46734 10558 46786 10610
rect 47070 10558 47122 10610
rect 47294 10558 47346 10610
rect 47742 10558 47794 10610
rect 47854 10558 47906 10610
rect 48134 10558 48186 10610
rect 4510 10446 4562 10498
rect 6974 10446 7026 10498
rect 2270 10334 2322 10386
rect 13358 10390 13410 10442
rect 14366 10446 14418 10498
rect 16718 10446 16770 10498
rect 19854 10446 19906 10498
rect 28814 10446 28866 10498
rect 30718 10446 30770 10498
rect 24446 10334 24498 10386
rect 27078 10334 27130 10386
rect 31278 10334 31330 10386
rect 36318 10334 36370 10386
rect 37662 10334 37714 10386
rect 46958 10390 47010 10442
rect 38334 10334 38386 10386
rect 39958 10334 40010 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 8206 9998 8258 10050
rect 13526 9998 13578 10050
rect 14366 9998 14418 10050
rect 39734 9998 39786 10050
rect 2382 9886 2434 9938
rect 7310 9886 7362 9938
rect 8878 9886 8930 9938
rect 10502 9886 10554 9938
rect 11398 9886 11450 9938
rect 16382 9886 16434 9938
rect 1598 9774 1650 9826
rect 4286 9774 4338 9826
rect 5182 9774 5234 9826
rect 5630 9774 5682 9826
rect 6302 9774 6354 9826
rect 6862 9774 6914 9826
rect 5966 9718 6018 9770
rect 7198 9730 7250 9782
rect 8542 9774 8594 9826
rect 8990 9730 9042 9782
rect 9214 9774 9266 9826
rect 10110 9774 10162 9826
rect 11846 9718 11898 9770
rect 12126 9741 12178 9793
rect 13806 9774 13858 9826
rect 12574 9718 12626 9770
rect 12910 9718 12962 9770
rect 14030 9774 14082 9826
rect 14926 9774 14978 9826
rect 15038 9774 15090 9826
rect 14758 9718 14810 9770
rect 15598 9774 15650 9826
rect 19574 9830 19626 9882
rect 20806 9830 20858 9882
rect 11678 9662 11730 9714
rect 5742 9606 5794 9658
rect 18286 9662 18338 9714
rect 18734 9718 18786 9770
rect 18846 9736 18898 9788
rect 20078 9736 20130 9788
rect 20414 9774 20466 9826
rect 22710 9830 22762 9882
rect 22430 9774 22482 9826
rect 22542 9774 22594 9826
rect 22878 9774 22930 9826
rect 23214 9774 23266 9826
rect 23382 9830 23434 9882
rect 27918 9886 27970 9938
rect 29822 9886 29874 9938
rect 23662 9774 23714 9826
rect 24222 9774 24274 9826
rect 25454 9774 25506 9826
rect 29150 9830 29202 9882
rect 29990 9830 30042 9882
rect 30550 9886 30602 9938
rect 32790 9886 32842 9938
rect 33238 9886 33290 9938
rect 34134 9886 34186 9938
rect 35086 9886 35138 9938
rect 36094 9886 36146 9938
rect 37606 9886 37658 9938
rect 38110 9886 38162 9938
rect 38558 9942 38610 9994
rect 43374 9998 43426 10050
rect 40910 9942 40962 9994
rect 41918 9942 41970 9994
rect 45054 9998 45106 10050
rect 42646 9886 42698 9938
rect 44102 9886 44154 9938
rect 46174 9886 46226 9938
rect 48078 9886 48130 9938
rect 27246 9774 27298 9826
rect 27358 9774 27410 9826
rect 31278 9774 31330 9826
rect 19406 9662 19458 9714
rect 20638 9662 20690 9714
rect 22150 9662 22202 9714
rect 23550 9662 23602 9714
rect 27524 9718 27576 9770
rect 29430 9718 29482 9770
rect 30942 9718 30994 9770
rect 23942 9662 23994 9714
rect 31502 9662 31554 9714
rect 31670 9718 31722 9770
rect 31838 9774 31890 9826
rect 34414 9774 34466 9826
rect 34526 9774 34578 9826
rect 34694 9774 34746 9826
rect 35646 9774 35698 9826
rect 35982 9759 36034 9811
rect 37774 9774 37826 9826
rect 38670 9774 38722 9826
rect 39006 9774 39058 9826
rect 39230 9774 39282 9826
rect 39454 9774 39506 9826
rect 40686 9774 40738 9826
rect 41022 9774 41074 9826
rect 41358 9774 41410 9826
rect 41694 9774 41746 9826
rect 42030 9774 42082 9826
rect 43710 9774 43762 9826
rect 44718 9774 44770 9826
rect 45390 9774 45442 9826
rect 4846 9550 4898 9602
rect 9774 9550 9826 9602
rect 21478 9550 21530 9602
rect 24558 9550 24610 9602
rect 25790 9550 25842 9602
rect 26518 9550 26570 9602
rect 26966 9550 27018 9602
rect 28646 9550 28698 9602
rect 32174 9550 32226 9602
rect 33686 9550 33738 9602
rect 37158 9550 37210 9602
rect 40350 9550 40402 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 10502 9214 10554 9266
rect 5742 9158 5794 9210
rect 8878 9158 8930 9210
rect 15038 9214 15090 9266
rect 15598 9214 15650 9266
rect 17670 9214 17722 9266
rect 18118 9214 18170 9266
rect 18678 9214 18730 9266
rect 22990 9214 23042 9266
rect 33686 9214 33738 9266
rect 34134 9214 34186 9266
rect 44550 9214 44602 9266
rect 47126 9214 47178 9266
rect 47574 9214 47626 9266
rect 48246 9214 48298 9266
rect 13358 9102 13410 9154
rect 1598 8990 1650 9042
rect 5462 9046 5514 9098
rect 16774 9102 16826 9154
rect 24334 9102 24386 9154
rect 36486 9102 36538 9154
rect 4286 8990 4338 9042
rect 5294 8990 5346 9042
rect 5854 8990 5906 9042
rect 6414 8990 6466 9042
rect 6750 9034 6802 9086
rect 7422 9005 7474 9057
rect 7758 8990 7810 9042
rect 8206 8990 8258 9042
rect 8430 9017 8482 9069
rect 8766 8990 8818 9042
rect 9438 8990 9490 9042
rect 10670 8990 10722 9042
rect 11454 8990 11506 9042
rect 13918 8990 13970 9042
rect 14254 8990 14306 9042
rect 14702 8990 14754 9042
rect 15934 8990 15986 9042
rect 18510 8990 18562 9042
rect 21198 8990 21250 9042
rect 21982 8990 22034 9042
rect 22374 8990 22426 9042
rect 22654 8990 22706 9042
rect 24502 9046 24554 9098
rect 39342 9102 39394 9154
rect 40294 9102 40346 9154
rect 41134 9102 41186 9154
rect 24222 8990 24274 9042
rect 24670 8990 24722 9042
rect 25790 8990 25842 9042
rect 26014 8990 26066 9042
rect 26462 8990 26514 9042
rect 26630 8990 26682 9042
rect 26798 8990 26850 9042
rect 26910 8990 26962 9042
rect 27806 8990 27858 9042
rect 30830 8990 30882 9042
rect 32232 8990 32284 9042
rect 32398 8990 32450 9042
rect 32510 8990 32562 9042
rect 33294 8990 33346 9042
rect 34638 8990 34690 9042
rect 34974 9034 35026 9086
rect 35310 8990 35362 9042
rect 35534 8990 35586 9042
rect 36654 8990 36706 9042
rect 39902 8990 39954 9042
rect 40014 8990 40066 9042
rect 43822 8990 43874 9042
rect 45278 8990 45330 9042
rect 45614 8990 45666 9042
rect 46286 8990 46338 9042
rect 46622 8990 46674 9042
rect 2382 8878 2434 8930
rect 4902 8878 4954 8930
rect 6862 8878 6914 8930
rect 7310 8878 7362 8930
rect 9774 8766 9826 8818
rect 13806 8822 13858 8874
rect 16326 8878 16378 8930
rect 19294 8878 19346 8930
rect 25398 8878 25450 8930
rect 28590 8878 28642 8930
rect 30494 8878 30546 8930
rect 31838 8878 31890 8930
rect 23942 8766 23994 8818
rect 25678 8822 25730 8874
rect 35086 8878 35138 8930
rect 37438 8878 37490 8930
rect 43038 8878 43090 8930
rect 45110 8878 45162 8930
rect 27190 8766 27242 8818
rect 31166 8766 31218 8818
rect 33126 8822 33178 8874
rect 46174 8822 46226 8874
rect 35814 8766 35866 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 2718 8430 2770 8482
rect 3558 8318 3610 8370
rect 4286 8318 4338 8370
rect 5070 8318 5122 8370
rect 6862 8318 6914 8370
rect 8654 8318 8706 8370
rect 11006 8318 11058 8370
rect 12182 8318 12234 8370
rect 13470 8374 13522 8426
rect 20470 8430 20522 8482
rect 27582 8430 27634 8482
rect 27806 8430 27858 8482
rect 14926 8318 14978 8370
rect 15542 8318 15594 8370
rect 18062 8318 18114 8370
rect 3054 8206 3106 8258
rect 3838 8206 3890 8258
rect 4622 8206 4674 8258
rect 4118 8150 4170 8202
rect 4958 8191 5010 8243
rect 5630 8206 5682 8258
rect 6078 8167 6130 8219
rect 6302 8206 6354 8258
rect 6974 8191 7026 8243
rect 7198 8206 7250 8258
rect 8206 8206 8258 8258
rect 8542 8162 8594 8214
rect 9102 8206 9154 8258
rect 11790 8206 11842 8258
rect 12518 8206 12570 8258
rect 12798 8206 12850 8258
rect 13022 8206 13074 8258
rect 13582 8206 13634 8258
rect 13806 8206 13858 8258
rect 14478 8206 14530 8258
rect 14814 8162 14866 8214
rect 18846 8206 18898 8258
rect 19238 8206 19290 8258
rect 19686 8206 19738 8258
rect 21254 8262 21306 8314
rect 20134 8206 20186 8258
rect 20302 8206 20354 8258
rect 21870 8178 21922 8230
rect 16158 8094 16210 8146
rect 5742 8038 5794 8090
rect 21422 8094 21474 8146
rect 22094 8150 22146 8202
rect 22318 8206 22370 8258
rect 23102 8206 23154 8258
rect 25454 8206 25506 8258
rect 25790 8206 25842 8258
rect 25902 8206 25954 8258
rect 25622 8150 25674 8202
rect 26574 8206 26626 8258
rect 26742 8262 26794 8314
rect 28478 8318 28530 8370
rect 30102 8318 30154 8370
rect 31502 8318 31554 8370
rect 35310 8318 35362 8370
rect 37158 8318 37210 8370
rect 38110 8318 38162 8370
rect 26910 8206 26962 8258
rect 27022 8206 27074 8258
rect 28142 8206 28194 8258
rect 29150 8206 29202 8258
rect 30718 8206 30770 8258
rect 34190 8206 34242 8258
rect 38278 8262 38330 8314
rect 39566 8318 39618 8370
rect 40014 8318 40066 8370
rect 41806 8318 41858 8370
rect 34414 8206 34466 8258
rect 34694 8206 34746 8258
rect 35422 8162 35474 8214
rect 35646 8206 35698 8258
rect 35982 8206 36034 8258
rect 37550 8168 37602 8220
rect 37886 8206 37938 8258
rect 41974 8262 42026 8314
rect 38894 8206 38946 8258
rect 39006 8206 39058 8258
rect 25006 8094 25058 8146
rect 26182 8094 26234 8146
rect 27302 8094 27354 8146
rect 30550 8094 30602 8146
rect 39172 8150 39224 8202
rect 40126 8162 40178 8214
rect 40462 8206 40514 8258
rect 41582 8206 41634 8258
rect 41414 8150 41466 8202
rect 43038 8150 43090 8202
rect 43318 8150 43370 8202
rect 43766 8150 43818 8202
rect 44132 8173 44184 8225
rect 44718 8206 44770 8258
rect 45502 8206 45554 8258
rect 48302 8206 48354 8258
rect 33406 8094 33458 8146
rect 44270 8094 44322 8146
rect 47406 8094 47458 8146
rect 27974 7982 28026 8034
rect 29486 7982 29538 8034
rect 34022 7982 34074 8034
rect 36318 7982 36370 8034
rect 42422 7982 42474 8034
rect 47966 7982 48018 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 12070 7646 12122 7698
rect 6974 7590 7026 7642
rect 7534 7590 7586 7642
rect 9774 7590 9826 7642
rect 17558 7646 17610 7698
rect 22150 7646 22202 7698
rect 23774 7646 23826 7698
rect 26742 7646 26794 7698
rect 30214 7646 30266 7698
rect 5966 7534 6018 7586
rect 3278 7422 3330 7474
rect 6750 7466 6802 7518
rect 7086 7422 7138 7474
rect 7646 7422 7698 7474
rect 7982 7449 8034 7501
rect 9886 7478 9938 7530
rect 8318 7422 8370 7474
rect 9550 7422 9602 7474
rect 10222 7422 10274 7474
rect 10894 7466 10946 7518
rect 11118 7422 11170 7474
rect 12686 7422 12738 7474
rect 12910 7422 12962 7474
rect 13470 7422 13522 7474
rect 13694 7422 13746 7474
rect 13862 7478 13914 7530
rect 14590 7478 14642 7530
rect 16158 7534 16210 7586
rect 33686 7534 33738 7586
rect 34750 7534 34802 7586
rect 14254 7422 14306 7474
rect 15038 7422 15090 7474
rect 15914 7422 15966 7474
rect 16942 7422 16994 7474
rect 18324 7459 18376 7511
rect 18510 7422 18562 7474
rect 18622 7422 18674 7474
rect 19182 7422 19234 7474
rect 21086 7422 21138 7474
rect 21870 7422 21922 7474
rect 21982 7442 22034 7494
rect 24110 7422 24162 7474
rect 25230 7422 25282 7474
rect 25342 7422 25394 7474
rect 25488 7460 25540 7512
rect 30774 7478 30826 7530
rect 26910 7422 26962 7474
rect 30942 7422 30994 7474
rect 31334 7422 31386 7474
rect 32140 7460 32192 7512
rect 32286 7422 32338 7474
rect 32398 7422 32450 7474
rect 33182 7422 33234 7474
rect 33406 7422 33458 7474
rect 34190 7460 34242 7512
rect 34918 7478 34970 7530
rect 38110 7534 38162 7586
rect 43430 7534 43482 7586
rect 34526 7422 34578 7474
rect 35422 7422 35474 7474
rect 39342 7422 39394 7474
rect 40014 7478 40066 7530
rect 39678 7422 39730 7474
rect 40350 7422 40402 7474
rect 41022 7422 41074 7474
rect 41134 7422 41186 7474
rect 41302 7422 41354 7474
rect 42254 7422 42306 7474
rect 42590 7422 42642 7474
rect 42926 7422 42978 7474
rect 43150 7422 43202 7474
rect 43934 7455 43986 7507
rect 44214 7478 44266 7530
rect 44662 7478 44714 7530
rect 44986 7462 45038 7514
rect 48302 7422 48354 7474
rect 4062 7310 4114 7362
rect 10782 7310 10834 7362
rect 14030 7310 14082 7362
rect 17950 7310 18002 7362
rect 24726 7310 24778 7362
rect 25902 7310 25954 7362
rect 27694 7310 27746 7362
rect 29598 7310 29650 7362
rect 31166 7310 31218 7362
rect 31726 7310 31778 7362
rect 36206 7310 36258 7362
rect 38726 7310 38778 7362
rect 40014 7310 40066 7362
rect 41694 7310 41746 7362
rect 45054 7310 45106 7362
rect 45614 7310 45666 7362
rect 47518 7310 47570 7362
rect 12406 7198 12458 7250
rect 13190 7198 13242 7250
rect 16774 7198 16826 7250
rect 42702 7254 42754 7306
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 4174 6862 4226 6914
rect 13918 6806 13970 6858
rect 25454 6862 25506 6914
rect 6526 6750 6578 6802
rect 10894 6750 10946 6802
rect 15150 6750 15202 6802
rect 18510 6750 18562 6802
rect 44046 6806 44098 6858
rect 47070 6806 47122 6858
rect 20022 6750 20074 6802
rect 4510 6638 4562 6690
rect 5182 6638 5234 6690
rect 5798 6638 5850 6690
rect 6078 6638 6130 6690
rect 6414 6594 6466 6646
rect 7086 6638 7138 6690
rect 7870 6638 7922 6690
rect 10110 6638 10162 6690
rect 12798 6638 12850 6690
rect 13806 6638 13858 6690
rect 14478 6638 14530 6690
rect 13582 6582 13634 6634
rect 14814 6638 14866 6690
rect 15038 6599 15090 6651
rect 15486 6638 15538 6690
rect 16158 6638 16210 6690
rect 15766 6582 15818 6634
rect 16382 6610 16434 6662
rect 17054 6638 17106 6690
rect 17390 6638 17442 6690
rect 17838 6638 17890 6690
rect 18174 6638 18226 6690
rect 18734 6638 18786 6690
rect 19630 6638 19682 6690
rect 9774 6526 9826 6578
rect 18510 6582 18562 6634
rect 20470 6638 20522 6690
rect 22374 6694 22426 6746
rect 25902 6750 25954 6802
rect 23942 6694 23994 6746
rect 21534 6582 21586 6634
rect 21758 6610 21810 6662
rect 23326 6610 23378 6662
rect 23550 6638 23602 6690
rect 27190 6694 27242 6746
rect 27358 6750 27410 6802
rect 31054 6750 31106 6802
rect 35422 6750 35474 6802
rect 41582 6750 41634 6802
rect 43038 6750 43090 6802
rect 24446 6638 24498 6690
rect 24782 6638 24834 6690
rect 24894 6638 24946 6690
rect 15934 6526 15986 6578
rect 22206 6526 22258 6578
rect 25062 6582 25114 6634
rect 26014 6594 26066 6646
rect 26238 6638 26290 6690
rect 27582 6638 27634 6690
rect 27806 6610 27858 6662
rect 28590 6638 28642 6690
rect 29374 6638 29426 6690
rect 29766 6638 29818 6690
rect 30270 6638 30322 6690
rect 36206 6638 36258 6690
rect 37270 6694 37322 6746
rect 37662 6638 37714 6690
rect 37998 6600 38050 6652
rect 38334 6638 38386 6690
rect 38670 6638 38722 6690
rect 39118 6638 39170 6690
rect 39454 6611 39506 6663
rect 39790 6638 39842 6690
rect 40238 6638 40290 6690
rect 23774 6526 23826 6578
rect 4846 6414 4898 6466
rect 19294 6414 19346 6466
rect 22822 6414 22874 6466
rect 24278 6470 24330 6522
rect 26854 6414 26906 6466
rect 28422 6414 28474 6466
rect 29206 6470 29258 6522
rect 32958 6526 33010 6578
rect 33518 6526 33570 6578
rect 41694 6594 41746 6646
rect 42030 6638 42082 6690
rect 42366 6638 42418 6690
rect 42478 6638 42530 6690
rect 43710 6638 43762 6690
rect 44046 6638 44098 6690
rect 44830 6638 44882 6690
rect 45390 6638 45442 6690
rect 42646 6582 42698 6634
rect 45614 6638 45666 6690
rect 46286 6638 46338 6690
rect 46398 6638 46450 6690
rect 46678 6638 46730 6690
rect 47182 6638 47234 6690
rect 47518 6638 47570 6690
rect 48134 6638 48186 6690
rect 37438 6526 37490 6578
rect 45894 6526 45946 6578
rect 39230 6470 39282 6522
rect 40574 6414 40626 6466
rect 41190 6414 41242 6466
rect 44998 6414 45050 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 8150 6078 8202 6130
rect 9662 6078 9714 6130
rect 10390 6078 10442 6130
rect 12070 6078 12122 6130
rect 32342 6078 32394 6130
rect 7534 5966 7586 6018
rect 12350 5966 12402 6018
rect 18398 6022 18450 6074
rect 14926 5966 14978 6018
rect 4846 5854 4898 5906
rect 5630 5854 5682 5906
rect 8710 5883 8762 5935
rect 8990 5854 9042 5906
rect 9998 5854 10050 5906
rect 12509 5887 12561 5939
rect 12798 5910 12850 5962
rect 13134 5910 13186 5962
rect 13470 5910 13522 5962
rect 24558 5966 24610 6018
rect 14814 5854 14866 5906
rect 8542 5742 8594 5794
rect 14198 5742 14250 5794
rect 15094 5798 15146 5850
rect 15262 5854 15314 5906
rect 15710 5854 15762 5906
rect 16046 5854 16098 5906
rect 16494 5869 16546 5921
rect 18062 5910 18114 5962
rect 29150 5966 29202 6018
rect 16830 5854 16882 5906
rect 17614 5854 17666 5906
rect 18286 5854 18338 5906
rect 20862 5854 20914 5906
rect 21646 5854 21698 5906
rect 21870 5854 21922 5906
rect 22654 5854 22706 5906
rect 25230 5854 25282 5906
rect 25342 5854 25394 5906
rect 25528 5891 25580 5943
rect 26462 5854 26514 5906
rect 29934 5910 29986 5962
rect 30046 5910 30098 5962
rect 37270 5966 37322 6018
rect 43990 5966 44042 6018
rect 45950 5966 46002 6018
rect 46902 5966 46954 6018
rect 30774 5854 30826 5906
rect 31166 5910 31218 5962
rect 31502 5854 31554 5906
rect 32510 5854 32562 5906
rect 33070 5854 33122 5906
rect 33182 5854 33234 5906
rect 33340 5904 33392 5956
rect 34526 5854 34578 5906
rect 16382 5742 16434 5794
rect 18958 5742 19010 5794
rect 27246 5742 27298 5794
rect 30606 5742 30658 5794
rect 14534 5630 14586 5682
rect 15598 5686 15650 5738
rect 31726 5742 31778 5794
rect 31894 5798 31946 5850
rect 34750 5854 34802 5906
rect 34974 5854 35026 5906
rect 35086 5854 35138 5906
rect 36206 5854 36258 5906
rect 36990 5854 37042 5906
rect 37550 5854 37602 5906
rect 37774 5854 37826 5906
rect 38054 5854 38106 5906
rect 38334 5854 38386 5906
rect 38446 5854 38498 5906
rect 39006 5854 39058 5906
rect 39118 5854 39170 5906
rect 39304 5892 39356 5944
rect 40014 5854 40066 5906
rect 40910 5854 40962 5906
rect 41246 5869 41298 5921
rect 41806 5854 41858 5906
rect 42142 5854 42194 5906
rect 43374 5854 43426 5906
rect 43598 5854 43650 5906
rect 44718 5910 44770 5962
rect 44998 5910 45050 5962
rect 45502 5910 45554 5962
rect 43710 5854 43762 5906
rect 45812 5887 45864 5939
rect 46398 5854 46450 5906
rect 46622 5854 46674 5906
rect 47406 5854 47458 5906
rect 47630 5854 47682 5906
rect 33742 5742 33794 5794
rect 35870 5742 35922 5794
rect 36654 5742 36706 5794
rect 39678 5742 39730 5794
rect 41358 5742 41410 5794
rect 42534 5742 42586 5794
rect 40182 5686 40234 5738
rect 25902 5630 25954 5682
rect 34246 5630 34298 5682
rect 35366 5630 35418 5682
rect 43038 5630 43090 5682
rect 47294 5686 47346 5738
rect 48246 5742 48298 5794
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 21366 5294 21418 5346
rect 12574 5238 12626 5290
rect 18510 5182 18562 5234
rect 19630 5182 19682 5234
rect 20806 5182 20858 5234
rect 21758 5238 21810 5290
rect 23214 5238 23266 5290
rect 32678 5294 32730 5346
rect 34302 5294 34354 5346
rect 12574 5070 12626 5122
rect 12798 5070 12850 5122
rect 13650 5030 13702 5082
rect 15262 5070 15314 5122
rect 16046 5070 16098 5122
rect 17950 5070 18002 5122
rect 13974 5014 14026 5066
rect 14422 5014 14474 5066
rect 14590 5014 14642 5066
rect 26854 5126 26906 5178
rect 27022 5182 27074 5234
rect 29318 5182 29370 5234
rect 32174 5182 32226 5234
rect 33350 5182 33402 5234
rect 34750 5238 34802 5290
rect 35534 5238 35586 5290
rect 41246 5294 41298 5346
rect 45054 5294 45106 5346
rect 27694 5126 27746 5178
rect 37662 5182 37714 5234
rect 18902 5070 18954 5122
rect 19070 5070 19122 5122
rect 19182 5070 19234 5122
rect 20190 5070 20242 5122
rect 20302 5070 20354 5122
rect 21198 5070 21250 5122
rect 21870 5070 21922 5122
rect 22206 5070 22258 5122
rect 22878 5070 22930 5122
rect 23102 5070 23154 5122
rect 23438 5070 23490 5122
rect 24222 5070 24274 5122
rect 20022 5014 20074 5066
rect 27470 5042 27522 5094
rect 27918 5070 27970 5122
rect 28254 5070 28306 5122
rect 29486 5070 29538 5122
rect 30270 5070 30322 5122
rect 32510 5070 32562 5122
rect 33630 5070 33682 5122
rect 33742 5070 33794 5122
rect 33910 5070 33962 5122
rect 34862 5070 34914 5122
rect 35198 5070 35250 5122
rect 35646 5070 35698 5122
rect 35982 5070 36034 5122
rect 36486 5070 36538 5122
rect 37102 5032 37154 5084
rect 37438 5070 37490 5122
rect 37830 5070 37882 5122
rect 13470 4958 13522 5010
rect 38558 5032 38610 5084
rect 38894 5070 38946 5122
rect 39118 5070 39170 5122
rect 39286 5126 39338 5178
rect 40462 5182 40514 5234
rect 43374 5182 43426 5234
rect 43822 5182 43874 5234
rect 45614 5182 45666 5234
rect 47518 5182 47570 5234
rect 39790 5070 39842 5122
rect 40126 5070 40178 5122
rect 40798 5070 40850 5122
rect 40350 5014 40402 5066
rect 41489 5039 41541 5091
rect 42366 5070 42418 5122
rect 42702 5070 42754 5122
rect 42814 5070 42866 5122
rect 42980 5070 43032 5122
rect 43934 5055 43986 5107
rect 44270 5070 44322 5122
rect 44718 5070 44770 5122
rect 48302 5070 48354 5122
rect 26126 4958 26178 5010
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 11734 4510 11786 4562
rect 14590 4398 14642 4450
rect 17446 4454 17498 4506
rect 30102 4510 30154 4562
rect 33238 4510 33290 4562
rect 47910 4510 47962 4562
rect 23158 4398 23210 4450
rect 25230 4398 25282 4450
rect 15374 4342 15426 4394
rect 15598 4342 15650 4394
rect 16046 4342 16098 4394
rect 29486 4398 29538 4450
rect 11902 4286 11954 4338
rect 12686 4286 12738 4338
rect 16356 4326 16408 4378
rect 17278 4286 17330 4338
rect 17950 4286 18002 4338
rect 18286 4330 18338 4382
rect 19070 4286 19122 4338
rect 19294 4286 19346 4338
rect 19630 4286 19682 4338
rect 22318 4286 22370 4338
rect 22654 4286 22706 4338
rect 22878 4286 22930 4338
rect 23438 4286 23490 4338
rect 24558 4286 24610 4338
rect 24782 4286 24834 4338
rect 25410 4319 25462 4371
rect 25566 4322 25618 4374
rect 26014 4342 26066 4394
rect 26350 4342 26402 4394
rect 36318 4398 36370 4450
rect 39342 4398 39394 4450
rect 45390 4398 45442 4450
rect 26798 4286 26850 4338
rect 31580 4324 31632 4376
rect 31726 4286 31778 4338
rect 31838 4286 31890 4338
rect 32398 4286 32450 4338
rect 33630 4286 33682 4338
rect 41414 4342 41466 4394
rect 41694 4342 41746 4394
rect 42198 4342 42250 4394
rect 42478 4342 42530 4394
rect 36654 4286 36706 4338
rect 39902 4286 39954 4338
rect 40238 4286 40290 4338
rect 42702 4286 42754 4338
rect 45726 4286 45778 4338
rect 45950 4286 46002 4338
rect 46734 4286 46786 4338
rect 47070 4286 47122 4338
rect 16382 4174 16434 4226
rect 18398 4174 18450 4226
rect 20414 4174 20466 4226
rect 24278 4174 24330 4226
rect 27582 4174 27634 4226
rect 30774 4174 30826 4226
rect 19182 4118 19234 4170
rect 31166 4174 31218 4226
rect 34414 4174 34466 4226
rect 37438 4174 37490 4226
rect 23774 4062 23826 4114
rect 32230 4118 32282 4170
rect 41358 4174 41410 4226
rect 43486 4174 43538 4226
rect 47462 4174 47514 4226
rect 39790 4118 39842 4170
rect 46230 4062 46282 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 13806 3670 13858 3722
rect 15038 3726 15090 3778
rect 16382 3670 16434 3722
rect 22430 3726 22482 3778
rect 38614 3726 38666 3778
rect 42198 3726 42250 3778
rect 17222 3614 17274 3666
rect 18398 3614 18450 3666
rect 23270 3614 23322 3666
rect 24838 3614 24890 3666
rect 25902 3670 25954 3722
rect 13358 3502 13410 3554
rect 13694 3502 13746 3554
rect 14198 3502 14250 3554
rect 14478 3502 14530 3554
rect 14702 3502 14754 3554
rect 15374 3502 15426 3554
rect 16046 3502 16098 3554
rect 16270 3502 16322 3554
rect 17558 3502 17610 3554
rect 17838 3502 17890 3554
rect 17950 3502 18002 3554
rect 18734 3502 18786 3554
rect 19798 3502 19850 3554
rect 20078 3502 20130 3554
rect 20302 3502 20354 3554
rect 20930 3469 20982 3521
rect 12630 3390 12682 3442
rect 21086 3446 21138 3498
rect 21534 3465 21586 3517
rect 21982 3469 22034 3521
rect 22766 3502 22818 3554
rect 25174 3502 25226 3554
rect 25454 3502 25506 3554
rect 26966 3558 27018 3610
rect 27134 3614 27186 3666
rect 29598 3614 29650 3666
rect 31502 3614 31554 3666
rect 32342 3614 32394 3666
rect 32790 3614 32842 3666
rect 33238 3614 33290 3666
rect 34638 3614 34690 3666
rect 35478 3614 35530 3666
rect 36374 3614 36426 3666
rect 37774 3614 37826 3666
rect 39174 3614 39226 3666
rect 41694 3670 41746 3722
rect 39958 3614 40010 3666
rect 43710 3670 43762 3722
rect 44830 3670 44882 3722
rect 25678 3502 25730 3554
rect 26014 3502 26066 3554
rect 26238 3502 26290 3554
rect 27694 3464 27746 3516
rect 20750 3390 20802 3442
rect 28590 3502 28642 3554
rect 28814 3502 28866 3554
rect 24054 3390 24106 3442
rect 27806 3446 27858 3498
rect 33630 3469 33682 3521
rect 33966 3465 34018 3517
rect 34246 3446 34298 3498
rect 34612 3462 34664 3514
rect 36766 3469 36818 3521
rect 37102 3465 37154 3517
rect 37438 3469 37490 3521
rect 37748 3462 37800 3514
rect 38222 3502 38274 3554
rect 38334 3502 38386 3554
rect 40294 3502 40346 3554
rect 40574 3502 40626 3554
rect 40854 3558 40906 3610
rect 43094 3614 43146 3666
rect 45334 3614 45386 3666
rect 45782 3614 45834 3666
rect 46678 3614 46730 3666
rect 47574 3614 47626 3666
rect 48022 3614 48074 3666
rect 41022 3502 41074 3554
rect 41470 3502 41522 3554
rect 41694 3502 41746 3554
rect 42478 3502 42530 3554
rect 42590 3502 42642 3554
rect 43710 3502 43762 3554
rect 44046 3502 44098 3554
rect 44494 3502 44546 3554
rect 44718 3502 44770 3554
rect 19462 3278 19514 3330
rect 28422 3334 28474 3386
rect 40686 3390 40738 3442
rect 46230 3278 46282 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 3584 49200 3696 50000
rect 5152 49200 5264 50000
rect 6720 49200 6832 50000
rect 8288 49200 8400 50000
rect 9856 49200 9968 50000
rect 11424 49200 11536 50000
rect 12992 49200 13104 50000
rect 14560 49200 14672 50000
rect 16128 49200 16240 50000
rect 17696 49200 17808 50000
rect 19264 49200 19376 50000
rect 20832 49200 20944 50000
rect 22400 49200 22512 50000
rect 23968 49200 24080 50000
rect 25536 49200 25648 50000
rect 27104 49200 27216 50000
rect 28672 49200 28784 50000
rect 28924 49308 29876 49364
rect 3612 46340 3668 49200
rect 3612 46284 3948 46340
rect 3892 45722 3948 46284
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 5180 46228 5236 49200
rect 6748 46340 6804 49200
rect 6748 46284 7084 46340
rect 5180 46172 5628 46228
rect 2380 45668 2436 45678
rect 2212 44996 2268 45006
rect 1708 44994 2268 44996
rect 1708 44942 2214 44994
rect 2266 44942 2268 44994
rect 1708 44940 2268 44942
rect 1708 43708 1764 44940
rect 2212 44930 2268 44940
rect 2268 44324 2324 44334
rect 2380 44324 2436 45612
rect 3108 45668 3164 45678
rect 3108 45574 3164 45612
rect 3556 45668 3612 45678
rect 3892 45670 3894 45722
rect 3946 45670 3948 45722
rect 5572 45722 5628 46172
rect 3556 45666 3780 45668
rect 3556 45614 3558 45666
rect 3610 45614 3780 45666
rect 3892 45658 3948 45670
rect 4564 45668 4620 45678
rect 3556 45612 3780 45614
rect 3556 45602 3612 45612
rect 2660 45220 2716 45230
rect 2660 45126 2716 45164
rect 3108 44996 3164 45006
rect 2268 44322 2436 44324
rect 2268 44270 2270 44322
rect 2322 44270 2436 44322
rect 2268 44268 2436 44270
rect 2940 44994 3164 44996
rect 2940 44942 3110 44994
rect 3162 44942 3164 44994
rect 2940 44940 3164 44942
rect 2100 44100 2156 44110
rect 1596 43652 1764 43708
rect 2044 44098 2156 44100
rect 2044 44046 2102 44098
rect 2154 44046 2156 44098
rect 2044 44034 2156 44046
rect 1596 42754 1652 43652
rect 1876 43428 1932 43438
rect 1876 43334 1932 43372
rect 1596 42702 1598 42754
rect 1650 42702 1652 42754
rect 1484 42532 1540 42542
rect 28 25284 84 25294
rect 28 8148 84 25228
rect 1484 21476 1540 42476
rect 1596 42196 1652 42702
rect 1932 42532 1988 42542
rect 1932 42438 1988 42476
rect 1596 42130 1652 42140
rect 2044 42084 2100 44034
rect 2268 43708 2324 44268
rect 2940 43708 2996 44940
rect 3108 44930 3164 44940
rect 3556 44994 3612 45006
rect 3556 44942 3558 44994
rect 3610 44942 3612 44994
rect 3556 44884 3612 44942
rect 3724 44996 3780 45612
rect 4564 45444 4620 45612
rect 4564 45378 4620 45388
rect 5012 45666 5068 45678
rect 5012 45614 5014 45666
rect 5066 45614 5068 45666
rect 5572 45670 5574 45722
rect 5626 45670 5628 45722
rect 6860 45892 6916 45902
rect 5572 45658 5628 45670
rect 6244 45668 6300 45678
rect 6692 45668 6748 45678
rect 6244 45666 6356 45668
rect 4452 45332 4508 45342
rect 3724 44930 3780 44940
rect 4004 44996 4060 45006
rect 4452 44996 4508 45276
rect 5012 45332 5068 45614
rect 6244 45614 6246 45666
rect 6298 45614 6356 45666
rect 6244 45602 6356 45614
rect 6300 45556 6356 45602
rect 6692 45574 6748 45612
rect 6300 45490 6356 45500
rect 5012 45266 5068 45276
rect 6188 45444 6244 45454
rect 5852 45106 5908 45118
rect 5852 45054 5854 45106
rect 5906 45054 5908 45106
rect 4004 44902 4060 44940
rect 4284 44994 4508 44996
rect 4284 44942 4454 44994
rect 4506 44942 4508 44994
rect 4284 44940 4508 44942
rect 3556 44818 3612 44828
rect 1708 42028 2100 42084
rect 2156 43652 2324 43708
rect 2604 43652 2996 43708
rect 3052 44322 3108 44334
rect 3052 44270 3054 44322
rect 3106 44270 3108 44322
rect 3052 43652 3108 44270
rect 4284 43988 4340 44940
rect 4452 44930 4508 44940
rect 4900 44996 4956 45006
rect 4900 44902 4956 44940
rect 5348 44994 5404 45006
rect 5348 44942 5350 44994
rect 5402 44942 5404 44994
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 5348 44436 5404 44942
rect 5684 44884 5740 44894
rect 5180 44380 5404 44436
rect 5516 44882 5740 44884
rect 5516 44830 5686 44882
rect 5738 44830 5740 44882
rect 5516 44828 5740 44830
rect 4956 44210 5012 44222
rect 4956 44158 4958 44210
rect 5010 44158 5012 44210
rect 4284 43922 4340 43932
rect 4732 44100 4788 44110
rect 1596 41972 1652 41982
rect 1708 41972 1764 42028
rect 1596 41970 1764 41972
rect 1596 41918 1598 41970
rect 1650 41918 1764 41970
rect 1596 41916 1764 41918
rect 1596 41906 1652 41916
rect 1820 40292 1876 42028
rect 1988 41300 2044 41310
rect 1988 41206 2044 41244
rect 1988 40516 2044 40526
rect 1988 40422 2044 40460
rect 1596 40236 1820 40292
rect 1596 39618 1652 40236
rect 1820 40226 1876 40236
rect 1596 39566 1598 39618
rect 1650 39566 1652 39618
rect 1596 39060 1652 39566
rect 1596 37266 1652 39004
rect 1596 37214 1598 37266
rect 1650 37214 1652 37266
rect 1596 35698 1652 37214
rect 1596 35646 1598 35698
rect 1650 35646 1652 35698
rect 1596 35634 1652 35646
rect 1596 33348 1652 33358
rect 1596 32788 1652 33292
rect 2156 33348 2212 43652
rect 2324 43428 2380 43438
rect 2604 43428 2660 43652
rect 3052 43586 3108 43596
rect 4060 43652 4116 43662
rect 4060 43558 4116 43596
rect 4396 43652 4452 43662
rect 4396 43538 4452 43596
rect 4396 43486 4398 43538
rect 4450 43486 4452 43538
rect 4396 43474 4452 43486
rect 4732 43538 4788 44044
rect 4956 43764 5012 44158
rect 4956 43698 5012 43708
rect 4732 43486 4734 43538
rect 4786 43486 4788 43538
rect 4732 43474 4788 43486
rect 4956 43553 5012 43565
rect 4956 43501 4958 43553
rect 5010 43501 5012 43553
rect 2324 43426 2660 43428
rect 2324 43374 2326 43426
rect 2378 43374 2660 43426
rect 2324 43372 2660 43374
rect 2324 43362 2380 43372
rect 2604 42980 2660 43372
rect 2604 42914 2660 42924
rect 2772 43426 2828 43438
rect 3220 43428 3276 43438
rect 2772 43374 2774 43426
rect 2826 43374 2828 43426
rect 2772 42980 2828 43374
rect 2772 42914 2828 42924
rect 2940 43426 3276 43428
rect 2940 43374 3222 43426
rect 3274 43374 3276 43426
rect 2940 43372 3276 43374
rect 2940 42756 2996 43372
rect 3220 43362 3276 43372
rect 3668 43426 3724 43438
rect 3668 43374 3670 43426
rect 3722 43374 3724 43426
rect 3668 43316 3724 43374
rect 3668 43250 3724 43260
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4956 43092 5012 43501
rect 5068 43540 5124 43550
rect 5068 43426 5124 43484
rect 5068 43374 5070 43426
rect 5122 43374 5124 43426
rect 5068 43362 5124 43374
rect 5180 43316 5236 44380
rect 5404 43540 5460 43550
rect 5516 43540 5572 44828
rect 5684 44818 5740 44828
rect 5852 43876 5908 45054
rect 6188 45106 6244 45388
rect 6188 45054 6190 45106
rect 6242 45054 6244 45106
rect 6188 45042 6244 45054
rect 6860 44558 6916 45836
rect 7028 45722 7084 46284
rect 7308 45892 7364 45902
rect 8316 45892 8372 49200
rect 9884 45892 9940 49200
rect 11452 46340 11508 49200
rect 13020 46788 13076 49200
rect 13020 46732 13412 46788
rect 11396 46284 11508 46340
rect 8316 45836 8652 45892
rect 9884 45836 10220 45892
rect 7308 45798 7364 45836
rect 7028 45670 7030 45722
rect 7082 45670 7084 45722
rect 8596 45722 8652 45836
rect 7028 45658 7084 45670
rect 7644 45668 7700 45678
rect 7196 45666 7700 45668
rect 7196 45614 7646 45666
rect 7698 45614 7700 45666
rect 7196 45612 7700 45614
rect 6972 45108 7028 45118
rect 7196 45108 7252 45612
rect 7644 45602 7700 45612
rect 8260 45666 8316 45678
rect 8260 45614 8262 45666
rect 8314 45614 8316 45666
rect 8596 45670 8598 45722
rect 8650 45670 8652 45722
rect 10164 45722 10220 45836
rect 8596 45658 8652 45670
rect 9212 45668 9268 45678
rect 8260 45556 8316 45614
rect 8260 45490 8316 45500
rect 6972 45106 7252 45108
rect 6972 45054 6974 45106
rect 7026 45054 7252 45106
rect 6972 45052 7252 45054
rect 9212 45108 9268 45612
rect 9828 45668 9884 45678
rect 10164 45670 10166 45722
rect 10218 45670 10220 45722
rect 10164 45658 10220 45670
rect 10556 45890 10612 45902
rect 10556 45838 10558 45890
rect 10610 45838 10612 45890
rect 9828 45574 9884 45612
rect 9772 45444 9828 45454
rect 9548 45108 9604 45118
rect 6972 45042 7028 45052
rect 5964 44492 6244 44548
rect 5964 44322 6020 44492
rect 5964 44270 5966 44322
rect 6018 44270 6020 44322
rect 5964 44100 6020 44270
rect 5964 44034 6020 44044
rect 6076 44322 6132 44334
rect 6076 44270 6078 44322
rect 6130 44270 6132 44322
rect 5852 43810 5908 43820
rect 5404 43538 5572 43540
rect 5404 43486 5406 43538
rect 5458 43486 5572 43538
rect 5404 43484 5572 43486
rect 5404 43474 5460 43484
rect 5180 43250 5236 43260
rect 4956 43026 5012 43036
rect 5684 43092 5740 43102
rect 6076 43092 6132 44270
rect 6188 43988 6244 44492
rect 6804 44546 6916 44558
rect 8876 44994 8932 45006
rect 8876 44942 8878 44994
rect 8930 44942 8932 44994
rect 6804 44494 6806 44546
rect 6858 44494 6916 44546
rect 6804 44492 6916 44494
rect 7980 44492 8316 44548
rect 6804 44482 6860 44492
rect 7084 44322 7140 44334
rect 7084 44270 7086 44322
rect 7138 44270 7140 44322
rect 6356 44212 6412 44222
rect 6356 44210 6692 44212
rect 6356 44158 6358 44210
rect 6410 44158 6692 44210
rect 6356 44156 6692 44158
rect 6356 44146 6412 44156
rect 6188 43932 6468 43988
rect 6412 43652 6468 43932
rect 6524 43652 6580 43662
rect 6412 43650 6580 43652
rect 6412 43598 6526 43650
rect 6578 43598 6580 43650
rect 6412 43596 6580 43598
rect 6524 43586 6580 43596
rect 6280 43540 6336 43550
rect 6280 43538 6356 43540
rect 6280 43486 6282 43538
rect 6334 43486 6356 43538
rect 6280 43474 6356 43486
rect 6300 43428 6356 43474
rect 6636 43428 6692 44156
rect 7084 44100 7140 44270
rect 7308 44324 7364 44334
rect 7588 44324 7644 44334
rect 7308 44322 7644 44324
rect 7308 44270 7310 44322
rect 7362 44270 7590 44322
rect 7642 44270 7644 44322
rect 7308 44268 7644 44270
rect 7308 44258 7364 44268
rect 7588 44258 7644 44268
rect 7868 44324 7924 44334
rect 7980 44324 8036 44492
rect 8260 44378 8316 44492
rect 8876 44436 8932 44942
rect 9100 44436 9156 44446
rect 8876 44380 9100 44436
rect 7868 44322 8036 44324
rect 7868 44270 7870 44322
rect 7922 44270 8036 44322
rect 7868 44268 8036 44270
rect 8092 44322 8148 44334
rect 8092 44270 8094 44322
rect 8146 44270 8148 44322
rect 8260 44326 8262 44378
rect 8314 44326 8316 44378
rect 9100 44378 9156 44380
rect 8260 44314 8316 44326
rect 8428 44324 8484 44334
rect 7084 44034 7140 44044
rect 7084 43706 7140 43718
rect 7084 43654 7086 43706
rect 7138 43654 7140 43706
rect 7084 43652 7140 43654
rect 7084 43586 7140 43596
rect 7420 43577 7476 43589
rect 7196 43538 7252 43550
rect 7196 43486 7198 43538
rect 7250 43486 7252 43538
rect 7196 43428 7252 43486
rect 7420 43540 7422 43577
rect 7474 43540 7476 43577
rect 7420 43474 7476 43484
rect 7756 43540 7812 43550
rect 7756 43446 7812 43484
rect 6300 43372 6580 43428
rect 5740 43036 6132 43092
rect 6412 43092 6468 43102
rect 3724 42924 4452 42980
rect 3724 42756 3780 42924
rect 2492 42700 2996 42756
rect 3612 42739 3780 42756
rect 2380 41858 2436 41870
rect 2380 41806 2382 41858
rect 2434 41806 2436 41858
rect 2380 41410 2436 41806
rect 2380 41358 2382 41410
rect 2434 41358 2436 41410
rect 2380 41346 2436 41358
rect 2492 40740 2548 42700
rect 3612 42687 3614 42739
rect 3666 42700 3780 42739
rect 3666 42687 3668 42700
rect 3612 42675 3668 42687
rect 3612 42586 3668 42598
rect 2772 42532 2828 42542
rect 2604 42530 2828 42532
rect 2604 42478 2774 42530
rect 2826 42478 2828 42530
rect 2604 42476 2828 42478
rect 2604 41860 2660 42476
rect 2772 42466 2828 42476
rect 3220 42530 3276 42542
rect 3220 42478 3222 42530
rect 3274 42478 3276 42530
rect 3220 42196 3276 42478
rect 3220 42130 3276 42140
rect 3612 42534 3614 42586
rect 3666 42534 3668 42586
rect 2604 41300 2660 41804
rect 2604 41234 2660 41244
rect 2716 41188 2772 41198
rect 2716 41094 2772 41132
rect 3276 41186 3332 41198
rect 3276 41134 3278 41186
rect 3330 41134 3332 41186
rect 2884 40740 2940 40750
rect 2492 40684 2884 40740
rect 2884 40626 2940 40684
rect 2884 40574 2886 40626
rect 2938 40574 2940 40626
rect 2884 40562 2940 40574
rect 3276 40628 3332 41134
rect 3388 41188 3444 41198
rect 3388 41018 3444 41132
rect 3612 41159 3668 42534
rect 3612 41107 3614 41159
rect 3666 41107 3668 41159
rect 3612 41095 3668 41107
rect 3388 40966 3390 41018
rect 3442 40966 3444 41018
rect 3388 40954 3444 40966
rect 3276 40572 3556 40628
rect 3388 40458 3444 40470
rect 2436 40402 2492 40414
rect 2436 40350 2438 40402
rect 2490 40350 2492 40402
rect 2436 40292 2492 40350
rect 2436 40226 2492 40236
rect 2604 40404 2660 40414
rect 2604 40068 2660 40348
rect 3388 40406 3390 40458
rect 3442 40406 3444 40458
rect 3388 40292 3444 40406
rect 3388 40226 3444 40236
rect 2492 40012 2660 40068
rect 3220 40178 3276 40190
rect 3220 40126 3222 40178
rect 3274 40126 3276 40178
rect 2380 39618 2436 39630
rect 2380 39566 2382 39618
rect 2434 39566 2436 39618
rect 2268 39060 2324 39070
rect 2380 39060 2436 39566
rect 2268 39058 2436 39060
rect 2268 39006 2270 39058
rect 2322 39006 2436 39058
rect 2268 39004 2436 39006
rect 2268 38994 2324 39004
rect 2492 38836 2548 40012
rect 3220 39956 3276 40126
rect 2604 39900 3276 39956
rect 2604 39396 2660 39900
rect 2604 39340 2996 39396
rect 2604 38836 2660 38846
rect 2492 38834 2660 38836
rect 2492 38782 2606 38834
rect 2658 38782 2660 38834
rect 2492 38780 2660 38782
rect 2604 38770 2660 38780
rect 2940 38834 2996 39340
rect 3500 39172 3556 40572
rect 3724 40178 3780 42700
rect 3948 42756 4004 42766
rect 4284 42756 4340 42766
rect 3948 42754 4340 42756
rect 3948 42702 3950 42754
rect 4002 42702 4286 42754
rect 4338 42702 4340 42754
rect 3948 42700 4340 42702
rect 3948 42690 4004 42700
rect 3948 42532 4004 42542
rect 3948 41186 4004 42476
rect 4284 42420 4340 42700
rect 4396 42754 4452 42924
rect 5684 42978 5740 43036
rect 5684 42926 5686 42978
rect 5738 42926 5740 42978
rect 5684 42914 5740 42926
rect 4396 42702 4398 42754
rect 4450 42702 4452 42754
rect 4396 42690 4452 42702
rect 5292 42868 5348 42878
rect 4676 42642 4732 42654
rect 4676 42590 4678 42642
rect 4730 42590 4732 42642
rect 4676 42532 4732 42590
rect 4676 42466 4732 42476
rect 4284 42364 4452 42420
rect 4396 42084 4452 42364
rect 4844 42084 4900 42094
rect 4396 42082 4900 42084
rect 4396 42030 4846 42082
rect 4898 42030 4900 42082
rect 4396 42028 4900 42030
rect 4844 42018 4900 42028
rect 4284 41972 4340 41982
rect 4284 41878 4340 41916
rect 5087 41970 5143 41982
rect 5087 41918 5089 41970
rect 5141 41918 5143 41970
rect 5087 41860 5143 41918
rect 5087 41794 5143 41804
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 5292 41524 5348 42812
rect 5964 42754 6020 42766
rect 5964 42702 5966 42754
rect 6018 42702 6020 42754
rect 5964 42532 6020 42702
rect 5964 42466 6020 42476
rect 6188 42754 6244 42766
rect 6188 42702 6190 42754
rect 6242 42702 6244 42754
rect 5964 41972 6020 41982
rect 5964 41878 6020 41916
rect 6188 41860 6244 42702
rect 6412 42754 6468 43036
rect 6412 42702 6414 42754
rect 6466 42702 6468 42754
rect 6412 42690 6468 42702
rect 6524 42868 6580 43372
rect 6524 42754 6580 42812
rect 6524 42702 6526 42754
rect 6578 42702 6580 42754
rect 6524 42690 6580 42702
rect 6636 43372 7252 43428
rect 6636 42766 6692 43372
rect 7084 43204 7140 43214
rect 7084 42978 7140 43148
rect 7868 43204 7924 44268
rect 7980 44100 8036 44110
rect 8092 44100 8148 44270
rect 9100 44326 9102 44378
rect 9154 44326 9156 44378
rect 9100 44314 9156 44326
rect 8428 44230 8484 44268
rect 8988 44266 9044 44278
rect 8988 44214 8990 44266
rect 9042 44214 9044 44266
rect 8092 44044 8484 44100
rect 7980 43652 8036 44044
rect 8428 43764 8484 44044
rect 8540 43764 8596 43774
rect 8428 43708 8540 43764
rect 8316 43652 8372 43662
rect 7980 43650 8372 43652
rect 7980 43598 8318 43650
rect 8370 43598 8372 43650
rect 7980 43596 8372 43598
rect 8316 43586 8372 43596
rect 8540 43538 8596 43708
rect 7868 43138 7924 43148
rect 8148 43482 8204 43494
rect 8148 43430 8150 43482
rect 8202 43430 8204 43482
rect 8540 43486 8542 43538
rect 8594 43486 8596 43538
rect 8540 43474 8596 43486
rect 8764 43566 8820 43578
rect 8764 43514 8766 43566
rect 8818 43514 8820 43566
rect 8148 42980 8204 43430
rect 8764 43204 8820 43514
rect 8764 43138 8820 43148
rect 8876 43540 8932 43550
rect 7084 42926 7086 42978
rect 7138 42926 7140 42978
rect 7084 42914 7140 42926
rect 7756 42924 8204 42980
rect 6636 42754 6746 42766
rect 7644 42756 7700 42766
rect 6636 42702 6692 42754
rect 6744 42702 6746 42754
rect 6636 42700 6746 42702
rect 6690 42690 6746 42700
rect 7420 42754 7700 42756
rect 7420 42702 7646 42754
rect 7698 42702 7700 42754
rect 7420 42700 7700 42702
rect 6300 41972 6356 41982
rect 6300 41878 6356 41916
rect 6860 41970 6916 41982
rect 6860 41918 6862 41970
rect 6914 41918 6916 41970
rect 6188 41794 6244 41804
rect 6860 41748 6916 41918
rect 7084 41860 7140 41870
rect 7084 41802 7140 41804
rect 7084 41750 7086 41802
rect 7138 41750 7140 41802
rect 7084 41738 7140 41750
rect 6860 41682 6916 41692
rect 6188 41636 6244 41646
rect 5292 41468 5684 41524
rect 3948 41134 3950 41186
rect 4002 41134 4004 41186
rect 3948 41122 4004 41134
rect 4172 41356 4676 41412
rect 3724 40126 3726 40178
rect 3778 40126 3780 40178
rect 3724 40114 3780 40126
rect 3836 40628 3892 40638
rect 3836 39508 3892 40572
rect 4172 40432 4228 41356
rect 4508 41186 4564 41198
rect 4508 41134 4510 41186
rect 4562 41134 4564 41186
rect 4172 40380 4174 40432
rect 4226 40380 4228 40432
rect 4396 40516 4452 40526
rect 4396 40458 4452 40460
rect 4396 40406 4398 40458
rect 4450 40406 4452 40458
rect 4396 40394 4452 40406
rect 4004 40346 4060 40358
rect 4004 40294 4006 40346
rect 4058 40294 4060 40346
rect 4004 40292 4060 40294
rect 4004 39844 4060 40236
rect 4172 40292 4228 40380
rect 4172 40226 4228 40236
rect 4508 40180 4564 41134
rect 4620 41186 4676 41356
rect 4620 41134 4622 41186
rect 4674 41134 4676 41186
rect 4620 41122 4676 41134
rect 5516 41186 5572 41198
rect 5516 41134 5518 41186
rect 5570 41134 5572 41186
rect 4900 41076 4956 41086
rect 4844 41074 4956 41076
rect 4844 41022 4902 41074
rect 4954 41022 4956 41074
rect 4844 41010 4956 41022
rect 4844 40402 4900 41010
rect 5180 40516 5236 40526
rect 4844 40350 4846 40402
rect 4898 40350 4900 40402
rect 4844 40338 4900 40350
rect 5068 40402 5124 40414
rect 5068 40350 5070 40402
rect 5122 40350 5124 40402
rect 4508 40124 4900 40180
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4004 39788 4340 39844
rect 4284 39730 4340 39788
rect 4284 39678 4286 39730
rect 4338 39678 4340 39730
rect 4284 39666 4340 39678
rect 3500 39106 3556 39116
rect 3816 39452 3892 39508
rect 4060 39620 4116 39630
rect 2940 38782 2942 38834
rect 2994 38782 2996 38834
rect 2940 38770 2996 38782
rect 3816 38890 3872 39452
rect 3816 38838 3818 38890
rect 3870 38838 3872 38890
rect 3816 38668 3872 38838
rect 3948 39172 4004 39182
rect 3816 38612 3892 38668
rect 3444 38276 3500 38286
rect 2996 38164 3052 38174
rect 2996 38070 3052 38108
rect 3444 38162 3500 38220
rect 3836 38276 3892 38612
rect 3836 38210 3892 38220
rect 3444 38110 3446 38162
rect 3498 38110 3500 38162
rect 3444 38098 3500 38110
rect 3948 38164 4004 39116
rect 4060 38946 4116 39564
rect 4844 39620 4900 40124
rect 5068 39732 5124 40350
rect 5068 39666 5124 39676
rect 4844 39554 4900 39564
rect 5180 39518 5236 40460
rect 5348 40404 5404 40414
rect 5348 40310 5404 40348
rect 5124 39506 5236 39518
rect 5124 39454 5126 39506
rect 5178 39454 5236 39506
rect 5124 39452 5236 39454
rect 5124 39442 5180 39452
rect 4060 38894 4062 38946
rect 4114 38894 4116 38946
rect 4060 38882 4116 38894
rect 4676 39060 4732 39070
rect 4676 38724 4732 39004
rect 5180 38948 5236 38958
rect 5180 38854 5236 38892
rect 4676 38658 4732 38668
rect 5516 38724 5572 41134
rect 5516 38658 5572 38668
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 2604 38052 2660 38062
rect 2604 37958 2660 37996
rect 3780 38052 3836 38062
rect 3780 37958 3836 37996
rect 2268 37826 2324 37838
rect 2268 37774 2270 37826
rect 2322 37774 2324 37826
rect 2268 37268 2324 37774
rect 3948 37828 4004 38108
rect 4060 38052 4116 38062
rect 4284 38052 4340 38062
rect 4564 38052 4620 38062
rect 4844 38052 4900 38062
rect 4060 38050 4228 38052
rect 4060 37998 4062 38050
rect 4114 37998 4228 38050
rect 4060 37996 4228 37998
rect 4060 37986 4116 37996
rect 3948 37772 4116 37828
rect 2380 37268 2436 37278
rect 2268 37266 2436 37268
rect 2268 37214 2382 37266
rect 2434 37214 2436 37266
rect 2268 37212 2436 37214
rect 2380 37202 2436 37212
rect 2604 36484 2660 36494
rect 2604 36390 2660 36428
rect 3500 36482 3556 36494
rect 3500 36430 3502 36482
rect 3554 36430 3556 36482
rect 2268 36258 2324 36270
rect 2268 36206 2270 36258
rect 2322 36206 2324 36258
rect 2268 35700 2324 36206
rect 2380 35700 2436 35710
rect 2268 35698 2436 35700
rect 2268 35646 2382 35698
rect 2434 35646 2436 35698
rect 2268 35644 2436 35646
rect 2380 35634 2436 35644
rect 2660 35364 2716 35374
rect 2660 35138 2716 35308
rect 3500 35364 3556 36430
rect 3612 36482 3668 36494
rect 3612 36430 3614 36482
rect 3666 36430 3668 36482
rect 3612 35812 3668 36430
rect 3892 36484 3948 36494
rect 3892 36390 3948 36428
rect 3612 35746 3668 35756
rect 3500 35298 3556 35308
rect 2660 35086 2662 35138
rect 2714 35086 2716 35138
rect 2660 35074 2716 35086
rect 2940 34914 2996 34926
rect 2940 34862 2942 34914
rect 2994 34862 2996 34914
rect 2604 34468 2660 34478
rect 2156 33282 2212 33292
rect 2380 33346 2436 33358
rect 2380 33294 2382 33346
rect 2434 33294 2436 33346
rect 1596 30994 1652 32732
rect 2268 32788 2324 32798
rect 2380 32788 2436 33294
rect 2268 32786 2436 32788
rect 2268 32734 2270 32786
rect 2322 32734 2436 32786
rect 2268 32732 2436 32734
rect 2268 32722 2324 32732
rect 2604 32562 2660 34412
rect 2940 34244 2996 34862
rect 3164 34916 3220 34926
rect 3164 34822 3220 34860
rect 3388 34914 3444 34926
rect 3388 34862 3390 34914
rect 3442 34862 3444 34914
rect 3388 34580 3444 34862
rect 4060 34916 4116 37772
rect 4172 36708 4228 37996
rect 4284 38050 4620 38052
rect 4284 37998 4286 38050
rect 4338 37998 4566 38050
rect 4618 37998 4620 38050
rect 4284 37996 4620 37998
rect 4284 37986 4340 37996
rect 4564 37986 4620 37996
rect 4732 38050 4900 38052
rect 4732 37998 4846 38050
rect 4898 37998 4900 38050
rect 4732 37996 4900 37998
rect 4284 37268 4340 37278
rect 4284 37174 4340 37212
rect 4732 37156 4788 37996
rect 4844 37986 4900 37996
rect 4956 38050 5012 38062
rect 4956 37998 4958 38050
rect 5010 37998 5012 38050
rect 4732 37090 4788 37100
rect 4844 37380 4900 37390
rect 4956 37380 5012 37998
rect 5628 37604 5684 41468
rect 6188 40964 6244 41580
rect 6300 41188 6356 41198
rect 6300 41186 6580 41188
rect 6300 41134 6302 41186
rect 6354 41134 6580 41186
rect 6300 41132 6580 41134
rect 6300 41122 6356 41132
rect 6188 40908 6468 40964
rect 6412 40740 6468 40908
rect 6244 40516 6300 40526
rect 6244 40422 6300 40460
rect 5852 40292 5908 40302
rect 5852 39844 5908 40236
rect 5852 39590 5908 39788
rect 6300 39732 6356 39742
rect 6300 39638 6356 39676
rect 5852 39538 5854 39590
rect 5906 39538 5908 39590
rect 5852 39526 5908 39538
rect 6076 39620 6132 39630
rect 6076 39526 6132 39564
rect 6412 39574 6468 40684
rect 6524 40628 6580 41132
rect 6972 40964 7028 40974
rect 7420 40964 7476 42700
rect 7644 42690 7700 42700
rect 7756 42532 7812 42924
rect 7532 42476 7812 42532
rect 7868 42754 7924 42766
rect 7868 42702 7870 42754
rect 7922 42702 7924 42754
rect 7532 41636 7588 42476
rect 7868 42082 7924 42702
rect 8148 42644 8204 42654
rect 7868 42030 7870 42082
rect 7922 42030 7924 42082
rect 7868 42018 7924 42030
rect 7980 42642 8204 42644
rect 7980 42590 8150 42642
rect 8202 42590 8204 42642
rect 7980 42588 8204 42590
rect 7700 41972 7756 41982
rect 7532 41570 7588 41580
rect 7644 41916 7700 41972
rect 7644 41878 7756 41916
rect 6636 40628 6692 40638
rect 6524 40626 6692 40628
rect 6524 40574 6638 40626
rect 6690 40574 6692 40626
rect 6524 40572 6692 40574
rect 6636 40562 6692 40572
rect 6972 40402 7028 40908
rect 7252 40908 7476 40964
rect 7252 40514 7308 40908
rect 7252 40462 7254 40514
rect 7306 40462 7308 40514
rect 7252 40450 7308 40462
rect 6972 40350 6974 40402
rect 7026 40350 7028 40402
rect 6972 40338 7028 40350
rect 7532 40404 7588 40414
rect 7532 40310 7588 40348
rect 7644 40180 7700 41878
rect 7980 41412 8036 42588
rect 8148 42578 8204 42588
rect 8876 42542 8932 43484
rect 8988 43092 9044 44214
rect 8988 43026 9044 43036
rect 9100 42756 9156 42766
rect 9212 42756 9268 45052
rect 9436 45106 9604 45108
rect 9436 45054 9550 45106
rect 9602 45054 9604 45106
rect 9436 45052 9604 45054
rect 9436 44436 9492 45052
rect 9548 45042 9604 45052
rect 9436 43538 9492 44380
rect 9660 44324 9716 44334
rect 9660 44230 9716 44268
rect 9772 44154 9828 45388
rect 10556 45444 10612 45838
rect 11396 45722 11452 46284
rect 12684 45892 12740 45902
rect 12684 45890 12852 45892
rect 12684 45838 12686 45890
rect 12738 45838 12852 45890
rect 12684 45836 12852 45838
rect 12684 45826 12740 45836
rect 10892 45668 10948 45678
rect 11396 45670 11398 45722
rect 11450 45670 11452 45722
rect 10892 45666 11172 45668
rect 10892 45614 10894 45666
rect 10946 45614 11172 45666
rect 11396 45658 11452 45670
rect 11844 45780 11900 45790
rect 11844 45722 11900 45724
rect 11844 45670 11846 45722
rect 11898 45670 11900 45722
rect 11844 45658 11900 45670
rect 12348 45666 12404 45678
rect 10892 45612 11172 45614
rect 10892 45602 10948 45612
rect 10556 45378 10612 45388
rect 9772 44102 9774 44154
rect 9826 44102 9828 44154
rect 9772 44090 9828 44102
rect 9884 45121 9940 45133
rect 9884 45069 9886 45121
rect 9938 45069 9940 45121
rect 9884 43988 9940 45069
rect 10332 45108 10388 45118
rect 10332 45014 10388 45052
rect 11116 45106 11172 45612
rect 12348 45614 12350 45666
rect 12402 45614 12404 45666
rect 11116 45054 11118 45106
rect 11170 45054 11172 45106
rect 11116 45042 11172 45054
rect 12236 45556 12292 45566
rect 9996 44994 10052 45006
rect 9996 44942 9998 44994
rect 10050 44942 10052 44994
rect 9996 44324 10052 44942
rect 10668 44434 10724 44446
rect 10668 44382 10670 44434
rect 10722 44382 10724 44434
rect 10220 44324 10276 44334
rect 9996 44243 9998 44268
rect 10050 44243 10052 44268
rect 9996 44230 10052 44243
rect 10108 44322 10276 44324
rect 10108 44270 10222 44322
rect 10274 44270 10276 44322
rect 10108 44268 10276 44270
rect 9436 43486 9438 43538
rect 9490 43486 9492 43538
rect 9436 43474 9492 43486
rect 9660 43932 9940 43988
rect 9996 43988 10052 43998
rect 9660 43538 9716 43932
rect 9996 43764 10052 43932
rect 9660 43486 9662 43538
rect 9714 43486 9716 43538
rect 9660 43092 9716 43486
rect 9884 43708 10052 43764
rect 9884 43438 9940 43708
rect 9884 43426 9996 43438
rect 9884 43374 9942 43426
rect 9994 43374 9996 43426
rect 9884 43372 9996 43374
rect 9940 43362 9996 43372
rect 9660 43026 9716 43036
rect 9996 43204 10052 43214
rect 9884 42756 9940 42766
rect 9100 42754 9268 42756
rect 9100 42702 9102 42754
rect 9154 42702 9268 42754
rect 9100 42700 9268 42702
rect 9100 42690 9156 42700
rect 8876 42530 8988 42542
rect 8876 42478 8934 42530
rect 8986 42478 8988 42530
rect 8876 42476 8988 42478
rect 8932 42084 8988 42476
rect 8932 42018 8988 42028
rect 8316 41998 8372 42010
rect 7868 41356 8036 41412
rect 8092 41970 8148 41982
rect 8092 41918 8094 41970
rect 8146 41918 8148 41970
rect 7868 41188 7924 41356
rect 7868 41122 7924 41132
rect 8092 41188 8148 41918
rect 8092 41122 8148 41132
rect 8204 41972 8260 41982
rect 7756 41076 7812 41086
rect 7756 40402 7812 41020
rect 8204 41074 8260 41916
rect 8204 41022 8206 41074
rect 8258 41022 8260 41074
rect 8204 40964 8260 41022
rect 7756 40350 7758 40402
rect 7810 40350 7812 40402
rect 7924 40908 8260 40964
rect 8316 41946 8318 41998
rect 8370 41946 8372 41998
rect 7924 40458 7980 40908
rect 7924 40406 7926 40458
rect 7978 40406 7980 40458
rect 7924 40394 7980 40406
rect 8092 40516 8148 40526
rect 8092 40458 8148 40460
rect 8092 40406 8094 40458
rect 8146 40406 8148 40458
rect 8092 40394 8148 40406
rect 8316 40458 8372 41946
rect 8764 41972 8820 41982
rect 8764 41878 8820 41916
rect 8932 41746 8988 41758
rect 8932 41694 8934 41746
rect 8986 41694 8988 41746
rect 8932 41412 8988 41694
rect 8932 41346 8988 41356
rect 9007 41130 9063 41142
rect 8764 41076 8820 41086
rect 8764 40982 8820 41020
rect 9007 41078 9009 41130
rect 9061 41078 9063 41130
rect 8316 40406 8318 40458
rect 8370 40406 8372 40458
rect 8876 40516 8932 40526
rect 9007 40516 9063 41078
rect 8876 40422 8932 40460
rect 8988 40460 9063 40516
rect 8316 40404 8372 40406
rect 7756 40338 7812 40350
rect 8204 40348 8316 40404
rect 7308 40124 7700 40180
rect 7308 39732 7364 40124
rect 8092 39844 8148 39854
rect 8204 39844 8260 40348
rect 8316 40328 8372 40348
rect 8988 40404 9044 40460
rect 8988 40338 9044 40348
rect 8092 39842 8260 39844
rect 8092 39790 8094 39842
rect 8146 39790 8260 39842
rect 8092 39788 8260 39790
rect 8092 39778 8148 39788
rect 7252 39676 7364 39732
rect 6972 39618 7028 39630
rect 6412 39562 6524 39574
rect 6412 39510 6470 39562
rect 6522 39510 6524 39562
rect 6412 39508 6524 39510
rect 6468 39396 6524 39508
rect 6972 39566 6974 39618
rect 7026 39566 7028 39618
rect 6972 39564 7028 39566
rect 7140 39564 7196 39574
rect 6972 39562 7196 39564
rect 6972 39510 7142 39562
rect 7194 39510 7196 39562
rect 6972 39508 7196 39510
rect 6468 39330 6524 39340
rect 6804 39396 6860 39406
rect 6804 39394 6916 39396
rect 6804 39342 6806 39394
rect 6858 39342 6916 39394
rect 6804 39330 6916 39342
rect 5964 38724 6020 38734
rect 5964 38276 6020 38668
rect 6860 38500 6916 39330
rect 6972 38948 7028 39508
rect 7140 39498 7196 39508
rect 7252 39396 7308 39676
rect 7420 39564 7476 39574
rect 7700 39564 7756 39574
rect 7420 39562 7588 39564
rect 7420 39510 7422 39562
rect 7474 39510 7588 39562
rect 7420 39508 7588 39510
rect 7420 39498 7476 39508
rect 7252 39340 7364 39396
rect 6972 38882 7028 38892
rect 7084 38836 7140 38846
rect 7084 38742 7140 38780
rect 6748 38444 6916 38500
rect 7308 38500 7364 39340
rect 7308 38444 7476 38500
rect 6748 38388 6804 38444
rect 6748 38322 6804 38332
rect 5964 38220 6524 38276
rect 6468 38162 6524 38220
rect 6468 38110 6470 38162
rect 6522 38110 6524 38162
rect 6468 38098 6524 38110
rect 6748 38052 6804 38062
rect 6748 37958 6804 37996
rect 4844 37378 5012 37380
rect 4844 37326 4846 37378
rect 4898 37326 5012 37378
rect 4844 37324 5012 37326
rect 5292 37548 5684 37604
rect 5796 37826 5852 37838
rect 5796 37774 5798 37826
rect 5850 37774 5852 37826
rect 5796 37604 5852 37774
rect 6860 37716 6916 37726
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4844 36708 4900 37324
rect 5087 37268 5143 37278
rect 5068 37266 5143 37268
rect 5068 37214 5089 37266
rect 5141 37214 5143 37266
rect 5068 37202 5143 37214
rect 4172 36652 4452 36708
rect 4396 36594 4452 36652
rect 4396 36542 4398 36594
rect 4450 36542 4452 36594
rect 4396 36530 4452 36542
rect 4620 36652 4900 36708
rect 4956 37156 5012 37166
rect 4228 36484 4284 36494
rect 4228 36390 4284 36428
rect 4620 36482 4676 36652
rect 4620 36430 4622 36482
rect 4674 36430 4676 36482
rect 4620 36418 4676 36430
rect 4956 36426 5012 37100
rect 4956 36374 4958 36426
rect 5010 36374 5012 36426
rect 4844 35736 4900 35748
rect 4844 35700 4846 35736
rect 4898 35700 4900 35736
rect 4844 35634 4900 35644
rect 4284 35586 4340 35598
rect 4284 35534 4286 35586
rect 4338 35534 4340 35586
rect 4284 35140 4340 35534
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4732 35140 4788 35150
rect 4284 35084 4452 35140
rect 4264 34916 4320 34926
rect 4060 34860 4172 34916
rect 4116 34804 4172 34860
rect 4264 34914 4340 34916
rect 4264 34862 4266 34914
rect 4318 34862 4340 34914
rect 4264 34850 4340 34862
rect 4284 34804 4340 34850
rect 4116 34748 4228 34804
rect 4060 34580 4116 34590
rect 3388 34524 3948 34580
rect 2940 34178 2996 34188
rect 3500 34356 3556 34366
rect 3220 32788 3276 32798
rect 3220 32694 3276 32732
rect 3500 32788 3556 34300
rect 3892 34186 3948 34524
rect 3892 34134 3894 34186
rect 3946 34134 3948 34186
rect 3668 34018 3724 34030
rect 3668 33966 3670 34018
rect 3722 33966 3724 34018
rect 3668 33908 3724 33966
rect 3892 34020 3948 34134
rect 4060 34186 4116 34524
rect 4172 34356 4228 34748
rect 4284 34738 4340 34748
rect 4172 34290 4228 34300
rect 4060 34134 4062 34186
rect 4114 34134 4116 34186
rect 4060 34122 4116 34134
rect 4284 34244 4340 34254
rect 4284 34186 4340 34188
rect 4284 34134 4286 34186
rect 4338 34134 4340 34186
rect 4284 34122 4340 34134
rect 4396 34020 4452 35084
rect 4508 34916 4564 34926
rect 4508 34822 4564 34860
rect 3892 33964 4452 34020
rect 4732 34020 4788 35084
rect 4956 34916 5012 36374
rect 5068 36372 5124 37202
rect 5068 36306 5124 36316
rect 5180 35700 5236 35710
rect 4900 34860 5012 34916
rect 5068 35698 5236 35700
rect 5068 35646 5182 35698
rect 5234 35646 5236 35698
rect 5068 35644 5236 35646
rect 5068 34916 5124 35644
rect 5180 35634 5236 35644
rect 5292 35588 5348 37548
rect 5796 37538 5852 37548
rect 6524 37604 6580 37614
rect 6244 37322 6300 37334
rect 5964 37268 6020 37278
rect 5964 37174 6020 37212
rect 6244 37270 6246 37322
rect 6298 37270 6300 37322
rect 6244 37268 6300 37270
rect 6244 37202 6300 37212
rect 6412 37296 6468 37308
rect 6412 37244 6414 37296
rect 6466 37244 6468 37296
rect 6244 36932 6300 36942
rect 5796 36596 5852 36606
rect 5628 36540 5796 36596
rect 5628 36484 5684 36540
rect 5796 36502 5852 36540
rect 6244 36594 6300 36876
rect 6244 36542 6246 36594
rect 6298 36542 6300 36594
rect 5628 36260 5684 36428
rect 5572 36204 5684 36260
rect 5908 36372 5964 36382
rect 5404 35812 5460 35822
rect 5404 35718 5460 35756
rect 5572 35754 5628 36204
rect 5908 35922 5964 36316
rect 5908 35870 5910 35922
rect 5962 35870 5964 35922
rect 5908 35858 5964 35870
rect 5572 35702 5574 35754
rect 5626 35702 5628 35754
rect 5572 35690 5628 35702
rect 6076 35718 6132 35730
rect 6076 35666 6078 35718
rect 6130 35666 6132 35718
rect 5292 35532 5460 35588
rect 4900 34804 4956 34860
rect 5068 34850 5124 34860
rect 5180 34914 5236 34926
rect 5180 34862 5182 34914
rect 5234 34862 5236 34914
rect 4844 34748 4956 34804
rect 5180 34804 5236 34862
rect 4844 34242 4900 34748
rect 5180 34738 5236 34748
rect 5012 34690 5068 34702
rect 5012 34638 5014 34690
rect 5066 34638 5068 34690
rect 5012 34580 5068 34638
rect 5012 34514 5068 34524
rect 4844 34190 4846 34242
rect 4898 34190 4900 34242
rect 4844 34178 4900 34190
rect 5292 34356 5348 34366
rect 4732 33954 4788 33964
rect 3668 33842 3724 33852
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4116 33348 4172 33358
rect 3668 32788 3724 32798
rect 3500 32786 3724 32788
rect 3500 32734 3670 32786
rect 3722 32734 3724 32786
rect 3500 32732 3724 32734
rect 2604 32510 2606 32562
rect 2658 32510 2660 32562
rect 2604 32498 2660 32510
rect 2940 31892 2996 31902
rect 2604 31780 2660 31790
rect 2604 31686 2660 31724
rect 2940 31778 2996 31836
rect 3500 31892 3556 32732
rect 3668 32722 3724 32732
rect 4116 32788 4172 33292
rect 5124 33348 5180 33358
rect 5124 33254 5180 33292
rect 4116 32694 4172 32732
rect 4284 33234 4340 33246
rect 4284 33182 4286 33234
rect 4338 33182 4340 33234
rect 4284 32564 4340 33182
rect 5292 32574 5348 34300
rect 4396 32564 4452 32574
rect 4172 32562 4452 32564
rect 4172 32510 4398 32562
rect 4450 32510 4452 32562
rect 4172 32508 4452 32510
rect 4172 32004 4228 32508
rect 4396 32498 4452 32508
rect 5272 32562 5348 32574
rect 5272 32510 5274 32562
rect 5326 32510 5348 32562
rect 5272 32498 5348 32510
rect 4172 31938 4228 31948
rect 4284 32228 4340 32238
rect 3500 31826 3556 31836
rect 2940 31726 2942 31778
rect 2994 31726 2996 31778
rect 2940 31714 2996 31726
rect 3052 31780 3108 31790
rect 3612 31778 3668 31790
rect 3052 31610 3108 31724
rect 1596 30942 1598 30994
rect 1650 30942 1652 30994
rect 1596 29764 1652 30942
rect 2268 31554 2324 31566
rect 2268 31502 2270 31554
rect 2322 31502 2324 31554
rect 3052 31558 3054 31610
rect 3106 31558 3108 31610
rect 3052 31546 3108 31558
rect 3276 31722 3332 31734
rect 3276 31670 3278 31722
rect 3330 31670 3332 31722
rect 2268 30996 2324 31502
rect 3276 31220 3332 31670
rect 3612 31726 3614 31778
rect 3666 31726 3668 31778
rect 3612 31668 3668 31726
rect 3612 31602 3668 31612
rect 4172 31778 4228 31790
rect 4172 31726 4174 31778
rect 4226 31726 4228 31778
rect 3276 31164 3556 31220
rect 2380 30996 2436 31006
rect 2268 30994 2436 30996
rect 2268 30942 2382 30994
rect 2434 30942 2436 30994
rect 2268 30940 2436 30942
rect 2380 30930 2436 30940
rect 2492 30660 2548 30670
rect 1596 29708 2156 29764
rect 1596 28644 1652 29708
rect 2100 29650 2156 29708
rect 2100 29598 2102 29650
rect 2154 29598 2156 29650
rect 2100 29586 2156 29598
rect 2492 29538 2548 30604
rect 3052 30660 3108 30670
rect 3500 30660 3556 31164
rect 2828 30210 2884 30222
rect 2828 30158 2830 30210
rect 2882 30158 2884 30210
rect 2828 30100 2884 30158
rect 3052 30195 3108 30604
rect 3164 30604 3556 30660
rect 4172 30996 4228 31726
rect 4284 31778 4340 32172
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4844 32004 4900 32014
rect 4844 31910 4900 31948
rect 4284 31726 4286 31778
rect 4338 31726 4340 31778
rect 5292 31780 5348 32498
rect 4284 31714 4340 31726
rect 4452 31722 4508 31734
rect 4452 31670 4454 31722
rect 4506 31670 4508 31722
rect 5292 31714 5348 31724
rect 4452 31668 4508 31670
rect 4452 31602 4508 31612
rect 5124 31668 5180 31678
rect 4732 31164 5012 31220
rect 4284 30996 4340 31006
rect 4172 30994 4340 30996
rect 4172 30942 4286 30994
rect 4338 30942 4340 30994
rect 4172 30940 4340 30942
rect 3164 30322 3220 30604
rect 3164 30270 3166 30322
rect 3218 30270 3220 30322
rect 3164 30258 3220 30270
rect 3052 30143 3054 30195
rect 3106 30143 3108 30195
rect 3052 30131 3108 30143
rect 3500 30212 3556 30222
rect 3500 30118 3556 30156
rect 4172 30212 4228 30940
rect 4284 30930 4340 30940
rect 4732 30994 4788 31164
rect 4732 30942 4734 30994
rect 4786 30942 4788 30994
rect 4732 30930 4788 30942
rect 4844 30994 4900 31006
rect 4844 30942 4846 30994
rect 4898 30942 4900 30994
rect 4844 30772 4900 30942
rect 4844 30706 4900 30716
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4172 30146 4228 30156
rect 4376 30436 4432 30446
rect 4376 30210 4432 30380
rect 4376 30158 4378 30210
rect 4430 30158 4432 30210
rect 4376 30146 4432 30158
rect 2828 30034 2884 30044
rect 4620 30100 4676 30110
rect 4620 30006 4676 30044
rect 4956 30100 5012 31164
rect 5124 31106 5180 31612
rect 5124 31054 5126 31106
rect 5178 31054 5180 31106
rect 5124 31042 5180 31054
rect 5404 30884 5460 35532
rect 6076 35476 6132 35666
rect 6244 35724 6300 36542
rect 6244 35672 6246 35724
rect 6298 35672 6300 35724
rect 6244 35660 6300 35672
rect 6076 35410 6132 35420
rect 6412 35476 6468 37244
rect 6524 36596 6580 37548
rect 6748 37296 6804 37308
rect 6748 37244 6750 37296
rect 6802 37244 6804 37296
rect 6748 37156 6804 37244
rect 6748 37090 6804 37100
rect 6524 36530 6580 36540
rect 6636 36260 6692 36270
rect 6636 36166 6692 36204
rect 6860 35588 6916 37660
rect 7420 37604 7476 38444
rect 7532 38164 7588 39508
rect 7700 39562 7812 39564
rect 7700 39510 7702 39562
rect 7754 39510 7812 39562
rect 7700 39498 7812 39510
rect 7756 39060 7812 39498
rect 9044 39396 9100 39406
rect 9212 39396 9268 42700
rect 9660 42754 9940 42756
rect 9660 42702 9886 42754
rect 9938 42702 9940 42754
rect 9660 42700 9940 42702
rect 9660 42194 9716 42700
rect 9884 42690 9940 42700
rect 9996 42532 10052 43148
rect 9660 42142 9662 42194
rect 9714 42142 9716 42194
rect 9660 42130 9716 42142
rect 9884 42476 10052 42532
rect 9884 41524 9940 42476
rect 10108 42420 10164 44268
rect 10220 44258 10276 44268
rect 10668 43764 10724 44382
rect 11004 44324 11060 44334
rect 10780 44278 10836 44290
rect 10780 44226 10782 44278
rect 10834 44226 10836 44278
rect 11004 44230 11060 44268
rect 11788 44324 11844 44334
rect 12236 44324 12292 45500
rect 12348 45108 12404 45614
rect 12348 45042 12404 45052
rect 12684 45444 12740 45454
rect 12684 44546 12740 45388
rect 12796 44884 12852 45836
rect 13132 45890 13188 45902
rect 13132 45838 13134 45890
rect 13186 45838 13188 45890
rect 13020 45220 13076 45230
rect 13132 45220 13188 45838
rect 13020 45218 13188 45220
rect 13020 45166 13022 45218
rect 13074 45166 13188 45218
rect 13020 45164 13188 45166
rect 13020 45154 13076 45164
rect 12796 44818 12852 44828
rect 12684 44494 12686 44546
rect 12738 44494 12740 44546
rect 12684 44482 12740 44494
rect 11788 44322 12292 44324
rect 11788 44270 11790 44322
rect 11842 44270 12292 44322
rect 11788 44268 12292 44270
rect 13020 44324 13076 44334
rect 10780 43988 10836 44226
rect 11620 44100 11676 44110
rect 11620 44098 11732 44100
rect 11620 44046 11622 44098
rect 11674 44046 11732 44098
rect 11620 44034 11732 44046
rect 10780 43922 10836 43932
rect 10668 43698 10724 43708
rect 10220 43540 10276 43550
rect 10220 43204 10276 43484
rect 11004 43540 11060 43578
rect 11004 43474 11060 43484
rect 10220 43138 10276 43148
rect 10556 43314 10612 43326
rect 10556 43262 10558 43314
rect 10610 43262 10612 43314
rect 10556 43092 10612 43262
rect 10556 43026 10612 43036
rect 10108 42354 10164 42364
rect 11340 42868 11396 42878
rect 9996 42140 10388 42196
rect 9996 41970 10052 42140
rect 10332 42138 10388 42140
rect 10332 42086 10334 42138
rect 10386 42086 10388 42138
rect 10332 42074 10388 42086
rect 10668 42009 10724 42021
rect 9996 41918 9998 41970
rect 10050 41918 10052 41970
rect 9996 41906 10052 41918
rect 10332 41972 10388 41982
rect 10332 41878 10388 41916
rect 10668 41957 10670 42009
rect 10722 41957 10724 42009
rect 10556 41860 10612 41870
rect 9884 41468 10164 41524
rect 9884 41188 9940 41198
rect 10108 41188 10164 41468
rect 9884 41094 9940 41132
rect 9996 41132 10164 41188
rect 9716 40628 9772 40638
rect 9716 40534 9772 40572
rect 9996 40404 10052 41132
rect 10556 41086 10612 41804
rect 10668 41300 10724 41957
rect 10892 41970 10948 41982
rect 10892 41918 10894 41970
rect 10946 41918 10948 41970
rect 10892 41636 10948 41918
rect 11340 41860 11396 42812
rect 11676 42868 11732 44034
rect 11788 43652 11844 44268
rect 13020 44230 13076 44268
rect 12124 44100 12180 44110
rect 12012 44098 12180 44100
rect 12012 44046 12126 44098
rect 12178 44046 12180 44098
rect 12012 44044 12180 44046
rect 13356 44100 13412 46732
rect 13916 45862 13972 45874
rect 13916 45810 13918 45862
rect 13970 45810 13972 45862
rect 13468 45666 13524 45678
rect 13468 45614 13470 45666
rect 13522 45614 13524 45666
rect 13468 44772 13524 45614
rect 13916 45444 13972 45810
rect 14588 45780 14644 49200
rect 16156 45890 16212 49200
rect 17724 46340 17780 49200
rect 17724 46284 17892 46340
rect 16156 45838 16158 45890
rect 16210 45838 16212 45890
rect 16156 45826 16212 45838
rect 17500 45890 17556 45902
rect 17500 45838 17502 45890
rect 17554 45838 17556 45890
rect 14588 45714 14644 45724
rect 17500 45780 17556 45838
rect 17500 45714 17556 45724
rect 17164 45668 17220 45678
rect 17164 45574 17220 45612
rect 13916 45378 13972 45388
rect 15484 45108 15540 45118
rect 15484 45014 15540 45052
rect 16268 45108 16324 45118
rect 16268 45014 16324 45052
rect 16940 45106 16996 45118
rect 16940 45054 16942 45106
rect 16994 45054 16996 45106
rect 13468 44706 13524 44716
rect 13580 44994 13636 45006
rect 13580 44942 13582 44994
rect 13634 44942 13636 44994
rect 13580 44324 13636 44942
rect 13580 44258 13636 44268
rect 13916 44996 13972 45006
rect 13524 44100 13580 44110
rect 13356 44098 13580 44100
rect 13356 44046 13526 44098
rect 13578 44046 13580 44098
rect 13356 44044 13580 44046
rect 13916 44100 13972 44940
rect 16940 44996 16996 45054
rect 16940 44930 16996 44940
rect 17500 45108 17556 45118
rect 15596 44884 15652 44894
rect 15148 44660 15204 44670
rect 14476 44436 14532 44446
rect 14476 44434 14644 44436
rect 14476 44382 14478 44434
rect 14530 44382 14644 44434
rect 14476 44380 14644 44382
rect 14476 44370 14532 44380
rect 14140 44322 14196 44334
rect 14140 44270 14142 44322
rect 14194 44270 14196 44322
rect 13916 44044 14084 44100
rect 11788 43596 11936 43652
rect 11880 43540 11936 43596
rect 11880 43538 11956 43540
rect 11880 43486 11882 43538
rect 11934 43486 11956 43538
rect 11880 43474 11956 43486
rect 11676 42802 11732 42812
rect 11788 42644 11844 42654
rect 11340 41794 11396 41804
rect 11676 42642 11844 42644
rect 11676 42590 11790 42642
rect 11842 42590 11844 42642
rect 11676 42588 11844 42590
rect 10892 41570 10948 41580
rect 11508 41746 11564 41758
rect 11508 41694 11510 41746
rect 11562 41694 11564 41746
rect 11508 41636 11564 41694
rect 11508 41570 11564 41580
rect 11676 41300 11732 42588
rect 11788 42578 11844 42588
rect 11788 41970 11844 41982
rect 11788 41918 11790 41970
rect 11842 41918 11844 41970
rect 11788 41412 11844 41918
rect 11900 41972 11956 43474
rect 12012 42756 12068 44044
rect 12124 44034 12180 44044
rect 13524 44034 13580 44044
rect 13580 43652 13636 43662
rect 12124 43540 12180 43550
rect 12572 43540 12628 43550
rect 12124 43538 12628 43540
rect 12124 43486 12126 43538
rect 12178 43486 12574 43538
rect 12626 43486 12628 43538
rect 12124 43484 12628 43486
rect 12124 43474 12180 43484
rect 12572 43474 12628 43484
rect 13448 43540 13504 43550
rect 13448 43446 13504 43484
rect 12460 42868 12516 42878
rect 12460 42774 12516 42812
rect 13580 42868 13636 43596
rect 13692 43314 13748 43326
rect 13692 43262 13694 43314
rect 13746 43262 13748 43314
rect 13692 43204 13748 43262
rect 13692 43138 13748 43148
rect 13916 43316 13972 43326
rect 13580 42802 13636 42812
rect 12012 42690 12068 42700
rect 12572 42756 12628 42766
rect 12572 42687 12574 42700
rect 12626 42687 12628 42700
rect 12572 42662 12628 42687
rect 12908 42756 12964 42766
rect 12908 42662 12964 42700
rect 13804 42756 13860 42766
rect 13804 42662 13860 42700
rect 13916 42754 13972 43260
rect 13916 42702 13918 42754
rect 13970 42702 13972 42754
rect 13916 42644 13972 42702
rect 13916 42578 13972 42588
rect 14028 42420 14084 44044
rect 14140 43652 14196 44270
rect 14140 43586 14196 43596
rect 14364 44278 14420 44290
rect 14364 44226 14366 44278
rect 14418 44226 14420 44278
rect 14252 43568 14308 43580
rect 14252 43516 14254 43568
rect 14306 43516 14308 43568
rect 14252 43316 14308 43516
rect 14252 43250 14308 43260
rect 14196 42980 14252 42990
rect 14364 42980 14420 44226
rect 14588 43652 14644 44380
rect 14924 44210 14980 44222
rect 14924 44158 14926 44210
rect 14978 44158 14980 44210
rect 14924 43876 14980 44158
rect 14924 43810 14980 43820
rect 14588 43596 14980 43652
rect 14196 42978 14420 42980
rect 14196 42926 14198 42978
rect 14250 42926 14420 42978
rect 14196 42924 14420 42926
rect 14476 43577 14532 43589
rect 14476 43540 14478 43577
rect 14530 43540 14532 43577
rect 14196 42914 14252 42924
rect 14028 42364 14308 42420
rect 11900 41906 11956 41916
rect 12012 41970 12068 41982
rect 12012 41918 12014 41970
rect 12066 41918 12068 41970
rect 11788 41346 11844 41356
rect 11900 41748 11956 41758
rect 10668 41234 10724 41244
rect 11564 41244 11732 41300
rect 10892 41188 10948 41198
rect 10892 41094 10948 41132
rect 11564 41188 11620 41244
rect 11732 41155 11824 41188
rect 11732 41132 11770 41155
rect 10556 41074 10668 41086
rect 10556 41022 10614 41074
rect 10666 41022 10668 41074
rect 10556 41020 10668 41022
rect 10612 41010 10668 41020
rect 11228 40740 11284 40750
rect 10164 40628 10220 40638
rect 10164 40534 10220 40572
rect 10892 40628 10948 40638
rect 9660 40348 10052 40404
rect 10612 40402 10668 40414
rect 10612 40350 10614 40402
rect 10666 40350 10668 40402
rect 9492 39396 9548 39406
rect 9044 39394 9156 39396
rect 9044 39342 9046 39394
rect 9098 39342 9156 39394
rect 9044 39330 9156 39342
rect 9212 39394 9548 39396
rect 9212 39342 9494 39394
rect 9546 39342 9548 39394
rect 9212 39340 9548 39342
rect 7756 39004 8148 39060
rect 7532 38108 7680 38164
rect 7624 38019 7680 38108
rect 7624 37967 7626 38019
rect 7678 37967 7680 38019
rect 7624 37604 7680 37967
rect 7420 37538 7476 37548
rect 7532 37548 7680 37604
rect 7196 37380 7252 37390
rect 7196 37286 7252 37324
rect 7532 36708 7588 37548
rect 7756 37492 7812 39004
rect 8092 38890 8148 39004
rect 7868 38834 7924 38846
rect 7868 38782 7870 38834
rect 7922 38782 7924 38834
rect 8092 38838 8094 38890
rect 8146 38838 8148 38890
rect 8092 38826 8148 38838
rect 8204 38872 8260 38884
rect 7868 38724 7924 38782
rect 8204 38820 8206 38872
rect 8258 38820 8260 38872
rect 8204 38668 8260 38820
rect 8764 38836 8820 38846
rect 8764 38742 8820 38780
rect 8932 38778 8988 38790
rect 8932 38726 8934 38778
rect 8986 38726 8988 38778
rect 8932 38668 8988 38726
rect 7868 38658 7924 38668
rect 7980 38612 8260 38668
rect 8652 38612 8988 38668
rect 7644 37436 7812 37492
rect 7868 38276 7924 38286
rect 7980 38276 8036 38612
rect 7868 38274 8036 38276
rect 7868 38222 7870 38274
rect 7922 38222 8036 38274
rect 7868 38220 8036 38222
rect 7644 37380 7700 37436
rect 7644 37266 7700 37324
rect 7644 37214 7646 37266
rect 7698 37214 7700 37266
rect 7644 37202 7700 37214
rect 7756 37268 7812 37278
rect 7868 37268 7924 38220
rect 8652 38218 8708 38612
rect 8652 38166 8654 38218
rect 8706 38166 8708 38218
rect 8652 38154 8708 38166
rect 8428 38050 8484 38062
rect 8428 37998 8430 38050
rect 8482 37998 8484 38050
rect 8036 37380 8092 37390
rect 8036 37286 8092 37324
rect 8428 37380 8484 37998
rect 8764 38050 8820 38062
rect 8764 37998 8766 38050
rect 8818 37998 8820 38050
rect 8764 37492 8820 37998
rect 9100 37502 9156 39330
rect 9436 39330 9548 39340
rect 8764 37426 8820 37436
rect 9044 37492 9156 37502
rect 9100 37436 9156 37492
rect 9212 39060 9268 39070
rect 9044 37398 9100 37436
rect 8428 37314 8484 37324
rect 7756 37266 7924 37268
rect 7756 37214 7758 37266
rect 7810 37214 7924 37266
rect 7756 37212 7924 37214
rect 7756 37202 7812 37212
rect 8596 37154 8652 37166
rect 8596 37102 8598 37154
rect 8650 37102 8652 37154
rect 8148 36932 8204 36942
rect 7532 36652 7700 36708
rect 6972 36484 7028 36494
rect 7252 36484 7308 36494
rect 7532 36484 7588 36494
rect 6972 36482 7308 36484
rect 6972 36430 6974 36482
rect 7026 36430 7254 36482
rect 7306 36430 7308 36482
rect 6972 36428 7308 36430
rect 6972 36418 7028 36428
rect 7252 36418 7308 36428
rect 7420 36482 7588 36484
rect 7420 36430 7534 36482
rect 7586 36430 7588 36482
rect 7420 36428 7588 36430
rect 6972 36260 7028 36270
rect 6972 35698 7028 36204
rect 7420 35924 7476 36428
rect 7532 36418 7588 36428
rect 7644 36148 7700 36652
rect 8148 36594 8204 36876
rect 8596 36932 8652 37102
rect 8596 36866 8652 36876
rect 9212 36596 9268 39004
rect 9436 38834 9492 39330
rect 9660 39060 9716 40348
rect 10612 40180 10668 40350
rect 10892 40402 10948 40572
rect 10892 40350 10894 40402
rect 10946 40350 10948 40402
rect 11228 40446 11284 40684
rect 11228 40394 11230 40446
rect 11282 40394 11284 40446
rect 11228 40382 11284 40394
rect 11452 40404 11508 40414
rect 10892 40338 10948 40350
rect 11564 40404 11620 41132
rect 11676 41103 11770 41132
rect 11822 41103 11824 41155
rect 11676 41091 11824 41103
rect 11676 41076 11788 41091
rect 11676 41010 11732 41020
rect 11900 40964 11956 41692
rect 12012 41410 12068 41918
rect 12460 41970 12516 41982
rect 13020 41972 13076 41982
rect 12460 41918 12462 41970
rect 12514 41918 12516 41970
rect 12292 41748 12348 41758
rect 12292 41654 12348 41692
rect 12460 41636 12516 41918
rect 12796 41970 13076 41972
rect 12796 41918 13022 41970
rect 13074 41918 13076 41970
rect 12796 41916 13076 41918
rect 12796 41860 12852 41916
rect 13020 41906 13076 41916
rect 13896 41972 13952 41982
rect 13896 41970 13972 41972
rect 13896 41918 13898 41970
rect 13950 41918 13972 41970
rect 13896 41906 13972 41918
rect 12796 41794 12852 41804
rect 13020 41636 13076 41646
rect 12460 41580 12964 41636
rect 12012 41358 12014 41410
rect 12066 41358 12068 41410
rect 12012 41300 12068 41358
rect 12348 41468 12852 41524
rect 12348 41300 12404 41468
rect 12012 41244 12404 41300
rect 12460 41300 12516 41310
rect 12684 41300 12740 41310
rect 12460 41206 12516 41244
rect 12572 41244 12684 41300
rect 12572 41142 12628 41244
rect 12684 41234 12740 41244
rect 12572 41090 12574 41142
rect 12626 41090 12628 41142
rect 12796 41186 12852 41468
rect 12796 41134 12798 41186
rect 12850 41134 12852 41186
rect 12796 41122 12852 41134
rect 11788 40908 11956 40964
rect 12012 41076 12068 41086
rect 11676 40404 11732 40414
rect 11564 40402 11732 40404
rect 11564 40350 11678 40402
rect 11730 40350 11732 40402
rect 11564 40348 11732 40350
rect 11340 40292 11396 40302
rect 11340 40198 11396 40236
rect 10444 40124 10668 40180
rect 11452 40180 11508 40348
rect 11676 40338 11732 40348
rect 11788 40402 11844 40908
rect 12012 40852 12068 41020
rect 11788 40350 11790 40402
rect 11842 40350 11844 40402
rect 11974 40796 12068 40852
rect 11974 40440 12030 40796
rect 11974 40388 11976 40440
rect 12028 40388 12030 40440
rect 11974 40376 12030 40388
rect 12348 40628 12404 40638
rect 11788 40338 11844 40350
rect 12124 40292 12180 40302
rect 11452 40124 11844 40180
rect 10332 39844 10388 39854
rect 10332 39750 10388 39788
rect 9996 39618 10052 39630
rect 9996 39566 9998 39618
rect 10050 39566 10052 39618
rect 9996 39508 10052 39566
rect 9996 39442 10052 39452
rect 9828 39396 9884 39406
rect 9828 39394 9940 39396
rect 9828 39342 9830 39394
rect 9882 39342 9940 39394
rect 9828 39330 9940 39342
rect 9660 38994 9716 39004
rect 9436 38782 9438 38834
rect 9490 38782 9492 38834
rect 9436 38724 9492 38782
rect 9436 38658 9492 38668
rect 9772 38218 9828 38230
rect 9772 38166 9774 38218
rect 9826 38166 9828 38218
rect 9436 38050 9492 38062
rect 9660 38052 9716 38062
rect 9436 37998 9438 38050
rect 9490 37998 9492 38050
rect 9436 37492 9492 37998
rect 9436 37426 9492 37436
rect 9548 38050 9716 38052
rect 9548 37998 9662 38050
rect 9714 37998 9716 38050
rect 9548 37996 9716 37998
rect 9548 36708 9604 37996
rect 9660 37986 9716 37996
rect 9660 37828 9716 37838
rect 9660 37166 9716 37772
rect 9772 37716 9828 38166
rect 9884 38052 9940 39330
rect 10332 39060 10388 39070
rect 10220 38722 10276 38734
rect 10220 38670 10222 38722
rect 10274 38670 10276 38722
rect 10220 38500 10276 38670
rect 10332 38668 10388 39004
rect 10444 38836 10500 40124
rect 10780 39562 10836 39574
rect 10780 39510 10782 39562
rect 10834 39510 10836 39562
rect 10780 39060 10836 39510
rect 11116 39562 11172 39574
rect 11116 39510 11118 39562
rect 11170 39510 11172 39562
rect 11116 39172 11172 39510
rect 11284 39562 11340 39574
rect 11284 39510 11286 39562
rect 11338 39510 11340 39562
rect 11284 39508 11340 39510
rect 11284 39442 11340 39452
rect 11788 39406 11844 40124
rect 12124 39618 12180 40236
rect 12348 40290 12404 40572
rect 12572 40516 12628 41090
rect 12572 40450 12628 40460
rect 12796 40852 12852 40862
rect 12796 40402 12852 40796
rect 12908 40740 12964 41580
rect 12908 40674 12964 40684
rect 12796 40350 12798 40402
rect 12850 40350 12852 40402
rect 12796 40338 12852 40350
rect 12908 40404 12964 40414
rect 12348 40238 12350 40290
rect 12402 40238 12404 40290
rect 12348 40226 12404 40238
rect 12908 39854 12964 40348
rect 12852 39842 12964 39854
rect 12852 39790 12854 39842
rect 12906 39790 12964 39842
rect 12852 39788 12964 39790
rect 12852 39778 12908 39788
rect 12124 39566 12126 39618
rect 12178 39566 12180 39618
rect 12012 39508 12068 39518
rect 11788 39396 11900 39406
rect 11788 39394 11956 39396
rect 11788 39342 11846 39394
rect 11898 39342 11956 39394
rect 11788 39340 11956 39342
rect 11844 39330 11956 39340
rect 11676 39284 11732 39294
rect 11116 39116 11508 39172
rect 10780 38994 10836 39004
rect 10444 38770 10500 38780
rect 10332 38612 10500 38668
rect 10444 38500 10500 38612
rect 10444 38444 10836 38500
rect 10220 38434 10276 38444
rect 10108 38052 10164 38062
rect 9884 38050 10164 38052
rect 9884 37998 10110 38050
rect 10162 37998 10164 38050
rect 9884 37996 10164 37998
rect 10108 37986 10164 37996
rect 10220 38052 10276 38062
rect 9772 37660 9996 37716
rect 9940 37322 9996 37660
rect 9940 37270 9942 37322
rect 9994 37270 9996 37322
rect 10108 37380 10164 37390
rect 10220 37380 10276 37996
rect 10780 37492 10836 38444
rect 10984 37994 11040 38006
rect 10984 37942 10986 37994
rect 11038 37942 11040 37994
rect 10984 37828 11040 37942
rect 11228 37940 11284 37950
rect 10984 37762 11040 37772
rect 11116 37938 11284 37940
rect 11116 37886 11230 37938
rect 11282 37886 11284 37938
rect 11116 37884 11284 37886
rect 10108 37378 10276 37380
rect 10108 37326 10110 37378
rect 10162 37326 10276 37378
rect 10108 37324 10276 37326
rect 10332 37436 10836 37492
rect 10108 37314 10164 37324
rect 9940 37258 9996 37270
rect 10332 37266 10388 37436
rect 10332 37214 10334 37266
rect 10386 37214 10388 37266
rect 10332 37202 10388 37214
rect 9660 37154 9772 37166
rect 9660 37102 9718 37154
rect 9770 37102 9772 37154
rect 9660 37100 9772 37102
rect 9716 37044 9772 37100
rect 10556 37044 10612 37436
rect 11116 37380 11172 37884
rect 11228 37874 11284 37884
rect 11452 37828 11508 39116
rect 11452 37762 11508 37772
rect 11564 38724 11620 38734
rect 10668 37324 11172 37380
rect 10668 37322 10724 37324
rect 10668 37270 10670 37322
rect 10722 37270 10724 37322
rect 10668 37258 10724 37270
rect 10556 36988 10724 37044
rect 9716 36978 9772 36988
rect 9548 36642 9604 36652
rect 10500 36708 10556 36718
rect 10500 36614 10556 36652
rect 8148 36542 8150 36594
rect 8202 36542 8204 36594
rect 8148 36530 8204 36542
rect 9100 36540 9268 36596
rect 7756 36484 7812 36494
rect 8316 36484 8372 36494
rect 7756 36482 8036 36484
rect 7756 36430 7758 36482
rect 7810 36430 8036 36482
rect 7756 36428 8036 36430
rect 7756 36418 7812 36428
rect 7644 36082 7700 36092
rect 6972 35646 6974 35698
rect 7026 35646 7028 35698
rect 6972 35634 7028 35646
rect 7084 35868 7476 35924
rect 7980 35924 8036 36428
rect 8204 36260 8260 36270
rect 7980 35868 8148 35924
rect 6412 35410 6468 35420
rect 6692 35532 6916 35588
rect 6692 35028 6748 35532
rect 6692 35026 6804 35028
rect 6692 34974 6694 35026
rect 6746 34974 6804 35026
rect 6692 34962 6804 34974
rect 7084 35026 7140 35868
rect 7084 34974 7086 35026
rect 7138 34974 7140 35026
rect 7084 34962 7140 34974
rect 7980 35364 8036 35374
rect 5964 34916 6020 34926
rect 5852 34914 6020 34916
rect 5852 34862 5966 34914
rect 6018 34862 6020 34914
rect 5852 34860 6020 34862
rect 5684 34802 5740 34814
rect 5684 34750 5686 34802
rect 5738 34750 5740 34802
rect 5572 34580 5628 34590
rect 5572 34186 5628 34524
rect 5684 34468 5740 34750
rect 5684 34402 5740 34412
rect 5572 34134 5574 34186
rect 5626 34134 5628 34186
rect 5740 34244 5796 34254
rect 5852 34244 5908 34860
rect 5964 34850 6020 34860
rect 6188 34914 6244 34926
rect 6188 34862 6190 34914
rect 6242 34862 6244 34914
rect 6188 34356 6244 34862
rect 6188 34290 6244 34300
rect 5740 34242 5908 34244
rect 5740 34190 5742 34242
rect 5794 34190 5908 34242
rect 5740 34188 5908 34190
rect 6300 34244 6356 34254
rect 5740 34178 5796 34188
rect 6300 34186 6356 34188
rect 5572 33908 5628 34134
rect 5964 34130 6020 34142
rect 5964 34078 5966 34130
rect 6018 34078 6020 34130
rect 6300 34134 6302 34186
rect 6354 34134 6356 34186
rect 6300 34122 6356 34134
rect 6636 34132 6692 34142
rect 6412 34130 6692 34132
rect 5964 34020 6020 34078
rect 6412 34078 6638 34130
rect 6690 34078 6692 34130
rect 6412 34076 6692 34078
rect 6412 34020 6468 34076
rect 6636 34066 6692 34076
rect 6748 34132 6804 34962
rect 7308 34916 7364 34926
rect 6916 34858 6972 34870
rect 6916 34806 6918 34858
rect 6970 34806 6972 34858
rect 7308 34822 7364 34860
rect 7532 34858 7588 34870
rect 6916 34580 6972 34806
rect 6916 34514 6972 34524
rect 7532 34806 7534 34858
rect 7586 34806 7588 34858
rect 7532 34804 7588 34806
rect 7140 34356 7196 34366
rect 6748 34066 6804 34076
rect 6860 34244 6916 34254
rect 6860 34130 6916 34188
rect 7140 34242 7196 34300
rect 7140 34190 7142 34242
rect 7194 34190 7196 34242
rect 7140 34178 7196 34190
rect 6860 34078 6862 34130
rect 6914 34078 6916 34130
rect 5964 33964 6468 34020
rect 5572 33842 5628 33852
rect 6188 33348 6244 33358
rect 6076 33290 6132 33302
rect 6076 33238 6078 33290
rect 6130 33238 6132 33290
rect 6188 33254 6244 33292
rect 6076 33236 6132 33238
rect 6076 33170 6132 33180
rect 5908 33124 5964 33134
rect 5740 33122 5964 33124
rect 5740 33070 5910 33122
rect 5962 33070 5964 33122
rect 5740 33068 5964 33070
rect 5516 32338 5572 32350
rect 5516 32286 5518 32338
rect 5570 32286 5572 32338
rect 5516 32116 5572 32286
rect 5740 32340 5796 33068
rect 5908 33058 5964 33068
rect 6300 32900 6356 33964
rect 5740 32274 5796 32284
rect 5964 32844 6356 32900
rect 6524 33908 6580 33918
rect 6860 33908 6916 34078
rect 5964 32562 6020 32844
rect 5964 32510 5966 32562
rect 6018 32510 6020 32562
rect 5964 32116 6020 32510
rect 5516 32060 6020 32116
rect 6076 32564 6132 32574
rect 6076 32004 6132 32508
rect 6242 32564 6298 32574
rect 6242 32562 6300 32564
rect 6242 32510 6244 32562
rect 6296 32510 6300 32562
rect 6242 32498 6300 32510
rect 6244 32116 6300 32498
rect 6524 32340 6580 33852
rect 6636 33852 6916 33908
rect 7532 33908 7588 34748
rect 7980 34356 8036 35308
rect 8092 35150 8148 35868
rect 8204 35364 8260 36204
rect 8204 35298 8260 35308
rect 8092 35138 8204 35150
rect 8092 35086 8150 35138
rect 8202 35086 8204 35138
rect 8092 35084 8204 35086
rect 8148 35074 8204 35084
rect 8092 34356 8148 34366
rect 7980 34354 8148 34356
rect 7980 34302 8094 34354
rect 8146 34302 8148 34354
rect 7980 34300 8148 34302
rect 8092 34290 8148 34300
rect 8092 34132 8148 34142
rect 6636 32564 6692 33852
rect 7532 33842 7588 33852
rect 7700 34018 7756 34030
rect 7700 33966 7702 34018
rect 7754 33966 7756 34018
rect 7700 33908 7756 33966
rect 6636 32498 6692 32508
rect 6748 33684 6804 33694
rect 6636 32340 6692 32350
rect 6524 32338 6692 32340
rect 6524 32286 6638 32338
rect 6690 32286 6692 32338
rect 6524 32284 6692 32286
rect 6636 32274 6692 32284
rect 6244 32060 6356 32116
rect 6076 31938 6132 31948
rect 5628 31892 5684 31902
rect 5628 31778 5684 31836
rect 5628 31726 5630 31778
rect 5682 31726 5684 31778
rect 5628 31714 5684 31726
rect 6076 31780 6132 31790
rect 6188 31780 6244 31790
rect 6132 31778 6244 31780
rect 6132 31726 6190 31778
rect 6242 31726 6244 31778
rect 6132 31724 6244 31726
rect 4956 30034 5012 30044
rect 5180 30828 5460 30884
rect 5908 30884 5964 30894
rect 2492 29486 2494 29538
rect 2546 29486 2548 29538
rect 2492 29474 2548 29486
rect 3052 29652 3108 29662
rect 3052 29482 3108 29596
rect 4956 29652 5012 29662
rect 3052 29430 3054 29482
rect 3106 29430 3108 29482
rect 2772 29370 2828 29382
rect 1820 29316 1876 29326
rect 1820 28754 1876 29260
rect 2772 29318 2774 29370
rect 2826 29318 2828 29370
rect 2772 29316 2828 29318
rect 2772 29250 2828 29260
rect 3052 28980 3108 29430
rect 3276 29540 3332 29550
rect 3276 29482 3332 29484
rect 3276 29430 3278 29482
rect 3330 29430 3332 29482
rect 3276 29418 3332 29430
rect 3724 29428 3780 29466
rect 3724 29362 3780 29372
rect 4600 29426 4656 29438
rect 4600 29374 4602 29426
rect 4654 29374 4656 29426
rect 4600 29316 4656 29374
rect 4600 29250 4656 29260
rect 4844 29202 4900 29214
rect 4844 29150 4846 29202
rect 4898 29150 4900 29202
rect 4476 29036 4740 29046
rect 1820 28702 1822 28754
rect 1874 28702 1876 28754
rect 1820 28690 1876 28702
rect 2604 28924 3108 28980
rect 4060 28980 4116 28990
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 1708 28644 1764 28654
rect 1596 28588 1708 28644
rect 1596 27858 1652 28588
rect 1708 28578 1764 28588
rect 1596 27806 1598 27858
rect 1650 27806 1652 27858
rect 1596 27794 1652 27806
rect 2380 27746 2436 27758
rect 2380 27694 2382 27746
rect 2434 27694 2436 27746
rect 2380 27188 2436 27694
rect 2604 27524 2660 28924
rect 3724 28756 3780 28766
rect 3724 28662 3780 28700
rect 2604 27468 3108 27524
rect 2828 27300 2884 27310
rect 2716 27188 2772 27198
rect 2380 27186 2772 27188
rect 2380 27134 2718 27186
rect 2770 27134 2772 27186
rect 2380 27132 2772 27134
rect 2716 27122 2772 27132
rect 2828 27059 2884 27244
rect 2828 27007 2830 27059
rect 2882 27007 2884 27059
rect 2828 26995 2884 27007
rect 3052 27076 3108 27468
rect 3052 26982 3108 27020
rect 3724 27074 3780 27086
rect 3724 27022 3726 27074
rect 3778 27022 3780 27074
rect 1596 26292 1652 26302
rect 3164 26292 3220 26302
rect 1596 26290 1764 26292
rect 1596 26238 1598 26290
rect 1650 26238 1764 26290
rect 1596 26236 1764 26238
rect 1596 26226 1652 26236
rect 1708 26180 1764 26236
rect 3052 26290 3220 26292
rect 3052 26238 3166 26290
rect 3218 26238 3220 26290
rect 3052 26236 3220 26238
rect 1708 24948 1764 26124
rect 2548 26180 2604 26190
rect 2548 26086 2604 26124
rect 1932 26068 1988 26078
rect 1932 25974 1988 26012
rect 2660 25732 2716 25742
rect 2660 25638 2716 25676
rect 2268 25506 2324 25518
rect 2268 25454 2270 25506
rect 2322 25454 2324 25506
rect 1708 24882 1764 24892
rect 2156 25396 2212 25406
rect 2156 24946 2212 25340
rect 2156 24894 2158 24946
rect 2210 24894 2212 24946
rect 2156 24882 2212 24894
rect 2268 24948 2324 25454
rect 2380 25506 2436 25518
rect 2380 25454 2382 25506
rect 2434 25454 2436 25506
rect 2380 25172 2436 25454
rect 3052 25172 3108 26236
rect 3164 26226 3220 26236
rect 3332 26234 3388 26246
rect 3332 26182 3334 26234
rect 3386 26182 3388 26234
rect 3332 25732 3388 26182
rect 3276 25676 3388 25732
rect 3276 25508 3332 25676
rect 3724 25618 3780 27022
rect 3948 27074 4004 27086
rect 3948 27022 3950 27074
rect 4002 27022 4004 27074
rect 3836 26964 3892 26974
rect 3836 26290 3892 26908
rect 3948 26908 4004 27022
rect 4060 27076 4116 28924
rect 4172 28868 4228 28878
rect 4172 27300 4228 28812
rect 4844 28868 4900 29150
rect 4844 28802 4900 28812
rect 4956 28654 5012 29596
rect 4508 28644 4564 28654
rect 4900 28644 5012 28654
rect 4564 28642 5012 28644
rect 4564 28590 4902 28642
rect 4954 28590 5012 28642
rect 4564 28588 5012 28590
rect 5068 29428 5124 29438
rect 4508 28550 4564 28588
rect 4900 28550 4956 28588
rect 4900 28026 4956 28038
rect 4900 27974 4902 28026
rect 4954 27974 4956 28026
rect 4900 27972 4956 27974
rect 4900 27906 4956 27916
rect 4284 27860 4340 27870
rect 4732 27860 4788 27870
rect 4284 27858 4788 27860
rect 4284 27806 4286 27858
rect 4338 27806 4734 27858
rect 4786 27806 4788 27858
rect 4284 27804 4788 27806
rect 4284 27794 4340 27804
rect 4732 27794 4788 27804
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 5068 27310 5124 29372
rect 5180 28420 5236 30828
rect 5908 30790 5964 30828
rect 5516 30210 5572 30222
rect 5516 30158 5518 30210
rect 5570 30158 5572 30210
rect 5516 29652 5572 30158
rect 5348 29594 5404 29606
rect 5348 29542 5350 29594
rect 5402 29542 5404 29594
rect 5516 29586 5572 29596
rect 5740 29764 5796 29774
rect 5348 29540 5404 29542
rect 5348 29474 5404 29484
rect 5628 29540 5684 29550
rect 5516 29426 5572 29438
rect 5516 29374 5518 29426
rect 5570 29374 5572 29426
rect 5516 29316 5572 29374
rect 5516 28980 5572 29260
rect 5516 28868 5572 28924
rect 5180 28354 5236 28364
rect 5292 28812 5572 28868
rect 5292 27748 5348 28812
rect 5628 28644 5684 29484
rect 5740 29316 5796 29708
rect 5852 29540 5908 29550
rect 5852 29470 5908 29484
rect 5852 29418 5854 29470
rect 5906 29418 5908 29470
rect 5852 29406 5908 29418
rect 5740 29314 6020 29316
rect 5740 29262 5742 29314
rect 5794 29262 6020 29314
rect 5740 29260 6020 29262
rect 5740 29250 5796 29260
rect 5460 27972 5516 27982
rect 5628 27972 5684 28588
rect 5740 28868 5796 28878
rect 5740 28604 5796 28812
rect 5740 28552 5742 28604
rect 5794 28552 5796 28604
rect 5964 28644 6020 29260
rect 6076 29204 6132 31724
rect 6188 31714 6244 31724
rect 6300 31610 6356 32060
rect 6300 31558 6302 31610
rect 6354 31558 6356 31610
rect 6300 31546 6356 31558
rect 6748 31556 6804 33628
rect 7700 33684 7756 33852
rect 7700 33618 7756 33628
rect 6972 33348 7028 33358
rect 6972 33346 7252 33348
rect 6972 33294 6974 33346
rect 7026 33294 7252 33346
rect 6972 33292 7252 33294
rect 6972 33282 7028 33292
rect 6580 31500 6804 31556
rect 7084 33124 7140 33134
rect 7084 32002 7140 33068
rect 7196 32786 7252 33292
rect 8092 32788 8148 34076
rect 8316 33460 8372 36428
rect 8428 36484 8484 36494
rect 8428 36482 8596 36484
rect 8428 36430 8430 36482
rect 8482 36430 8596 36482
rect 8428 36428 8596 36430
rect 8428 36418 8484 36428
rect 8428 35252 8484 35262
rect 8428 34914 8484 35196
rect 8428 34862 8430 34914
rect 8482 34862 8484 34914
rect 8428 34804 8484 34862
rect 8428 34738 8484 34748
rect 8428 34130 8484 34142
rect 8428 34078 8430 34130
rect 8482 34078 8484 34130
rect 8428 33796 8484 34078
rect 8428 33730 8484 33740
rect 8540 33684 8596 36428
rect 8988 36148 9044 36158
rect 8876 35812 8932 35822
rect 8876 35718 8932 35756
rect 8652 34916 8708 34926
rect 8652 34822 8708 34860
rect 8988 34356 9044 36092
rect 9100 36036 9156 36540
rect 9548 36484 9604 36494
rect 9304 36426 9360 36438
rect 9304 36374 9306 36426
rect 9358 36374 9360 36426
rect 9548 36390 9604 36428
rect 9884 36482 9940 36494
rect 9884 36430 9886 36482
rect 9938 36430 9940 36482
rect 9304 36372 9360 36374
rect 9304 36306 9360 36316
rect 9100 35980 9380 36036
rect 9212 34916 9268 34926
rect 9212 34822 9268 34860
rect 8988 34290 9044 34300
rect 9100 34804 9156 34814
rect 9100 34130 9156 34748
rect 9324 34692 9380 35980
rect 9884 35924 9940 36430
rect 10052 36260 10108 36270
rect 10668 36260 10724 36988
rect 10780 36482 10836 37324
rect 11284 37156 11340 37166
rect 11284 36596 11340 37100
rect 11116 36540 11340 36596
rect 11452 36820 11508 36830
rect 10780 36430 10782 36482
rect 10834 36430 10836 36482
rect 10780 36418 10836 36430
rect 10892 36482 10948 36494
rect 10892 36430 10894 36482
rect 10946 36430 10948 36482
rect 10892 36260 10948 36430
rect 10052 36258 10388 36260
rect 10052 36206 10054 36258
rect 10106 36206 10388 36258
rect 10052 36204 10388 36206
rect 10052 36194 10108 36204
rect 9548 35868 9940 35924
rect 9548 35822 9604 35868
rect 9492 35812 9604 35822
rect 9548 35756 9604 35812
rect 9492 35754 9548 35756
rect 9492 35702 9494 35754
rect 9546 35702 9548 35754
rect 9492 35690 9548 35702
rect 9660 35728 9716 35740
rect 9660 35676 9662 35728
rect 9714 35676 9716 35728
rect 9455 34916 9511 34926
rect 9455 34822 9511 34860
rect 9660 34916 9716 35676
rect 9884 35737 9940 35749
rect 9884 35685 9886 35737
rect 9938 35685 9940 35737
rect 9884 35364 9940 35685
rect 9884 35298 9940 35308
rect 10332 35252 10388 36204
rect 10444 36204 10948 36260
rect 10444 35810 10500 36204
rect 10444 35758 10446 35810
rect 10498 35758 10500 35810
rect 10444 35746 10500 35758
rect 11116 35812 11172 36540
rect 11452 36482 11508 36764
rect 11452 36430 11454 36482
rect 11506 36430 11508 36482
rect 11452 36148 11508 36430
rect 11452 36082 11508 36092
rect 11564 36036 11620 38668
rect 11676 38052 11732 39228
rect 11900 38052 11956 39330
rect 12012 38836 12068 39452
rect 12124 39060 12180 39566
rect 12292 39620 12348 39630
rect 12292 39526 12348 39564
rect 12572 39618 12628 39630
rect 12572 39566 12574 39618
rect 12626 39566 12628 39618
rect 12460 39508 12516 39518
rect 12460 39414 12516 39452
rect 12124 38994 12180 39004
rect 12012 38780 12180 38836
rect 12124 38722 12180 38780
rect 12124 38670 12126 38722
rect 12178 38670 12180 38722
rect 12124 38658 12180 38670
rect 12124 38218 12180 38230
rect 12124 38166 12126 38218
rect 12178 38166 12180 38218
rect 12012 38052 12068 38062
rect 11900 38050 12068 38052
rect 11900 37998 12014 38050
rect 12066 37998 12068 38050
rect 11900 37996 12068 37998
rect 11676 37986 11732 37996
rect 12012 37940 12068 37996
rect 12124 38052 12180 38166
rect 12572 38218 12628 39566
rect 12728 39060 12784 39070
rect 12728 38872 12784 39004
rect 12728 38820 12730 38872
rect 12782 38820 12784 38872
rect 12728 38808 12784 38820
rect 12572 38166 12574 38218
rect 12626 38166 12628 38218
rect 12572 38154 12628 38166
rect 12124 37986 12180 37996
rect 12572 38052 12628 38062
rect 12572 37958 12628 37996
rect 12796 38050 12852 38062
rect 12796 37998 12798 38050
rect 12850 37998 12852 38050
rect 12012 37874 12068 37884
rect 11676 37828 11732 37838
rect 11676 37266 11732 37772
rect 12796 37390 12852 37998
rect 12460 37380 12516 37390
rect 12796 37378 12908 37390
rect 12796 37326 12854 37378
rect 12906 37326 12908 37378
rect 12796 37324 12908 37326
rect 11676 37214 11678 37266
rect 11730 37214 11732 37266
rect 11676 36484 11732 37214
rect 12012 37281 12068 37293
rect 12012 37229 12014 37281
rect 12066 37229 12068 37281
rect 12012 36820 12068 37229
rect 12348 37266 12404 37278
rect 12348 37214 12350 37266
rect 12402 37214 12404 37266
rect 12124 37156 12180 37166
rect 12348 37156 12404 37214
rect 12124 37154 12348 37156
rect 12124 37102 12126 37154
rect 12178 37102 12348 37154
rect 12124 37100 12348 37102
rect 12124 37090 12180 37100
rect 12348 37062 12404 37100
rect 12012 36754 12068 36764
rect 12460 36708 12516 37324
rect 12852 37314 12908 37324
rect 12572 37268 12628 37278
rect 12572 37156 12628 37212
rect 12572 37100 12740 37156
rect 12124 36652 12516 36708
rect 11788 36484 11844 36494
rect 11676 36482 11844 36484
rect 11676 36430 11790 36482
rect 11842 36430 11844 36482
rect 11676 36428 11844 36430
rect 11788 36260 11844 36428
rect 11788 36194 11844 36204
rect 11564 35980 11732 36036
rect 11116 35746 11172 35756
rect 11004 35700 11060 35710
rect 10668 35698 11060 35700
rect 10668 35646 11006 35698
rect 11058 35646 11060 35698
rect 10668 35644 11060 35646
rect 10332 35196 10612 35252
rect 9324 34636 9492 34692
rect 9100 34078 9102 34130
rect 9154 34078 9156 34130
rect 9100 34066 9156 34078
rect 8764 33908 8820 33918
rect 8764 33906 9156 33908
rect 8764 33854 8766 33906
rect 8818 33854 9156 33906
rect 8764 33852 9156 33854
rect 8764 33842 8820 33852
rect 8540 33628 9044 33684
rect 7196 32734 7198 32786
rect 7250 32734 7252 32786
rect 7196 32722 7252 32734
rect 7532 32732 7924 32788
rect 7532 32562 7588 32732
rect 7868 32730 7924 32732
rect 7868 32678 7870 32730
rect 7922 32678 7924 32730
rect 7868 32666 7924 32678
rect 7980 32732 8148 32788
rect 8204 33404 8372 33460
rect 7532 32510 7534 32562
rect 7586 32510 7588 32562
rect 7532 32498 7588 32510
rect 7868 32564 7924 32574
rect 7980 32564 8036 32732
rect 7868 32562 8036 32564
rect 7868 32510 7870 32562
rect 7922 32510 8036 32562
rect 7868 32508 8036 32510
rect 8092 32589 8148 32601
rect 8092 32537 8094 32589
rect 8146 32537 8148 32589
rect 7868 32498 7924 32508
rect 7084 31950 7086 32002
rect 7138 31950 7140 32002
rect 6412 31108 6468 31118
rect 6188 30996 6244 31006
rect 6188 30902 6244 30940
rect 6412 30994 6468 31052
rect 6412 30942 6414 30994
rect 6466 30942 6468 30994
rect 6580 31050 6636 31500
rect 6580 30998 6582 31050
rect 6634 30998 6636 31050
rect 6580 30986 6636 30998
rect 6748 30996 6804 31006
rect 6412 30930 6468 30942
rect 6748 30902 6804 30940
rect 6972 30996 7028 31006
rect 6972 30902 7028 30940
rect 7084 30548 7140 31950
rect 7756 32004 7812 32014
rect 7420 31780 7476 31790
rect 7196 31778 7476 31780
rect 7196 31726 7422 31778
rect 7474 31726 7476 31778
rect 7196 31724 7476 31726
rect 7196 30772 7252 31724
rect 7420 31714 7476 31724
rect 7756 31778 7812 31948
rect 8092 31890 8148 32537
rect 8092 31838 8094 31890
rect 8146 31838 8148 31890
rect 8092 31826 8148 31838
rect 7756 31726 7758 31778
rect 7810 31726 7812 31778
rect 7756 31714 7812 31726
rect 7980 31780 8036 31790
rect 7980 31711 7982 31724
rect 8034 31711 8036 31724
rect 7980 31686 8036 31711
rect 8204 31556 8260 33404
rect 8316 33236 8372 33246
rect 8316 32004 8372 33180
rect 8876 33236 8932 33246
rect 8876 33142 8932 33180
rect 8316 31778 8372 31948
rect 8316 31726 8318 31778
rect 8370 31726 8372 31778
rect 8316 31714 8372 31726
rect 8428 32562 8484 32574
rect 8428 32510 8430 32562
rect 8482 32510 8484 32562
rect 8428 31556 8484 32510
rect 8540 31780 8596 31790
rect 8540 31686 8596 31724
rect 8988 31724 9044 33628
rect 9100 33460 9156 33852
rect 9100 33394 9156 33404
rect 9324 33572 9380 33582
rect 9212 33346 9268 33358
rect 9212 33294 9214 33346
rect 9266 33294 9268 33346
rect 9212 32788 9268 33294
rect 9212 32722 9268 32732
rect 9324 31902 9380 33516
rect 9436 33348 9492 34636
rect 9660 34580 9716 34860
rect 10332 34916 10388 34926
rect 10556 34916 10612 35196
rect 10332 34914 10612 34916
rect 10332 34862 10334 34914
rect 10386 34862 10612 34914
rect 10332 34860 10612 34862
rect 10332 34850 10388 34860
rect 9660 34524 9828 34580
rect 9660 34356 9716 34366
rect 9660 34262 9716 34300
rect 9436 33292 9716 33348
rect 9268 31890 9380 31902
rect 9268 31838 9270 31890
rect 9322 31838 9380 31890
rect 9268 31836 9380 31838
rect 9436 32562 9492 32574
rect 9436 32510 9438 32562
rect 9490 32510 9492 32562
rect 9268 31826 9324 31836
rect 9436 31724 9492 32510
rect 8820 31666 8876 31678
rect 8988 31668 9492 31724
rect 9548 31780 9604 31790
rect 9548 31686 9604 31724
rect 8820 31614 8822 31666
rect 8874 31614 8876 31666
rect 8820 31556 8876 31614
rect 8204 31500 8372 31556
rect 8428 31500 8876 31556
rect 7812 31108 7868 31118
rect 7308 31032 7364 31044
rect 7308 30980 7310 31032
rect 7362 30980 7364 31032
rect 7812 31014 7868 31052
rect 8092 30996 8148 31006
rect 7308 30884 7364 30980
rect 7980 30994 8148 30996
rect 7980 30942 8094 30994
rect 8146 30942 8148 30994
rect 7980 30940 8148 30942
rect 7980 30884 8036 30940
rect 8092 30930 8148 30940
rect 8204 30996 8260 31006
rect 8204 30902 8260 30940
rect 7308 30828 8036 30884
rect 7196 30716 7476 30772
rect 7084 30482 7140 30492
rect 6300 30324 6356 30334
rect 6300 30230 6356 30268
rect 7420 29988 7476 30716
rect 7420 29876 7476 29932
rect 7196 29820 7476 29876
rect 7756 30660 7812 30670
rect 6076 29138 6132 29148
rect 6188 29426 6244 29438
rect 6188 29374 6190 29426
rect 6242 29374 6244 29426
rect 6076 28644 6132 28654
rect 5964 28642 6132 28644
rect 5964 28590 6078 28642
rect 6130 28590 6132 28642
rect 5964 28588 6132 28590
rect 6076 28578 6132 28588
rect 5740 28540 5796 28552
rect 5460 27970 5684 27972
rect 5460 27918 5462 27970
rect 5514 27918 5684 27970
rect 5460 27916 5684 27918
rect 6076 28420 6132 28430
rect 5460 27906 5516 27916
rect 5740 27858 5796 27870
rect 5740 27806 5742 27858
rect 5794 27806 5796 27858
rect 5292 27692 5460 27748
rect 4172 27244 4788 27300
rect 4228 27076 4284 27086
rect 4060 27074 4284 27076
rect 4060 27022 4230 27074
rect 4282 27022 4284 27074
rect 4060 27020 4284 27022
rect 4228 27010 4284 27020
rect 4508 27076 4564 27086
rect 4508 26982 4564 27020
rect 4732 27074 4788 27244
rect 5012 27298 5124 27310
rect 5012 27246 5014 27298
rect 5066 27246 5124 27298
rect 5012 27244 5124 27246
rect 5292 27524 5348 27534
rect 5012 27234 5068 27244
rect 4732 27022 4734 27074
rect 4786 27022 4788 27074
rect 4732 27010 4788 27022
rect 4844 27076 4900 27086
rect 4844 26908 4900 27020
rect 3948 26852 4116 26908
rect 4844 26852 5012 26908
rect 4060 26414 4116 26852
rect 4060 26402 4134 26414
rect 4060 26350 4080 26402
rect 4132 26350 4134 26402
rect 4060 26348 4134 26350
rect 4078 26338 4134 26348
rect 3836 26238 3838 26290
rect 3890 26238 3892 26290
rect 3836 26226 3892 26238
rect 4844 26290 4900 26302
rect 4844 26238 4846 26290
rect 4898 26238 4900 26290
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 3724 25566 3726 25618
rect 3778 25566 3780 25618
rect 4844 25674 4900 26238
rect 4956 26292 5012 26852
rect 5180 26292 5236 26302
rect 4956 26236 5124 26292
rect 5068 25956 5124 26236
rect 5180 26198 5236 26236
rect 5292 26122 5348 27468
rect 5292 26070 5294 26122
rect 5346 26070 5348 26122
rect 5292 26058 5348 26070
rect 4844 25622 4846 25674
rect 4898 25622 4900 25674
rect 4844 25610 4900 25622
rect 4956 25900 5124 25956
rect 3724 25554 3780 25566
rect 3500 25508 3556 25518
rect 3276 25506 3556 25508
rect 3164 25450 3220 25462
rect 3164 25398 3166 25450
rect 3218 25398 3220 25450
rect 3164 25396 3220 25398
rect 3164 25330 3220 25340
rect 3276 25454 3502 25506
rect 3554 25454 3556 25506
rect 4844 25506 4900 25518
rect 4104 25468 4160 25480
rect 3276 25452 3556 25454
rect 3892 25452 3948 25462
rect 2380 25116 3108 25172
rect 2268 24892 2660 24948
rect 2492 24724 2548 24734
rect 2268 24668 2492 24724
rect 2044 23714 2100 23726
rect 2044 23662 2046 23714
rect 2098 23662 2100 23714
rect 2044 23492 2100 23662
rect 2044 23426 2100 23436
rect 1484 21410 1540 21420
rect 1596 23154 1652 23166
rect 1596 23102 1598 23154
rect 1650 23102 1652 23154
rect 1596 20802 1652 23102
rect 2156 22370 2212 22382
rect 2156 22318 2158 22370
rect 2210 22318 2212 22370
rect 2156 21812 2212 22318
rect 2268 22202 2324 24668
rect 2492 24630 2548 24668
rect 2380 23940 2436 23950
rect 2604 23940 2660 24892
rect 2828 24500 2884 25116
rect 3276 25060 3332 25452
rect 3500 25442 3556 25452
rect 3836 25450 3948 25452
rect 3836 25398 3894 25450
rect 3946 25398 3948 25450
rect 3836 25386 3948 25398
rect 4104 25416 4106 25468
rect 4158 25416 4160 25468
rect 2828 24406 2884 24444
rect 3052 25004 3332 25060
rect 3388 25172 3444 25182
rect 2380 23938 2660 23940
rect 2380 23886 2382 23938
rect 2434 23900 2660 23938
rect 2434 23886 2602 23900
rect 2380 23884 2602 23886
rect 2380 23874 2436 23884
rect 2600 23848 2602 23884
rect 2654 23884 2660 23900
rect 2654 23848 2656 23884
rect 2600 23604 2656 23848
rect 2600 23538 2656 23548
rect 3052 23492 3108 25004
rect 3052 23426 3108 23436
rect 3164 24836 3220 24846
rect 3164 24722 3220 24780
rect 3164 24670 3166 24722
rect 3218 24670 3220 24722
rect 3164 23380 3220 24670
rect 3388 24722 3444 25116
rect 3388 24670 3390 24722
rect 3442 24670 3444 24722
rect 3388 24106 3444 24670
rect 3556 24724 3612 24734
rect 3556 24630 3612 24668
rect 3388 24054 3390 24106
rect 3442 24054 3444 24106
rect 3276 23938 3332 23950
rect 3276 23886 3278 23938
rect 3330 23886 3332 23938
rect 3276 23380 3332 23886
rect 3388 23828 3444 24054
rect 3836 23828 3892 25386
rect 4104 24948 4160 25416
rect 4844 25454 4846 25506
rect 4898 25454 4900 25506
rect 4844 25172 4900 25454
rect 4844 25106 4900 25116
rect 3948 24892 4160 24948
rect 3948 24500 4004 24892
rect 4844 24778 4900 24790
rect 4060 24724 4116 24734
rect 4844 24726 4846 24778
rect 4898 24726 4900 24778
rect 4060 24722 4228 24724
rect 4060 24670 4062 24722
rect 4114 24670 4228 24722
rect 4060 24668 4228 24670
rect 4060 24658 4116 24668
rect 3948 23910 4004 24444
rect 3948 23858 3950 23910
rect 4002 23858 4004 23910
rect 3948 23846 4004 23858
rect 4172 23940 4228 24668
rect 4302 24612 4358 24622
rect 4302 24518 4358 24556
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4396 24052 4452 24062
rect 4396 23958 4452 23996
rect 3388 23772 3780 23828
rect 3276 23324 3556 23380
rect 3164 23314 3220 23324
rect 2268 22150 2270 22202
rect 2322 22150 2324 22202
rect 2268 22138 2324 22150
rect 2380 23042 2436 23054
rect 2380 22990 2382 23042
rect 2434 22990 2436 23042
rect 2156 21746 2212 21756
rect 2268 21812 2324 21822
rect 2380 21812 2436 22990
rect 3164 22820 3220 22830
rect 2828 22484 2884 22494
rect 2828 22370 2884 22428
rect 2828 22318 2830 22370
rect 2882 22318 2884 22370
rect 2828 22306 2884 22318
rect 3164 22370 3220 22764
rect 3164 22318 3166 22370
rect 3218 22318 3220 22370
rect 3332 22820 3388 22830
rect 3332 22426 3388 22764
rect 3332 22374 3334 22426
rect 3386 22374 3388 22426
rect 3500 22484 3556 23324
rect 3500 22418 3556 22428
rect 3332 22362 3388 22374
rect 3612 22370 3668 22382
rect 3164 22306 3220 22318
rect 3612 22318 3614 22370
rect 3666 22318 3668 22370
rect 3500 22258 3556 22270
rect 3500 22206 3502 22258
rect 3554 22206 3556 22258
rect 2268 21810 2436 21812
rect 2268 21758 2270 21810
rect 2322 21758 2436 21810
rect 2268 21756 2436 21758
rect 3276 21812 3332 21822
rect 2268 21746 2324 21756
rect 2604 21588 2660 21598
rect 2604 21494 2660 21532
rect 3276 21586 3332 21756
rect 3500 21812 3556 22206
rect 3612 21924 3668 22318
rect 3724 22260 3780 23772
rect 3836 23762 3892 23772
rect 3892 23156 3948 23166
rect 3892 22594 3948 23100
rect 3892 22542 3894 22594
rect 3946 22542 3948 22594
rect 3892 22530 3948 22542
rect 3724 22194 3780 22204
rect 3612 21868 3892 21924
rect 3500 21746 3556 21756
rect 3612 21700 3668 21710
rect 3612 21606 3668 21644
rect 3276 21534 3278 21586
rect 3330 21534 3332 21586
rect 3276 21522 3332 21534
rect 2380 20804 2436 20814
rect 1596 20750 1598 20802
rect 1650 20750 1652 20802
rect 1596 20020 1652 20750
rect 1820 20802 2436 20804
rect 1820 20750 2382 20802
rect 2434 20750 2436 20802
rect 1820 20748 2436 20750
rect 1820 20242 1876 20748
rect 2380 20738 2436 20748
rect 1820 20190 1822 20242
rect 1874 20190 1876 20242
rect 1820 20178 1876 20190
rect 3836 20244 3892 21868
rect 4056 21812 4112 21822
rect 4056 21626 4112 21756
rect 4172 21700 4228 23884
rect 4564 23882 4620 23894
rect 4564 23830 4566 23882
rect 4618 23830 4620 23882
rect 4564 23828 4620 23830
rect 4564 23762 4620 23772
rect 4284 23604 4340 23614
rect 4284 23268 4340 23548
rect 4284 23266 4676 23268
rect 4284 23214 4286 23266
rect 4338 23214 4676 23266
rect 4284 23212 4676 23214
rect 4284 23202 4340 23212
rect 4620 23154 4676 23212
rect 4620 23102 4622 23154
rect 4674 23102 4676 23154
rect 4620 23090 4676 23102
rect 4844 23156 4900 24726
rect 4844 23090 4900 23100
rect 4788 22932 4844 22970
rect 4788 22866 4844 22876
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4620 22484 4676 22494
rect 4508 22314 4564 22326
rect 4508 22262 4510 22314
rect 4562 22262 4564 22314
rect 4508 22260 4564 22262
rect 4508 22194 4564 22204
rect 4172 21634 4228 21644
rect 4508 22036 4564 22046
rect 4056 21624 4116 21626
rect 4056 21572 4058 21624
rect 4110 21572 4116 21624
rect 4056 21560 4116 21572
rect 4060 20916 4116 21560
rect 4508 21418 4564 21980
rect 4620 21924 4676 22428
rect 4956 22482 5012 25900
rect 5404 24834 5460 27692
rect 5740 27524 5796 27806
rect 5964 27860 6020 27870
rect 5964 27766 6020 27804
rect 5740 27458 5796 27468
rect 5628 27076 5684 27086
rect 5628 26982 5684 27020
rect 6076 26906 6132 28364
rect 6188 27972 6244 29374
rect 6636 29428 6692 29438
rect 6636 29334 6692 29372
rect 6860 29426 6916 29438
rect 6860 29374 6862 29426
rect 6914 29374 6916 29426
rect 6524 29258 6580 29270
rect 6524 29206 6526 29258
rect 6578 29206 6580 29258
rect 6524 28980 6580 29206
rect 6468 28924 6580 28980
rect 6300 28756 6356 28766
rect 6300 28662 6356 28700
rect 6468 28698 6524 28924
rect 6468 28646 6470 28698
rect 6522 28646 6524 28698
rect 6468 28634 6524 28646
rect 6188 27906 6244 27916
rect 6412 28420 6468 28430
rect 6244 27634 6300 27646
rect 6244 27582 6246 27634
rect 6298 27582 6300 27634
rect 6244 27300 6300 27582
rect 6244 27234 6300 27244
rect 5852 26852 5908 26862
rect 6076 26854 6078 26906
rect 6130 26854 6132 26906
rect 6076 26842 6132 26854
rect 6188 27074 6244 27086
rect 6188 27022 6190 27074
rect 6242 27022 6244 27074
rect 5740 26290 5796 26302
rect 5740 26238 5742 26290
rect 5794 26238 5796 26290
rect 5404 24782 5406 24834
rect 5458 24782 5460 24834
rect 5404 24770 5460 24782
rect 5516 25506 5572 25518
rect 5516 25454 5518 25506
rect 5570 25454 5572 25506
rect 5516 24836 5572 25454
rect 5516 24388 5572 24780
rect 5516 24322 5572 24332
rect 5628 24722 5684 24734
rect 5628 24670 5630 24722
rect 5682 24670 5684 24722
rect 5628 24052 5684 24670
rect 5628 23986 5684 23996
rect 5292 23828 5348 23838
rect 5180 23380 5236 23390
rect 5180 22484 5236 23324
rect 4956 22430 4958 22482
rect 5010 22430 5012 22482
rect 4956 22418 5012 22430
rect 5124 22428 5236 22484
rect 5124 22426 5180 22428
rect 4732 22372 4788 22382
rect 5124 22374 5126 22426
rect 5178 22374 5180 22426
rect 5124 22362 5180 22374
rect 4732 22036 4788 22316
rect 5292 22148 5348 23772
rect 5740 23716 5796 26238
rect 5852 25730 5908 26796
rect 6188 26404 6244 27022
rect 5852 25678 5854 25730
rect 5906 25678 5908 25730
rect 5852 25666 5908 25678
rect 5964 26348 6244 26404
rect 5964 26305 6020 26348
rect 5964 26253 5966 26305
rect 6018 26253 6020 26305
rect 5964 25732 6020 26253
rect 5964 25666 6020 25676
rect 6076 26178 6132 26190
rect 6076 26126 6078 26178
rect 6130 26126 6132 26178
rect 6076 25508 6132 26126
rect 6076 25442 6132 25452
rect 6300 25506 6356 25518
rect 6300 25454 6302 25506
rect 6354 25454 6356 25506
rect 6300 25396 6356 25454
rect 6300 25330 6356 25340
rect 6188 24724 6244 24734
rect 5740 23660 5908 23716
rect 5740 23492 5796 23502
rect 5628 23268 5684 23278
rect 5516 23156 5572 23166
rect 5404 23154 5572 23156
rect 5404 23102 5518 23154
rect 5570 23102 5572 23154
rect 5404 23100 5572 23102
rect 5404 22372 5460 23100
rect 5516 23090 5572 23100
rect 5404 22306 5460 22316
rect 5516 22932 5572 22942
rect 5516 22370 5572 22876
rect 5516 22318 5518 22370
rect 5570 22318 5572 22370
rect 5516 22306 5572 22318
rect 4732 21970 4788 21980
rect 5068 22092 5348 22148
rect 4620 21588 4676 21868
rect 4732 21588 4788 21598
rect 4620 21586 4788 21588
rect 4620 21534 4734 21586
rect 4786 21534 4788 21586
rect 4620 21532 4788 21534
rect 4508 21366 4510 21418
rect 4562 21366 4564 21418
rect 4508 21354 4564 21366
rect 4732 21364 4788 21532
rect 4732 21308 4900 21364
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4844 21026 4900 21308
rect 4844 20974 4846 21026
rect 4898 20974 4900 21026
rect 4844 20962 4900 20974
rect 4284 20916 4340 20926
rect 4060 20914 4340 20916
rect 4060 20862 4286 20914
rect 4338 20862 4340 20914
rect 4060 20860 4340 20862
rect 4284 20850 4340 20860
rect 3836 20188 4340 20244
rect 1596 19954 1652 19964
rect 2156 20018 2212 20030
rect 2156 19966 2158 20018
rect 2210 19966 2212 20018
rect 2156 19796 2212 19966
rect 2156 19730 2212 19740
rect 2268 20020 2324 20030
rect 2268 18452 2324 19964
rect 3052 19908 3108 19918
rect 3052 19814 3108 19852
rect 4284 19234 4340 20188
rect 4956 19906 5012 19918
rect 4956 19854 4958 19906
rect 5010 19854 5012 19906
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4284 19182 4286 19234
rect 4338 19182 4340 19234
rect 4004 19010 4060 19022
rect 4004 18958 4006 19010
rect 4058 18958 4060 19010
rect 4004 18788 4060 18958
rect 4284 19012 4340 19182
rect 4956 19236 5012 19854
rect 5068 19402 5124 22092
rect 5404 21924 5460 21934
rect 5404 21586 5460 21868
rect 5404 21534 5406 21586
rect 5458 21534 5460 21586
rect 5404 21522 5460 21534
rect 5628 21474 5684 23212
rect 5740 23210 5796 23436
rect 5740 23158 5742 23210
rect 5794 23158 5796 23210
rect 5852 23268 5908 23660
rect 6076 23380 6132 23390
rect 5852 23202 5908 23212
rect 5964 23322 6020 23334
rect 5964 23270 5966 23322
rect 6018 23270 6020 23322
rect 5740 21924 5796 23158
rect 5964 23156 6020 23270
rect 5964 23090 6020 23100
rect 6076 23154 6132 23324
rect 6076 23102 6078 23154
rect 6130 23102 6132 23154
rect 6076 23090 6132 23102
rect 6188 22932 6244 24668
rect 5852 22876 6244 22932
rect 5852 22594 5908 22876
rect 6412 22596 6468 28364
rect 6860 28420 6916 29374
rect 7196 28644 7252 29820
rect 7476 29652 7532 29662
rect 7476 29558 7532 29596
rect 7756 29316 7812 30604
rect 7868 29540 7924 29550
rect 7980 29540 8036 30828
rect 8316 30660 8372 31500
rect 8428 30994 8484 31006
rect 8428 30942 8430 30994
rect 8482 30942 8484 30994
rect 8428 30884 8484 30942
rect 8540 30996 8596 31500
rect 8540 30930 8596 30940
rect 8428 30818 8484 30828
rect 8316 30594 8372 30604
rect 8764 30770 8820 30782
rect 8764 30718 8766 30770
rect 8818 30718 8820 30770
rect 8764 30324 8820 30718
rect 9212 30436 9268 31668
rect 9660 31444 9716 33292
rect 9772 32786 9828 34524
rect 10332 34168 10388 34180
rect 9996 34132 10052 34142
rect 10332 34116 10334 34168
rect 10386 34116 10388 34168
rect 9996 34038 10052 34076
rect 10220 34074 10276 34086
rect 10220 34022 10222 34074
rect 10274 34022 10276 34074
rect 10220 33796 10276 34022
rect 10108 33740 10276 33796
rect 9996 33460 10052 33470
rect 9996 33366 10052 33404
rect 9772 32734 9774 32786
rect 9826 32734 9828 32786
rect 9772 32722 9828 32734
rect 10108 31892 10164 33740
rect 10332 33684 10388 34116
rect 10668 33796 10724 35644
rect 11004 35634 11060 35644
rect 11116 35252 11172 35262
rect 10668 33730 10724 33740
rect 10780 34914 10836 34926
rect 11004 34916 11060 34926
rect 10780 34862 10782 34914
rect 10834 34862 10836 34914
rect 9996 31836 10164 31892
rect 10220 33628 10388 33684
rect 10780 33684 10836 34862
rect 10892 34914 11060 34916
rect 10892 34862 11006 34914
rect 11058 34862 11060 34914
rect 10892 34860 11060 34862
rect 10892 34242 10948 34860
rect 11004 34850 11060 34860
rect 11116 34692 11172 35196
rect 11284 34804 11340 34814
rect 11284 34710 11340 34748
rect 10892 34190 10894 34242
rect 10946 34190 10948 34242
rect 10892 34178 10948 34190
rect 11060 34636 11172 34692
rect 11060 34468 11116 34636
rect 11060 34074 11116 34412
rect 11060 34022 11062 34074
rect 11114 34022 11116 34074
rect 11060 33908 11116 34022
rect 11228 34580 11284 34590
rect 11228 33908 11284 34524
rect 11340 34132 11396 34142
rect 11676 34132 11732 35980
rect 12124 35924 12180 36652
rect 12684 36594 12740 37100
rect 12684 36542 12686 36594
rect 12738 36542 12740 36594
rect 12684 36530 12740 36542
rect 12012 35868 12180 35924
rect 12236 36482 12292 36494
rect 12572 36484 12628 36494
rect 12236 36430 12238 36482
rect 12290 36430 12292 36482
rect 11880 35698 11936 35710
rect 11880 35646 11882 35698
rect 11934 35646 11936 35698
rect 11880 35140 11936 35646
rect 12012 35252 12068 35868
rect 12124 35700 12180 35710
rect 12124 35606 12180 35644
rect 12236 35476 12292 36430
rect 12460 36482 12628 36484
rect 12460 36430 12574 36482
rect 12626 36430 12628 36482
rect 12460 36428 12628 36430
rect 12460 35812 12516 36428
rect 12572 36418 12628 36428
rect 13020 36036 13076 41580
rect 13580 41524 13636 41534
rect 13580 41156 13636 41468
rect 13412 41130 13468 41142
rect 13412 41078 13414 41130
rect 13466 41078 13468 41130
rect 13580 41104 13582 41156
rect 13634 41104 13636 41156
rect 13580 41092 13636 41104
rect 13916 41130 13972 41906
rect 13132 40740 13188 40750
rect 13132 40402 13188 40684
rect 13412 40516 13468 41078
rect 13916 41078 13918 41130
rect 13970 41078 13972 41130
rect 13916 41076 13972 41078
rect 13916 41010 13972 41020
rect 14140 41746 14196 41758
rect 14140 41694 14142 41746
rect 14194 41694 14196 41746
rect 14140 40740 14196 41694
rect 14140 40674 14196 40684
rect 13412 40460 13636 40516
rect 13132 40350 13134 40402
rect 13186 40350 13188 40402
rect 13132 37380 13188 40350
rect 13580 40404 13636 40460
rect 13580 40338 13636 40348
rect 13244 40234 13300 40246
rect 13244 40182 13246 40234
rect 13298 40182 13300 40234
rect 13244 39508 13300 40182
rect 14252 39956 14308 42364
rect 14364 41412 14420 41422
rect 14476 41412 14532 43484
rect 14756 43482 14812 43494
rect 14364 41410 14532 41412
rect 14364 41358 14366 41410
rect 14418 41358 14532 41410
rect 14364 41356 14532 41358
rect 14588 43428 14644 43438
rect 14364 41346 14420 41356
rect 14588 40964 14644 43372
rect 14756 43430 14758 43482
rect 14810 43430 14812 43482
rect 14756 43092 14812 43430
rect 14756 43026 14812 43036
rect 14924 42868 14980 43596
rect 15036 43540 15092 43578
rect 15036 43474 15092 43484
rect 14924 42802 14980 42812
rect 15036 43092 15092 43102
rect 15036 42756 15092 43036
rect 14700 42698 14756 42710
rect 14700 42646 14702 42698
rect 14754 42646 14756 42698
rect 15036 42662 15092 42700
rect 14700 42644 14756 42646
rect 14700 42578 14756 42588
rect 15148 42196 15204 44604
rect 15596 43706 15652 44828
rect 16604 44884 16660 44894
rect 16604 44790 16660 44828
rect 16828 44324 16884 44334
rect 17500 44324 17556 45052
rect 17668 44994 17724 45006
rect 17668 44942 17670 44994
rect 17722 44942 17724 44994
rect 17668 44772 17724 44942
rect 17668 44706 17724 44716
rect 17612 44324 17668 44334
rect 17724 44324 17780 44334
rect 16828 44322 17108 44324
rect 16828 44270 16830 44322
rect 16882 44270 17108 44322
rect 16828 44268 17108 44270
rect 16828 44258 16884 44268
rect 15596 43654 15598 43706
rect 15650 43654 15652 43706
rect 15596 43642 15652 43654
rect 15932 43652 15988 43662
rect 15932 43594 15988 43596
rect 15708 43540 15764 43550
rect 15260 43538 15764 43540
rect 15260 43486 15710 43538
rect 15762 43486 15764 43538
rect 15932 43542 15934 43594
rect 15986 43542 15988 43594
rect 15932 43530 15988 43542
rect 16380 43540 16436 43550
rect 15260 43484 15764 43486
rect 15260 42866 15316 43484
rect 15708 43474 15764 43484
rect 16380 43446 16436 43484
rect 16716 43540 16772 43550
rect 15260 42814 15262 42866
rect 15314 42814 15316 42866
rect 15260 42802 15316 42814
rect 16156 42868 16212 42878
rect 16156 42754 16212 42812
rect 15428 42698 15484 42710
rect 15428 42646 15430 42698
rect 15482 42646 15484 42698
rect 15428 42644 15484 42646
rect 15428 42578 15484 42588
rect 15932 42698 15988 42710
rect 15932 42646 15934 42698
rect 15986 42646 15988 42698
rect 16156 42702 16158 42754
rect 16210 42702 16212 42754
rect 16156 42690 16212 42702
rect 16380 42756 16436 42766
rect 16380 42662 16436 42700
rect 16548 42698 16604 42710
rect 15932 42644 15988 42646
rect 15932 42578 15988 42588
rect 16268 42644 16324 42654
rect 15148 42140 15316 42196
rect 14868 41972 14924 41982
rect 14868 41878 14924 41916
rect 15148 41970 15204 41982
rect 15148 41918 15150 41970
rect 15202 41918 15204 41970
rect 15148 41636 15204 41918
rect 15260 41748 15316 42140
rect 15894 42007 15950 42019
rect 15260 41682 15316 41692
rect 15372 41970 15428 41982
rect 15372 41918 15374 41970
rect 15426 41918 15428 41970
rect 15148 41570 15204 41580
rect 15372 41636 15428 41918
rect 15372 41570 15428 41580
rect 15596 41970 15652 41982
rect 15596 41918 15598 41970
rect 15650 41918 15652 41970
rect 14924 41188 14980 41198
rect 15596 41188 15652 41918
rect 15708 41970 15764 41982
rect 15708 41918 15710 41970
rect 15762 41918 15764 41970
rect 15708 41524 15764 41918
rect 15894 41972 15896 42007
rect 15948 41972 15950 42007
rect 15894 41748 15950 41916
rect 16268 41858 16324 42588
rect 16548 42646 16550 42698
rect 16602 42646 16604 42698
rect 16548 42196 16604 42646
rect 16548 42140 16660 42196
rect 16268 41806 16270 41858
rect 16322 41806 16324 41858
rect 16268 41794 16324 41806
rect 16492 41972 16548 41982
rect 15894 41692 16212 41748
rect 16044 41524 16100 41534
rect 15708 41468 15856 41524
rect 14924 41186 15092 41188
rect 14924 41134 14926 41186
rect 14978 41134 15092 41186
rect 14924 41132 15092 41134
rect 14924 41122 14980 41132
rect 14588 40908 14980 40964
rect 14456 40740 14512 40750
rect 14456 40458 14512 40684
rect 14456 40406 14458 40458
rect 14510 40406 14512 40458
rect 14700 40740 14756 40750
rect 14700 40514 14756 40684
rect 14700 40462 14702 40514
rect 14754 40462 14756 40514
rect 14700 40450 14756 40462
rect 14456 40394 14512 40406
rect 14252 39890 14308 39900
rect 13916 39732 13972 39742
rect 13524 39620 13580 39630
rect 13804 39620 13860 39630
rect 13524 39526 13580 39564
rect 13692 39618 13860 39620
rect 13692 39566 13806 39618
rect 13858 39566 13860 39618
rect 13692 39564 13860 39566
rect 13244 38836 13300 39452
rect 13468 38836 13524 38846
rect 13244 38834 13524 38836
rect 13244 38782 13470 38834
rect 13522 38782 13524 38834
rect 13244 38780 13524 38782
rect 13468 38770 13524 38780
rect 13580 38836 13636 38846
rect 13580 38666 13636 38780
rect 13580 38614 13582 38666
rect 13634 38614 13636 38666
rect 13580 38602 13636 38614
rect 13132 37314 13188 37324
rect 13356 38164 13412 38174
rect 13356 37378 13412 38108
rect 13356 37326 13358 37378
rect 13410 37326 13412 37378
rect 13356 37314 13412 37326
rect 13692 37940 13748 39564
rect 13804 39554 13860 39564
rect 13916 39618 13972 39676
rect 13916 39566 13918 39618
rect 13970 39566 13972 39618
rect 13916 39284 13972 39566
rect 13916 39218 13972 39228
rect 14252 39618 14308 39630
rect 14252 39566 14254 39618
rect 14306 39566 14308 39618
rect 14252 38836 14308 39566
rect 14364 39620 14420 39630
rect 14364 39172 14420 39564
rect 14924 39508 14980 40908
rect 15036 40740 15092 41132
rect 15036 40684 15372 40740
rect 15316 40626 15372 40684
rect 15316 40574 15318 40626
rect 15370 40574 15372 40626
rect 15316 40562 15372 40574
rect 15484 40404 15540 40414
rect 15596 40404 15652 41132
rect 15800 41130 15856 41468
rect 16044 41412 16100 41468
rect 15800 41078 15802 41130
rect 15854 41078 15856 41130
rect 15800 41076 15856 41078
rect 15800 40852 15856 41020
rect 15484 40402 15652 40404
rect 15484 40350 15486 40402
rect 15538 40350 15652 40402
rect 15484 40348 15652 40350
rect 15708 40796 15856 40852
rect 15932 41410 16100 41412
rect 15932 41358 16046 41410
rect 16098 41358 16100 41410
rect 15932 41356 16100 41358
rect 15484 40338 15540 40348
rect 14924 39442 14980 39452
rect 15128 39562 15184 39574
rect 15128 39510 15130 39562
rect 15182 39510 15184 39562
rect 15128 39172 15184 39510
rect 15372 39506 15428 39518
rect 15372 39454 15374 39506
rect 15426 39454 15428 39506
rect 15372 39396 15428 39454
rect 15372 39330 15428 39340
rect 15708 39284 15764 40796
rect 15820 40628 15876 40638
rect 15820 39396 15876 40572
rect 15932 39618 15988 41356
rect 16044 41346 16100 41356
rect 16044 40404 16100 40414
rect 16156 40404 16212 41692
rect 16492 40740 16548 41916
rect 16604 41860 16660 42140
rect 16716 42084 16772 43484
rect 16884 43540 16940 43550
rect 16884 43446 16940 43484
rect 16716 42018 16772 42028
rect 16884 42642 16940 42654
rect 16884 42590 16886 42642
rect 16938 42590 16940 42642
rect 16884 42084 16940 42590
rect 16884 42018 16940 42028
rect 16884 41860 16940 41870
rect 16604 41858 16940 41860
rect 16604 41806 16886 41858
rect 16938 41806 16940 41858
rect 16604 41804 16940 41806
rect 16604 40852 16660 41804
rect 16884 41794 16940 41804
rect 17052 41636 17108 44268
rect 17500 44322 17780 44324
rect 17500 44270 17614 44322
rect 17666 44270 17726 44322
rect 17778 44270 17780 44322
rect 17500 44268 17780 44270
rect 17500 43204 17556 44268
rect 17612 44258 17668 44268
rect 17724 44258 17780 44268
rect 17836 43764 17892 46284
rect 19180 46116 19236 46126
rect 19292 46116 19348 49200
rect 19180 46114 19348 46116
rect 19180 46062 19182 46114
rect 19234 46062 19348 46114
rect 19180 46060 19348 46062
rect 19180 46050 19236 46060
rect 20076 45892 20132 45902
rect 20748 45892 20804 45902
rect 20076 45810 20078 45836
rect 20130 45810 20132 45836
rect 20076 45798 20132 45810
rect 20636 45890 20804 45892
rect 20636 45838 20750 45890
rect 20802 45838 20804 45890
rect 20636 45836 20804 45838
rect 18508 45668 18564 45678
rect 18060 44996 18116 45006
rect 18060 44902 18116 44940
rect 17836 43698 17892 43708
rect 17948 44660 18004 44670
rect 17668 43652 17724 43662
rect 17668 43558 17724 43596
rect 17948 43565 18004 44604
rect 18508 44434 18564 45612
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 19964 44996 20020 45006
rect 19964 44902 20020 44940
rect 18508 44382 18510 44434
rect 18562 44382 18564 44434
rect 18508 44370 18564 44382
rect 20412 44212 20468 44222
rect 20636 44212 20692 45836
rect 20748 45826 20804 45836
rect 20748 45108 20804 45118
rect 20748 45014 20804 45052
rect 20860 44548 20916 49200
rect 22428 46116 22484 49200
rect 22540 46116 22596 46126
rect 22428 46114 22596 46116
rect 22428 46062 22542 46114
rect 22594 46062 22596 46114
rect 22428 46060 22596 46062
rect 22540 46050 22596 46060
rect 21532 45862 21588 45874
rect 21532 45810 21534 45862
rect 21586 45810 21588 45862
rect 21084 45780 21140 45790
rect 21532 45780 21588 45810
rect 21084 45778 21588 45780
rect 21084 45726 21086 45778
rect 21138 45726 21588 45778
rect 21084 45724 21588 45726
rect 21084 45714 21140 45724
rect 20860 44482 20916 44492
rect 20972 45106 21028 45118
rect 20972 45054 20974 45106
rect 21026 45054 21028 45106
rect 20188 44210 20468 44212
rect 20188 44158 20414 44210
rect 20466 44158 20468 44210
rect 20188 44156 20468 44158
rect 19404 44100 19460 44110
rect 19292 43764 19348 43774
rect 19292 43670 19348 43708
rect 17948 43513 17950 43565
rect 18002 43513 18004 43565
rect 17948 43501 18004 43513
rect 17500 43148 17668 43204
rect 17500 42868 17556 42878
rect 17164 42756 17220 42766
rect 17164 42662 17220 42700
rect 17388 42756 17444 42766
rect 17388 42662 17444 42700
rect 17500 42754 17556 42812
rect 17500 42702 17502 42754
rect 17554 42702 17556 42754
rect 17500 42690 17556 42702
rect 16828 41580 17108 41636
rect 17164 42084 17220 42094
rect 16716 41188 16772 41198
rect 16716 41094 16772 41132
rect 16604 40796 16772 40852
rect 16492 40684 16660 40740
rect 16492 40570 16548 40582
rect 16492 40518 16494 40570
rect 16546 40518 16548 40570
rect 16044 40402 16212 40404
rect 16044 40350 16046 40402
rect 16098 40350 16212 40402
rect 16044 40348 16212 40350
rect 16268 40441 16324 40453
rect 16268 40389 16270 40441
rect 16322 40389 16324 40441
rect 16044 40338 16100 40348
rect 16268 39730 16324 40389
rect 16492 40404 16548 40518
rect 16492 40338 16548 40348
rect 16604 40516 16660 40684
rect 16604 40402 16660 40460
rect 16604 40350 16606 40402
rect 16658 40350 16660 40402
rect 16268 39678 16270 39730
rect 16322 39678 16324 39730
rect 16268 39666 16324 39678
rect 15932 39566 15934 39618
rect 15986 39566 15988 39618
rect 15932 39554 15988 39566
rect 16100 39562 16156 39574
rect 16100 39510 16102 39562
rect 16154 39510 16156 39562
rect 16100 39508 16156 39510
rect 16044 39452 16156 39508
rect 16044 39396 16100 39452
rect 15820 39340 16100 39396
rect 15708 39228 16212 39284
rect 14364 39116 14532 39172
rect 14252 38770 14308 38780
rect 14364 38872 14420 38884
rect 14364 38820 14366 38872
rect 14418 38820 14420 38872
rect 13804 38724 13860 38734
rect 13804 38174 13860 38668
rect 14364 38612 14420 38820
rect 13804 38164 13916 38174
rect 14364 38164 14420 38556
rect 13804 38162 14196 38164
rect 13804 38110 13862 38162
rect 13914 38110 14196 38162
rect 13804 38108 14196 38110
rect 13860 38098 13916 38108
rect 13580 37266 13636 37278
rect 13188 37210 13244 37222
rect 13188 37158 13190 37210
rect 13242 37158 13244 37210
rect 13188 37156 13244 37158
rect 13188 37090 13244 37100
rect 13580 37214 13582 37266
rect 13634 37214 13636 37266
rect 13580 36650 13636 37214
rect 13692 37156 13748 37884
rect 13804 37294 13860 37306
rect 13804 37268 13806 37294
rect 13858 37268 13860 37294
rect 13804 37202 13860 37212
rect 13692 36708 13748 37100
rect 14140 37044 14196 38108
rect 14364 38098 14420 38108
rect 14476 38836 14532 39116
rect 14924 39116 15184 39172
rect 15596 39172 15652 39182
rect 14924 38946 14980 39116
rect 15596 39058 15652 39116
rect 15596 39006 15598 39058
rect 15650 39006 15652 39058
rect 15596 38994 15652 39006
rect 14924 38894 14926 38946
rect 14978 38894 14980 38946
rect 14924 38882 14980 38894
rect 14700 38836 14756 38846
rect 14476 38834 14756 38836
rect 14476 38782 14702 38834
rect 14754 38782 14756 38834
rect 15932 38836 15988 38846
rect 14476 38780 14756 38782
rect 14252 38052 14308 38062
rect 14252 37268 14308 37996
rect 14476 38050 14532 38780
rect 14700 38770 14756 38780
rect 15092 38778 15148 38790
rect 15092 38726 15094 38778
rect 15146 38726 15148 38778
rect 15932 38742 15988 38780
rect 15092 38668 15148 38726
rect 14700 38612 15148 38668
rect 15800 38612 15856 38622
rect 14476 37998 14478 38050
rect 14530 37998 14532 38050
rect 14476 37986 14532 37998
rect 14588 38218 14644 38230
rect 14588 38166 14590 38218
rect 14642 38166 14644 38218
rect 14588 38052 14644 38166
rect 14588 37986 14644 37996
rect 14700 37502 14756 38612
rect 14924 38052 14980 38062
rect 14924 37958 14980 37996
rect 15800 38050 15856 38556
rect 15800 37998 15802 38050
rect 15854 37998 15856 38050
rect 15800 37986 15856 37998
rect 16044 38052 16100 38062
rect 16044 37958 16100 37996
rect 14644 37490 14756 37502
rect 14644 37438 14646 37490
rect 14698 37438 14756 37490
rect 14644 37436 14756 37438
rect 14644 37426 14700 37436
rect 14476 37268 14532 37278
rect 14252 37266 14532 37268
rect 14252 37214 14478 37266
rect 14530 37214 14532 37266
rect 14252 37212 14532 37214
rect 14476 37202 14532 37212
rect 15204 37156 15260 37166
rect 15204 37062 15260 37100
rect 15988 37156 16044 37166
rect 15988 37154 16100 37156
rect 15988 37102 15990 37154
rect 16042 37102 16100 37154
rect 15988 37090 16100 37102
rect 14028 36988 14476 37044
rect 13692 36652 13972 36708
rect 13580 36598 13582 36650
rect 13634 36598 13636 36650
rect 13580 36586 13636 36598
rect 13580 36482 13636 36494
rect 13580 36430 13582 36482
rect 13634 36430 13636 36482
rect 13020 35980 13300 36036
rect 12236 35410 12292 35420
rect 12348 35756 12516 35812
rect 12348 35364 12404 35756
rect 12572 35700 12628 35738
rect 12572 35634 12628 35644
rect 12348 35308 12572 35364
rect 12012 35196 12292 35252
rect 11880 35084 12180 35140
rect 11788 35028 11844 35038
rect 11788 34804 11844 34972
rect 12012 34858 12068 34870
rect 12012 34806 12014 34858
rect 12066 34806 12068 34858
rect 12012 34804 12068 34806
rect 11788 34748 12068 34804
rect 11340 34130 11732 34132
rect 11340 34078 11342 34130
rect 11394 34078 11732 34130
rect 11340 34076 11732 34078
rect 11340 34066 11396 34076
rect 11228 33852 11396 33908
rect 11060 33842 11116 33852
rect 9772 31778 9828 31790
rect 9772 31726 9774 31778
rect 9826 31726 9828 31778
rect 9772 31668 9828 31726
rect 9772 31602 9828 31612
rect 9996 31668 10052 31836
rect 10220 31780 10276 33628
rect 10780 33618 10836 33628
rect 11228 33236 11284 33246
rect 11004 32788 11060 32798
rect 10780 32730 10836 32742
rect 10780 32678 10782 32730
rect 10834 32678 10836 32730
rect 10332 32564 10388 32574
rect 10332 32562 10724 32564
rect 10332 32510 10334 32562
rect 10386 32510 10724 32562
rect 10332 32508 10724 32510
rect 10332 32498 10388 32508
rect 10500 31724 10556 31734
rect 10220 31722 10556 31724
rect 9996 31602 10052 31612
rect 10108 31666 10164 31678
rect 10220 31670 10502 31722
rect 10554 31670 10556 31722
rect 10220 31668 10556 31670
rect 10108 31614 10110 31666
rect 10162 31614 10164 31666
rect 10108 31444 10164 31614
rect 9660 31388 9828 31444
rect 9492 31050 9548 31062
rect 9492 30998 9494 31050
rect 9546 30998 9548 31050
rect 9492 30548 9548 30998
rect 9212 30370 9268 30380
rect 9324 30492 9548 30548
rect 9660 31024 9716 31036
rect 9660 30972 9662 31024
rect 9714 30972 9716 31024
rect 8764 30258 8820 30268
rect 9324 30324 9380 30492
rect 9660 30324 9716 30972
rect 9324 30258 9380 30268
rect 9436 30268 9716 30324
rect 8204 30212 8260 30222
rect 8260 30156 8372 30212
rect 8204 30118 8260 30156
rect 7868 29538 8036 29540
rect 7868 29486 7870 29538
rect 7922 29486 8036 29538
rect 7868 29484 8036 29486
rect 8092 30100 8148 30110
rect 8092 29494 8148 30044
rect 7868 29474 7924 29484
rect 8092 29482 8167 29494
rect 8092 29430 8113 29482
rect 8165 29430 8167 29482
rect 8092 29428 8167 29430
rect 8111 29418 8167 29428
rect 8316 29428 8372 30156
rect 8988 30210 9044 30222
rect 8988 30158 8990 30210
rect 9042 30158 9044 30210
rect 8820 30100 8876 30110
rect 8820 29986 8876 30044
rect 8820 29934 8822 29986
rect 8874 29934 8876 29986
rect 8820 29922 8876 29934
rect 8988 29652 9044 30158
rect 9156 30154 9212 30166
rect 9156 30102 9158 30154
rect 9210 30102 9212 30154
rect 9156 30100 9212 30102
rect 9156 30034 9212 30044
rect 9324 30154 9380 30166
rect 9324 30102 9326 30154
rect 9378 30102 9380 30154
rect 9324 30100 9380 30102
rect 9324 30034 9380 30044
rect 9436 29652 9492 30268
rect 8988 29596 9492 29652
rect 9548 30154 9604 30166
rect 9548 30102 9550 30154
rect 9602 30102 9604 30154
rect 8316 29362 8372 29372
rect 8988 29428 9044 29466
rect 8988 29362 9044 29372
rect 7756 29260 8148 29316
rect 7420 28644 7476 28654
rect 7196 28588 7364 28644
rect 6860 28354 6916 28364
rect 7140 28420 7196 28430
rect 7140 28326 7196 28364
rect 6972 28084 7028 28094
rect 6804 27972 6860 27982
rect 6804 27914 6860 27916
rect 6524 27858 6580 27870
rect 6524 27806 6526 27858
rect 6578 27806 6580 27858
rect 6524 27524 6580 27806
rect 6524 27458 6580 27468
rect 6636 27860 6692 27870
rect 6804 27862 6806 27914
rect 6858 27862 6860 27914
rect 6804 27850 6860 27862
rect 6972 27858 7028 28028
rect 6636 26908 6692 27804
rect 6972 27806 6974 27858
rect 7026 27806 7028 27858
rect 6972 27794 7028 27806
rect 7080 27076 7136 27086
rect 7080 26984 7082 27020
rect 7134 26984 7136 27020
rect 7080 26972 7136 26984
rect 7308 26908 7364 28588
rect 7420 28550 7476 28588
rect 8092 28532 8148 29260
rect 9212 29092 9268 29596
rect 9548 29428 9604 30102
rect 9772 29764 9828 31388
rect 10108 31378 10164 31388
rect 10444 31658 10556 31668
rect 10444 31106 10500 31658
rect 10444 31054 10446 31106
rect 10498 31054 10500 31106
rect 9884 31033 9940 31045
rect 10444 31042 10500 31054
rect 10556 31556 10612 31566
rect 9884 30996 9886 31033
rect 9938 30996 9940 31033
rect 9884 30930 9940 30940
rect 10108 30996 10164 31006
rect 10108 30434 10164 30940
rect 10108 30382 10110 30434
rect 10162 30382 10164 30434
rect 10108 30370 10164 30382
rect 8988 29036 9268 29092
rect 9324 29426 9604 29428
rect 9324 29374 9550 29426
rect 9602 29374 9604 29426
rect 9324 29372 9604 29374
rect 9324 29092 9380 29372
rect 9548 29362 9604 29372
rect 9660 29708 9828 29764
rect 9660 29428 9716 29708
rect 9660 29362 9716 29372
rect 10424 29426 10480 29438
rect 10424 29374 10426 29426
rect 10478 29374 10480 29426
rect 8428 28980 8484 28990
rect 8988 28980 9044 29036
rect 9324 29026 9380 29036
rect 8296 28644 8352 28682
rect 8296 28578 8352 28588
rect 8092 28476 8260 28532
rect 7476 28084 7532 28094
rect 7532 28028 7700 28084
rect 7476 27990 7532 28028
rect 7532 27242 7588 27254
rect 7532 27190 7534 27242
rect 7586 27190 7588 27242
rect 7532 26908 7588 27190
rect 7644 27188 7700 28028
rect 7756 27860 7812 27870
rect 7756 27766 7812 27804
rect 7868 27858 7924 27870
rect 7868 27806 7870 27858
rect 7922 27806 7924 27858
rect 7868 27524 7924 27806
rect 8036 27860 8092 27870
rect 8036 27766 8092 27804
rect 7868 27458 7924 27468
rect 8204 27188 8260 28476
rect 8428 27746 8484 28924
rect 8764 28924 9044 28980
rect 9660 28980 9716 28990
rect 8764 28644 8820 28924
rect 8988 28644 9044 28654
rect 8764 28642 9044 28644
rect 8764 28590 8990 28642
rect 9042 28590 9044 28642
rect 8764 28588 9044 28590
rect 8540 28532 8596 28542
rect 8540 28530 8820 28532
rect 8540 28478 8542 28530
rect 8594 28478 8820 28530
rect 8540 28476 8820 28478
rect 8540 28466 8596 28476
rect 8428 27694 8430 27746
rect 8482 27694 8484 27746
rect 8428 27682 8484 27694
rect 8764 27188 8820 28476
rect 8988 28308 9044 28588
rect 9660 28420 9716 28924
rect 9864 28868 9920 28878
rect 9864 28642 9920 28812
rect 10108 28868 10164 28878
rect 10424 28868 10480 29374
rect 10108 28866 10480 28868
rect 10108 28814 10110 28866
rect 10162 28814 10480 28866
rect 10108 28812 10480 28814
rect 10108 28802 10164 28812
rect 9864 28590 9866 28642
rect 9918 28590 9920 28642
rect 9864 28578 9920 28590
rect 10556 28654 10612 31500
rect 10668 30772 10724 32508
rect 10780 31722 10836 32678
rect 10892 32564 10948 32574
rect 10892 32470 10948 32508
rect 11004 31892 11060 32732
rect 11228 32116 11284 33180
rect 11340 32900 11396 33852
rect 11340 32834 11396 32844
rect 11676 32788 11732 34076
rect 11900 33572 11956 34748
rect 12124 34692 12180 35084
rect 11900 33506 11956 33516
rect 12012 34636 12180 34692
rect 12012 34132 12068 34636
rect 11900 33236 11956 33246
rect 11900 33142 11956 33180
rect 11676 32722 11732 32732
rect 11676 32589 11732 32601
rect 11676 32537 11678 32589
rect 11730 32537 11732 32589
rect 11676 32228 11732 32537
rect 11676 32162 11732 32172
rect 10780 31670 10782 31722
rect 10834 31670 10836 31722
rect 10780 30996 10836 31670
rect 10892 31836 11060 31892
rect 11116 32060 11284 32116
rect 10892 31220 10948 31836
rect 11116 31780 11172 32060
rect 11340 31780 11396 31790
rect 11116 31778 11396 31780
rect 11116 31734 11342 31778
rect 11060 31726 11342 31734
rect 11394 31726 11396 31778
rect 11060 31724 11396 31726
rect 11060 31722 11172 31724
rect 11060 31670 11062 31722
rect 11114 31670 11172 31722
rect 11340 31714 11396 31724
rect 11452 31780 11508 31790
rect 11060 31668 11172 31670
rect 11060 31658 11116 31668
rect 11060 31220 11116 31230
rect 10892 31218 11116 31220
rect 10892 31166 11062 31218
rect 11114 31166 11116 31218
rect 10892 31164 11116 31166
rect 11060 31154 11116 31164
rect 11452 31021 11508 31724
rect 10780 30940 11060 30996
rect 11452 30969 11454 31021
rect 11506 30969 11508 31021
rect 11452 30957 11508 30969
rect 10668 30716 10948 30772
rect 10780 30548 10836 30558
rect 10668 29540 10724 29550
rect 10668 29446 10724 29484
rect 10556 28644 10668 28654
rect 10556 28588 10612 28644
rect 10612 28550 10668 28588
rect 10780 28420 10836 30492
rect 10892 30378 10948 30716
rect 10892 30326 10894 30378
rect 10946 30326 10948 30378
rect 11004 30436 11060 30940
rect 11004 30370 11060 30380
rect 11788 30436 11844 30446
rect 12012 30436 12068 34076
rect 12236 32228 12292 35196
rect 12348 35140 12404 35150
rect 12348 34858 12404 35084
rect 12348 34806 12350 34858
rect 12402 34806 12404 34858
rect 12516 34970 12572 35308
rect 12796 35252 12852 35262
rect 12796 35138 12852 35196
rect 12796 35086 12798 35138
rect 12850 35086 12852 35138
rect 12796 35074 12852 35086
rect 12516 34918 12518 34970
rect 12570 34918 12572 34970
rect 12516 34916 12572 34918
rect 12516 34840 12572 34860
rect 12348 33796 12404 34806
rect 12684 34692 12740 34702
rect 12460 34356 12516 34366
rect 12460 34130 12516 34300
rect 12460 34078 12462 34130
rect 12514 34078 12516 34130
rect 12460 33908 12516 34078
rect 12684 34356 12740 34636
rect 12684 34130 12740 34300
rect 12964 34244 13020 34254
rect 12964 34150 13020 34188
rect 12684 34078 12686 34130
rect 12738 34078 12740 34130
rect 12684 34066 12740 34078
rect 12460 33842 12516 33852
rect 12348 33730 12404 33740
rect 12124 32172 12292 32228
rect 12348 33572 12404 33582
rect 12124 31892 12180 32172
rect 12124 31826 12180 31836
rect 12236 32004 12292 32014
rect 12236 31734 12292 31948
rect 12216 31722 12292 31734
rect 12216 31670 12218 31722
rect 12270 31670 12292 31722
rect 12216 31668 12292 31670
rect 12216 31658 12272 31668
rect 11788 30434 12068 30436
rect 11788 30382 11790 30434
rect 11842 30382 12068 30434
rect 11788 30380 12068 30382
rect 12124 31556 12180 31566
rect 12348 31556 12404 33516
rect 12852 33572 12908 33582
rect 12852 33478 12908 33516
rect 12460 33346 12516 33358
rect 12460 33294 12462 33346
rect 12514 33294 12516 33346
rect 12460 32004 12516 33294
rect 12572 33348 12628 33358
rect 12572 32676 12628 33292
rect 12796 32788 12852 32798
rect 12796 32694 12852 32732
rect 12572 32610 12628 32620
rect 12460 31938 12516 31948
rect 12460 31668 12516 31678
rect 12460 31574 12516 31612
rect 11788 30370 11844 30380
rect 10892 29988 10948 30326
rect 12124 30324 12180 31500
rect 11900 30268 12180 30324
rect 12236 31500 12404 31556
rect 11004 30212 11060 30222
rect 11004 30118 11060 30156
rect 11340 30212 11396 30222
rect 11340 30210 11508 30212
rect 11340 30158 11342 30210
rect 11394 30158 11508 30210
rect 11340 30156 11508 30158
rect 11340 30146 11396 30156
rect 10892 29932 11396 29988
rect 11340 29482 11396 29932
rect 11340 29430 11342 29482
rect 11394 29430 11396 29482
rect 11340 29418 11396 29430
rect 11452 29092 11508 30156
rect 11900 29316 11956 30268
rect 12031 30154 12087 30166
rect 12031 30102 12033 30154
rect 12085 30102 12087 30154
rect 12031 29540 12087 30102
rect 12236 29876 12292 31500
rect 13244 31220 13300 35980
rect 13448 35698 13504 35710
rect 13448 35646 13450 35698
rect 13502 35646 13504 35698
rect 13448 35364 13504 35646
rect 13448 35298 13504 35308
rect 13580 35140 13636 36430
rect 13804 36484 13860 36494
rect 13692 35588 13748 35598
rect 13692 35494 13748 35532
rect 13580 35074 13636 35084
rect 13804 34916 13860 36428
rect 13916 35252 13972 36652
rect 14028 35698 14084 36988
rect 14420 36594 14476 36988
rect 14420 36542 14422 36594
rect 14474 36542 14476 36594
rect 14420 36530 14476 36542
rect 15596 36932 15652 36942
rect 15484 36482 15540 36494
rect 15484 36430 15486 36482
rect 15538 36430 15540 36482
rect 15148 36260 15204 36270
rect 14028 35646 14030 35698
rect 14082 35646 14084 35698
rect 14028 35634 14084 35646
rect 14812 36258 15204 36260
rect 14812 36206 15150 36258
rect 15202 36206 15204 36258
rect 14812 36204 15204 36206
rect 14812 35698 14868 36204
rect 15148 36194 15204 36204
rect 15484 35924 15540 36430
rect 15596 36482 15652 36876
rect 15596 36430 15598 36482
rect 15650 36430 15652 36482
rect 15596 36418 15652 36430
rect 15484 35858 15540 35868
rect 14812 35646 14814 35698
rect 14866 35646 14868 35698
rect 14812 35634 14868 35646
rect 13916 35186 13972 35196
rect 15596 35364 15652 35374
rect 15148 35140 15204 35150
rect 15148 35046 15204 35084
rect 14028 34916 14084 34926
rect 13804 34914 14084 34916
rect 13804 34862 14030 34914
rect 14082 34862 14084 34914
rect 13804 34860 14084 34862
rect 14028 34850 14084 34860
rect 14904 34858 14960 34870
rect 14904 34806 14906 34858
rect 14958 34806 14960 34858
rect 13748 34692 13804 34702
rect 13748 34690 13860 34692
rect 13748 34638 13750 34690
rect 13802 34638 13860 34690
rect 13748 34626 13860 34638
rect 13636 34020 13692 34030
rect 13244 31154 13300 31164
rect 13468 34018 13692 34020
rect 13468 33966 13638 34018
rect 13690 33966 13692 34018
rect 13468 33964 13692 33966
rect 13468 31780 13524 33964
rect 13636 33954 13692 33964
rect 13804 33908 13860 34626
rect 14904 34356 14960 34806
rect 14644 34300 14960 34356
rect 14364 34244 14420 34254
rect 13916 34132 13972 34142
rect 14252 34130 14308 34142
rect 13916 34038 13972 34076
rect 14084 34074 14140 34086
rect 14084 34022 14086 34074
rect 14138 34022 14140 34074
rect 13804 33852 13972 33908
rect 13580 33796 13636 33806
rect 13580 33458 13636 33740
rect 13580 33406 13582 33458
rect 13634 33406 13636 33458
rect 13580 33394 13636 33406
rect 13692 33684 13748 33694
rect 13692 33318 13748 33628
rect 13648 33306 13748 33318
rect 13648 33254 13650 33306
rect 13702 33254 13748 33306
rect 13648 33180 13748 33254
rect 13804 33348 13860 33358
rect 13804 33257 13806 33292
rect 13858 33257 13860 33292
rect 13804 33245 13860 33257
rect 13916 32228 13972 33852
rect 14084 33572 14140 34022
rect 14084 33506 14140 33516
rect 14252 34078 14254 34130
rect 14306 34078 14308 34130
rect 14252 33290 14308 34078
rect 14252 33238 14254 33290
rect 14306 33238 14308 33290
rect 14364 34130 14420 34188
rect 14644 34242 14700 34300
rect 14644 34190 14646 34242
rect 14698 34190 14700 34242
rect 14644 34178 14700 34190
rect 14364 34078 14366 34130
rect 14418 34078 14420 34130
rect 14364 33348 14420 34078
rect 14812 34132 14868 34142
rect 14364 33282 14420 33292
rect 14588 33572 14644 33582
rect 14588 33313 14644 33516
rect 14588 33261 14590 33313
rect 14642 33261 14644 33313
rect 14588 33249 14644 33261
rect 14252 32900 14308 33238
rect 14252 32844 14644 32900
rect 14364 32676 14420 32686
rect 14364 32618 14420 32620
rect 13916 32162 13972 32172
rect 14028 32564 14084 32574
rect 14364 32566 14366 32618
rect 14418 32566 14420 32618
rect 14364 32554 14420 32566
rect 14588 32601 14644 32844
rect 14812 32676 14868 34076
rect 14924 34130 14980 34142
rect 14924 34078 14926 34130
rect 14978 34078 14980 34130
rect 14924 33908 14980 34078
rect 15148 34132 15204 34142
rect 15148 34038 15204 34076
rect 14924 33842 14980 33852
rect 15036 34020 15092 34030
rect 15036 33908 15092 33964
rect 15428 33908 15484 33918
rect 15036 33906 15484 33908
rect 15036 33854 15430 33906
rect 15482 33854 15484 33906
rect 15036 33852 15484 33854
rect 15036 33694 15092 33852
rect 15428 33842 15484 33852
rect 15032 33684 15092 33694
rect 15596 33684 15652 35308
rect 16044 34914 16100 37090
rect 16044 34862 16046 34914
rect 16098 34862 16100 34914
rect 15708 34692 15764 34702
rect 15708 34598 15764 34636
rect 15088 33628 15092 33684
rect 15148 33628 15652 33684
rect 15032 33308 15088 33628
rect 15032 33256 15034 33308
rect 15086 33256 15088 33308
rect 15032 33244 15088 33256
rect 14812 32620 15092 32676
rect 13580 32004 13636 32014
rect 13580 31910 13636 31948
rect 14028 31734 14084 32508
rect 14588 32549 14590 32601
rect 14642 32549 14644 32601
rect 13356 30996 13412 31006
rect 13468 30996 13524 31724
rect 13974 31722 14084 31734
rect 13974 31670 13976 31722
rect 14028 31670 14084 31722
rect 13974 31668 14084 31670
rect 14140 31778 14196 31790
rect 14140 31726 14142 31778
rect 14194 31726 14196 31778
rect 13974 31556 14030 31668
rect 13974 31490 14030 31500
rect 14140 31332 14196 31726
rect 13244 30994 13524 30996
rect 13244 30942 13358 30994
rect 13410 30942 13524 30994
rect 13244 30940 13524 30942
rect 13804 31276 14196 31332
rect 14252 31778 14308 31790
rect 14252 31726 14254 31778
rect 14306 31726 14308 31778
rect 12908 30212 12964 30222
rect 12796 30210 12964 30212
rect 12796 30158 12910 30210
rect 12962 30158 12964 30210
rect 12796 30156 12964 30158
rect 12236 29820 12516 29876
rect 12031 29484 12180 29540
rect 12012 29316 12068 29326
rect 11900 29314 12068 29316
rect 11900 29262 12014 29314
rect 12066 29262 12068 29314
rect 11900 29260 12068 29262
rect 12012 29250 12068 29260
rect 12124 29092 12180 29484
rect 11452 29026 11508 29036
rect 12012 29036 12180 29092
rect 12236 29426 12292 29438
rect 12236 29374 12238 29426
rect 12290 29374 12292 29426
rect 11340 28868 11396 28878
rect 11340 28614 11396 28812
rect 9660 28364 9940 28420
rect 8988 28252 9772 28308
rect 8932 28026 8988 28038
rect 8932 27974 8934 28026
rect 8986 27974 8988 28026
rect 8932 27972 8988 27974
rect 8932 27906 8988 27916
rect 9716 27970 9772 28252
rect 9716 27918 9718 27970
rect 9770 27918 9772 27970
rect 9716 27906 9772 27918
rect 9100 27858 9156 27870
rect 9100 27806 9102 27858
rect 9154 27806 9156 27858
rect 9100 27748 9156 27806
rect 9100 27682 9156 27692
rect 9324 27860 9380 27870
rect 8204 27132 8484 27188
rect 8764 27132 8932 27188
rect 7644 27122 7700 27132
rect 7756 27074 7812 27086
rect 7756 27022 7758 27074
rect 7810 27022 7812 27074
rect 7756 26908 7812 27022
rect 8260 26962 8316 26974
rect 8260 26910 8262 26962
rect 8314 26910 8316 26962
rect 8260 26908 8316 26910
rect 6636 26852 6804 26908
rect 6524 26180 6580 26190
rect 6524 24778 6580 26124
rect 6636 25732 6692 25742
rect 6636 25506 6692 25676
rect 6636 25454 6638 25506
rect 6690 25454 6692 25506
rect 6636 25442 6692 25454
rect 6748 24948 6804 26852
rect 6860 26852 7364 26908
rect 7420 26852 7588 26908
rect 7644 26852 7812 26908
rect 7868 26852 7924 26862
rect 6860 25618 6916 26852
rect 6972 26346 7028 26358
rect 6972 26294 6974 26346
rect 7026 26294 7028 26346
rect 6972 25844 7028 26294
rect 6972 25788 7252 25844
rect 6860 25566 6862 25618
rect 6914 25566 6916 25618
rect 6860 25554 6916 25566
rect 6972 25620 7028 25630
rect 6748 24892 6916 24948
rect 6524 24726 6526 24778
rect 6578 24726 6580 24778
rect 6524 23770 6580 24726
rect 6860 24612 6916 24892
rect 6748 24556 6916 24612
rect 6972 24778 7028 25564
rect 7084 25508 7140 25518
rect 7084 25414 7140 25452
rect 6972 24726 6974 24778
rect 7026 24726 7028 24778
rect 6972 24724 7028 24726
rect 6524 23718 6526 23770
rect 6578 23718 6580 23770
rect 6524 23706 6580 23718
rect 6636 23940 6692 23960
rect 6636 23882 6692 23884
rect 6636 23830 6638 23882
rect 6690 23830 6692 23882
rect 6524 23268 6580 23278
rect 6524 23154 6580 23212
rect 6524 23102 6526 23154
rect 6578 23102 6580 23154
rect 6524 23090 6580 23102
rect 6636 22820 6692 23830
rect 6748 23042 6804 24556
rect 6860 24388 6916 24398
rect 6860 23882 6916 24332
rect 6860 23830 6862 23882
rect 6914 23830 6916 23882
rect 6972 23940 7028 24668
rect 6972 23874 7028 23884
rect 6860 23716 6916 23830
rect 6860 23660 7028 23716
rect 6748 22990 6750 23042
rect 6802 22990 6804 23042
rect 6748 22978 6804 22990
rect 6860 23181 6916 23193
rect 6860 23129 6862 23181
rect 6914 23129 6916 23181
rect 6860 23044 6916 23129
rect 6860 22978 6916 22988
rect 6972 22820 7028 23660
rect 7196 23380 7252 25788
rect 7420 25732 7476 26852
rect 7532 26516 7588 26526
rect 7532 26346 7588 26460
rect 7532 26294 7534 26346
rect 7586 26294 7588 26346
rect 7532 26282 7588 26294
rect 7532 25732 7588 25742
rect 7420 25676 7532 25732
rect 7532 25506 7588 25676
rect 7532 25454 7534 25506
rect 7586 25454 7588 25506
rect 7532 25442 7588 25454
rect 7644 24612 7700 26852
rect 7644 24546 7700 24556
rect 7756 25396 7812 25406
rect 7756 24724 7812 25340
rect 7756 24164 7812 24668
rect 7868 24500 7924 26796
rect 8092 26852 8316 26908
rect 8092 26516 8148 26852
rect 8428 26740 8484 27132
rect 8540 27076 8596 27086
rect 8540 26982 8596 27020
rect 8652 27074 8708 27086
rect 8652 27022 8654 27074
rect 8706 27022 8708 27074
rect 8652 26740 8708 27022
rect 8092 26450 8148 26460
rect 8316 26684 8484 26740
rect 8540 26684 8708 26740
rect 8764 26964 8820 26974
rect 8316 26402 8372 26684
rect 8540 26628 8596 26684
rect 8316 26350 8318 26402
rect 8370 26350 8372 26402
rect 8316 26338 8372 26350
rect 8428 26572 8596 26628
rect 8092 26292 8148 26302
rect 8092 26198 8148 26236
rect 8428 25620 8484 26572
rect 8652 26516 8708 26526
rect 8540 26346 8596 26358
rect 8540 26294 8542 26346
rect 8594 26294 8596 26346
rect 8540 25732 8596 26294
rect 8540 25666 8596 25676
rect 8428 25554 8484 25564
rect 8092 25506 8148 25518
rect 8092 25454 8094 25506
rect 8146 25454 8148 25506
rect 8540 25506 8596 25518
rect 7980 25172 8036 25182
rect 7980 24778 8036 25116
rect 7980 24726 7982 24778
rect 8034 24726 8036 24778
rect 8092 24836 8148 25454
rect 8260 25450 8316 25462
rect 8260 25398 8262 25450
rect 8314 25398 8316 25450
rect 8540 25454 8542 25506
rect 8594 25454 8596 25506
rect 8260 24948 8316 25398
rect 8428 25396 8484 25406
rect 8428 25302 8484 25340
rect 8540 25172 8596 25454
rect 8540 25106 8596 25116
rect 8652 24948 8708 26460
rect 8764 25742 8820 26908
rect 8876 26516 8932 27132
rect 9324 27186 9380 27804
rect 9324 27134 9326 27186
rect 9378 27134 9380 27186
rect 9324 27122 9380 27134
rect 9772 27412 9828 27422
rect 9548 27076 9604 27086
rect 9548 26982 9604 27020
rect 9772 27074 9828 27356
rect 9772 27022 9774 27074
rect 9826 27022 9828 27074
rect 9772 27010 9828 27022
rect 8876 26450 8932 26460
rect 9436 26292 9492 26302
rect 9436 26198 9492 26236
rect 9604 26068 9660 26078
rect 8988 26066 9660 26068
rect 8988 26014 9606 26066
rect 9658 26014 9660 26066
rect 8988 26012 9660 26014
rect 8764 25730 8876 25742
rect 8764 25678 8822 25730
rect 8874 25678 8876 25730
rect 8764 25676 8876 25678
rect 8820 25666 8876 25676
rect 8260 24892 8484 24948
rect 8652 24892 8932 24948
rect 8092 24770 8148 24780
rect 7980 24714 8036 24726
rect 8316 24724 8372 24734
rect 8316 24630 8372 24668
rect 7868 24444 8090 24500
rect 7756 24108 7924 24164
rect 7756 23940 7812 23950
rect 7196 23314 7252 23324
rect 7308 23882 7364 23894
rect 7308 23830 7310 23882
rect 7362 23830 7364 23882
rect 7756 23846 7812 23884
rect 7868 23938 7924 24108
rect 7868 23886 7870 23938
rect 7922 23886 7924 23938
rect 7868 23874 7924 23886
rect 8034 23940 8090 24444
rect 8428 24162 8484 24892
rect 8540 24836 8596 24846
rect 8540 24742 8596 24780
rect 8708 24724 8764 24734
rect 8708 24630 8764 24668
rect 8876 24164 8932 24892
rect 8988 24724 9044 26012
rect 9604 26002 9660 26012
rect 9884 25620 9940 28364
rect 10668 28364 10836 28420
rect 10892 28586 10948 28598
rect 10892 28534 10894 28586
rect 10946 28534 10948 28586
rect 10220 28084 10276 28094
rect 10220 27914 10276 28028
rect 9996 27886 10052 27898
rect 9996 27834 9998 27886
rect 10050 27834 10052 27886
rect 9996 27524 10052 27834
rect 10220 27862 10222 27914
rect 10274 27862 10276 27914
rect 9996 27468 10164 27524
rect 9996 27188 10052 27198
rect 9996 26740 10052 27132
rect 10108 26964 10164 27468
rect 10220 27412 10276 27862
rect 10444 27886 10500 27898
rect 10444 27860 10446 27886
rect 10498 27860 10500 27886
rect 10444 27794 10500 27804
rect 10556 27893 10612 27905
rect 10556 27841 10558 27893
rect 10610 27841 10612 27893
rect 10556 27636 10612 27841
rect 10556 27570 10612 27580
rect 10668 27412 10724 28364
rect 10892 28196 10948 28534
rect 11116 28586 11172 28598
rect 11116 28534 11118 28586
rect 11170 28534 11172 28586
rect 10220 27346 10276 27356
rect 10556 27356 10724 27412
rect 10780 28140 10948 28196
rect 11004 28420 11060 28430
rect 10780 27860 10836 28140
rect 10892 27972 10948 27982
rect 10892 27914 10948 27916
rect 10892 27862 10894 27914
rect 10946 27862 10948 27914
rect 10892 27850 10948 27862
rect 11004 27914 11060 28364
rect 11004 27862 11006 27914
rect 11058 27862 11060 27914
rect 11004 27850 11060 27862
rect 10332 27188 10388 27198
rect 10332 27074 10388 27132
rect 10332 27022 10334 27074
rect 10386 27022 10388 27074
rect 10332 27010 10388 27022
rect 10220 26964 10276 26974
rect 10108 26908 10220 26964
rect 9996 26684 10164 26740
rect 9884 25554 9940 25564
rect 10108 25620 10164 26684
rect 10220 26526 10276 26908
rect 10220 26514 10332 26526
rect 10220 26462 10278 26514
rect 10330 26462 10332 26514
rect 10220 26460 10332 26462
rect 10276 26450 10332 26460
rect 10444 26290 10500 26302
rect 10444 26238 10446 26290
rect 10498 26238 10500 26290
rect 10444 26180 10500 26238
rect 10108 25554 10164 25564
rect 10220 26124 10500 26180
rect 8988 24658 9044 24668
rect 9100 25508 9156 25518
rect 8428 24110 8430 24162
rect 8482 24110 8484 24162
rect 8428 24098 8484 24110
rect 8540 24108 8932 24164
rect 8034 23846 8090 23884
rect 7308 23268 7364 23830
rect 6636 22764 6804 22820
rect 5852 22542 5854 22594
rect 5906 22542 5908 22594
rect 5852 22530 5908 22542
rect 6076 22540 6468 22596
rect 5740 21858 5796 21868
rect 5628 21422 5630 21474
rect 5682 21422 5684 21474
rect 5628 21410 5684 21422
rect 5852 21588 5908 21598
rect 5852 21026 5908 21532
rect 5852 20974 5854 21026
rect 5906 20974 5908 21026
rect 5852 20962 5908 20974
rect 5180 20804 5236 20814
rect 5180 20710 5236 20748
rect 5516 20804 5572 20814
rect 6076 20804 6132 22540
rect 6300 22372 6356 22382
rect 6300 22278 6356 22316
rect 6412 22370 6468 22382
rect 6412 22318 6414 22370
rect 6466 22318 6468 22370
rect 6412 22260 6468 22318
rect 6580 22372 6636 22382
rect 6580 22278 6636 22316
rect 6412 22194 6468 22204
rect 6524 21924 6580 21934
rect 5068 19350 5070 19402
rect 5122 19350 5124 19402
rect 5068 19338 5124 19350
rect 4956 19142 5012 19180
rect 4284 18946 4340 18956
rect 5404 19012 5460 19022
rect 4004 18722 4060 18732
rect 2268 18386 2324 18396
rect 3052 18452 3108 18462
rect 3052 18358 3108 18396
rect 5292 18452 5348 18462
rect 3836 18340 3892 18350
rect 3836 18246 3892 18284
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 5124 17780 5180 17790
rect 5124 17686 5180 17724
rect 5292 17668 5348 18396
rect 5404 17668 5460 18956
rect 5516 18452 5572 20748
rect 5852 20748 6132 20804
rect 6412 20802 6468 20814
rect 5684 19908 5740 19918
rect 5516 18386 5572 18396
rect 5628 19906 5740 19908
rect 5628 19854 5686 19906
rect 5738 19854 5740 19906
rect 5628 19842 5740 19854
rect 5516 17668 5572 17678
rect 5404 17666 5572 17668
rect 5404 17614 5518 17666
rect 5570 17614 5572 17666
rect 5404 17612 5572 17614
rect 4228 17556 4284 17566
rect 4228 17462 4284 17500
rect 4676 17556 4732 17566
rect 4676 17462 4732 17500
rect 4340 17108 4396 17118
rect 4340 17014 4396 17052
rect 5068 16882 5124 16894
rect 5068 16830 5070 16882
rect 5122 16830 5124 16882
rect 3892 16770 3948 16782
rect 3892 16718 3894 16770
rect 3946 16718 3948 16770
rect 2268 16658 2324 16670
rect 2268 16606 2270 16658
rect 2322 16606 2324 16658
rect 2268 16100 2324 16606
rect 3052 16660 3108 16670
rect 3892 16660 3948 16718
rect 4732 16772 4788 16782
rect 4732 16678 4788 16716
rect 3052 16658 3948 16660
rect 3052 16606 3054 16658
rect 3106 16606 3948 16658
rect 3052 16604 3948 16606
rect 3052 16594 3108 16604
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 5068 16324 5124 16830
rect 5180 16884 5236 16894
rect 5292 16884 5348 17612
rect 5516 17602 5572 17612
rect 5628 17108 5684 19842
rect 5740 18452 5796 18462
rect 5740 18358 5796 18396
rect 5740 17666 5796 17678
rect 5740 17614 5742 17666
rect 5794 17614 5796 17666
rect 5740 17556 5796 17614
rect 5740 17490 5796 17500
rect 5628 17042 5684 17052
rect 5180 16882 5348 16884
rect 5180 16830 5182 16882
rect 5234 16830 5348 16882
rect 5180 16828 5348 16830
rect 5180 16818 5236 16828
rect 5852 16548 5908 20748
rect 6246 20746 6302 20758
rect 6246 20694 6248 20746
rect 6300 20694 6302 20746
rect 6246 20468 6302 20694
rect 6246 20402 6302 20412
rect 6412 20750 6414 20802
rect 6466 20750 6468 20802
rect 6412 20244 6468 20750
rect 6524 20802 6580 21868
rect 6748 21812 6804 22764
rect 6860 22764 7028 22820
rect 7196 23154 7252 23166
rect 7196 23102 7198 23154
rect 7250 23102 7252 23154
rect 7196 22932 7252 23102
rect 6860 22372 6916 22764
rect 6972 22596 7028 22606
rect 7196 22596 7252 22876
rect 6972 22594 7252 22596
rect 6972 22542 6974 22594
rect 7026 22542 7252 22594
rect 6972 22540 7252 22542
rect 6972 22530 7028 22540
rect 7196 22372 7252 22382
rect 6860 22316 7028 22372
rect 6748 21756 6916 21812
rect 6639 21625 6695 21637
rect 6639 21573 6641 21625
rect 6693 21573 6695 21625
rect 6639 21140 6695 21573
rect 6524 20750 6526 20802
rect 6578 20750 6580 20802
rect 6524 20738 6580 20750
rect 6636 21084 6695 21140
rect 6636 20580 6692 21084
rect 6636 20514 6692 20524
rect 6412 20188 6692 20244
rect 6636 20132 6692 20188
rect 6490 20055 6546 20067
rect 6490 20003 6492 20055
rect 6544 20030 6546 20055
rect 6544 20020 6580 20030
rect 6490 19964 6524 20003
rect 6524 19954 6580 19964
rect 6636 20018 6692 20076
rect 6636 19966 6638 20018
rect 6690 19966 6692 20018
rect 6636 19954 6692 19966
rect 6748 20020 6804 20030
rect 6860 20020 6916 21756
rect 6972 21754 7028 22316
rect 6972 21702 6974 21754
rect 7026 21702 7028 21754
rect 6972 21690 7028 21702
rect 7196 21586 7252 22316
rect 7308 22370 7364 23212
rect 7308 22318 7310 22370
rect 7362 22318 7364 22370
rect 7308 22306 7364 22318
rect 7532 23380 7588 23390
rect 7532 22260 7588 23324
rect 8540 23278 8596 24108
rect 8876 23938 8932 23950
rect 8876 23886 8878 23938
rect 8930 23886 8932 23938
rect 8876 23828 8932 23886
rect 8876 23762 8932 23772
rect 8484 23266 8596 23278
rect 8484 23214 8486 23266
rect 8538 23214 8596 23266
rect 8484 23212 8596 23214
rect 8484 23202 8540 23212
rect 7756 23156 7812 23166
rect 8092 23156 8148 23166
rect 7756 23062 7812 23100
rect 7924 23098 7980 23110
rect 7924 23046 7926 23098
rect 7978 23046 7980 23098
rect 8092 23062 8148 23100
rect 8204 23154 8260 23166
rect 8204 23102 8206 23154
rect 8258 23102 8260 23154
rect 7924 22820 7980 23046
rect 8204 22932 8260 23102
rect 8204 22866 8260 22876
rect 7644 22764 7980 22820
rect 7644 22594 7700 22764
rect 7644 22542 7646 22594
rect 7698 22542 7700 22594
rect 7644 22530 7700 22542
rect 7924 22596 7980 22764
rect 7924 22530 7980 22540
rect 9100 22482 9156 25452
rect 9212 25506 9268 25518
rect 9212 25454 9214 25506
rect 9266 25454 9268 25506
rect 9212 25172 9268 25454
rect 10088 25452 10144 25462
rect 9940 25450 10144 25452
rect 9324 25396 9380 25406
rect 9324 25172 9380 25340
rect 9940 25398 10090 25450
rect 10142 25398 10144 25450
rect 9940 25396 10144 25398
rect 9324 25116 9716 25172
rect 9212 24106 9268 25116
rect 9436 24722 9492 24734
rect 9436 24670 9438 24722
rect 9490 24670 9492 24722
rect 9436 24612 9492 24670
rect 9436 24546 9492 24556
rect 9660 24722 9716 25116
rect 9940 24834 9996 25396
rect 10088 25386 10144 25396
rect 10220 25172 10276 26124
rect 10556 26068 10612 27356
rect 10668 27076 10724 27086
rect 10780 27076 10836 27804
rect 11116 27748 11172 28534
rect 11340 28562 11342 28614
rect 11394 28562 11396 28614
rect 11676 28642 11732 28654
rect 11900 28644 11956 28654
rect 11340 28084 11396 28562
rect 11452 28586 11508 28598
rect 11452 28534 11454 28586
rect 11506 28534 11508 28586
rect 11452 28084 11508 28534
rect 11676 28590 11678 28642
rect 11730 28590 11732 28642
rect 11452 28028 11620 28084
rect 11340 28018 11396 28028
rect 11228 27972 11284 27982
rect 11228 27914 11284 27916
rect 11228 27862 11230 27914
rect 11282 27862 11284 27914
rect 11228 27850 11284 27862
rect 11452 27886 11508 27898
rect 11452 27834 11454 27886
rect 11506 27834 11508 27886
rect 11452 27748 11508 27834
rect 11116 27692 11508 27748
rect 11116 27188 11172 27692
rect 11116 27094 11172 27132
rect 11564 27188 11620 28028
rect 11564 27122 11620 27132
rect 10668 27074 10836 27076
rect 10668 27022 10670 27074
rect 10722 27022 10836 27074
rect 11340 27074 11396 27086
rect 10668 27020 10836 27022
rect 10668 27010 10724 27020
rect 10948 27018 11004 27030
rect 10948 26966 10950 27018
rect 11002 26966 11004 27018
rect 10948 26908 11004 26966
rect 11340 27022 11342 27074
rect 11394 27022 11396 27074
rect 11340 26964 11396 27022
rect 11508 27018 11564 27030
rect 11508 26966 11510 27018
rect 11562 26966 11564 27018
rect 11508 26964 11564 26966
rect 10948 26852 11060 26908
rect 11004 26740 11060 26852
rect 10780 26684 11004 26740
rect 10780 26514 10836 26684
rect 11004 26674 11060 26684
rect 11228 26852 11396 26908
rect 11452 26908 11564 26964
rect 11676 26964 11732 28590
rect 10780 26462 10782 26514
rect 10834 26462 10836 26514
rect 10780 26450 10836 26462
rect 10332 26012 10612 26068
rect 11116 26290 11172 26302
rect 11116 26238 11118 26290
rect 11170 26238 11172 26290
rect 10332 25730 10388 26012
rect 10332 25678 10334 25730
rect 10386 25678 10388 25730
rect 10332 25666 10388 25678
rect 10220 25106 10276 25116
rect 10332 25508 10388 25518
rect 9940 24782 9942 24834
rect 9994 24782 9996 24834
rect 9940 24770 9996 24782
rect 9660 24670 9662 24722
rect 9714 24670 9716 24722
rect 9212 24054 9214 24106
rect 9266 24054 9268 24106
rect 9212 24042 9268 24054
rect 9212 23940 9268 23950
rect 9212 23846 9268 23884
rect 9436 23156 9492 23166
rect 9436 23154 9604 23156
rect 9436 23102 9438 23154
rect 9490 23102 9604 23154
rect 9436 23100 9604 23102
rect 9436 23090 9492 23100
rect 9100 22430 9102 22482
rect 9154 22430 9156 22482
rect 9100 22418 9156 22430
rect 9212 22596 9268 22606
rect 9212 22355 9268 22540
rect 9212 22303 9214 22355
rect 9266 22303 9268 22355
rect 9212 22291 9268 22303
rect 9436 22372 9492 22382
rect 9436 22278 9492 22316
rect 7532 22204 7924 22260
rect 7756 21588 7812 21598
rect 7196 21534 7198 21586
rect 7250 21534 7252 21586
rect 6972 20916 7028 20926
rect 7196 20916 7252 21534
rect 6972 20914 7252 20916
rect 6972 20862 6974 20914
rect 7026 20862 7252 20914
rect 6972 20860 7252 20862
rect 7644 21586 7812 21588
rect 7644 21534 7758 21586
rect 7810 21534 7812 21586
rect 7644 21532 7812 21534
rect 6972 20850 7028 20860
rect 7644 20804 7700 21532
rect 7756 21522 7812 21532
rect 7868 21364 7924 22204
rect 8764 21588 8820 21598
rect 9548 21588 9604 23100
rect 9660 22596 9716 24670
rect 10108 23938 10164 23950
rect 10108 23886 10110 23938
rect 10162 23886 10164 23938
rect 9772 23714 9828 23726
rect 9772 23662 9774 23714
rect 9826 23662 9828 23714
rect 9772 23156 9828 23662
rect 9772 23090 9828 23100
rect 9660 22530 9716 22540
rect 10108 22596 10164 23886
rect 10220 23156 10276 23166
rect 10220 23062 10276 23100
rect 10108 22530 10164 22540
rect 9884 22372 9940 22382
rect 9660 21588 9716 21598
rect 9548 21586 9716 21588
rect 9548 21534 9662 21586
rect 9714 21534 9716 21586
rect 9548 21532 9716 21534
rect 8764 21494 8820 21532
rect 6748 20018 6916 20020
rect 6748 19966 6750 20018
rect 6802 19966 6916 20018
rect 6748 19964 6916 19966
rect 6972 20132 7028 20142
rect 6748 19954 6804 19964
rect 6076 19796 6132 19806
rect 6076 19702 6132 19740
rect 6636 19796 6692 19806
rect 6188 19402 6244 19414
rect 6188 19350 6190 19402
rect 6242 19350 6244 19402
rect 6076 19236 6132 19246
rect 5964 19234 6132 19236
rect 5964 19182 6078 19234
rect 6130 19182 6132 19234
rect 5964 19180 6132 19182
rect 5964 17902 6020 19180
rect 6076 19170 6132 19180
rect 6188 18900 6244 19350
rect 6132 18844 6244 18900
rect 6412 19234 6468 19246
rect 6412 19182 6414 19234
rect 6466 19182 6468 19234
rect 6132 18506 6188 18844
rect 6412 18788 6468 19182
rect 6636 19236 6692 19740
rect 6972 19796 7028 20076
rect 7532 20020 7588 20030
rect 7532 19926 7588 19964
rect 7196 19908 7252 19918
rect 7196 19814 7252 19852
rect 6972 19730 7028 19740
rect 6972 19460 7028 19470
rect 6972 19366 7028 19404
rect 7644 19236 7700 20748
rect 7756 21308 7924 21364
rect 8428 21364 8484 21374
rect 8428 21362 8932 21364
rect 8428 21310 8430 21362
rect 8482 21310 8932 21362
rect 8428 21308 8932 21310
rect 7756 20018 7812 21308
rect 8428 21298 8484 21308
rect 8876 20914 8932 21308
rect 8876 20862 8878 20914
rect 8930 20862 8932 20914
rect 8876 20850 8932 20862
rect 9324 20916 9380 20926
rect 7756 19966 7758 20018
rect 7810 19966 7812 20018
rect 7756 19460 7812 19966
rect 7868 20018 7924 20030
rect 7868 19966 7870 20018
rect 7922 19966 7924 20018
rect 7868 19908 7924 19966
rect 7868 19842 7924 19852
rect 8036 20018 8092 20030
rect 8036 19966 8038 20018
rect 8090 19966 8092 20018
rect 8036 19684 8092 19966
rect 8428 20020 8484 20030
rect 8428 19906 8484 19964
rect 8428 19854 8430 19906
rect 8482 19854 8484 19906
rect 8428 19842 8484 19854
rect 9044 19906 9100 19918
rect 9044 19854 9046 19906
rect 9098 19854 9100 19906
rect 9044 19796 9100 19854
rect 9044 19730 9100 19740
rect 9212 19796 9268 19806
rect 8036 19618 8092 19628
rect 7756 19394 7812 19404
rect 8988 19460 9044 19470
rect 8988 19366 9044 19404
rect 7868 19236 7924 19246
rect 7644 19234 7924 19236
rect 7644 19182 7870 19234
rect 7922 19182 7924 19234
rect 7644 19180 7924 19182
rect 6636 19142 6692 19180
rect 7868 19170 7924 19180
rect 6412 18722 6468 18732
rect 6524 19012 6580 19022
rect 6132 18454 6134 18506
rect 6186 18454 6188 18506
rect 6132 18442 6188 18454
rect 6524 18450 6580 18956
rect 7532 19012 7588 19022
rect 7532 18918 7588 18956
rect 8596 19012 8652 19022
rect 8596 19010 8820 19012
rect 8596 18958 8598 19010
rect 8650 18958 8820 19010
rect 8596 18956 8820 18958
rect 8596 18946 8652 18956
rect 6524 18398 6526 18450
rect 6578 18398 6580 18450
rect 6524 18386 6580 18398
rect 6860 18488 6916 18500
rect 6860 18436 6862 18488
rect 6914 18436 6916 18488
rect 8316 18465 8372 18477
rect 6300 18340 6356 18350
rect 6300 18246 6356 18284
rect 5964 17890 6076 17902
rect 5964 17838 6022 17890
rect 6074 17838 6076 17890
rect 5964 17836 6076 17838
rect 6020 17826 6076 17836
rect 6412 17668 6468 17678
rect 6412 17574 6468 17612
rect 6860 17556 6916 18436
rect 7924 18452 7980 18462
rect 7924 18358 7980 18396
rect 8316 18413 8318 18465
rect 8370 18413 8372 18465
rect 7476 18338 7532 18350
rect 7476 18286 7478 18338
rect 7530 18286 7532 18338
rect 7476 18228 7532 18286
rect 7476 18162 7532 18172
rect 8204 18338 8260 18350
rect 8204 18286 8206 18338
rect 8258 18286 8260 18338
rect 8204 18004 8260 18286
rect 7196 17948 8260 18004
rect 7196 17778 7252 17948
rect 7196 17726 7198 17778
rect 7250 17726 7252 17778
rect 7196 17714 7252 17726
rect 8316 17892 8372 18413
rect 6916 17500 7140 17556
rect 6860 17462 6916 17500
rect 5964 16772 6020 16782
rect 5964 16678 6020 16716
rect 7084 16548 7140 17500
rect 8316 17108 8372 17836
rect 8540 18450 8596 18462
rect 8540 18398 8542 18450
rect 8594 18398 8596 18450
rect 8540 18340 8596 18398
rect 8540 17780 8596 18284
rect 8540 17714 8596 17724
rect 8652 17892 8708 17902
rect 7868 16772 7924 16782
rect 5852 16492 6356 16548
rect 5068 16268 6132 16324
rect 2044 16098 2324 16100
rect 2044 16046 2270 16098
rect 2322 16046 2324 16098
rect 2044 16044 2324 16046
rect 2044 14530 2100 16044
rect 2268 16034 2324 16044
rect 3052 16098 3108 16110
rect 3052 16046 3054 16098
rect 3106 16046 3108 16098
rect 3052 15540 3108 16046
rect 5964 16098 6020 16110
rect 5964 16046 5966 16098
rect 6018 16046 6020 16098
rect 4284 15988 4340 15998
rect 3052 15474 3108 15484
rect 3500 15540 3556 15550
rect 3500 15446 3556 15484
rect 3836 15316 3892 15326
rect 3836 15222 3892 15260
rect 4284 15314 4340 15932
rect 4956 15988 5012 15998
rect 4956 15894 5012 15932
rect 4284 15262 4286 15314
rect 4338 15262 4340 15314
rect 4508 15876 4564 15886
rect 4508 15358 4564 15820
rect 5068 15482 5124 15494
rect 4508 15306 4510 15358
rect 4562 15306 4564 15358
rect 4508 15294 4564 15306
rect 4956 15428 5012 15438
rect 4956 15314 5012 15372
rect 4284 15250 4340 15262
rect 4956 15262 4958 15314
rect 5010 15262 5012 15314
rect 4956 15250 5012 15262
rect 5068 15430 5070 15482
rect 5122 15430 5124 15482
rect 5068 15316 5124 15430
rect 5404 15428 5460 15438
rect 5068 15250 5124 15260
rect 5292 15341 5348 15353
rect 5292 15289 5294 15341
rect 5346 15289 5348 15341
rect 4620 15204 4676 15242
rect 4620 15138 4676 15148
rect 5292 15204 5348 15289
rect 5292 15138 5348 15148
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 2044 14478 2046 14530
rect 2098 14478 2100 14530
rect 2044 13972 2100 14478
rect 2828 14532 2884 14542
rect 4732 14532 4788 14542
rect 2828 14530 3108 14532
rect 2828 14478 2830 14530
rect 2882 14478 3108 14530
rect 2828 14476 3108 14478
rect 2828 14466 2884 14476
rect 3052 13972 3108 14476
rect 4732 14438 4788 14476
rect 5068 14308 5124 14318
rect 3164 13972 3220 13982
rect 3052 13970 3220 13972
rect 3052 13918 3166 13970
rect 3218 13918 3220 13970
rect 3052 13916 3220 13918
rect 2044 13906 2100 13916
rect 3164 13906 3220 13916
rect 3388 13972 3444 13982
rect 3388 11732 3444 13916
rect 4900 13972 4956 13982
rect 4900 13878 4956 13916
rect 3500 13748 3556 13758
rect 3500 13654 3556 13692
rect 5068 13746 5124 14252
rect 5404 13972 5460 15372
rect 5964 15428 6020 16046
rect 6076 15930 6132 16268
rect 6076 15878 6078 15930
rect 6130 15878 6132 15930
rect 6076 15866 6132 15878
rect 6188 15988 6244 15998
rect 5964 15362 6020 15372
rect 5628 15314 5684 15326
rect 5628 15262 5630 15314
rect 5682 15262 5684 15314
rect 5628 15148 5684 15262
rect 6188 15314 6244 15932
rect 6188 15262 6190 15314
rect 6242 15262 6244 15314
rect 6188 15250 6244 15262
rect 6300 15148 6356 16492
rect 6860 16492 7140 16548
rect 7644 16770 7924 16772
rect 7644 16718 7870 16770
rect 7922 16718 7924 16770
rect 7644 16716 7924 16718
rect 6412 16212 6468 16222
rect 6412 16059 6468 16156
rect 6412 16007 6414 16059
rect 6466 16007 6468 16059
rect 6412 15995 6468 16007
rect 6636 16098 6692 16110
rect 6636 16046 6638 16098
rect 6690 16046 6692 16098
rect 6524 15329 6580 15341
rect 6524 15277 6526 15329
rect 6578 15277 6580 15329
rect 5628 15092 5796 15148
rect 6300 15092 6468 15148
rect 5740 14642 5796 15092
rect 5740 14590 5742 14642
rect 5794 14590 5796 14642
rect 5740 14578 5796 14590
rect 5852 14980 5908 14990
rect 5852 14515 5908 14924
rect 5852 14463 5854 14515
rect 5906 14463 5908 14515
rect 5852 14451 5908 14463
rect 6076 14532 6132 14542
rect 6076 14438 6132 14476
rect 5404 13970 5908 13972
rect 5404 13918 5406 13970
rect 5458 13918 5908 13970
rect 5404 13916 5908 13918
rect 5404 13906 5460 13916
rect 5068 13694 5070 13746
rect 5122 13694 5124 13746
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4844 12738 4900 12750
rect 4844 12686 4846 12738
rect 4898 12686 4900 12738
rect 3388 11666 3444 11676
rect 3948 12178 4004 12190
rect 3948 12126 3950 12178
rect 4002 12126 4004 12178
rect 3948 11732 4004 12126
rect 4732 12180 4788 12190
rect 4844 12180 4900 12686
rect 5068 12404 5124 13694
rect 5180 12962 5236 12974
rect 5180 12910 5182 12962
rect 5234 12910 5236 12962
rect 5180 12740 5236 12910
rect 5628 12962 5684 13916
rect 5852 13746 5908 13916
rect 5852 13694 5854 13746
rect 5906 13694 5908 13746
rect 5852 13682 5908 13694
rect 5964 13914 6020 13926
rect 5964 13862 5966 13914
rect 6018 13862 6020 13914
rect 5964 13748 6020 13862
rect 5964 13682 6020 13692
rect 6300 13785 6356 13797
rect 6300 13733 6302 13785
rect 6354 13733 6356 13785
rect 6300 13412 6356 13733
rect 6300 13346 6356 13356
rect 5628 12910 5630 12962
rect 5682 12910 5684 12962
rect 6300 13076 6356 13086
rect 6300 12962 6356 13020
rect 5628 12898 5684 12910
rect 6076 12906 6132 12918
rect 6076 12854 6078 12906
rect 6130 12854 6132 12906
rect 6300 12910 6302 12962
rect 6354 12910 6356 12962
rect 6300 12898 6356 12910
rect 5740 12794 5796 12806
rect 5740 12742 5742 12794
rect 5794 12742 5796 12794
rect 5740 12740 5796 12742
rect 5180 12684 5796 12740
rect 4732 12178 4900 12180
rect 4732 12126 4734 12178
rect 4786 12126 4900 12178
rect 4732 12124 4900 12126
rect 4956 12348 5124 12404
rect 4732 12114 4788 12124
rect 4956 11844 5012 12348
rect 4476 11788 4740 11798
rect 4956 11788 5348 11844
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 1820 11508 1876 11518
rect 1820 11396 1876 11452
rect 1708 11394 1876 11396
rect 1708 11342 1822 11394
rect 1874 11342 1876 11394
rect 1708 11340 1876 11342
rect 1596 9828 1652 9838
rect 1708 9828 1764 11340
rect 1820 11330 1876 11340
rect 2604 11396 2660 11406
rect 2604 11394 2884 11396
rect 2604 11342 2606 11394
rect 2658 11342 2884 11394
rect 2604 11340 2884 11342
rect 2604 11330 2660 11340
rect 2828 10836 2884 11340
rect 2940 10836 2996 10846
rect 2828 10834 2996 10836
rect 2828 10782 2942 10834
rect 2994 10782 2996 10834
rect 2828 10780 2996 10782
rect 2940 10770 2996 10780
rect 3276 10836 3332 10846
rect 2604 10610 2660 10622
rect 2604 10558 2606 10610
rect 2658 10558 2660 10610
rect 2268 10388 2324 10398
rect 2268 10386 2436 10388
rect 2268 10334 2270 10386
rect 2322 10334 2436 10386
rect 2268 10332 2436 10334
rect 2268 10322 2324 10332
rect 2380 9938 2436 10332
rect 2604 10052 2660 10558
rect 3276 10610 3332 10780
rect 3276 10558 3278 10610
rect 3330 10558 3332 10610
rect 3276 10546 3332 10558
rect 2604 9986 2660 9996
rect 2380 9886 2382 9938
rect 2434 9886 2436 9938
rect 2380 9874 2436 9886
rect 1596 9826 1764 9828
rect 1596 9774 1598 9826
rect 1650 9774 1764 9826
rect 1596 9772 1764 9774
rect 1596 9042 1652 9772
rect 1596 8990 1598 9042
rect 1650 8990 1652 9042
rect 1596 8708 1652 8990
rect 2380 8932 2436 8942
rect 3556 8932 3612 8942
rect 2380 8930 2660 8932
rect 2380 8878 2382 8930
rect 2434 8878 2660 8930
rect 2380 8876 2660 8878
rect 2380 8866 2436 8876
rect 1596 8642 1652 8652
rect 2604 8484 2660 8876
rect 3556 8708 3612 8876
rect 2716 8484 2772 8494
rect 2604 8482 2772 8484
rect 2604 8430 2718 8482
rect 2770 8430 2772 8482
rect 2604 8428 2772 8430
rect 2716 8418 2772 8428
rect 3052 8484 3108 8494
rect 3052 8258 3108 8428
rect 3556 8372 3612 8652
rect 3052 8206 3054 8258
rect 3106 8206 3108 8258
rect 3052 8194 3108 8206
rect 3276 8370 3612 8372
rect 3276 8318 3558 8370
rect 3610 8318 3612 8370
rect 3276 8316 3612 8318
rect 28 8082 84 8092
rect 3276 7474 3332 8316
rect 3556 8306 3612 8316
rect 3836 8260 3892 8270
rect 3836 8166 3892 8204
rect 3276 7422 3278 7474
rect 3330 7422 3332 7474
rect 3276 7410 3332 7422
rect 3948 6692 4004 11676
rect 5124 11620 5180 11630
rect 5124 11506 5180 11564
rect 5124 11454 5126 11506
rect 5178 11454 5180 11506
rect 5124 11442 5180 11454
rect 4508 11396 4564 11406
rect 4508 11302 4564 11340
rect 4396 11284 4452 11294
rect 4396 10836 4452 11228
rect 5292 11172 5348 11788
rect 4060 10780 4452 10836
rect 4060 8214 4116 10780
rect 4396 10654 4452 10780
rect 5068 10836 5124 10846
rect 5068 10778 5124 10780
rect 5068 10726 5070 10778
rect 5122 10726 5124 10778
rect 5068 10714 5124 10726
rect 4172 10612 4228 10622
rect 4172 10610 4340 10612
rect 4172 10558 4174 10610
rect 4226 10558 4340 10610
rect 4396 10602 4398 10654
rect 4450 10602 4452 10654
rect 5180 10637 5236 10649
rect 4396 10590 4452 10602
rect 4844 10610 4900 10622
rect 4172 10556 4340 10558
rect 4172 10546 4228 10556
rect 4284 9828 4340 10556
rect 4844 10558 4846 10610
rect 4898 10558 4900 10610
rect 4508 10500 4564 10510
rect 4508 10406 4564 10444
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4284 9734 4340 9772
rect 4396 9716 4452 9726
rect 4284 9044 4340 9054
rect 4172 9042 4340 9044
rect 4172 8990 4286 9042
rect 4338 8990 4340 9042
rect 4172 8988 4340 8990
rect 4172 8372 4228 8988
rect 4284 8978 4340 8988
rect 4396 8820 4452 9660
rect 4844 9604 4900 10558
rect 5180 10585 5182 10637
rect 5234 10585 5236 10637
rect 5180 10500 5236 10585
rect 5180 10434 5236 10444
rect 5180 9828 5236 9838
rect 5292 9828 5348 11116
rect 5516 11508 5572 11518
rect 5516 10610 5572 11452
rect 6076 11506 6132 12854
rect 6412 12516 6468 15092
rect 6524 14980 6580 15277
rect 6636 15202 6692 16046
rect 6636 15150 6638 15202
rect 6690 15150 6692 15202
rect 6636 15138 6692 15150
rect 6860 15148 6916 16492
rect 7196 16212 7252 16222
rect 7196 16118 7252 16156
rect 7644 16098 7700 16716
rect 7868 16706 7924 16716
rect 8316 16436 8372 17052
rect 8652 16884 8708 17836
rect 8764 17108 8820 18956
rect 9212 18340 9268 19740
rect 9324 19234 9380 20860
rect 9660 20802 9716 21532
rect 9660 20750 9662 20802
rect 9714 20750 9716 20802
rect 9660 20018 9716 20750
rect 9884 20802 9940 22316
rect 9884 20750 9886 20802
rect 9938 20750 9940 20802
rect 9884 20738 9940 20750
rect 9996 20802 10052 20814
rect 9996 20750 9998 20802
rect 10050 20750 10052 20802
rect 9660 19966 9662 20018
rect 9714 19966 9716 20018
rect 9324 19182 9326 19234
rect 9378 19182 9380 19234
rect 9324 19170 9380 19182
rect 9436 19236 9492 19246
rect 9660 19236 9716 19966
rect 9436 19234 9716 19236
rect 9436 19182 9438 19234
rect 9490 19182 9716 19234
rect 9436 19180 9716 19182
rect 9996 19908 10052 20750
rect 10162 20746 10218 20758
rect 10162 20694 10164 20746
rect 10216 20694 10218 20746
rect 10162 20244 10218 20694
rect 10108 20188 10218 20244
rect 10108 20132 10164 20188
rect 10108 20066 10164 20076
rect 9436 18452 9492 19180
rect 9996 19012 10052 19852
rect 9996 18946 10052 18956
rect 10220 19234 10276 19246
rect 10220 19182 10222 19234
rect 10274 19182 10276 19234
rect 9772 18452 9828 18462
rect 9436 18450 9828 18452
rect 9436 18398 9774 18450
rect 9826 18398 9828 18450
rect 9436 18396 9828 18398
rect 9772 18340 9828 18396
rect 9212 18284 9716 18340
rect 9772 18284 10164 18340
rect 9212 17892 9268 17902
rect 8764 17042 8820 17052
rect 9100 17554 9156 17566
rect 9100 17502 9102 17554
rect 9154 17502 9156 17554
rect 8764 16884 8820 16894
rect 8988 16884 9044 16894
rect 9100 16884 9156 17502
rect 8652 16882 8820 16884
rect 8652 16830 8766 16882
rect 8818 16830 8820 16882
rect 8652 16828 8820 16830
rect 8764 16818 8820 16828
rect 8876 16882 9156 16884
rect 8876 16830 8990 16882
rect 9042 16830 9156 16882
rect 8876 16828 9156 16830
rect 8484 16660 8540 16670
rect 8484 16658 8708 16660
rect 8484 16606 8486 16658
rect 8538 16606 8708 16658
rect 8484 16604 8708 16606
rect 8484 16594 8540 16604
rect 8316 16380 8484 16436
rect 7308 16054 7364 16066
rect 7308 16002 7310 16054
rect 7362 16002 7364 16054
rect 6972 15876 7028 15886
rect 6972 15316 7028 15820
rect 7308 15876 7364 16002
rect 7308 15810 7364 15820
rect 7644 16046 7646 16098
rect 7698 16046 7700 16098
rect 7140 15652 7196 15662
rect 7644 15652 7700 16046
rect 8316 16210 8372 16222
rect 8316 16158 8318 16210
rect 8370 16158 8372 16210
rect 7140 15538 7196 15596
rect 7140 15486 7142 15538
rect 7194 15486 7196 15538
rect 7140 15474 7196 15486
rect 7308 15596 7700 15652
rect 8204 15652 8260 15662
rect 6972 15260 7252 15316
rect 6860 15092 7028 15148
rect 6524 14914 6580 14924
rect 6524 14532 6580 14542
rect 6524 14438 6580 14476
rect 6804 14474 6860 14486
rect 6804 14422 6806 14474
rect 6858 14422 6860 14474
rect 6804 14420 6860 14422
rect 6636 14362 6692 14374
rect 6636 14310 6638 14362
rect 6690 14310 6692 14362
rect 6524 13748 6580 13758
rect 6636 13748 6692 14310
rect 6524 13746 6692 13748
rect 6524 13694 6526 13746
rect 6578 13694 6692 13746
rect 6524 13692 6692 13694
rect 6748 14364 6860 14420
rect 6524 13682 6580 13692
rect 6412 12450 6468 12460
rect 6748 13524 6804 14364
rect 6972 14196 7028 15092
rect 6972 14130 7028 14140
rect 7196 13972 7252 15260
rect 7308 15314 7364 15596
rect 7308 15262 7310 15314
rect 7362 15262 7364 15314
rect 7308 15250 7364 15262
rect 7420 15316 7476 15326
rect 7420 15222 7476 15260
rect 7756 15316 7812 15326
rect 7756 15222 7812 15260
rect 8204 15314 8260 15596
rect 8316 15540 8372 16158
rect 8428 16083 8484 16380
rect 8428 16031 8430 16083
rect 8482 16031 8484 16083
rect 8428 16019 8484 16031
rect 8316 15474 8372 15484
rect 8204 15262 8206 15314
rect 8258 15262 8260 15314
rect 8204 15250 8260 15262
rect 8316 15316 8372 15326
rect 8092 15204 8148 15214
rect 8092 14530 8148 15148
rect 8092 14478 8094 14530
rect 8146 14478 8148 14530
rect 7756 14306 7812 14318
rect 7756 14254 7758 14306
rect 7810 14254 7812 14306
rect 7756 13972 7812 14254
rect 6636 12292 6692 12302
rect 6636 12198 6692 12236
rect 6076 11454 6078 11506
rect 6130 11454 6132 11506
rect 6076 11442 6132 11454
rect 6188 11620 6244 11630
rect 5628 11396 5684 11406
rect 5628 11302 5684 11340
rect 5964 11350 6020 11362
rect 5964 11298 5966 11350
rect 6018 11298 6020 11350
rect 5964 11284 6020 11298
rect 5964 11218 6020 11228
rect 5516 10558 5518 10610
rect 5570 10558 5572 10610
rect 5516 10546 5572 10558
rect 6188 10610 6244 11564
rect 6412 11396 6468 11406
rect 6412 11302 6468 11340
rect 6748 11379 6804 13468
rect 7084 13916 7812 13972
rect 6860 13412 6916 13422
rect 6860 13074 6916 13356
rect 6860 13022 6862 13074
rect 6914 13022 6916 13074
rect 6860 13010 6916 13022
rect 6972 12918 7028 12930
rect 6972 12866 6974 12918
rect 7026 12866 7028 12918
rect 6972 12852 7028 12866
rect 6972 12786 7028 12796
rect 6860 11508 6916 11518
rect 6860 11414 6916 11452
rect 6748 11327 6750 11379
rect 6802 11327 6804 11379
rect 6748 11315 6804 11327
rect 6188 10558 6190 10610
rect 6242 10558 6244 10610
rect 6188 10546 6244 10558
rect 6860 11284 6916 11294
rect 5740 10052 5796 10062
rect 6860 10052 6916 11228
rect 6972 10500 7028 10510
rect 6972 10406 7028 10444
rect 6860 9996 7028 10052
rect 5180 9826 5348 9828
rect 5180 9774 5182 9826
rect 5234 9774 5348 9826
rect 5180 9772 5348 9774
rect 5628 9826 5684 9838
rect 5628 9774 5630 9826
rect 5682 9774 5684 9826
rect 5180 9762 5236 9772
rect 4844 9510 4900 9548
rect 5628 9604 5684 9774
rect 5740 9658 5796 9996
rect 6300 9940 6356 9950
rect 6300 9826 6356 9884
rect 5740 9606 5742 9658
rect 5794 9606 5796 9658
rect 5964 9770 6020 9782
rect 5964 9718 5966 9770
rect 6018 9718 6020 9770
rect 6300 9774 6302 9826
rect 6354 9774 6356 9826
rect 6300 9762 6356 9774
rect 6860 9828 6916 9838
rect 6860 9734 6916 9772
rect 5964 9716 6020 9718
rect 5964 9650 6020 9660
rect 6748 9716 6804 9726
rect 5740 9594 5796 9606
rect 5460 9098 5516 9110
rect 5292 9044 5348 9054
rect 5460 9046 5462 9098
rect 5514 9046 5516 9098
rect 5460 9044 5516 9046
rect 5292 8950 5348 8988
rect 5404 8988 5516 9044
rect 5628 9044 5684 9548
rect 4900 8932 4956 8942
rect 4900 8838 4956 8876
rect 5404 8820 5460 8988
rect 4340 8764 4452 8820
rect 5068 8764 5460 8820
rect 4340 8708 4396 8764
rect 4172 8306 4228 8316
rect 4284 8652 4396 8708
rect 4956 8708 5012 8718
rect 4476 8652 4740 8662
rect 4284 8370 4340 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4284 8318 4286 8370
rect 4338 8318 4340 8370
rect 4284 8306 4340 8318
rect 4620 8260 4676 8270
rect 4060 8202 4172 8214
rect 4060 8150 4118 8202
rect 4170 8150 4172 8202
rect 4620 8166 4676 8204
rect 4956 8243 5012 8652
rect 5068 8370 5124 8764
rect 5068 8318 5070 8370
rect 5122 8318 5124 8370
rect 5068 8306 5124 8318
rect 4956 8191 4958 8243
rect 5010 8191 5012 8243
rect 5628 8258 5684 8988
rect 5740 9210 5796 9222
rect 5740 9158 5742 9210
rect 5794 9158 5796 9210
rect 5740 8484 5796 9158
rect 6748 9086 6804 9660
rect 5852 9042 5908 9054
rect 6412 9044 6468 9054
rect 5852 8990 5854 9042
rect 5906 8990 5908 9042
rect 5852 8932 5908 8990
rect 5852 8866 5908 8876
rect 5964 9042 6468 9044
rect 5964 8990 6414 9042
rect 6466 8990 6468 9042
rect 6748 9034 6750 9086
rect 6802 9034 6804 9086
rect 6748 9022 6804 9034
rect 5964 8988 6468 8990
rect 5740 8418 5796 8428
rect 5628 8206 5630 8258
rect 5682 8206 5684 8258
rect 5628 8194 5684 8206
rect 4956 8179 5012 8191
rect 4060 8092 4172 8150
rect 5740 8090 5796 8102
rect 5740 8038 5742 8090
rect 5794 8038 5796 8090
rect 5180 7700 5236 7710
rect 4060 7362 4116 7374
rect 4060 7310 4062 7362
rect 4114 7310 4116 7362
rect 4060 6916 4116 7310
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4172 6916 4228 6926
rect 4060 6914 4228 6916
rect 4060 6862 4174 6914
rect 4226 6862 4228 6914
rect 4060 6860 4228 6862
rect 4172 6850 4228 6860
rect 4508 6916 4564 6926
rect 3948 6626 4004 6636
rect 4508 6690 4564 6860
rect 4508 6638 4510 6690
rect 4562 6638 4564 6690
rect 4508 6626 4564 6638
rect 4956 6692 5012 6702
rect 4844 6468 4900 6478
rect 4844 6374 4900 6412
rect 4844 5908 4900 5918
rect 4956 5908 5012 6636
rect 5180 6690 5236 7644
rect 5740 6916 5796 8038
rect 5740 6850 5796 6860
rect 5964 7586 6020 8988
rect 6412 8978 6468 8988
rect 6860 8932 6916 8942
rect 6860 8838 6916 8876
rect 6076 8372 6132 8382
rect 6076 8219 6132 8316
rect 6860 8372 6916 8382
rect 6860 8278 6916 8316
rect 6076 8167 6078 8219
rect 6130 8167 6132 8219
rect 6076 8155 6132 8167
rect 6300 8258 6356 8270
rect 6300 8206 6302 8258
rect 6354 8206 6356 8258
rect 5964 7534 5966 7586
rect 6018 7534 6020 7586
rect 5180 6638 5182 6690
rect 5234 6638 5236 6690
rect 5180 6626 5236 6638
rect 5796 6692 5852 6702
rect 5964 6692 6020 7534
rect 6300 6804 6356 8206
rect 6748 8260 6804 8270
rect 6748 7518 6804 8204
rect 6972 8243 7028 9996
rect 7084 8708 7140 13916
rect 7756 13748 7812 13758
rect 8092 13748 8148 14478
rect 8316 14420 8372 15260
rect 8484 15314 8540 15326
rect 8484 15262 8486 15314
rect 8538 15262 8540 15314
rect 8484 15148 8540 15262
rect 8484 15092 8596 15148
rect 8540 14868 8596 15092
rect 8540 14802 8596 14812
rect 8316 14354 8372 14364
rect 8428 14308 8484 14318
rect 8428 14214 8484 14252
rect 8652 13972 8708 16604
rect 8764 16100 8820 16110
rect 8876 16100 8932 16828
rect 8988 16818 9044 16828
rect 8764 16098 8932 16100
rect 8764 16046 8766 16098
rect 8818 16046 8932 16098
rect 8764 16044 8932 16046
rect 8764 16034 8820 16044
rect 8876 15316 8932 15326
rect 8876 15202 8932 15260
rect 8876 15150 8878 15202
rect 8930 15150 8932 15202
rect 8876 15138 8932 15150
rect 9212 15148 9268 17836
rect 9660 17890 9716 18284
rect 9660 17838 9662 17890
rect 9714 17838 9716 17890
rect 9660 17826 9716 17838
rect 9996 18116 10052 18126
rect 9996 17666 10052 18060
rect 9996 17614 9998 17666
rect 10050 17614 10052 17666
rect 9436 17108 9492 17118
rect 9324 16884 9380 16894
rect 9324 16098 9380 16828
rect 9436 16882 9492 17052
rect 9996 16996 10052 17614
rect 9996 16930 10052 16940
rect 10108 17668 10164 18284
rect 10220 18004 10276 19182
rect 10220 17938 10276 17948
rect 9436 16830 9438 16882
rect 9490 16830 9492 16882
rect 9436 16818 9492 16830
rect 10108 16884 10164 17612
rect 10108 16818 10164 16828
rect 10220 16770 10276 16782
rect 10220 16718 10222 16770
rect 10274 16718 10276 16770
rect 10108 16100 10164 16110
rect 9324 16046 9326 16098
rect 9378 16046 9380 16098
rect 9324 16034 9380 16046
rect 9660 16098 10164 16100
rect 9660 16046 10110 16098
rect 10162 16046 10164 16098
rect 9660 16044 10164 16046
rect 9660 15426 9716 16044
rect 10108 16034 10164 16044
rect 9660 15374 9662 15426
rect 9714 15374 9716 15426
rect 9660 15362 9716 15374
rect 10108 15342 10164 15354
rect 9492 15316 9548 15326
rect 9492 15222 9548 15260
rect 10108 15290 10110 15342
rect 10162 15290 10164 15342
rect 9660 15204 9716 15214
rect 9212 15092 9380 15148
rect 8764 14868 8820 14878
rect 8764 14530 8820 14812
rect 8764 14478 8766 14530
rect 8818 14478 8820 14530
rect 8764 14466 8820 14478
rect 9100 14474 9156 14486
rect 7756 13746 8148 13748
rect 7756 13694 7758 13746
rect 7810 13694 8148 13746
rect 7756 13692 8148 13694
rect 8428 13916 8708 13972
rect 9100 14422 9102 14474
rect 9154 14422 9156 14474
rect 8428 13746 8484 13916
rect 8428 13694 8430 13746
rect 8482 13694 8484 13746
rect 7756 13682 7812 13692
rect 7420 13524 7476 13534
rect 7420 13430 7476 13468
rect 7980 13524 8036 13534
rect 7196 12964 7252 12974
rect 7644 12964 7700 12974
rect 7196 12962 7700 12964
rect 7196 12910 7198 12962
rect 7250 12910 7646 12962
rect 7698 12910 7700 12962
rect 7196 12908 7700 12910
rect 7196 12292 7252 12908
rect 7644 12898 7700 12908
rect 7980 12947 8036 13468
rect 8092 13522 8148 13534
rect 8092 13470 8094 13522
rect 8146 13470 8148 13522
rect 8092 13412 8148 13470
rect 8092 13346 8148 13356
rect 8092 13076 8148 13086
rect 8092 12982 8148 13020
rect 8428 12964 8484 13694
rect 7980 12895 7982 12947
rect 8034 12895 8036 12947
rect 7980 12883 8036 12895
rect 8204 12962 8484 12964
rect 8204 12910 8430 12962
rect 8482 12910 8484 12962
rect 8204 12908 8484 12910
rect 7196 12226 7252 12236
rect 8092 12180 8148 12190
rect 8204 12180 8260 12908
rect 8428 12898 8484 12908
rect 8540 13748 8596 13758
rect 8092 12178 8260 12180
rect 8092 12126 8094 12178
rect 8146 12126 8260 12178
rect 8092 12124 8260 12126
rect 8428 12740 8484 12750
rect 8540 12740 8596 13692
rect 8876 13636 8932 13646
rect 8876 13542 8932 13580
rect 9100 13524 9156 14422
rect 9100 13458 9156 13468
rect 8484 12684 8596 12740
rect 8652 13412 8708 13422
rect 8652 12852 8708 13356
rect 8092 12114 8148 12124
rect 7252 12066 7308 12078
rect 7252 12014 7254 12066
rect 7306 12014 7308 12066
rect 7252 11844 7308 12014
rect 7252 11778 7308 11788
rect 7756 11954 7812 11966
rect 7756 11902 7758 11954
rect 7810 11902 7812 11954
rect 7532 11394 7588 11406
rect 7532 11342 7534 11394
rect 7586 11342 7588 11394
rect 7532 11172 7588 11342
rect 7756 11284 7812 11902
rect 7868 11396 7924 11406
rect 7868 11302 7924 11340
rect 8316 11396 8372 11406
rect 7756 11218 7812 11228
rect 7532 11106 7588 11116
rect 8204 10500 8260 10510
rect 8204 10050 8260 10444
rect 8204 9998 8206 10050
rect 8258 9998 8260 10050
rect 8204 9986 8260 9998
rect 7308 9940 7364 9950
rect 7308 9846 7364 9884
rect 7084 8642 7140 8652
rect 7196 9782 7252 9794
rect 7196 9730 7198 9782
rect 7250 9730 7252 9782
rect 7196 8484 7252 9730
rect 7420 9057 7476 9069
rect 7420 9005 7422 9057
rect 7474 9005 7476 9057
rect 7308 8932 7364 8942
rect 7308 8838 7364 8876
rect 7420 8708 7476 9005
rect 7420 8642 7476 8652
rect 7756 9042 7812 9054
rect 7756 8990 7758 9042
rect 7810 8990 7812 9042
rect 7196 8428 7364 8484
rect 7308 8372 7364 8428
rect 7308 8306 7364 8316
rect 6972 8191 6974 8243
rect 7026 8191 7028 8243
rect 6972 8179 7028 8191
rect 7196 8258 7252 8270
rect 7196 8206 7198 8258
rect 7250 8206 7252 8258
rect 6748 7466 6750 7518
rect 6802 7466 6804 7518
rect 6748 7252 6804 7466
rect 6972 7642 7028 7654
rect 6972 7590 6974 7642
rect 7026 7590 7028 7642
rect 6972 7476 7028 7590
rect 6972 7410 7028 7420
rect 7084 7476 7140 7486
rect 7196 7476 7252 8206
rect 7756 8260 7812 8990
rect 8204 9044 8260 9054
rect 8316 9044 8372 11340
rect 8428 9604 8484 12684
rect 8652 12193 8708 12796
rect 8764 12740 8820 12750
rect 8764 12646 8820 12684
rect 8652 12141 8654 12193
rect 8706 12141 8708 12193
rect 8540 12066 8596 12078
rect 8540 12014 8542 12066
rect 8594 12014 8596 12066
rect 8540 11394 8596 12014
rect 8540 11342 8542 11394
rect 8594 11342 8596 11394
rect 8540 11330 8596 11342
rect 8540 11226 8596 11238
rect 8540 11174 8542 11226
rect 8594 11174 8596 11226
rect 8540 9826 8596 11174
rect 8540 9774 8542 9826
rect 8594 9774 8596 9826
rect 8540 9762 8596 9774
rect 8652 9716 8708 12141
rect 8988 12180 9044 12190
rect 8988 12086 9044 12124
rect 9324 11956 9380 15092
rect 9436 15092 9492 15102
rect 9436 14530 9492 15036
rect 9436 14478 9438 14530
rect 9490 14478 9492 14530
rect 9436 14466 9492 14478
rect 9548 14980 9604 14990
rect 9548 13636 9604 14924
rect 9660 14642 9716 15148
rect 10108 14980 10164 15290
rect 10220 15204 10276 16718
rect 10332 15428 10388 25452
rect 10892 25396 10948 25406
rect 10780 25172 10836 25182
rect 10780 24722 10836 25116
rect 10780 24670 10782 24722
rect 10834 24670 10836 24722
rect 10780 24658 10836 24670
rect 10892 24554 10948 25340
rect 11116 24948 11172 26238
rect 11228 26290 11284 26852
rect 11228 26238 11230 26290
rect 11282 26238 11284 26290
rect 11228 26226 11284 26238
rect 11340 26292 11396 26302
rect 11116 24882 11172 24892
rect 11004 24724 11060 24734
rect 11340 24724 11396 26236
rect 11452 26290 11508 26908
rect 11676 26898 11732 26908
rect 11788 28642 11956 28644
rect 11788 28590 11902 28642
rect 11954 28590 11956 28642
rect 11788 28588 11956 28590
rect 11788 26740 11844 28588
rect 11900 28578 11956 28588
rect 12012 28196 12068 29036
rect 12236 28868 12292 29374
rect 12236 28802 12292 28812
rect 12348 29428 12404 29438
rect 12180 28642 12236 28654
rect 12180 28590 12182 28642
rect 12234 28590 12236 28642
rect 12180 28420 12236 28590
rect 12180 28354 12236 28364
rect 12012 28140 12180 28196
rect 11788 26674 11844 26684
rect 11900 28084 11956 28094
rect 11676 26628 11732 26638
rect 11676 26516 11732 26572
rect 11676 26460 11788 26516
rect 11732 26402 11788 26460
rect 11732 26350 11734 26402
rect 11786 26350 11788 26402
rect 11732 26338 11788 26350
rect 11452 26238 11454 26290
rect 11506 26238 11508 26290
rect 11452 25452 11508 26238
rect 11452 25450 11620 25452
rect 11452 25398 11454 25450
rect 11506 25398 11620 25450
rect 11452 25396 11620 25398
rect 11452 25386 11508 25396
rect 11452 24724 11508 24734
rect 11004 24722 11172 24724
rect 11004 24670 11006 24722
rect 11058 24670 11172 24722
rect 11004 24668 11172 24670
rect 11004 24658 11060 24668
rect 10892 24502 10894 24554
rect 10946 24502 10948 24554
rect 10892 24490 10948 24502
rect 11116 23938 11172 24668
rect 11116 23886 11118 23938
rect 11170 23886 11172 23938
rect 11116 23380 11172 23886
rect 11340 24722 11508 24724
rect 11340 24670 11454 24722
rect 11506 24670 11508 24722
rect 11340 24668 11508 24670
rect 11340 23940 11396 24668
rect 11452 24658 11508 24668
rect 11564 24724 11620 25396
rect 11900 25338 11956 28028
rect 12012 27897 12068 27909
rect 12012 27860 12014 27897
rect 12066 27860 12068 27897
rect 12012 27794 12068 27804
rect 12124 27412 12180 28140
rect 12124 27346 12180 27356
rect 12348 26628 12404 29372
rect 12460 27860 12516 29820
rect 12796 29482 12852 30156
rect 12908 30146 12964 30156
rect 13244 29652 13300 30940
rect 13356 30930 13412 30940
rect 13804 30660 13860 31276
rect 14252 31220 14308 31726
rect 14476 31780 14532 31790
rect 14476 31686 14532 31724
rect 14588 31332 14644 32549
rect 14868 32506 14924 32518
rect 14868 32454 14870 32506
rect 14922 32454 14924 32506
rect 14868 32004 14924 32454
rect 14868 31938 14924 31948
rect 14588 31266 14644 31276
rect 13916 31164 14308 31220
rect 15036 31220 15092 32620
rect 15148 32674 15204 33628
rect 15820 33572 15876 33582
rect 15820 33514 15876 33516
rect 15820 33462 15822 33514
rect 15874 33462 15876 33514
rect 15820 33450 15876 33462
rect 15708 33348 15764 33358
rect 15708 33254 15764 33292
rect 16044 33012 16100 34862
rect 15148 32622 15150 32674
rect 15202 32622 15204 32674
rect 15148 32610 15204 32622
rect 15484 32956 16100 33012
rect 15036 31164 15204 31220
rect 13916 30660 13972 31164
rect 14140 30996 14196 31006
rect 15016 30996 15072 31006
rect 14140 30902 14196 30940
rect 14812 30994 15072 30996
rect 14812 30942 15018 30994
rect 15070 30942 15072 30994
rect 14812 30940 15072 30942
rect 13916 30604 14196 30660
rect 13804 30594 13860 30604
rect 13468 30212 13524 30222
rect 13468 30118 13524 30156
rect 13244 29586 13300 29596
rect 13356 30100 13412 30110
rect 12796 29430 12798 29482
rect 12850 29430 12852 29482
rect 12796 29428 12852 29430
rect 12796 29362 12852 29372
rect 12684 29092 12740 29102
rect 12684 28866 12740 29036
rect 12684 28814 12686 28866
rect 12738 28814 12740 28866
rect 12684 28802 12740 28814
rect 13020 28644 13076 28654
rect 13020 28642 13300 28644
rect 13020 28590 13022 28642
rect 13074 28590 13300 28642
rect 13020 28588 13300 28590
rect 13020 28578 13076 28588
rect 13020 27886 13076 27898
rect 12684 27860 12740 27870
rect 12460 27794 12516 27804
rect 12572 27804 12684 27860
rect 12460 27242 12516 27254
rect 12460 27190 12462 27242
rect 12514 27190 12516 27242
rect 12460 27076 12516 27190
rect 12460 27010 12516 27020
rect 12572 27074 12628 27804
rect 12684 27794 12740 27804
rect 13020 27860 13022 27886
rect 13074 27860 13076 27886
rect 13020 27794 13076 27804
rect 13244 27858 13300 28588
rect 13244 27806 13246 27858
rect 13298 27806 13300 27858
rect 13244 27188 13300 27806
rect 12572 27022 12574 27074
rect 12626 27022 12628 27074
rect 12572 27010 12628 27022
rect 12908 27132 13300 27188
rect 12908 27074 12964 27132
rect 12908 27022 12910 27074
rect 12962 27022 12964 27074
rect 12908 27010 12964 27022
rect 13244 27076 13300 27132
rect 13244 27010 13300 27020
rect 13356 26908 13412 30044
rect 13804 29482 13860 29494
rect 13804 29430 13806 29482
rect 13858 29430 13860 29482
rect 13804 28868 13860 29430
rect 14140 29092 14196 30604
rect 14812 30548 14868 30940
rect 15016 30930 15072 30940
rect 15148 30772 15204 31164
rect 14588 30492 14868 30548
rect 14924 30716 15204 30772
rect 15260 30770 15316 30782
rect 15260 30718 15262 30770
rect 15314 30718 15316 30770
rect 14588 30434 14644 30492
rect 14588 30382 14590 30434
rect 14642 30382 14644 30434
rect 14588 30370 14644 30382
rect 14344 30212 14400 30222
rect 14344 30118 14400 30156
rect 14140 29026 14196 29036
rect 14252 29988 14308 29998
rect 14924 29988 14980 30716
rect 15260 30436 15316 30718
rect 15260 30370 15316 30380
rect 15484 30660 15540 32956
rect 13804 28812 14196 28868
rect 14028 28642 14084 28654
rect 13636 28586 13692 28598
rect 13636 28534 13638 28586
rect 13690 28534 13692 28586
rect 14028 28590 14030 28642
rect 14082 28590 14084 28642
rect 13468 27972 13524 27982
rect 13468 27878 13524 27916
rect 13636 27914 13692 28534
rect 13636 27862 13638 27914
rect 13690 27862 13692 27914
rect 13804 28530 13860 28542
rect 13804 28478 13806 28530
rect 13858 28478 13860 28530
rect 13804 27972 13860 28478
rect 14028 28532 14084 28590
rect 14028 28466 14084 28476
rect 13804 27906 13860 27916
rect 13636 27300 13692 27862
rect 14028 27896 14084 27908
rect 14028 27860 14030 27896
rect 14082 27860 14084 27896
rect 14028 27794 14084 27804
rect 14140 27748 14196 28812
rect 14140 27682 14196 27692
rect 14252 27524 14308 29932
rect 14364 29932 14980 29988
rect 15036 30212 15092 30222
rect 14364 29314 14420 29932
rect 15036 29652 15092 30156
rect 15484 29652 15540 30604
rect 15036 29596 15316 29652
rect 14750 29451 14806 29463
rect 14364 29262 14366 29314
rect 14418 29262 14420 29314
rect 14364 29250 14420 29262
rect 14588 29428 14644 29438
rect 14750 29399 14752 29451
rect 14804 29428 14806 29451
rect 14924 29428 14980 29438
rect 14804 29399 14812 29428
rect 14750 29372 14812 29399
rect 14364 28644 14420 28654
rect 14364 28552 14366 28588
rect 14418 28552 14420 28588
rect 14364 28540 14420 28552
rect 14476 27972 14532 27982
rect 14364 27858 14420 27870
rect 14364 27806 14366 27858
rect 14418 27806 14420 27858
rect 14364 27636 14420 27806
rect 14476 27748 14532 27916
rect 14588 27970 14644 29372
rect 14756 28822 14812 29372
rect 14924 29334 14980 29372
rect 15036 29426 15092 29438
rect 15036 29374 15038 29426
rect 15090 29374 15092 29426
rect 15036 29092 15092 29374
rect 15036 29026 15092 29036
rect 14756 28810 14868 28822
rect 14756 28758 14814 28810
rect 14866 28758 14868 28810
rect 14756 28756 14868 28758
rect 14812 28746 14868 28756
rect 14588 27918 14590 27970
rect 14642 27918 14644 27970
rect 14588 27906 14644 27918
rect 14924 28642 14980 28654
rect 15148 28644 15204 28654
rect 14924 28590 14926 28642
rect 14978 28590 14980 28642
rect 14756 27860 14812 27870
rect 14756 27766 14812 27804
rect 14476 27692 14644 27748
rect 14364 27570 14420 27580
rect 13636 27234 13692 27244
rect 14028 27468 14308 27524
rect 12348 26562 12404 26572
rect 13132 26852 13412 26908
rect 13468 27076 13524 27086
rect 12292 26319 12348 26331
rect 12292 26267 12294 26319
rect 12346 26292 12348 26319
rect 12840 26328 12896 26340
rect 12460 26292 12516 26302
rect 12346 26267 12404 26292
rect 12292 26236 12404 26267
rect 12124 26180 12180 26190
rect 12124 26086 12180 26124
rect 11900 25286 11902 25338
rect 11954 25286 11956 25338
rect 11900 25274 11956 25286
rect 12012 25732 12068 25742
rect 11452 24164 11508 24174
rect 11564 24164 11620 24668
rect 11452 24162 11620 24164
rect 11452 24110 11454 24162
rect 11506 24110 11620 24162
rect 11452 24108 11620 24110
rect 11676 25172 11732 25182
rect 11452 24098 11508 24108
rect 11340 23884 11508 23940
rect 11116 23324 11396 23380
rect 11228 22708 11284 22718
rect 11228 22594 11284 22652
rect 11228 22542 11230 22594
rect 11282 22542 11284 22594
rect 11228 22530 11284 22542
rect 10892 22370 10948 22382
rect 10892 22318 10894 22370
rect 10946 22318 10948 22370
rect 10556 22146 10612 22158
rect 10556 22094 10558 22146
rect 10610 22094 10612 22146
rect 10444 21588 10500 21598
rect 10556 21588 10612 22094
rect 10892 21812 10948 22318
rect 11340 22148 11396 23324
rect 11452 22148 11508 23884
rect 11676 23604 11732 25116
rect 11788 24948 11844 24958
rect 11788 24722 11844 24892
rect 11788 24670 11790 24722
rect 11842 24670 11844 24722
rect 11788 24658 11844 24670
rect 12012 24174 12068 25676
rect 12236 25620 12292 25630
rect 12124 25452 12180 25462
rect 12236 25452 12292 25564
rect 12124 25450 12292 25452
rect 12124 25398 12126 25450
rect 12178 25398 12292 25450
rect 12124 25396 12292 25398
rect 12348 25452 12404 26236
rect 12460 26198 12516 26236
rect 12840 26292 12842 26328
rect 12894 26292 12896 26328
rect 12840 26226 12896 26236
rect 13132 25732 13188 26852
rect 13468 26122 13524 27020
rect 13860 27076 13916 27114
rect 13860 27010 13916 27020
rect 14028 26908 14084 27468
rect 14420 27188 14476 27198
rect 14420 27130 14476 27132
rect 14140 27076 14196 27086
rect 14140 26982 14196 27020
rect 14420 27078 14422 27130
rect 14474 27078 14476 27130
rect 13916 26852 14084 26908
rect 14252 26964 14308 27002
rect 14420 26908 14476 27078
rect 14588 27074 14644 27692
rect 14924 27636 14980 28590
rect 15036 28642 15204 28644
rect 15036 28590 15150 28642
rect 15202 28590 15204 28642
rect 15036 28588 15204 28590
rect 15036 28532 15092 28588
rect 15148 28578 15204 28588
rect 15036 27748 15092 28476
rect 15148 28420 15204 28430
rect 15148 27858 15204 28364
rect 15260 28308 15316 29596
rect 15484 29586 15540 29596
rect 15596 32788 15652 32798
rect 15372 29426 15428 29438
rect 15372 29374 15374 29426
rect 15426 29374 15428 29426
rect 15372 28868 15428 29374
rect 15484 29428 15540 29438
rect 15596 29428 15652 32732
rect 15951 32788 16007 32798
rect 15951 32618 16007 32732
rect 15951 32566 15953 32618
rect 16005 32566 16007 32618
rect 15951 32554 16007 32566
rect 15708 32338 15764 32350
rect 15708 32286 15710 32338
rect 15762 32286 15764 32338
rect 15708 31892 15764 32286
rect 16156 31892 16212 39228
rect 16604 39060 16660 40350
rect 16268 39058 16660 39060
rect 16268 39006 16606 39058
rect 16658 39006 16660 39058
rect 16268 39004 16660 39006
rect 16268 35252 16324 39004
rect 16604 38994 16660 39004
rect 16716 38668 16772 40796
rect 16828 39842 16884 41580
rect 16828 39790 16830 39842
rect 16882 39790 16884 39842
rect 16828 39778 16884 39790
rect 17164 39618 17220 42028
rect 17612 41972 17668 43148
rect 17724 42754 17780 42766
rect 17724 42702 17726 42754
rect 17778 42702 17780 42754
rect 17724 42644 17780 42702
rect 18004 42756 18060 42766
rect 18004 42662 18060 42700
rect 19180 42756 19236 42766
rect 19180 42754 19348 42756
rect 19180 42702 19182 42754
rect 19234 42702 19348 42754
rect 19180 42700 19348 42702
rect 19180 42690 19236 42700
rect 17724 42578 17780 42588
rect 18844 42532 18900 42542
rect 17500 41970 17668 41972
rect 17500 41918 17614 41970
rect 17666 41918 17668 41970
rect 17500 41916 17668 41918
rect 17500 41188 17556 41916
rect 17612 41906 17668 41916
rect 18396 42530 18900 42532
rect 18396 42478 18846 42530
rect 18898 42478 18900 42530
rect 18396 42476 18900 42478
rect 18396 41970 18452 42476
rect 18844 42466 18900 42476
rect 19292 42196 19348 42700
rect 19404 42308 19460 44044
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 20188 43764 20244 44156
rect 20412 44146 20468 44156
rect 20524 44156 20636 44212
rect 19964 43708 20244 43764
rect 20412 43876 20468 43886
rect 19740 42756 19796 42766
rect 19740 42662 19796 42700
rect 19964 42756 20020 43708
rect 20244 43092 20300 43102
rect 19964 42662 20020 42700
rect 20076 42980 20132 42990
rect 20076 42754 20132 42924
rect 20076 42702 20078 42754
rect 20130 42702 20132 42754
rect 20076 42690 20132 42702
rect 20244 42754 20300 43036
rect 20244 42702 20246 42754
rect 20298 42702 20300 42754
rect 20244 42690 20300 42702
rect 19572 42644 19628 42654
rect 19572 42586 19628 42588
rect 19572 42534 19574 42586
rect 19626 42534 19628 42586
rect 19572 42522 19628 42534
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19404 42252 19684 42308
rect 19836 42298 20100 42308
rect 19292 42140 19572 42196
rect 18396 41918 18398 41970
rect 18450 41918 18452 41970
rect 18396 41906 18452 41918
rect 19516 41524 19572 42140
rect 19516 41458 19572 41468
rect 17500 41122 17556 41132
rect 18620 41186 18676 41198
rect 18620 41134 18622 41186
rect 18674 41134 18676 41186
rect 17836 40964 17892 40974
rect 17612 40628 17668 40638
rect 17612 40534 17668 40572
rect 17276 40404 17332 40414
rect 17276 40310 17332 40348
rect 17556 39732 17612 39742
rect 17556 39638 17612 39676
rect 17164 39566 17166 39618
rect 17218 39566 17220 39618
rect 17164 39554 17220 39566
rect 17836 39618 17892 40908
rect 18620 40628 18676 41134
rect 19404 41188 19460 41198
rect 19404 41094 19460 41132
rect 19628 40628 19684 42252
rect 20412 42196 20468 43820
rect 20524 43764 20580 44156
rect 20636 44146 20692 44156
rect 20972 43988 21028 45054
rect 20524 43698 20580 43708
rect 20636 43932 21028 43988
rect 21196 45106 21252 45118
rect 21196 45054 21198 45106
rect 21250 45054 21252 45106
rect 20524 43540 20580 43550
rect 20524 42644 20580 43484
rect 20636 42978 20692 43932
rect 21196 43876 21252 45054
rect 21756 45108 21812 45118
rect 21308 44884 21364 44894
rect 21308 44294 21364 44828
rect 21476 44884 21532 44894
rect 21476 44882 21700 44884
rect 21476 44830 21478 44882
rect 21530 44830 21700 44882
rect 21476 44828 21700 44830
rect 21476 44818 21532 44828
rect 21308 44242 21310 44294
rect 21362 44242 21364 44294
rect 21308 44230 21364 44242
rect 21644 43876 21700 44828
rect 21196 43820 21588 43876
rect 20860 43540 20916 43578
rect 20860 43474 20916 43484
rect 20636 42926 20638 42978
rect 20690 42926 20692 42978
rect 20636 42914 20692 42926
rect 21420 42980 21476 42990
rect 20524 42578 20580 42588
rect 20076 42140 20468 42196
rect 19740 41412 19796 41422
rect 19740 41318 19796 41356
rect 20076 41186 20132 42140
rect 20748 41972 20804 41982
rect 20524 41970 20804 41972
rect 20524 41918 20750 41970
rect 20802 41918 20804 41970
rect 20524 41916 20804 41918
rect 20300 41860 20356 41870
rect 20524 41860 20580 41916
rect 20748 41906 20804 41916
rect 20300 41858 20580 41860
rect 20300 41806 20302 41858
rect 20354 41806 20580 41858
rect 20300 41804 20580 41806
rect 20300 41794 20356 41804
rect 20524 41524 20580 41804
rect 20524 41468 21308 41524
rect 20412 41412 20468 41422
rect 20412 41354 20468 41356
rect 20412 41302 20414 41354
rect 20466 41302 20468 41354
rect 20412 41290 20468 41302
rect 20076 41134 20078 41186
rect 20130 41134 20132 41186
rect 20076 41122 20132 41134
rect 20412 41186 20468 41198
rect 20412 41134 20414 41186
rect 20466 41134 20468 41186
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19796 40628 19852 40638
rect 19628 40626 19852 40628
rect 19628 40574 19798 40626
rect 19850 40574 19852 40626
rect 19628 40572 19852 40574
rect 18620 40562 18676 40572
rect 19796 40562 19852 40572
rect 18228 40516 18284 40526
rect 18228 40422 18284 40460
rect 19292 40402 19348 40414
rect 19292 40350 19294 40402
rect 19346 40350 19348 40402
rect 18956 40180 19012 40190
rect 18620 40178 19012 40180
rect 18620 40126 18958 40178
rect 19010 40126 19012 40178
rect 18620 40124 19012 40126
rect 17836 39566 17838 39618
rect 17890 39566 17892 39618
rect 16380 38612 16772 38668
rect 16940 38836 16996 38846
rect 16380 37380 16436 38612
rect 16940 38164 16996 38780
rect 17500 38834 17556 38846
rect 17500 38782 17502 38834
rect 17554 38782 17556 38834
rect 17500 38668 17556 38782
rect 17836 38668 17892 39566
rect 18396 39956 18452 39966
rect 18284 38722 18340 38734
rect 18284 38670 18286 38722
rect 18338 38670 18340 38722
rect 17500 38612 18116 38668
rect 16940 38050 16996 38108
rect 16940 37998 16942 38050
rect 16994 37998 16996 38050
rect 16940 37986 16996 37998
rect 16604 37826 16660 37838
rect 16604 37774 16606 37826
rect 16658 37774 16660 37826
rect 16604 37716 16660 37774
rect 16604 37650 16660 37660
rect 17332 37828 17388 37838
rect 17780 37828 17836 37838
rect 17332 37826 17836 37828
rect 17332 37774 17334 37826
rect 17386 37774 17782 37826
rect 17834 37774 17836 37826
rect 17332 37772 17836 37774
rect 16380 37286 16436 37324
rect 16716 37268 16772 37278
rect 16716 37174 16772 37212
rect 17332 37268 17388 37772
rect 17780 37380 17836 37772
rect 17780 37324 18004 37380
rect 17332 37202 17388 37212
rect 16492 37156 16548 37166
rect 16380 36596 16436 36606
rect 16492 36596 16548 37100
rect 17780 37154 17836 37166
rect 17780 37102 17782 37154
rect 17834 37102 17836 37154
rect 17780 36932 17836 37102
rect 17780 36866 17836 36876
rect 16380 36594 16548 36596
rect 16380 36542 16382 36594
rect 16434 36542 16548 36594
rect 16380 36540 16548 36542
rect 16380 36530 16436 36540
rect 17948 36484 18004 37324
rect 17836 36428 18004 36484
rect 17836 36372 17892 36428
rect 17836 35698 17892 36316
rect 17836 35646 17838 35698
rect 17890 35646 17892 35698
rect 16268 35186 16324 35196
rect 16716 35586 16772 35598
rect 16716 35534 16718 35586
rect 16770 35534 16772 35586
rect 16716 35028 16772 35534
rect 17500 35476 17556 35486
rect 17836 35476 17892 35646
rect 17500 35474 17668 35476
rect 17500 35422 17502 35474
rect 17554 35422 17668 35474
rect 17500 35420 17668 35422
rect 17500 35410 17556 35420
rect 16716 34962 16772 34972
rect 17220 35028 17276 35038
rect 16268 34914 16324 34926
rect 16268 34862 16270 34914
rect 16322 34862 16324 34914
rect 16268 33460 16324 34862
rect 16268 33402 16324 33404
rect 16268 33350 16270 33402
rect 16322 33350 16324 33402
rect 16268 33338 16324 33350
rect 16492 34914 16548 34926
rect 16492 34862 16494 34914
rect 16546 34862 16548 34914
rect 16492 33290 16548 34862
rect 17052 34916 17108 34926
rect 16772 34804 16828 34814
rect 16772 34710 16828 34748
rect 16940 34132 16996 34142
rect 16940 34038 16996 34076
rect 17052 33908 17108 34860
rect 17220 34860 17276 34972
rect 17220 34858 17332 34860
rect 17220 34806 17222 34858
rect 17274 34806 17332 34858
rect 17220 34794 17332 34806
rect 17276 34130 17332 34794
rect 17500 34858 17556 34870
rect 17500 34806 17502 34858
rect 17554 34806 17556 34858
rect 17500 34468 17556 34806
rect 17500 34402 17556 34412
rect 17276 34078 17278 34130
rect 17330 34078 17332 34130
rect 17276 34066 17332 34078
rect 17444 33908 17500 33918
rect 16940 33852 17108 33908
rect 17164 33906 17500 33908
rect 17164 33854 17446 33906
rect 17498 33854 17500 33906
rect 17164 33852 17500 33854
rect 16940 33458 16996 33852
rect 16940 33406 16942 33458
rect 16994 33406 16996 33458
rect 16940 33394 16996 33406
rect 17052 33684 17108 33694
rect 17052 33348 17108 33628
rect 17164 33460 17220 33852
rect 17444 33842 17500 33852
rect 17612 33796 17668 35420
rect 17836 35410 17892 35420
rect 17948 35698 18004 35710
rect 17948 35646 17950 35698
rect 18002 35646 18004 35698
rect 17780 34860 17836 34870
rect 17780 34858 17892 34860
rect 17780 34806 17782 34858
rect 17834 34806 17892 34858
rect 17780 34794 17892 34806
rect 17836 33908 17892 34794
rect 17948 34804 18004 35646
rect 17948 34738 18004 34748
rect 18060 34132 18116 38612
rect 18284 38276 18340 38670
rect 18284 38210 18340 38220
rect 18228 37828 18284 37838
rect 18228 37734 18284 37772
rect 18396 37828 18452 39900
rect 18620 39730 18676 40124
rect 18956 40114 19012 40124
rect 19292 40180 19348 40350
rect 20300 40404 20356 40414
rect 20300 40310 20356 40348
rect 20412 40402 20468 41134
rect 20636 41186 20692 41198
rect 20636 41134 20638 41186
rect 20690 41134 20692 41186
rect 20412 40350 20414 40402
rect 20466 40350 20468 40402
rect 19292 40114 19348 40124
rect 20132 40178 20188 40190
rect 20132 40126 20134 40178
rect 20186 40126 20188 40178
rect 18620 39678 18622 39730
rect 18674 39678 18676 39730
rect 18620 39666 18676 39678
rect 20132 39620 20188 40126
rect 20132 39554 20188 39564
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 20188 38722 20244 38734
rect 20188 38670 20190 38722
rect 20242 38670 20244 38722
rect 20188 38388 20244 38670
rect 20188 38322 20244 38332
rect 18620 38276 18676 38286
rect 18620 38182 18676 38220
rect 20412 38276 20468 40350
rect 20524 40404 20580 40414
rect 20524 39730 20580 40348
rect 20524 39678 20526 39730
rect 20578 39678 20580 39730
rect 20524 39666 20580 39678
rect 20636 40402 20692 41134
rect 21252 41130 21308 41468
rect 21252 41078 21254 41130
rect 21306 41078 21308 41130
rect 21252 41066 21308 41078
rect 21420 40964 21476 42924
rect 21532 42868 21588 43820
rect 21644 43810 21700 43820
rect 21756 43764 21812 45052
rect 22540 44994 22596 45006
rect 22540 44942 22542 44994
rect 22594 44942 22596 44994
rect 22316 44548 22372 44558
rect 22316 44454 22372 44492
rect 22540 44548 22596 44942
rect 23996 44548 24052 49200
rect 25564 46340 25620 49200
rect 25396 46284 25620 46340
rect 24444 45890 24500 45902
rect 24444 45838 24446 45890
rect 24498 45838 24500 45890
rect 22540 44482 22596 44492
rect 23772 44492 24052 44548
rect 24332 45780 24388 45790
rect 23100 44324 23156 44334
rect 21756 43708 21924 43764
rect 21736 43540 21792 43550
rect 21868 43540 21924 43708
rect 23100 43650 23156 44268
rect 23100 43598 23102 43650
rect 23154 43598 23156 43650
rect 23100 43586 23156 43598
rect 22652 43566 22708 43578
rect 21736 43538 21812 43540
rect 21736 43486 21738 43538
rect 21790 43486 21812 43538
rect 21736 43474 21812 43486
rect 21868 43484 22484 43540
rect 21756 42980 21812 43474
rect 21980 43316 22036 43326
rect 21980 43222 22036 43260
rect 21756 42914 21812 42924
rect 21868 43092 21924 43102
rect 21532 42802 21588 42812
rect 21756 42754 21812 42766
rect 21532 42698 21588 42710
rect 21532 42646 21534 42698
rect 21586 42646 21588 42698
rect 21532 42532 21588 42646
rect 21756 42702 21758 42754
rect 21810 42702 21812 42754
rect 21756 42644 21812 42702
rect 21756 42578 21812 42588
rect 21868 42532 21924 43036
rect 22316 42980 22372 42990
rect 21980 42868 22036 42878
rect 21980 42774 22036 42812
rect 22148 42756 22204 42766
rect 22148 42662 22204 42700
rect 22316 42754 22372 42924
rect 22316 42702 22318 42754
rect 22370 42702 22372 42754
rect 22316 42690 22372 42702
rect 22428 42756 22484 43484
rect 22652 43514 22654 43566
rect 22706 43514 22708 43566
rect 22652 43092 22708 43514
rect 22876 43538 22932 43550
rect 22876 43486 22878 43538
rect 22930 43486 22932 43538
rect 22876 43316 22932 43486
rect 22876 43250 22932 43260
rect 22988 43540 23044 43550
rect 23436 43538 23492 43550
rect 22652 43026 22708 43036
rect 22764 42756 22820 42766
rect 22428 42754 22932 42756
rect 22428 42702 22766 42754
rect 22818 42702 22932 42754
rect 22428 42700 22932 42702
rect 22764 42690 22820 42700
rect 22484 42532 22540 42542
rect 21868 42476 22260 42532
rect 21532 42466 21588 42476
rect 21624 41972 21680 41982
rect 21868 41972 21924 41982
rect 21624 41970 21700 41972
rect 21624 41918 21626 41970
rect 21678 41918 21700 41970
rect 21624 41906 21700 41918
rect 20636 40350 20638 40402
rect 20690 40350 20692 40402
rect 20636 38668 20692 40350
rect 20412 38210 20468 38220
rect 20524 38612 20692 38668
rect 20748 40908 21476 40964
rect 21532 41636 21588 41646
rect 21532 41147 21588 41580
rect 21644 41412 21700 41906
rect 21868 41878 21924 41916
rect 21644 41346 21700 41356
rect 22204 41410 22260 42476
rect 22484 42438 22540 42476
rect 22204 41358 22206 41410
rect 22258 41358 22260 41410
rect 22204 41346 22260 41358
rect 22428 42008 22484 42020
rect 22428 41956 22430 42008
rect 22482 41956 22484 42008
rect 21532 41095 21534 41147
rect 21586 41095 21588 41147
rect 18956 38052 19012 38062
rect 20524 38052 20580 38612
rect 18956 38050 19236 38052
rect 18956 37998 18958 38050
rect 19010 37998 19236 38050
rect 18956 37996 19236 37998
rect 18956 37986 19012 37996
rect 18396 37762 18452 37772
rect 18508 37380 18564 37390
rect 18284 37294 18340 37306
rect 18284 37268 18286 37294
rect 18338 37268 18340 37294
rect 18284 37202 18340 37212
rect 18508 37266 18564 37324
rect 19068 37380 19124 37390
rect 18508 37214 18510 37266
rect 18562 37214 18564 37266
rect 18284 36370 18340 36382
rect 18284 36318 18286 36370
rect 18338 36318 18340 36370
rect 18284 35812 18340 36318
rect 18508 36260 18564 37214
rect 18620 37268 18676 37278
rect 19068 37266 19124 37324
rect 18620 36932 18676 37212
rect 18900 37210 18956 37222
rect 18732 37156 18788 37166
rect 18732 37062 18788 37100
rect 18900 37158 18902 37210
rect 18954 37158 18956 37210
rect 19068 37214 19070 37266
rect 19122 37214 19124 37266
rect 19068 37202 19124 37214
rect 18900 37156 18956 37158
rect 18900 37090 18956 37100
rect 18620 36876 18900 36932
rect 18844 36706 18900 36876
rect 18844 36654 18846 36706
rect 18898 36654 18900 36706
rect 18844 36642 18900 36654
rect 19180 36708 19236 37996
rect 20412 37996 20580 38052
rect 19684 37940 19740 37950
rect 19684 37846 19740 37884
rect 20132 37828 20188 37838
rect 20132 37826 20244 37828
rect 20132 37774 20134 37826
rect 20186 37774 20244 37826
rect 20132 37762 20244 37774
rect 20188 37716 20244 37762
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20188 37650 20244 37660
rect 20412 37716 20468 37996
rect 20412 37650 20468 37660
rect 20580 37826 20636 37838
rect 20580 37774 20582 37826
rect 20634 37774 20636 37826
rect 20580 37716 20636 37774
rect 20580 37650 20636 37660
rect 19836 37594 20100 37604
rect 20244 37492 20300 37502
rect 20244 37490 20692 37492
rect 20244 37438 20246 37490
rect 20298 37438 20692 37490
rect 20244 37436 20692 37438
rect 20244 37426 20300 37436
rect 19292 37268 19348 37278
rect 19292 37174 19348 37212
rect 20300 37268 20356 37278
rect 20076 37156 20132 37166
rect 19572 37044 19628 37054
rect 19180 36642 19236 36652
rect 19292 37042 19628 37044
rect 19292 36990 19574 37042
rect 19626 36990 19628 37042
rect 19292 36988 19628 36990
rect 19292 36596 19348 36988
rect 19572 36978 19628 36988
rect 20076 36820 20132 37100
rect 20300 36932 20356 37212
rect 20412 37266 20468 37278
rect 20412 37214 20414 37266
rect 20466 37214 20468 37266
rect 20412 37156 20468 37214
rect 20636 37266 20692 37436
rect 20636 37214 20638 37266
rect 20690 37214 20692 37266
rect 20636 37202 20692 37214
rect 20748 37268 20804 40908
rect 20916 40628 20972 40638
rect 20916 40514 20972 40572
rect 21532 40628 21588 41095
rect 21812 41130 21868 41142
rect 21812 41078 21814 41130
rect 21866 41078 21868 41130
rect 21812 41076 21868 41078
rect 21980 41076 22036 41086
rect 21812 41020 21980 41076
rect 21532 40562 21588 40572
rect 20916 40462 20918 40514
rect 20970 40462 20972 40514
rect 20916 40450 20972 40462
rect 21308 40404 21364 40414
rect 21308 40310 21364 40348
rect 21420 40402 21476 40414
rect 21420 40350 21422 40402
rect 21474 40350 21476 40402
rect 21420 40292 21476 40350
rect 21588 40404 21644 40414
rect 21588 40310 21644 40348
rect 21420 40226 21476 40236
rect 21980 40290 22036 41020
rect 22428 41076 22484 41956
rect 22764 41972 22820 41982
rect 22764 41878 22820 41916
rect 22708 41524 22764 41534
rect 22708 41410 22764 41468
rect 22708 41358 22710 41410
rect 22762 41358 22764 41410
rect 22708 41346 22764 41358
rect 22428 41010 22484 41020
rect 22876 41188 22932 42700
rect 22988 42532 23044 43484
rect 23268 43482 23324 43494
rect 23268 43430 23270 43482
rect 23322 43430 23324 43482
rect 23268 42868 23324 43430
rect 23436 43486 23438 43538
rect 23490 43486 23492 43538
rect 23436 43316 23492 43486
rect 23660 43538 23716 43550
rect 23660 43486 23662 43538
rect 23714 43486 23716 43538
rect 23436 43250 23492 43260
rect 23548 43428 23604 43438
rect 23212 42812 23324 42868
rect 23548 42866 23604 43372
rect 23660 43092 23716 43486
rect 23660 43026 23716 43036
rect 23548 42814 23550 42866
rect 23602 42814 23604 42866
rect 23212 42756 23268 42812
rect 23548 42802 23604 42814
rect 23212 42532 23268 42700
rect 22988 42466 23044 42476
rect 23156 42476 23268 42532
rect 23156 41914 23212 42476
rect 23772 42196 23828 44492
rect 23996 44322 24052 44334
rect 23996 44270 23998 44322
rect 24050 44270 24052 44322
rect 23996 43662 24052 44270
rect 24220 44324 24276 44334
rect 24220 44230 24276 44268
rect 24332 44212 24388 45724
rect 24444 45218 24500 45838
rect 24780 45892 24836 45902
rect 24780 45798 24836 45836
rect 25396 45722 25452 46284
rect 25844 46116 25900 46126
rect 25844 46114 26516 46116
rect 25844 46062 25846 46114
rect 25898 46062 26516 46114
rect 25844 46060 26516 46062
rect 25844 46050 25900 46060
rect 26124 45892 26180 45902
rect 25396 45670 25398 45722
rect 25450 45670 25452 45722
rect 25396 45658 25452 45670
rect 25676 45890 26180 45892
rect 25676 45838 26126 45890
rect 26178 45838 26180 45890
rect 25676 45836 26180 45838
rect 24444 45166 24446 45218
rect 24498 45166 24500 45218
rect 24444 45154 24500 45166
rect 25228 45108 25284 45118
rect 25004 44548 25060 44558
rect 25004 44454 25060 44492
rect 24500 44212 24556 44222
rect 24332 44210 24556 44212
rect 24332 44158 24502 44210
rect 24554 44158 24556 44210
rect 24332 44156 24556 44158
rect 24500 44146 24556 44156
rect 25228 44100 25284 45052
rect 25676 44434 25732 45836
rect 26124 45826 26180 45836
rect 26236 45890 26292 45902
rect 26236 45838 26238 45890
rect 26290 45838 26292 45890
rect 26012 45668 26068 45678
rect 26012 45106 26068 45612
rect 26012 45054 26014 45106
rect 26066 45054 26068 45106
rect 26012 45042 26068 45054
rect 26236 44772 26292 45838
rect 26460 45890 26516 46060
rect 26460 45838 26462 45890
rect 26514 45838 26516 45890
rect 26460 45826 26516 45838
rect 27132 45780 27188 49200
rect 28700 49140 28756 49200
rect 28924 49140 28980 49308
rect 28700 49084 28980 49140
rect 28812 46058 28868 46070
rect 28812 46006 28814 46058
rect 28866 46006 28868 46058
rect 28812 46004 28868 46006
rect 28812 45948 29428 46004
rect 27916 45892 27972 45902
rect 28364 45892 28420 45902
rect 27132 45714 27188 45724
rect 27804 45890 27972 45892
rect 27804 45838 27918 45890
rect 27970 45838 27972 45890
rect 27804 45836 27972 45838
rect 26796 45668 26852 45678
rect 26796 45574 26852 45612
rect 27580 45666 27636 45678
rect 27580 45614 27582 45666
rect 27634 45614 27636 45666
rect 27244 45556 27300 45566
rect 26908 44772 26964 44782
rect 26236 44716 26796 44772
rect 26236 44548 26292 44558
rect 25676 44382 25678 44434
rect 25730 44382 25732 44434
rect 25676 44370 25732 44382
rect 25900 44436 25956 44446
rect 25340 44324 25396 44334
rect 25900 44322 25956 44380
rect 25340 44230 25396 44268
rect 25508 44266 25564 44278
rect 25228 44034 25284 44044
rect 25508 44214 25510 44266
rect 25562 44214 25564 44266
rect 25900 44270 25902 44322
rect 25954 44270 25956 44322
rect 25900 44258 25956 44270
rect 26236 44266 26292 44492
rect 26740 44546 26796 44716
rect 26740 44494 26742 44546
rect 26794 44494 26796 44546
rect 26740 44482 26796 44494
rect 25508 43764 25564 44214
rect 26236 44214 26238 44266
rect 26290 44214 26292 44266
rect 26236 43876 26292 44214
rect 26236 43820 26628 43876
rect 25508 43708 25620 43764
rect 23940 43650 24052 43662
rect 23940 43598 23942 43650
rect 23994 43598 24052 43650
rect 23940 43596 24052 43598
rect 23940 43586 23996 43596
rect 24220 43540 24276 43550
rect 24220 43538 24724 43540
rect 24220 43486 24222 43538
rect 24274 43486 24724 43538
rect 24220 43484 24724 43486
rect 24220 43474 24276 43484
rect 24556 43316 24612 43326
rect 24556 43222 24612 43260
rect 24668 42532 24724 43484
rect 25452 43538 25508 43550
rect 25452 43486 25454 43538
rect 25506 43486 25508 43538
rect 25284 43316 25340 43326
rect 24556 42476 24724 42532
rect 25228 43314 25340 43316
rect 25228 43262 25286 43314
rect 25338 43262 25340 43314
rect 25228 43250 25340 43262
rect 23772 42140 24164 42196
rect 22876 40964 22932 41132
rect 22988 41858 23044 41870
rect 22988 41806 22990 41858
rect 23042 41806 23044 41858
rect 22988 41186 23044 41806
rect 23156 41862 23158 41914
rect 23210 41862 23212 41914
rect 23156 41748 23212 41862
rect 22988 41134 22990 41186
rect 23042 41134 23044 41186
rect 22988 41122 23044 41134
rect 23100 41692 23212 41748
rect 23324 41972 23380 41982
rect 23772 41972 23828 41982
rect 22876 40908 23044 40964
rect 21980 40238 21982 40290
rect 22034 40238 22036 40290
rect 21980 40226 22036 40238
rect 22092 40404 22148 40414
rect 22092 39844 22148 40348
rect 22428 40402 22484 40414
rect 22428 40350 22430 40402
rect 22482 40350 22484 40402
rect 21980 39788 22148 39844
rect 22204 40292 22260 40302
rect 21308 39620 21364 39630
rect 21308 39526 21364 39564
rect 21980 39284 22036 39788
rect 22204 39732 22260 40236
rect 21756 39228 22036 39284
rect 22184 39676 22260 39732
rect 22316 40180 22372 40190
rect 22184 39620 22240 39676
rect 22184 39562 22240 39564
rect 22184 39510 22186 39562
rect 22238 39510 22240 39562
rect 21084 38948 21140 38958
rect 21084 38878 21140 38892
rect 20860 38836 20916 38846
rect 21084 38826 21086 38878
rect 21138 38826 21140 38878
rect 21084 38814 21140 38826
rect 21756 38834 21812 39228
rect 22184 39060 22240 39510
rect 22184 38994 22240 39004
rect 22316 39002 22372 40124
rect 22316 38950 22318 39002
rect 22370 38950 22372 39002
rect 22316 38938 22372 38950
rect 22428 39506 22484 40350
rect 22428 39454 22430 39506
rect 22482 39454 22484 39506
rect 20860 38742 20916 38780
rect 21756 38782 21758 38834
rect 21810 38782 21812 38834
rect 21756 38770 21812 38782
rect 21980 38873 22036 38885
rect 21980 38821 21982 38873
rect 22034 38821 22036 38873
rect 22316 38836 22372 38846
rect 21196 38724 21252 38762
rect 21196 38658 21252 38668
rect 21980 38724 22036 38821
rect 21980 38658 22036 38668
rect 22092 38834 22372 38836
rect 22092 38782 22318 38834
rect 22370 38782 22372 38834
rect 22092 38780 22372 38782
rect 22092 38612 22148 38780
rect 22316 38770 22372 38780
rect 22428 38836 22484 39454
rect 22428 38770 22484 38780
rect 22540 40402 22596 40414
rect 22540 40350 22542 40402
rect 22594 40350 22596 40402
rect 22540 38948 22596 40350
rect 22820 40404 22876 40414
rect 22820 40310 22876 40348
rect 22092 38546 22148 38556
rect 21084 38388 21140 38398
rect 21084 37940 21140 38332
rect 22204 38276 22260 38286
rect 22540 38276 22596 38892
rect 22764 39620 22820 39630
rect 22988 39620 23044 40908
rect 22764 39618 23044 39620
rect 22764 39566 22766 39618
rect 22818 39566 23044 39618
rect 22764 39564 23044 39566
rect 22764 38668 22820 39564
rect 22204 38274 22596 38276
rect 22204 38222 22206 38274
rect 22258 38222 22596 38274
rect 22204 38220 22596 38222
rect 22652 38612 22820 38668
rect 22932 38724 22988 38762
rect 22932 38658 22988 38668
rect 22204 38210 22260 38220
rect 21252 37994 21308 38006
rect 21252 37942 21254 37994
rect 21306 37942 21308 37994
rect 21252 37940 21308 37942
rect 21084 37884 21308 37940
rect 21476 37994 21532 38006
rect 21476 37942 21478 37994
rect 21530 37942 21532 37994
rect 21476 37940 21532 37942
rect 21644 37994 21700 38006
rect 21644 37942 21646 37994
rect 21698 37942 21700 37994
rect 21476 37884 21568 37940
rect 21084 37604 21140 37884
rect 21084 37538 21140 37548
rect 21308 37716 21364 37726
rect 20748 37202 20804 37212
rect 20412 37090 20468 37100
rect 20300 36876 20580 36932
rect 20076 36764 20356 36820
rect 20300 36650 20356 36764
rect 20300 36598 20302 36650
rect 20354 36598 20356 36650
rect 20300 36586 20356 36598
rect 20412 36596 20468 36606
rect 19292 36530 19348 36540
rect 19964 36482 20020 36494
rect 19087 36428 19143 36438
rect 19964 36430 19966 36482
rect 20018 36430 20020 36482
rect 19068 36426 19348 36428
rect 19068 36374 19089 36426
rect 19141 36374 19348 36426
rect 19068 36372 19348 36374
rect 19068 36362 19143 36372
rect 18508 36204 18676 36260
rect 18284 35746 18340 35756
rect 18452 35924 18508 35934
rect 18452 35810 18508 35868
rect 18452 35758 18454 35810
rect 18506 35758 18508 35810
rect 18452 35746 18508 35758
rect 18172 35698 18228 35710
rect 18172 35646 18174 35698
rect 18226 35646 18228 35698
rect 18172 35028 18228 35646
rect 18620 35588 18676 36204
rect 18788 35812 18844 35822
rect 19068 35812 19124 36362
rect 18788 35754 18844 35756
rect 18788 35702 18790 35754
rect 18842 35702 18844 35754
rect 18788 35690 18844 35702
rect 19012 35756 19124 35812
rect 19012 35754 19068 35756
rect 19012 35702 19014 35754
rect 19066 35702 19068 35754
rect 19012 35690 19068 35702
rect 19180 35737 19236 35749
rect 19180 35685 19182 35737
rect 19234 35685 19236 35737
rect 19180 35588 19236 35685
rect 18620 35532 19236 35588
rect 18172 34962 18228 34972
rect 18284 35476 18340 35486
rect 18172 34804 18228 34842
rect 18172 34738 18228 34748
rect 18284 34692 18340 35420
rect 19068 34916 19124 34926
rect 19068 34822 19124 34860
rect 18788 34802 18844 34814
rect 18788 34750 18790 34802
rect 18842 34750 18844 34802
rect 18284 34636 18452 34692
rect 18060 34038 18116 34076
rect 18284 34468 18340 34478
rect 17836 33852 18116 33908
rect 17612 33730 17668 33740
rect 17164 33404 17276 33460
rect 17220 33348 17276 33404
rect 17388 33348 17444 33358
rect 17052 33292 17164 33348
rect 17220 33346 17444 33348
rect 17220 33294 17390 33346
rect 17442 33294 17444 33346
rect 17220 33292 17444 33294
rect 16492 33238 16494 33290
rect 16546 33238 16548 33290
rect 16492 33236 16548 33238
rect 16492 33170 16548 33180
rect 17108 33290 17164 33292
rect 17108 33238 17110 33290
rect 17162 33238 17164 33290
rect 17388 33282 17444 33292
rect 17108 32788 17164 33238
rect 17500 33236 17556 33246
rect 17108 32732 17220 32788
rect 16828 32564 16884 32602
rect 16828 32498 16884 32508
rect 17164 32228 17220 32732
rect 17500 32674 17556 33180
rect 18060 33236 18116 33852
rect 18284 33358 18340 34412
rect 18264 33348 18340 33358
rect 18320 33292 18340 33348
rect 18264 33263 18266 33292
rect 18318 33263 18320 33292
rect 18264 33251 18320 33263
rect 18060 33170 18116 33180
rect 18396 33124 18452 34636
rect 18788 34244 18844 34750
rect 19180 34804 19236 35532
rect 19292 35476 19348 36372
rect 19964 36260 20020 36430
rect 20412 36482 20468 36540
rect 20412 36430 20414 36482
rect 20466 36430 20468 36482
rect 20412 36418 20468 36430
rect 20524 36260 20580 36876
rect 20748 36820 20804 36830
rect 21308 36820 21364 37660
rect 21512 37492 21568 37884
rect 21512 37322 21568 37436
rect 21512 37270 21514 37322
rect 21566 37270 21568 37322
rect 21512 37258 21568 37270
rect 21644 37380 21700 37942
rect 22540 37940 22596 37950
rect 22428 37492 22484 37502
rect 20748 36482 20804 36764
rect 20748 36430 20750 36482
rect 20802 36430 20804 36482
rect 20524 36204 20692 36260
rect 19964 36194 20020 36204
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19740 35924 19796 35934
rect 19740 35810 19796 35868
rect 19740 35758 19742 35810
rect 19794 35758 19796 35810
rect 19740 35746 19796 35758
rect 20468 35727 20524 35739
rect 20188 35700 20244 35710
rect 20468 35700 20470 35727
rect 20188 35606 20244 35644
rect 20412 35675 20470 35700
rect 20522 35675 20524 35727
rect 20412 35644 20524 35675
rect 19292 35410 19348 35420
rect 19628 35476 19684 35486
rect 19516 35252 19572 35262
rect 19180 34738 19236 34748
rect 19292 34914 19348 34926
rect 19292 34862 19294 34914
rect 19346 34862 19348 34914
rect 18788 34178 18844 34188
rect 18620 33796 18676 33806
rect 18508 33460 18564 33470
rect 18508 33366 18564 33404
rect 17500 32622 17502 32674
rect 17554 32622 17556 32674
rect 17500 32610 17556 32622
rect 18172 33068 18452 33124
rect 18060 32601 18116 32613
rect 18060 32549 18062 32601
rect 18114 32549 18116 32601
rect 17780 32506 17836 32518
rect 17780 32454 17782 32506
rect 17834 32454 17836 32506
rect 17780 32452 17836 32454
rect 17164 32162 17220 32172
rect 17612 32228 17668 32238
rect 15708 31826 15764 31836
rect 16044 31836 16212 31892
rect 16268 32116 16324 32126
rect 15876 31780 15932 31790
rect 15876 31686 15932 31724
rect 16044 31108 16100 31836
rect 16268 31678 16324 32060
rect 16828 31892 16884 31902
rect 16212 31666 16324 31678
rect 16212 31614 16214 31666
rect 16266 31614 16324 31666
rect 16212 31612 16324 31614
rect 16492 31778 16548 31790
rect 16492 31726 16494 31778
rect 16546 31726 16548 31778
rect 16212 31602 16268 31612
rect 16492 31220 16548 31726
rect 16492 31154 16548 31164
rect 16604 31778 16660 31790
rect 16604 31726 16606 31778
rect 16658 31726 16660 31778
rect 15932 31052 16100 31108
rect 16604 31108 16660 31726
rect 15820 30770 15876 30782
rect 15820 30718 15822 30770
rect 15874 30718 15876 30770
rect 15820 30322 15876 30718
rect 15820 30270 15822 30322
rect 15874 30270 15876 30322
rect 15820 30258 15876 30270
rect 15764 29540 15820 29550
rect 15932 29540 15988 31052
rect 16604 31042 16660 31052
rect 16716 31556 16772 31566
rect 16156 30996 16212 31006
rect 15764 29538 15988 29540
rect 15764 29486 15766 29538
rect 15818 29486 15988 29538
rect 15764 29484 15988 29486
rect 16044 30994 16212 30996
rect 16044 30942 16158 30994
rect 16210 30942 16212 30994
rect 16044 30940 16212 30942
rect 16044 29540 16100 30940
rect 16156 30930 16212 30940
rect 16716 30994 16772 31500
rect 16716 30942 16718 30994
rect 16770 30942 16772 30994
rect 16716 30930 16772 30942
rect 16828 30994 16884 31836
rect 17388 31892 17444 31902
rect 17612 31892 17668 32172
rect 17780 32004 17836 32396
rect 17780 31948 18004 32004
rect 17612 31836 17836 31892
rect 17388 31778 17444 31836
rect 17164 31722 17220 31734
rect 17164 31670 17166 31722
rect 17218 31670 17220 31722
rect 17388 31726 17390 31778
rect 17442 31726 17444 31778
rect 17780 31834 17836 31836
rect 17780 31782 17782 31834
rect 17834 31782 17836 31834
rect 17780 31770 17836 31782
rect 17388 31714 17444 31726
rect 17164 31556 17220 31670
rect 17612 31668 17668 31678
rect 17164 31490 17220 31500
rect 17500 31666 17668 31668
rect 17500 31614 17614 31666
rect 17666 31614 17668 31666
rect 17500 31612 17668 31614
rect 16828 30942 16830 30994
rect 16882 30942 16884 30994
rect 16828 30930 16884 30942
rect 16436 30772 16492 30782
rect 16436 30770 16772 30772
rect 16436 30718 16438 30770
rect 16490 30718 16772 30770
rect 16436 30716 16772 30718
rect 16436 30706 16492 30716
rect 16716 30548 16772 30716
rect 16716 30492 16996 30548
rect 16492 29988 16548 29998
rect 16940 29988 16996 30492
rect 16380 29652 16436 29662
rect 16212 29540 16268 29550
rect 16044 29538 16268 29540
rect 16044 29486 16214 29538
rect 16266 29486 16268 29538
rect 16044 29484 16268 29486
rect 15764 29474 15820 29484
rect 16212 29474 16268 29484
rect 15596 29372 15708 29428
rect 15484 29334 15540 29372
rect 15652 29316 15708 29372
rect 15652 29260 15764 29316
rect 15596 29092 15652 29102
rect 15372 28812 15540 28868
rect 15260 28242 15316 28252
rect 15372 28644 15428 28654
rect 15372 28084 15428 28588
rect 15484 28532 15540 28812
rect 15484 28466 15540 28476
rect 15148 27806 15150 27858
rect 15202 27806 15204 27858
rect 15148 27794 15204 27806
rect 15260 28028 15428 28084
rect 15484 28308 15540 28318
rect 15036 27682 15092 27692
rect 15260 27690 15316 28028
rect 15372 27860 15428 27898
rect 15372 27794 15428 27804
rect 14588 27022 14590 27074
rect 14642 27022 14644 27074
rect 14588 27010 14644 27022
rect 14700 27580 14980 27636
rect 15260 27638 15262 27690
rect 15314 27638 15316 27690
rect 15260 27626 15316 27638
rect 15372 27636 15428 27646
rect 14252 26898 14308 26908
rect 14364 26852 14476 26908
rect 13580 26292 13636 26302
rect 13580 26290 13748 26292
rect 13580 26238 13582 26290
rect 13634 26238 13748 26290
rect 13580 26236 13748 26238
rect 13580 26226 13636 26236
rect 13468 26070 13470 26122
rect 13522 26070 13524 26122
rect 13468 26058 13524 26070
rect 13132 25666 13188 25676
rect 13562 25844 13618 25854
rect 13562 25730 13618 25788
rect 13562 25678 13564 25730
rect 13616 25678 13618 25730
rect 13562 25666 13618 25678
rect 12684 25508 12740 25528
rect 12348 25450 12740 25452
rect 12348 25398 12686 25450
rect 12738 25398 12740 25450
rect 12348 25396 12740 25398
rect 12124 25386 12180 25396
rect 12236 24948 12292 25396
rect 12684 25386 12740 25396
rect 13580 25508 13636 25518
rect 13132 25060 13188 25070
rect 12684 24948 12740 24958
rect 12236 24892 12628 24948
rect 12124 24836 12180 24846
rect 12124 24742 12180 24780
rect 12236 24724 12292 24734
rect 12236 24630 12292 24668
rect 12572 24722 12628 24892
rect 12572 24670 12574 24722
rect 12626 24670 12628 24722
rect 11994 24162 12068 24174
rect 11994 24110 11996 24162
rect 12048 24110 12068 24162
rect 11994 24108 12068 24110
rect 11994 24098 12050 24108
rect 11676 22708 11732 23548
rect 12236 23938 12292 23950
rect 12236 23886 12238 23938
rect 12290 23886 12292 23938
rect 12236 23156 12292 23886
rect 12572 23380 12628 24670
rect 12572 23314 12628 23324
rect 12684 23960 12740 24892
rect 12684 23938 12796 23960
rect 12684 23886 12742 23938
rect 12794 23886 12796 23938
rect 12684 23874 12796 23886
rect 12908 23940 12964 23950
rect 12684 23322 12740 23874
rect 12684 23270 12686 23322
rect 12738 23270 12740 23322
rect 12684 23258 12740 23270
rect 12684 23156 12740 23166
rect 12236 23154 12740 23156
rect 12236 23102 12686 23154
rect 12738 23102 12740 23154
rect 12236 23100 12740 23102
rect 12124 23044 12180 23054
rect 11676 22642 11732 22652
rect 11788 23042 12180 23044
rect 11788 22990 12126 23042
rect 12178 22990 12180 23042
rect 11788 22988 12180 22990
rect 11788 22596 11844 22988
rect 12124 22978 12180 22988
rect 11784 22540 11844 22596
rect 11564 22372 11620 22382
rect 11784 22372 11840 22540
rect 11564 22370 11840 22372
rect 11564 22318 11566 22370
rect 11618 22332 11840 22370
rect 11618 22318 11786 22332
rect 11564 22316 11786 22318
rect 11564 22306 11620 22316
rect 11784 22280 11786 22316
rect 11838 22280 11840 22332
rect 11784 22268 11840 22280
rect 11788 22148 11844 22158
rect 11452 22092 11620 22148
rect 11340 22082 11396 22092
rect 10892 21746 10948 21756
rect 10444 21586 10612 21588
rect 10444 21534 10446 21586
rect 10498 21534 10612 21586
rect 10444 21532 10612 21534
rect 10444 21522 10500 21532
rect 10556 21364 10612 21374
rect 10556 21026 10612 21308
rect 10556 20974 10558 21026
rect 10610 20974 10612 21026
rect 10556 20962 10612 20974
rect 11228 21028 11284 21038
rect 11228 20934 11284 20972
rect 11564 21028 11620 22092
rect 11564 20962 11620 20972
rect 11788 20970 11844 22092
rect 12348 21700 12404 23100
rect 12684 23090 12740 23100
rect 12908 22708 12964 23884
rect 12572 22652 12964 22708
rect 13020 23380 13076 23390
rect 12572 22538 12628 22652
rect 12572 22486 12574 22538
rect 12626 22486 12628 22538
rect 12572 22474 12628 22486
rect 12460 22372 12516 22382
rect 12460 22278 12516 22316
rect 13020 21810 13076 23324
rect 13020 21758 13022 21810
rect 13074 21758 13076 21810
rect 13020 21746 13076 21758
rect 12348 21698 12740 21700
rect 12348 21646 12350 21698
rect 12402 21646 12740 21698
rect 12348 21644 12740 21646
rect 12348 21634 12404 21644
rect 12684 21586 12740 21644
rect 12684 21534 12686 21586
rect 12738 21534 12740 21586
rect 12684 21522 12740 21534
rect 11788 20918 11790 20970
rect 11842 20918 11844 20970
rect 11788 20906 11844 20918
rect 11564 20804 11620 20814
rect 12012 20804 12068 20814
rect 11564 20802 12068 20804
rect 11564 20750 11566 20802
rect 11618 20750 12014 20802
rect 12066 20750 12068 20802
rect 11564 20748 12068 20750
rect 11564 20738 11620 20748
rect 11676 20468 11732 20478
rect 10444 19906 10500 19918
rect 10444 19854 10446 19906
rect 10498 19854 10500 19906
rect 10444 19460 10500 19854
rect 10444 19394 10500 19404
rect 11676 19124 11732 20412
rect 12012 20132 12068 20748
rect 12572 20802 12628 20814
rect 12572 20750 12574 20802
rect 12626 20750 12628 20802
rect 12348 20132 12404 20142
rect 12012 20130 12404 20132
rect 12012 20078 12350 20130
rect 12402 20078 12404 20130
rect 12012 20076 12404 20078
rect 12348 20066 12404 20076
rect 12124 19236 12180 19246
rect 12460 19236 12516 19246
rect 12572 19236 12628 20750
rect 13020 20020 13076 20030
rect 13132 20020 13188 25004
rect 13580 24554 13636 25452
rect 13580 24502 13582 24554
rect 13634 24502 13636 24554
rect 13580 24490 13636 24502
rect 13692 24722 13748 26236
rect 13916 25844 13972 26852
rect 14140 26740 14196 26750
rect 14364 26740 14420 26852
rect 13916 25778 13972 25788
rect 14028 26290 14084 26302
rect 14028 26238 14030 26290
rect 14082 26238 14084 26290
rect 13804 25620 13860 25630
rect 13804 25506 13860 25564
rect 13804 25454 13806 25506
rect 13858 25454 13860 25506
rect 13804 25442 13860 25454
rect 14028 25172 14084 26238
rect 14140 26290 14196 26684
rect 14140 26238 14142 26290
rect 14194 26238 14196 26290
rect 14140 26226 14196 26238
rect 14286 26684 14420 26740
rect 14286 26327 14342 26684
rect 14286 26275 14288 26327
rect 14340 26275 14342 26327
rect 14286 25844 14342 26275
rect 14700 26178 14756 27580
rect 14980 27412 15036 27422
rect 14980 27298 15036 27356
rect 14980 27246 14982 27298
rect 15034 27246 15036 27298
rect 14980 27234 15036 27246
rect 14812 27076 14868 27114
rect 14812 27010 14868 27020
rect 15372 26964 15428 27580
rect 14700 26126 14702 26178
rect 14754 26126 14756 26178
rect 14700 26114 14756 26126
rect 14812 26852 14868 26862
rect 14140 25788 14342 25844
rect 14140 25284 14196 25788
rect 14812 25674 14868 26796
rect 15372 26514 15428 26908
rect 15372 26462 15374 26514
rect 15426 26462 15428 26514
rect 15372 26450 15428 26462
rect 15484 27074 15540 28252
rect 15596 27860 15652 29036
rect 15708 28868 15764 29260
rect 15932 28868 15988 28878
rect 15708 28866 15988 28868
rect 15708 28814 15934 28866
rect 15986 28814 15988 28866
rect 15708 28812 15988 28814
rect 15932 28802 15988 28812
rect 16268 28644 16324 28654
rect 16380 28644 16436 29596
rect 16492 29426 16548 29932
rect 16492 29374 16494 29426
rect 16546 29374 16548 29426
rect 16492 29362 16548 29374
rect 16716 29932 16996 29988
rect 17500 29988 17556 31612
rect 17612 31602 17668 31612
rect 17948 31556 18004 31948
rect 17836 31500 18004 31556
rect 18060 31556 18116 32549
rect 17668 30996 17724 31006
rect 17668 30902 17724 30940
rect 17724 30324 17780 30334
rect 17836 30324 17892 31500
rect 18060 31490 18116 31500
rect 17724 30322 17892 30324
rect 17724 30270 17726 30322
rect 17778 30270 17892 30322
rect 17724 30268 17892 30270
rect 17948 31108 18004 31118
rect 17948 30994 18004 31052
rect 17948 30942 17950 30994
rect 18002 30942 18004 30994
rect 17948 30324 18004 30942
rect 17724 30258 17780 30268
rect 17948 30258 18004 30268
rect 18172 30100 18228 33068
rect 18284 32788 18340 32798
rect 18620 32788 18676 33740
rect 18284 32618 18340 32732
rect 18284 32566 18286 32618
rect 18338 32566 18340 32618
rect 18284 32554 18340 32566
rect 18508 32732 18676 32788
rect 18508 31892 18564 32732
rect 18620 32562 18676 32574
rect 18620 32510 18622 32562
rect 18674 32510 18676 32562
rect 18620 32452 18676 32510
rect 18620 32386 18676 32396
rect 18788 32564 18844 32574
rect 18788 32394 18844 32508
rect 18788 32342 18790 32394
rect 18842 32342 18844 32394
rect 18788 32330 18844 32342
rect 19292 32564 19348 34862
rect 19516 33460 19572 35196
rect 19628 35138 19684 35420
rect 20412 35364 20468 35644
rect 20636 35586 20692 36204
rect 20748 36148 20804 36430
rect 21196 36764 21364 36820
rect 21532 37156 21588 37166
rect 20748 36082 20804 36092
rect 20860 36372 20916 36382
rect 20860 36036 20916 36316
rect 20860 35970 20916 35980
rect 21028 36260 21084 36270
rect 21028 35922 21084 36204
rect 21028 35870 21030 35922
rect 21082 35870 21084 35922
rect 21028 35858 21084 35870
rect 20860 35812 20916 35822
rect 20860 35698 20916 35756
rect 20860 35646 20862 35698
rect 20914 35646 20916 35698
rect 20860 35634 20916 35646
rect 20636 35534 20638 35586
rect 20690 35534 20692 35586
rect 20636 35522 20692 35534
rect 19628 35086 19630 35138
rect 19682 35086 19684 35138
rect 19628 35074 19684 35086
rect 20076 35308 20468 35364
rect 19871 34860 19927 34870
rect 19628 34858 19927 34860
rect 19628 34806 19873 34858
rect 19925 34806 19927 34858
rect 19628 34804 19927 34806
rect 19628 34356 19684 34804
rect 19871 34794 19927 34804
rect 20076 34804 20132 35308
rect 20076 34738 20132 34748
rect 20748 34914 20804 34926
rect 20748 34862 20750 34914
rect 20802 34862 20804 34914
rect 20300 34580 20356 34590
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19964 34356 20020 34366
rect 19628 34300 19796 34356
rect 19516 33404 19684 33460
rect 19404 33348 19460 33358
rect 19404 33346 19572 33348
rect 19404 33294 19406 33346
rect 19458 33294 19572 33346
rect 19404 33292 19572 33294
rect 19404 33282 19460 33292
rect 18396 31836 18564 31892
rect 18956 32004 19012 32014
rect 18284 31220 18340 31230
rect 18284 31038 18340 31164
rect 18284 30986 18286 31038
rect 18338 30986 18340 31038
rect 18284 30974 18340 30986
rect 18396 30884 18452 31836
rect 18620 31780 18676 31790
rect 18620 31698 18622 31724
rect 18674 31698 18676 31724
rect 18620 31686 18676 31698
rect 18620 30996 18676 31006
rect 18396 30790 18452 30828
rect 18508 30940 18620 30996
rect 18508 30660 18564 30940
rect 18620 30902 18676 30940
rect 18340 30604 18564 30660
rect 18732 30884 18788 30894
rect 18340 30322 18396 30604
rect 18340 30270 18342 30322
rect 18394 30270 18396 30322
rect 18340 30212 18396 30270
rect 18340 30146 18396 30156
rect 18508 30324 18564 30334
rect 16716 29426 16772 29932
rect 17500 29922 17556 29932
rect 17836 30044 18228 30100
rect 16716 29374 16718 29426
rect 16770 29374 16772 29426
rect 16716 29362 16772 29374
rect 17556 29314 17612 29326
rect 17556 29262 17558 29314
rect 17610 29262 17612 29314
rect 17556 29204 17612 29262
rect 17444 29148 17556 29204
rect 17444 28756 17500 29148
rect 17556 29138 17612 29148
rect 17388 28754 17500 28756
rect 17388 28702 17446 28754
rect 17498 28702 17500 28754
rect 17388 28690 17500 28702
rect 16268 28642 16492 28644
rect 16268 28590 16270 28642
rect 16322 28590 16492 28642
rect 16268 28588 16492 28590
rect 16268 28578 16324 28588
rect 16436 28084 16492 28588
rect 16996 28420 17052 28430
rect 15596 27794 15652 27804
rect 15820 28082 16492 28084
rect 15820 28030 16438 28082
rect 16490 28030 16492 28082
rect 15820 28028 16492 28030
rect 15484 27022 15486 27074
rect 15538 27022 15540 27074
rect 14812 25622 14814 25674
rect 14866 25622 14868 25674
rect 14812 25610 14868 25622
rect 15036 26290 15092 26302
rect 15036 26238 15038 26290
rect 15090 26238 15092 26290
rect 14308 25508 14364 25518
rect 14308 25414 14364 25452
rect 14924 25508 14980 25518
rect 14924 25414 14980 25452
rect 14476 25396 14532 25406
rect 14476 25302 14532 25340
rect 15036 25396 15092 26238
rect 15484 26180 15540 27022
rect 15372 26068 15428 26078
rect 15148 25844 15204 25854
rect 15148 25506 15204 25788
rect 15148 25454 15150 25506
rect 15202 25454 15204 25506
rect 15148 25442 15204 25454
rect 15036 25330 15092 25340
rect 14140 25228 14308 25284
rect 14028 25106 14084 25116
rect 13692 24670 13694 24722
rect 13746 24670 13748 24722
rect 13468 23940 13524 23950
rect 13356 23938 13524 23940
rect 13356 23886 13470 23938
rect 13522 23886 13524 23938
rect 13356 23884 13524 23886
rect 13356 23154 13412 23884
rect 13468 23874 13524 23884
rect 13356 23102 13358 23154
rect 13410 23102 13412 23154
rect 13356 22372 13412 23102
rect 13356 20804 13412 22316
rect 13468 23604 13524 23614
rect 13468 22370 13524 23548
rect 13692 22932 13748 24670
rect 14252 24106 14308 25228
rect 14368 24760 14424 24772
rect 14368 24708 14370 24760
rect 14422 24708 14424 24760
rect 14368 24276 14424 24708
rect 14252 24054 14254 24106
rect 14306 24054 14308 24106
rect 14252 24042 14308 24054
rect 14364 24220 14424 24276
rect 15148 24722 15204 24734
rect 15148 24670 15150 24722
rect 15202 24670 15204 24722
rect 14140 23940 14196 23950
rect 14140 23846 14196 23884
rect 14364 23940 14420 24220
rect 14364 23874 14420 23884
rect 15148 24050 15204 24670
rect 15372 24724 15428 26012
rect 15484 25508 15540 26124
rect 15484 25442 15540 25452
rect 15596 27524 15652 27534
rect 15484 24948 15540 24958
rect 15596 24948 15652 27468
rect 15708 25508 15764 25518
rect 15708 25414 15764 25452
rect 15484 24946 15764 24948
rect 15484 24894 15486 24946
rect 15538 24894 15764 24946
rect 15484 24892 15764 24894
rect 15484 24882 15540 24892
rect 15372 24668 15652 24724
rect 15148 23998 15150 24050
rect 15202 23998 15204 24050
rect 15148 23940 15204 23998
rect 15148 23874 15204 23884
rect 13916 23380 13972 23390
rect 13916 23154 13972 23324
rect 13916 23102 13918 23154
rect 13970 23102 13972 23154
rect 13916 23090 13972 23102
rect 14028 23154 14084 23166
rect 14028 23102 14030 23154
rect 14082 23102 14084 23154
rect 13692 22876 13972 22932
rect 13748 22708 13804 22718
rect 13468 22318 13470 22370
rect 13522 22318 13524 22370
rect 13468 22306 13524 22318
rect 13580 22370 13636 22382
rect 13580 22318 13582 22370
rect 13634 22318 13636 22370
rect 13580 21924 13636 22318
rect 13748 22372 13804 22652
rect 13748 22370 13860 22372
rect 13748 22318 13750 22370
rect 13802 22318 13860 22370
rect 13748 22306 13860 22318
rect 13692 21924 13748 21934
rect 13580 21868 13692 21924
rect 13580 21586 13636 21598
rect 13580 21534 13582 21586
rect 13634 21534 13636 21586
rect 13580 21028 13636 21534
rect 13692 21586 13748 21868
rect 13692 21534 13694 21586
rect 13746 21534 13748 21586
rect 13804 21636 13860 22306
rect 13916 21812 13972 22876
rect 14028 22036 14084 23102
rect 14196 23154 14252 23166
rect 14196 23102 14198 23154
rect 14250 23102 14252 23154
rect 14196 22932 14252 23102
rect 14196 22866 14252 22876
rect 14588 22930 14644 22942
rect 14588 22878 14590 22930
rect 14642 22878 14644 22930
rect 14140 22482 14196 22494
rect 14140 22430 14142 22482
rect 14194 22430 14196 22482
rect 14140 22372 14196 22430
rect 14140 22306 14196 22316
rect 14028 21970 14084 21980
rect 13916 21756 14028 21812
rect 13972 21700 14028 21756
rect 14588 21700 14644 22878
rect 14700 22596 14756 22606
rect 14700 22502 14756 22540
rect 15372 22484 15428 22494
rect 15092 22372 15148 22382
rect 15092 22278 15148 22316
rect 15260 22370 15316 22382
rect 15260 22318 15262 22370
rect 15314 22318 15316 22370
rect 13972 21644 14084 21700
rect 13804 21624 13894 21636
rect 13804 21572 13840 21624
rect 13892 21572 13894 21624
rect 13804 21570 13894 21572
rect 13838 21560 13894 21570
rect 13692 21522 13748 21534
rect 14028 21364 14084 21644
rect 14588 21634 14644 21644
rect 14700 22148 14756 22158
rect 14700 21476 14756 22092
rect 15260 21924 15316 22318
rect 15372 22370 15428 22428
rect 15372 22318 15374 22370
rect 15426 22318 15428 22370
rect 15372 22148 15428 22318
rect 15372 22082 15428 22092
rect 15260 21868 15428 21924
rect 14588 21420 14756 21476
rect 14812 21812 14868 21822
rect 14812 21474 14868 21756
rect 15186 21700 15242 21710
rect 15186 21624 15242 21644
rect 15186 21572 15188 21624
rect 15240 21572 15242 21624
rect 15186 21560 15242 21572
rect 15372 21586 15428 21868
rect 15596 21700 15652 24668
rect 15708 22370 15764 24892
rect 15820 22596 15876 28028
rect 16436 28018 16492 28028
rect 16940 28418 17052 28420
rect 16940 28366 16998 28418
rect 17050 28366 17052 28418
rect 16940 28354 17052 28366
rect 16940 27860 16996 28354
rect 16940 27758 16996 27804
rect 16884 27746 16996 27758
rect 16884 27694 16886 27746
rect 16938 27694 16996 27746
rect 16884 27692 16996 27694
rect 16884 27412 16940 27692
rect 16492 27356 16940 27412
rect 16492 27300 16548 27356
rect 16156 27244 16548 27300
rect 16156 26908 16212 27244
rect 16268 27076 16324 27086
rect 16268 27074 16548 27076
rect 16268 27022 16270 27074
rect 16322 27022 16548 27074
rect 16268 27020 16548 27022
rect 16268 27010 16324 27020
rect 16156 26852 16268 26908
rect 16212 26178 16268 26852
rect 16492 26516 16548 27020
rect 17388 26908 17444 28690
rect 17720 28604 17776 28616
rect 17720 28552 17722 28604
rect 17774 28552 17776 28604
rect 17720 28532 17776 28552
rect 17720 28466 17776 28476
rect 17612 27634 17668 27646
rect 17612 27582 17614 27634
rect 17666 27582 17668 27634
rect 17612 27076 17668 27582
rect 17612 27010 17668 27020
rect 16828 26852 17444 26908
rect 16604 26516 16660 26526
rect 16492 26514 16660 26516
rect 16492 26462 16606 26514
rect 16658 26462 16660 26514
rect 16492 26460 16660 26462
rect 16604 26450 16660 26460
rect 16212 26126 16214 26178
rect 16266 26126 16268 26178
rect 16212 26068 16268 26126
rect 16212 26002 16268 26012
rect 16604 25956 16660 25966
rect 16492 25506 16548 25518
rect 16492 25454 16494 25506
rect 16546 25454 16548 25506
rect 16492 24948 16548 25454
rect 16492 24882 16548 24892
rect 16044 24724 16100 24734
rect 15932 24722 16100 24724
rect 15932 24670 16046 24722
rect 16098 24670 16100 24722
rect 15932 24668 16100 24670
rect 15932 23044 15988 24668
rect 16044 24658 16100 24668
rect 16380 24500 16436 24510
rect 16380 24406 16436 24444
rect 16604 24388 16660 25900
rect 16828 25844 16884 26852
rect 16940 26292 16996 26302
rect 16940 26198 16996 26236
rect 17556 26180 17612 26190
rect 17556 26086 17612 26124
rect 16716 25788 16884 25844
rect 16716 25060 16772 25788
rect 17836 25172 17892 30044
rect 17948 29652 18004 29662
rect 17948 29428 18004 29596
rect 18172 29428 18228 29438
rect 17948 29426 18116 29428
rect 17948 29374 17950 29426
rect 18002 29374 18116 29426
rect 17948 29372 18116 29374
rect 17948 29362 18004 29372
rect 18060 28644 18116 29372
rect 18172 29426 18340 29428
rect 18172 29374 18174 29426
rect 18226 29374 18340 29426
rect 18172 29372 18340 29374
rect 18172 29362 18228 29372
rect 18172 29258 18228 29270
rect 18172 29206 18174 29258
rect 18226 29206 18228 29258
rect 18172 28980 18228 29206
rect 18172 28914 18228 28924
rect 18284 28810 18340 29372
rect 18284 28758 18286 28810
rect 18338 28758 18340 28810
rect 18060 28588 18228 28644
rect 17948 28532 18004 28542
rect 17948 27858 18004 28476
rect 17948 27806 17950 27858
rect 18002 27806 18004 27858
rect 17948 27188 18004 27806
rect 18172 27690 18228 28588
rect 18284 28532 18340 28758
rect 18284 28466 18340 28476
rect 18396 28642 18452 28654
rect 18396 28590 18398 28642
rect 18450 28590 18452 28642
rect 18172 27638 18174 27690
rect 18226 27638 18228 27690
rect 18172 27626 18228 27638
rect 18284 27860 18340 27870
rect 18396 27860 18452 28590
rect 18340 27804 18452 27860
rect 18172 27188 18228 27198
rect 17948 27186 18228 27188
rect 17948 27134 18174 27186
rect 18226 27134 18228 27186
rect 17948 27132 18228 27134
rect 18172 27122 18228 27132
rect 18284 26908 18340 27804
rect 18508 27188 18564 30268
rect 18732 30210 18788 30828
rect 18732 30158 18734 30210
rect 18786 30158 18788 30210
rect 18732 30146 18788 30158
rect 18844 30548 18900 30558
rect 18844 30210 18900 30492
rect 18844 30158 18846 30210
rect 18898 30158 18900 30210
rect 18844 30146 18900 30158
rect 18844 29764 18900 29774
rect 18956 29764 19012 31948
rect 19124 30436 19180 30446
rect 19292 30436 19348 32508
rect 19404 33124 19460 33134
rect 19404 32618 19460 33068
rect 19404 32566 19406 32618
rect 19458 32566 19460 32618
rect 19404 32116 19460 32566
rect 19404 32050 19460 32060
rect 19124 30434 19348 30436
rect 19124 30382 19126 30434
rect 19178 30382 19348 30434
rect 19124 30380 19348 30382
rect 19404 31108 19460 31118
rect 19124 30370 19180 30380
rect 18956 29708 19236 29764
rect 18844 29540 18900 29708
rect 18956 29540 19012 29550
rect 18844 29538 19012 29540
rect 18844 29486 18958 29538
rect 19010 29486 19012 29538
rect 18844 29484 19012 29486
rect 18956 29474 19012 29484
rect 18620 29426 18676 29438
rect 18620 29374 18622 29426
rect 18674 29374 18676 29426
rect 19068 29426 19124 29438
rect 18620 28980 18676 29374
rect 18620 28914 18676 28924
rect 18788 29370 18844 29382
rect 18788 29318 18790 29370
rect 18842 29318 18844 29370
rect 18788 28868 18844 29318
rect 19068 29374 19070 29426
rect 19122 29374 19124 29426
rect 19068 29316 19124 29374
rect 18956 29260 19124 29316
rect 18956 29204 19012 29260
rect 19180 29204 19236 29708
rect 19404 29550 19460 31052
rect 19516 30884 19572 33292
rect 19628 33307 19684 33404
rect 19740 33458 19796 34300
rect 19740 33406 19742 33458
rect 19794 33406 19796 33458
rect 19740 33394 19796 33406
rect 19964 34157 20020 34300
rect 19964 34105 19966 34157
rect 20018 34105 20020 34157
rect 19628 33255 19630 33307
rect 19682 33255 19684 33307
rect 19628 33243 19684 33255
rect 19964 33124 20020 34105
rect 20076 33460 20132 33470
rect 20076 33346 20132 33404
rect 20076 33294 20078 33346
rect 20130 33294 20132 33346
rect 20076 33282 20132 33294
rect 19628 33068 20020 33124
rect 19628 31780 19684 33068
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19628 31714 19684 31724
rect 20188 32618 20244 32630
rect 20188 32566 20190 32618
rect 20242 32566 20244 32618
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 20188 31108 20244 32566
rect 20188 31042 20244 31052
rect 19516 30818 19572 30828
rect 20132 30884 20188 30894
rect 20132 30790 20188 30828
rect 20076 30548 20132 30558
rect 19516 30324 19572 30334
rect 19516 30177 19572 30268
rect 19516 30125 19518 30177
rect 19570 30125 19572 30177
rect 19516 30113 19572 30125
rect 19796 30154 19852 30166
rect 19796 30102 19798 30154
rect 19850 30102 19852 30154
rect 19796 30100 19852 30102
rect 19348 29538 19460 29550
rect 19348 29486 19350 29538
rect 19402 29486 19460 29538
rect 19348 29484 19460 29486
rect 19628 30044 19852 30100
rect 19628 29764 19684 30044
rect 20076 29988 20132 30492
rect 20300 30324 20356 34524
rect 20748 34186 20804 34862
rect 21084 34916 21140 34926
rect 21084 34356 21140 34860
rect 20580 34146 20636 34158
rect 20580 34132 20582 34146
rect 20412 34094 20582 34132
rect 20634 34094 20636 34146
rect 20412 34076 20636 34094
rect 20748 34134 20750 34186
rect 20802 34134 20804 34186
rect 20412 32004 20468 34076
rect 20748 33796 20804 34134
rect 20748 33730 20804 33740
rect 20860 34300 21140 34356
rect 21196 34356 21252 36764
rect 21364 36484 21420 36494
rect 21364 36390 21420 36428
rect 21308 36036 21364 36046
rect 21308 35588 21364 35980
rect 21532 35812 21588 37100
rect 21644 36482 21700 37324
rect 22316 37380 22372 37390
rect 22316 37322 22372 37324
rect 21756 37268 21812 37278
rect 22316 37270 22318 37322
rect 22370 37270 22372 37322
rect 21812 37212 21924 37268
rect 22316 37258 22372 37270
rect 21756 37174 21812 37212
rect 21644 36430 21646 36482
rect 21698 36430 21700 36482
rect 21644 36036 21700 36430
rect 21644 35970 21700 35980
rect 21756 37044 21812 37054
rect 21308 35522 21364 35532
rect 21420 35756 21588 35812
rect 21308 34356 21364 34366
rect 21196 34300 21308 34356
rect 20860 33684 20916 34300
rect 21084 34244 21140 34300
rect 21308 34290 21364 34300
rect 21084 34188 21252 34244
rect 21196 34186 21252 34188
rect 20972 34158 21028 34170
rect 20972 34132 20974 34158
rect 21026 34132 21028 34158
rect 21196 34134 21198 34186
rect 21250 34134 21252 34186
rect 21196 34122 21252 34134
rect 21420 34142 21476 35756
rect 21756 35698 21812 36988
rect 21868 36482 21924 37212
rect 22204 37156 22260 37166
rect 21868 36430 21870 36482
rect 21922 36430 21924 36482
rect 21868 36418 21924 36430
rect 21980 36484 22036 36494
rect 21980 36390 22036 36428
rect 22204 36482 22260 37100
rect 22428 36932 22484 37436
rect 22204 36430 22206 36482
rect 22258 36430 22260 36482
rect 22204 36418 22260 36430
rect 22316 36876 22484 36932
rect 22540 36932 22596 37884
rect 22652 37604 22708 38612
rect 22820 38276 22876 38286
rect 22820 38162 22876 38220
rect 22820 38110 22822 38162
rect 22874 38110 22876 38162
rect 22820 38098 22876 38110
rect 22652 37548 22820 37604
rect 22652 37268 22708 37278
rect 22652 37174 22708 37212
rect 22540 36876 22708 36932
rect 21756 35646 21758 35698
rect 21810 35646 21812 35698
rect 21588 35588 21644 35598
rect 21588 35494 21644 35532
rect 21756 35140 21812 35646
rect 21868 36036 21924 36046
rect 21868 35364 21924 35980
rect 21868 35298 21924 35308
rect 21980 35252 22036 35262
rect 21644 35082 21700 35094
rect 21756 35084 21924 35140
rect 21644 35030 21646 35082
rect 21698 35030 21700 35082
rect 21420 34130 21532 34142
rect 21420 34078 21478 34130
rect 21530 34078 21532 34130
rect 21420 34076 21532 34078
rect 20972 34066 21028 34076
rect 21476 34066 21532 34076
rect 21644 34132 21700 35030
rect 21756 34916 21812 34926
rect 21756 34822 21812 34860
rect 21868 34692 21924 35084
rect 21980 34914 22036 35196
rect 21980 34862 21982 34914
rect 22034 34862 22036 34914
rect 21980 34850 22036 34862
rect 21644 34066 21700 34076
rect 21756 34636 21924 34692
rect 21532 33908 21588 33918
rect 21364 33796 21420 33806
rect 20860 33628 21028 33684
rect 20804 33122 20860 33134
rect 20804 33070 20806 33122
rect 20858 33070 20860 33122
rect 20804 33012 20860 33070
rect 20412 31938 20468 31948
rect 20524 32956 20804 33012
rect 20524 31780 20580 32956
rect 20804 32946 20860 32956
rect 20748 32564 20804 32574
rect 20748 32470 20804 32508
rect 20524 31778 20692 31780
rect 20524 31726 20526 31778
rect 20578 31726 20692 31778
rect 20524 31724 20692 31726
rect 20524 31714 20580 31724
rect 20412 31108 20468 31118
rect 20412 30994 20468 31052
rect 20412 30942 20414 30994
rect 20466 30942 20468 30994
rect 20412 30930 20468 30942
rect 20524 30994 20580 31006
rect 20524 30942 20526 30994
rect 20578 30942 20580 30994
rect 20524 30772 20580 30942
rect 20524 30706 20580 30716
rect 20636 30996 20692 31724
rect 20636 30324 20692 30940
rect 20300 30268 20580 30324
rect 20524 30182 20580 30268
rect 20748 31220 20804 31230
rect 20972 31220 21028 33628
rect 21364 33178 21420 33740
rect 21364 33126 21366 33178
rect 21418 33126 21420 33178
rect 21364 33114 21420 33126
rect 21532 33346 21588 33852
rect 21756 33348 21812 34636
rect 22316 34468 22372 36876
rect 22484 36708 22540 36718
rect 22484 36614 22540 36652
rect 22428 35588 22484 35598
rect 22428 35364 22484 35532
rect 22428 35298 22484 35308
rect 22540 35586 22596 35598
rect 22540 35534 22542 35586
rect 22594 35534 22596 35586
rect 22428 35140 22484 35150
rect 22428 34692 22484 35084
rect 22540 34916 22596 35534
rect 22540 34850 22596 34860
rect 22652 34860 22708 36876
rect 22764 36484 22820 37548
rect 23100 37268 23156 41692
rect 23212 41188 23268 41198
rect 23212 41094 23268 41132
rect 23324 41186 23380 41916
rect 23660 41970 23828 41972
rect 23660 41918 23774 41970
rect 23826 41918 23828 41970
rect 23660 41916 23828 41918
rect 23324 41134 23326 41186
rect 23378 41134 23380 41186
rect 23324 41122 23380 41134
rect 23436 41748 23492 41758
rect 23436 40964 23492 41692
rect 23548 41186 23604 41198
rect 23548 41134 23550 41186
rect 23602 41134 23604 41186
rect 23548 41076 23604 41134
rect 23548 41010 23604 41020
rect 23324 40908 23492 40964
rect 23324 40740 23380 40908
rect 23324 38276 23380 40684
rect 23492 40292 23548 40302
rect 23660 40292 23716 41916
rect 23772 41906 23828 41916
rect 23996 41300 24052 41310
rect 23828 41188 23884 41198
rect 23828 41094 23884 41132
rect 23436 40290 23716 40292
rect 23436 40238 23494 40290
rect 23546 40238 23716 40290
rect 23436 40236 23716 40238
rect 23436 40226 23548 40236
rect 23436 39182 23492 40226
rect 23884 40180 23940 40190
rect 23660 40178 23940 40180
rect 23660 40126 23886 40178
rect 23938 40126 23940 40178
rect 23660 40124 23940 40126
rect 23548 39732 23604 39742
rect 23660 39732 23716 40124
rect 23884 40114 23940 40124
rect 23996 39956 24052 41244
rect 24108 41188 24164 42140
rect 24556 42138 24612 42476
rect 24556 42086 24558 42138
rect 24610 42086 24612 42138
rect 24556 42074 24612 42086
rect 24892 42308 24948 42318
rect 24220 42009 24276 42021
rect 24220 41957 24222 42009
rect 24274 41957 24276 42009
rect 24220 41300 24276 41957
rect 24444 41972 24500 41982
rect 24444 41878 24500 41916
rect 24780 41636 24836 41646
rect 24668 41300 24724 41310
rect 24220 41298 24724 41300
rect 24220 41246 24670 41298
rect 24722 41246 24724 41298
rect 24220 41244 24724 41246
rect 24668 41234 24724 41244
rect 24108 41132 24332 41188
rect 24276 41018 24332 41132
rect 24780 41171 24836 41580
rect 24780 41119 24782 41171
rect 24834 41119 24836 41171
rect 24780 41107 24836 41119
rect 24276 40966 24278 41018
rect 24330 40966 24332 41018
rect 24276 40954 24332 40966
rect 24724 40628 24780 40638
rect 24780 40572 24836 40628
rect 24724 40534 24836 40572
rect 23548 39730 23716 39732
rect 23548 39678 23550 39730
rect 23602 39678 23716 39730
rect 23548 39676 23716 39678
rect 23772 39900 24052 39956
rect 24220 40402 24276 40414
rect 24220 40350 24222 40402
rect 24274 40350 24276 40402
rect 24220 39956 24276 40350
rect 24220 39900 24724 39956
rect 23548 39666 23604 39676
rect 23660 39508 23716 39518
rect 23660 39284 23716 39452
rect 23772 39396 23828 39900
rect 24668 39396 24724 39900
rect 23772 39340 23940 39396
rect 23660 39218 23716 39228
rect 23436 39172 23548 39182
rect 23436 39116 23492 39172
rect 23492 39060 23548 39116
rect 23492 39058 23828 39060
rect 23492 39006 23494 39058
rect 23546 39006 23828 39058
rect 23492 39004 23828 39006
rect 23492 38994 23548 39004
rect 23772 38834 23828 39004
rect 23884 38948 23940 39340
rect 24556 39340 24724 39396
rect 24444 39284 24500 39294
rect 23884 38892 24108 38948
rect 23772 38782 23774 38834
rect 23826 38782 23828 38834
rect 24052 38890 24108 38892
rect 24052 38838 24054 38890
rect 24106 38838 24108 38890
rect 24052 38826 24108 38838
rect 24444 38834 24500 39228
rect 24556 39002 24612 39340
rect 24556 38950 24558 39002
rect 24610 38950 24612 39002
rect 24556 38938 24612 38950
rect 23772 38770 23828 38782
rect 24444 38782 24446 38834
rect 24498 38782 24500 38834
rect 24444 38770 24500 38782
rect 23996 38724 24052 38734
rect 23212 38164 23268 38174
rect 23212 38070 23268 38108
rect 23044 37212 23156 37268
rect 23044 37210 23100 37212
rect 22876 37156 22932 37166
rect 22876 37062 22932 37100
rect 23044 37158 23046 37210
rect 23098 37158 23100 37210
rect 23044 36932 23100 37158
rect 22988 36876 23100 36932
rect 22876 36484 22932 36494
rect 22764 36482 22932 36484
rect 22764 36430 22878 36482
rect 22930 36430 22932 36482
rect 22764 36428 22932 36430
rect 22876 36418 22932 36428
rect 22988 36260 23044 36876
rect 23324 36820 23380 38220
rect 23548 38500 23604 38510
rect 23548 38050 23604 38444
rect 23548 37998 23550 38050
rect 23602 37998 23604 38050
rect 23548 37986 23604 37998
rect 23660 38164 23716 38174
rect 23660 38050 23716 38108
rect 23660 37998 23662 38050
rect 23714 37998 23716 38050
rect 23660 37986 23716 37998
rect 23996 37826 24052 38668
rect 24612 38500 24668 38510
rect 24612 38162 24668 38444
rect 24612 38110 24614 38162
rect 24666 38110 24668 38162
rect 24612 38098 24668 38110
rect 23996 37774 23998 37826
rect 24050 37774 24052 37826
rect 23492 37154 23548 37166
rect 23884 37156 23940 37166
rect 23492 37102 23494 37154
rect 23546 37102 23548 37154
rect 23492 37044 23548 37102
rect 23492 36978 23548 36988
rect 23660 37154 23940 37156
rect 23660 37102 23886 37154
rect 23938 37102 23940 37154
rect 23660 37100 23940 37102
rect 23324 36764 23604 36820
rect 22764 36204 23044 36260
rect 22764 35140 22820 36204
rect 23548 35924 23604 36764
rect 23660 36594 23716 37100
rect 23884 37090 23940 37100
rect 23996 36932 24052 37774
rect 24220 37940 24276 37950
rect 24220 37266 24276 37884
rect 24780 37380 24836 40534
rect 24780 37314 24836 37324
rect 24220 37214 24222 37266
rect 24274 37214 24276 37266
rect 24220 37202 24276 37214
rect 23660 36542 23662 36594
rect 23714 36542 23716 36594
rect 23660 36530 23716 36542
rect 23772 36876 24052 36932
rect 24724 37156 24780 37166
rect 24892 37156 24948 42252
rect 25228 41970 25284 43250
rect 25452 42866 25508 43486
rect 25452 42814 25454 42866
rect 25506 42814 25508 42866
rect 25452 42756 25508 42814
rect 25452 42690 25508 42700
rect 25564 42308 25620 43708
rect 25900 43540 25956 43578
rect 25900 43474 25956 43484
rect 26572 42978 26628 43820
rect 26776 43550 26832 43596
rect 26776 43540 26852 43550
rect 26776 43538 26796 43540
rect 26776 43486 26778 43538
rect 26776 43484 26796 43486
rect 26776 43474 26852 43484
rect 26572 42926 26574 42978
rect 26626 42926 26628 42978
rect 26572 42914 26628 42926
rect 25900 42756 25956 42766
rect 25900 42662 25956 42700
rect 26012 42754 26068 42766
rect 26012 42702 26014 42754
rect 26066 42702 26068 42754
rect 25564 42252 25956 42308
rect 25228 41918 25230 41970
rect 25282 41918 25284 41970
rect 25228 41906 25284 41918
rect 25900 41412 25956 42252
rect 26012 42196 26068 42702
rect 26178 42698 26236 42756
rect 26178 42646 26180 42698
rect 26232 42646 26236 42698
rect 26178 42634 26236 42646
rect 26180 42308 26236 42634
rect 26180 42252 26292 42308
rect 26012 42140 26160 42196
rect 26104 41970 26160 42140
rect 26104 41918 26106 41970
rect 26158 41918 26160 41970
rect 26104 41860 26160 41918
rect 26236 41972 26292 42252
rect 26796 42084 26852 43474
rect 26908 43092 26964 44716
rect 27020 44660 27076 44670
rect 27020 44322 27076 44604
rect 27020 44270 27022 44322
rect 27074 44270 27076 44322
rect 27020 44258 27076 44270
rect 27244 44436 27300 45500
rect 27580 45220 27636 45614
rect 27580 45154 27636 45164
rect 27804 44772 27860 45836
rect 27916 45826 27972 45836
rect 28252 45890 28420 45892
rect 28252 45838 28366 45890
rect 28418 45838 28420 45890
rect 28252 45836 28420 45838
rect 27916 44996 27972 45006
rect 27916 44902 27972 44940
rect 28252 44996 28308 45836
rect 28364 45826 28420 45836
rect 28700 45892 28756 45902
rect 29372 45892 29428 45948
rect 29484 45892 29540 45902
rect 29708 45892 29764 45902
rect 28700 45890 29092 45892
rect 28700 45838 28702 45890
rect 28754 45838 29092 45890
rect 28700 45836 29092 45838
rect 29372 45890 29540 45892
rect 29372 45838 29486 45890
rect 29538 45838 29540 45890
rect 29372 45836 29540 45838
rect 28700 45826 28756 45836
rect 28252 44930 28308 44940
rect 28364 45444 28420 45454
rect 27804 44706 27860 44716
rect 27244 44322 27300 44380
rect 27244 44270 27246 44322
rect 27298 44270 27300 44322
rect 27244 44258 27300 44270
rect 27916 44322 27972 44334
rect 27916 44270 27918 44322
rect 27970 44270 27972 44322
rect 27804 44212 27860 44222
rect 27580 44098 27636 44110
rect 27580 44046 27582 44098
rect 27634 44046 27636 44098
rect 27580 43876 27636 44046
rect 27580 43810 27636 43820
rect 27804 43652 27860 44156
rect 27916 44100 27972 44270
rect 28196 44324 28252 44334
rect 28364 44324 28420 45388
rect 28868 45106 28924 45118
rect 28868 45054 28870 45106
rect 28922 45054 28924 45106
rect 28476 44884 28532 44894
rect 28476 44882 28644 44884
rect 28476 44830 28478 44882
rect 28530 44830 28644 44882
rect 28476 44828 28644 44830
rect 28476 44818 28532 44828
rect 28476 44324 28532 44334
rect 28364 44322 28532 44324
rect 28364 44270 28478 44322
rect 28530 44270 28532 44322
rect 28364 44268 28532 44270
rect 28196 44230 28252 44268
rect 28476 44258 28532 44268
rect 28588 44322 28644 44828
rect 28868 44660 28924 45054
rect 28868 44594 28924 44604
rect 29036 45106 29092 45836
rect 29484 45826 29540 45836
rect 29596 45836 29708 45892
rect 29204 45778 29260 45790
rect 29204 45726 29206 45778
rect 29258 45726 29260 45778
rect 29204 45556 29260 45726
rect 29204 45490 29260 45500
rect 29036 45054 29038 45106
rect 29090 45054 29092 45106
rect 28588 44270 28590 44322
rect 28642 44270 28644 44322
rect 28588 44258 28644 44270
rect 27916 44034 27972 44044
rect 28364 44100 28420 44110
rect 29036 44100 29092 45054
rect 29148 45106 29204 45118
rect 29148 45054 29150 45106
rect 29202 45054 29204 45106
rect 29148 44996 29204 45054
rect 29148 44322 29204 44940
rect 29596 44558 29652 45836
rect 29708 45798 29764 45836
rect 29708 45108 29764 45118
rect 29708 45014 29764 45052
rect 29820 44772 29876 49308
rect 30240 49200 30352 50000
rect 31808 49200 31920 50000
rect 33376 49200 33488 50000
rect 34944 49200 35056 50000
rect 36512 49200 36624 50000
rect 38080 49200 38192 50000
rect 39648 49200 39760 50000
rect 41216 49200 41328 50000
rect 42784 49200 42896 50000
rect 44352 49200 44464 50000
rect 45920 49200 46032 50000
rect 30156 47012 30212 47022
rect 29988 45778 30044 45790
rect 29988 45726 29990 45778
rect 30042 45726 30044 45778
rect 29988 45444 30044 45726
rect 29988 45378 30044 45388
rect 29820 44716 30044 44772
rect 29540 44546 29652 44558
rect 29540 44494 29542 44546
rect 29594 44494 29652 44546
rect 29540 44492 29652 44494
rect 29540 44482 29596 44492
rect 29148 44270 29150 44322
rect 29202 44270 29204 44322
rect 29148 44258 29204 44270
rect 29260 44322 29316 44334
rect 29260 44270 29262 44322
rect 29314 44270 29316 44322
rect 29260 44100 29316 44270
rect 29036 44044 29316 44100
rect 29988 44154 30044 44716
rect 29988 44102 29990 44154
rect 30042 44102 30044 44154
rect 29988 44090 30044 44102
rect 27804 43586 27860 43596
rect 28084 43594 28140 43606
rect 27356 43540 27412 43550
rect 27356 43446 27412 43484
rect 27692 43540 27748 43550
rect 27692 43446 27748 43484
rect 28084 43542 28086 43594
rect 28138 43542 28140 43594
rect 27020 43316 27076 43326
rect 27020 43314 27188 43316
rect 27020 43262 27022 43314
rect 27074 43262 27188 43314
rect 27020 43260 27188 43262
rect 27020 43250 27076 43260
rect 26908 43036 27076 43092
rect 26796 42018 26852 42028
rect 26236 41906 26292 41916
rect 26684 41970 26740 41982
rect 26684 41918 26686 41970
rect 26738 41918 26740 41970
rect 26104 41794 26160 41804
rect 26348 41748 26404 41758
rect 26684 41748 26740 41918
rect 26348 41746 26740 41748
rect 26348 41694 26350 41746
rect 26402 41694 26740 41746
rect 26348 41692 26740 41694
rect 26908 41970 26964 41982
rect 26908 41918 26910 41970
rect 26962 41918 26964 41970
rect 25788 41356 25956 41412
rect 26124 41636 26180 41646
rect 25452 41300 25508 41310
rect 25452 41206 25508 41244
rect 25116 41188 25172 41198
rect 25116 41094 25172 41132
rect 25564 41142 25620 41154
rect 25564 41090 25566 41142
rect 25618 41090 25620 41142
rect 25564 40628 25620 41090
rect 25340 40572 25620 40628
rect 25788 40628 25844 41356
rect 25340 40180 25396 40572
rect 25788 40562 25844 40572
rect 25900 41186 25956 41198
rect 25900 41134 25902 41186
rect 25954 41134 25956 41186
rect 25710 40439 25766 40451
rect 25340 40114 25396 40124
rect 25452 40402 25508 40414
rect 25452 40350 25454 40402
rect 25506 40350 25508 40402
rect 25452 39732 25508 40350
rect 25228 39730 25508 39732
rect 25228 39678 25454 39730
rect 25506 39678 25508 39730
rect 25228 39676 25508 39678
rect 25004 38948 25060 38958
rect 25004 38276 25060 38892
rect 25228 38834 25284 39676
rect 25452 39666 25508 39676
rect 25564 40402 25620 40414
rect 25710 40404 25712 40439
rect 25564 40350 25566 40402
rect 25618 40350 25620 40402
rect 25564 39172 25620 40350
rect 25676 40387 25712 40404
rect 25764 40387 25766 40439
rect 25676 40348 25766 40387
rect 25676 40292 25732 40348
rect 25676 39284 25732 40236
rect 25788 40180 25844 40190
rect 25788 39844 25844 40124
rect 25900 39956 25956 41134
rect 26124 40290 26180 41580
rect 26348 41188 26404 41692
rect 26908 41636 26964 41918
rect 27020 41748 27076 43036
rect 27132 42756 27188 43260
rect 28084 43204 28140 43542
rect 28252 43568 28308 43580
rect 28252 43540 28254 43568
rect 28306 43540 28308 43568
rect 28252 43474 28308 43484
rect 28084 43138 28140 43148
rect 28232 43316 28288 43326
rect 27356 42756 27412 42766
rect 27132 42754 27412 42756
rect 27132 42702 27358 42754
rect 27410 42702 27412 42754
rect 27132 42700 27412 42702
rect 27356 42690 27412 42700
rect 28232 42754 28288 43260
rect 28232 42702 28234 42754
rect 28286 42702 28288 42754
rect 28232 42690 28288 42702
rect 27636 42026 27692 42038
rect 27188 41972 27244 41982
rect 27188 41878 27244 41916
rect 27636 41974 27638 42026
rect 27690 41974 27692 42026
rect 27468 41860 27524 41870
rect 27468 41748 27524 41804
rect 27020 41692 27300 41748
rect 26908 41570 26964 41580
rect 26348 41122 26404 41132
rect 26572 41188 26628 41198
rect 26572 41094 26628 41132
rect 27132 40740 27188 40750
rect 26460 40402 26516 40414
rect 26460 40350 26462 40402
rect 26514 40350 26516 40402
rect 26460 40292 26516 40350
rect 26124 40238 26126 40290
rect 26178 40238 26180 40290
rect 26124 40226 26180 40238
rect 26236 40236 26516 40292
rect 26684 40402 26740 40414
rect 26684 40350 26686 40402
rect 26738 40350 26740 40402
rect 26236 39956 26292 40236
rect 26684 40180 26740 40350
rect 26964 40292 27020 40302
rect 26964 40198 27020 40236
rect 26684 40114 26740 40124
rect 27132 40068 27188 40684
rect 25900 39900 26292 39956
rect 26908 40012 27188 40068
rect 25788 39788 25956 39844
rect 25676 39218 25732 39228
rect 25564 39106 25620 39116
rect 25228 38782 25230 38834
rect 25282 38782 25284 38834
rect 25228 38770 25284 38782
rect 25452 38388 25508 38398
rect 25340 38276 25396 38286
rect 25004 38220 25228 38276
rect 25172 38164 25228 38220
rect 25172 38162 25284 38164
rect 25172 38110 25174 38162
rect 25226 38110 25284 38162
rect 25172 38098 25284 38110
rect 24724 37154 24948 37156
rect 24724 37102 24726 37154
rect 24778 37102 24948 37154
rect 24724 37100 24948 37102
rect 23548 35868 23716 35924
rect 22764 35074 22820 35084
rect 22876 35364 22932 35374
rect 22876 34914 22932 35308
rect 23324 35252 23380 35262
rect 23324 35138 23380 35196
rect 23324 35086 23326 35138
rect 23378 35086 23380 35138
rect 23324 35074 23380 35086
rect 22876 34862 22878 34914
rect 22930 34862 22932 34914
rect 22652 34748 22722 34860
rect 22876 34850 22932 34862
rect 22988 34914 23044 34926
rect 22988 34862 22990 34914
rect 23042 34862 23044 34914
rect 22540 34692 22596 34702
rect 22428 34690 22596 34692
rect 22428 34638 22542 34690
rect 22594 34638 22596 34690
rect 22428 34636 22596 34638
rect 22540 34626 22596 34636
rect 22652 34580 22708 34748
rect 22652 34524 22820 34580
rect 22316 34412 22652 34468
rect 21868 34244 21924 34254
rect 21868 34130 21924 34188
rect 22596 34242 22652 34412
rect 22596 34190 22598 34242
rect 22650 34190 22652 34242
rect 22596 34178 22652 34190
rect 21868 34078 21870 34130
rect 21922 34078 21924 34130
rect 22204 34130 22260 34142
rect 21868 34066 21924 34078
rect 22036 34074 22092 34086
rect 22036 34022 22038 34074
rect 22090 34022 22092 34074
rect 22036 34020 22092 34022
rect 21980 33964 22036 34020
rect 21980 33954 22092 33964
rect 22204 34078 22206 34130
rect 22258 34078 22260 34130
rect 21532 33294 21534 33346
rect 21586 33294 21588 33346
rect 21196 32788 21252 32798
rect 21196 32674 21252 32732
rect 21532 32676 21588 33294
rect 21644 33346 21812 33348
rect 21644 33294 21758 33346
rect 21810 33294 21812 33346
rect 21644 33292 21812 33294
rect 21644 33012 21700 33292
rect 21756 33282 21812 33292
rect 21868 33908 21924 33918
rect 21868 33348 21924 33852
rect 21868 33282 21924 33292
rect 21644 32946 21700 32956
rect 21196 32622 21198 32674
rect 21250 32622 21252 32674
rect 21196 32610 21252 32622
rect 21420 32620 21588 32676
rect 21868 32620 21924 32630
rect 21980 32620 22036 33954
rect 22204 33908 22260 34078
rect 22204 33842 22260 33852
rect 22316 34130 22372 34142
rect 22316 34078 22318 34130
rect 22370 34078 22372 34130
rect 22316 33796 22372 34078
rect 22316 33730 22372 33740
rect 22428 34132 22484 34142
rect 21308 31778 21364 31790
rect 21308 31726 21310 31778
rect 21362 31726 21364 31778
rect 21308 31668 21364 31726
rect 21308 31602 21364 31612
rect 21420 31778 21476 32620
rect 21868 32618 22036 32620
rect 21868 32566 21870 32618
rect 21922 32566 22036 32618
rect 21868 32564 22036 32566
rect 21868 32554 21924 32564
rect 21980 32116 22036 32564
rect 21980 32050 22036 32060
rect 22204 33684 22260 33694
rect 21980 31892 22036 31902
rect 21980 31798 22036 31836
rect 21420 31726 21422 31778
rect 21474 31726 21476 31778
rect 21420 31444 21476 31726
rect 20748 30994 20804 31164
rect 20748 30942 20750 30994
rect 20802 30942 20804 30994
rect 20748 30324 20804 30942
rect 20860 31164 21028 31220
rect 21252 31388 21476 31444
rect 21586 31722 21642 31734
rect 21586 31670 21588 31722
rect 21640 31670 21642 31722
rect 20860 30660 20916 31164
rect 21252 31106 21308 31388
rect 21586 31108 21642 31670
rect 22204 31668 22260 33628
rect 22428 32676 22484 34076
rect 22540 33908 22596 33918
rect 22540 33458 22596 33852
rect 22540 33406 22542 33458
rect 22594 33406 22596 33458
rect 22540 33394 22596 33406
rect 22764 33012 22820 34524
rect 22988 33684 23044 34862
rect 23660 34468 23716 35868
rect 23660 34402 23716 34412
rect 23772 34356 23828 36876
rect 24724 36820 24780 37100
rect 23772 34290 23828 34300
rect 23884 36764 24780 36820
rect 23660 34130 23716 34142
rect 23660 34078 23662 34130
rect 23714 34078 23716 34130
rect 23548 34020 23604 34030
rect 23324 33908 23380 33918
rect 23324 33814 23380 33852
rect 23548 33796 23604 33964
rect 23660 33908 23716 34078
rect 23772 34132 23828 34142
rect 23772 34038 23828 34076
rect 23772 33908 23828 33918
rect 23660 33852 23772 33908
rect 23772 33842 23828 33852
rect 23884 33796 23940 36764
rect 24444 35588 24500 35598
rect 24332 35532 24444 35588
rect 24332 34914 24388 35532
rect 24444 35494 24500 35532
rect 24332 34862 24334 34914
rect 24386 34862 24388 34914
rect 24332 34850 24388 34862
rect 24556 34914 24612 34926
rect 24556 34862 24558 34914
rect 24610 34862 24612 34914
rect 24164 34692 24220 34702
rect 24556 34692 24612 34862
rect 24164 34690 24612 34692
rect 24164 34638 24166 34690
rect 24218 34638 24612 34690
rect 24164 34636 24612 34638
rect 24164 34626 24220 34636
rect 25116 34468 25172 34478
rect 23996 34132 24052 34142
rect 23996 34130 25060 34132
rect 23996 34078 23998 34130
rect 24050 34078 25060 34130
rect 23996 34076 25060 34078
rect 23996 34066 24052 34076
rect 24276 33908 24332 33918
rect 24276 33814 24332 33852
rect 23548 33740 23716 33796
rect 23884 33740 24052 33796
rect 22988 33618 23044 33628
rect 22764 32956 23156 33012
rect 22708 32676 22764 32686
rect 22428 32674 22764 32676
rect 22428 32622 22710 32674
rect 22762 32622 22764 32674
rect 22428 32620 22764 32622
rect 22708 32610 22764 32620
rect 22988 32562 23044 32574
rect 22988 32510 22990 32562
rect 23042 32510 23044 32562
rect 22372 32452 22428 32462
rect 22372 32450 22484 32452
rect 22372 32398 22374 32450
rect 22426 32398 22484 32450
rect 22372 32386 22484 32398
rect 22092 31612 22204 31668
rect 21252 31054 21254 31106
rect 21306 31054 21308 31106
rect 21252 31042 21308 31054
rect 21532 31052 21642 31108
rect 21756 31108 21812 31118
rect 20972 30994 21028 31006
rect 20972 30942 20974 30994
rect 21026 30942 21028 30994
rect 20972 30884 21028 30942
rect 21532 30884 21588 31052
rect 20972 30818 21028 30828
rect 21084 30828 21588 30884
rect 21756 30994 21812 31052
rect 21756 30942 21758 30994
rect 21810 30942 21812 30994
rect 20860 30594 20916 30604
rect 20748 30268 20916 30324
rect 20636 30258 20692 30268
rect 20524 30170 20624 30182
rect 20412 30154 20468 30166
rect 20412 30102 20414 30154
rect 20466 30102 20468 30154
rect 20412 30100 20468 30102
rect 20300 30044 20412 30100
rect 20524 30118 20570 30170
rect 20622 30118 20624 30170
rect 20524 30100 20624 30118
rect 20524 30044 20692 30100
rect 20076 29932 20244 29988
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19348 29474 19404 29484
rect 18956 29138 19012 29148
rect 19068 29148 19236 29204
rect 19404 29204 19460 29214
rect 18900 28868 18956 28878
rect 18788 28866 18956 28868
rect 18788 28814 18902 28866
rect 18954 28814 18956 28866
rect 18788 28812 18956 28814
rect 18900 28802 18956 28812
rect 19068 28756 19124 29148
rect 19068 28700 19348 28756
rect 19068 28642 19124 28700
rect 19068 28590 19070 28642
rect 19122 28590 19124 28642
rect 19068 28578 19124 28590
rect 19180 28532 19236 28542
rect 18960 27896 19016 27908
rect 18960 27844 18962 27896
rect 19014 27844 19016 27896
rect 18960 27412 19016 27844
rect 19180 27858 19236 28476
rect 19180 27806 19182 27858
rect 19234 27806 19236 27858
rect 19180 27794 19236 27806
rect 18508 27122 18564 27132
rect 18620 27356 19016 27412
rect 18620 27074 18676 27356
rect 18620 27022 18622 27074
rect 18674 27022 18676 27074
rect 18620 27010 18676 27022
rect 18508 26964 18564 26974
rect 18284 26852 18452 26908
rect 18508 26852 18676 26908
rect 18396 26628 18452 26852
rect 18396 26562 18452 26572
rect 18322 26327 18378 26339
rect 17948 26292 18004 26302
rect 17948 26178 18004 26236
rect 17948 26126 17950 26178
rect 18002 26126 18004 26178
rect 17948 26114 18004 26126
rect 18322 26275 18324 26327
rect 18376 26275 18378 26327
rect 18322 25844 18378 26275
rect 16716 24994 16772 25004
rect 17388 25116 17892 25172
rect 18284 25788 18378 25844
rect 18508 26290 18564 26302
rect 18508 26238 18510 26290
rect 18562 26238 18564 26290
rect 16604 24322 16660 24332
rect 17052 24500 17108 24510
rect 17052 24050 17108 24444
rect 17052 23998 17054 24050
rect 17106 23998 17108 24050
rect 17052 23986 17108 23998
rect 16438 23156 16494 23166
rect 16436 23154 16494 23156
rect 16436 23102 16440 23154
rect 16492 23102 16494 23154
rect 16436 23090 16494 23102
rect 16604 23154 16660 23166
rect 16604 23102 16606 23154
rect 16658 23102 16660 23154
rect 16044 23044 16100 23054
rect 15932 23042 16100 23044
rect 15932 22990 16046 23042
rect 16098 22990 16100 23042
rect 15932 22988 16100 22990
rect 16044 22978 16100 22988
rect 16436 22606 16492 23090
rect 15820 22540 16324 22596
rect 15708 22318 15710 22370
rect 15762 22318 15764 22370
rect 15708 22306 15764 22318
rect 15820 22370 15876 22382
rect 15820 22318 15822 22370
rect 15874 22318 15876 22370
rect 15820 22260 15876 22318
rect 15988 22372 16044 22382
rect 15988 22278 16044 22316
rect 15820 21924 15876 22204
rect 15820 21858 15876 21868
rect 16156 21812 16212 21822
rect 15596 21644 15876 21700
rect 15372 21534 15374 21586
rect 15426 21534 15428 21586
rect 15372 21476 15428 21534
rect 14812 21422 14814 21474
rect 14866 21422 14868 21474
rect 13580 20962 13636 20972
rect 13692 21308 14084 21364
rect 14252 21362 14308 21374
rect 14252 21310 14254 21362
rect 14306 21310 14308 21362
rect 13020 20018 13188 20020
rect 13020 19966 13022 20018
rect 13074 19966 13188 20018
rect 13020 19964 13188 19966
rect 13244 20802 13412 20804
rect 13244 20750 13358 20802
rect 13410 20750 13412 20802
rect 13244 20748 13412 20750
rect 12852 19796 12908 19806
rect 12124 19234 12628 19236
rect 12124 19182 12126 19234
rect 12178 19182 12462 19234
rect 12514 19182 12628 19234
rect 12124 19180 12628 19182
rect 12684 19794 12908 19796
rect 12684 19742 12854 19794
rect 12906 19742 12908 19794
rect 12684 19740 12908 19742
rect 12124 19170 12180 19180
rect 12460 19170 12516 19180
rect 11676 19058 11732 19068
rect 12236 18676 12292 18686
rect 12124 18228 12180 18238
rect 12012 18226 12180 18228
rect 12012 18174 12126 18226
rect 12178 18174 12180 18226
rect 12012 18172 12180 18174
rect 10892 17668 10948 17678
rect 10892 17666 11172 17668
rect 10892 17614 10894 17666
rect 10946 17614 11172 17666
rect 10892 17612 11172 17614
rect 10892 17602 10948 17612
rect 11116 17108 11172 17612
rect 11116 17052 11396 17108
rect 11340 15540 11396 17052
rect 11788 16884 11844 16894
rect 11340 15474 11396 15484
rect 11564 16660 11620 16670
rect 10332 15362 10388 15372
rect 10220 15138 10276 15148
rect 10332 15258 10388 15270
rect 10332 15206 10334 15258
rect 10386 15206 10388 15258
rect 10332 15092 10388 15206
rect 10332 15026 10388 15036
rect 10108 14914 10164 14924
rect 10614 14868 10670 14878
rect 10220 14644 10276 14654
rect 9660 14590 9662 14642
rect 9714 14590 9716 14642
rect 9660 14578 9716 14590
rect 9996 14642 10276 14644
rect 9996 14590 10222 14642
rect 10274 14590 10276 14642
rect 9996 14588 10276 14590
rect 9828 14474 9884 14486
rect 9828 14422 9830 14474
rect 9882 14422 9884 14474
rect 9828 13972 9884 14422
rect 9996 13972 10052 14588
rect 10220 14578 10276 14588
rect 10332 14532 10388 14542
rect 9772 13916 9884 13972
rect 9940 13916 10052 13972
rect 10108 14308 10164 14318
rect 9548 13412 9604 13580
rect 9660 13636 9716 13646
rect 9772 13636 9828 13916
rect 9940 13860 9996 13916
rect 10108 13860 10164 14252
rect 9660 13634 9828 13636
rect 9660 13582 9662 13634
rect 9714 13582 9828 13634
rect 9660 13580 9828 13582
rect 9884 13804 9996 13860
rect 10074 13804 10164 13860
rect 9660 13570 9716 13580
rect 9548 13356 9716 13412
rect 9436 12850 9492 12862
rect 9436 12798 9438 12850
rect 9490 12798 9492 12850
rect 9436 12180 9492 12798
rect 9548 12180 9604 12190
rect 9492 12178 9604 12180
rect 9492 12126 9550 12178
rect 9602 12126 9604 12178
rect 9492 12124 9604 12126
rect 9436 12086 9492 12124
rect 9548 12114 9604 12124
rect 9660 12178 9716 13356
rect 9884 12740 9940 13804
rect 10074 13784 10130 13804
rect 10074 13732 10076 13784
rect 10128 13732 10130 13784
rect 10074 13720 10130 13732
rect 10220 13748 10276 13758
rect 10220 13654 10276 13692
rect 10332 13746 10388 14476
rect 10614 14530 10670 14812
rect 11340 14756 11396 14766
rect 10614 14478 10616 14530
rect 10668 14478 10670 14530
rect 10614 14466 10670 14478
rect 10780 14754 11396 14756
rect 10780 14702 11342 14754
rect 11394 14702 11396 14754
rect 10780 14700 11396 14702
rect 10780 14530 10836 14700
rect 11340 14690 11396 14700
rect 11564 14542 11620 16604
rect 11788 15538 11844 16828
rect 12012 16660 12068 18172
rect 12124 18162 12180 18172
rect 12236 17892 12292 18620
rect 12684 18228 12740 19740
rect 12852 19730 12908 19740
rect 13020 19796 13076 19964
rect 13020 19730 13076 19740
rect 12796 19460 12852 19470
rect 13244 19460 13300 20748
rect 13356 20738 13412 20748
rect 13692 20580 13748 21308
rect 14252 20804 14308 21310
rect 14364 20916 14420 20926
rect 14364 20822 14420 20860
rect 14252 20738 14308 20748
rect 13580 20578 13748 20580
rect 13580 20526 13694 20578
rect 13746 20526 13748 20578
rect 13580 20524 13748 20526
rect 13412 20132 13468 20142
rect 13412 20038 13468 20076
rect 12796 19458 13300 19460
rect 12796 19406 12798 19458
rect 12850 19406 13300 19458
rect 12796 19404 13300 19406
rect 12796 19394 12852 19404
rect 12236 17826 12292 17836
rect 12348 18172 12740 18228
rect 13132 18477 13188 18490
rect 13132 18452 13134 18477
rect 13186 18452 13188 18477
rect 12124 16996 12180 17006
rect 12124 16902 12180 16940
rect 11788 15486 11790 15538
rect 11842 15486 11844 15538
rect 11788 15474 11844 15486
rect 11900 16604 12068 16660
rect 11900 15148 11956 16604
rect 12012 15988 12068 15998
rect 12012 15894 12068 15932
rect 11788 15092 11956 15148
rect 10780 14478 10782 14530
rect 10834 14478 10836 14530
rect 10780 14466 10836 14478
rect 10892 14530 10948 14542
rect 10892 14478 10894 14530
rect 10946 14478 10948 14530
rect 10332 13694 10334 13746
rect 10386 13694 10388 13746
rect 10332 13682 10388 13694
rect 10444 14420 10500 14430
rect 10444 13412 10500 14364
rect 10892 14420 10948 14478
rect 11564 14530 11639 14542
rect 11564 14478 11585 14530
rect 11637 14478 11639 14530
rect 11564 14476 11639 14478
rect 11583 14466 11639 14476
rect 10892 14354 10948 14364
rect 9660 12126 9662 12178
rect 9714 12126 9716 12178
rect 9846 12684 9940 12740
rect 10108 13356 10500 13412
rect 10556 13746 10612 13758
rect 10556 13694 10558 13746
rect 10610 13694 10612 13746
rect 9846 12216 9902 12684
rect 9846 12164 9848 12216
rect 9900 12164 9902 12216
rect 9846 12152 9902 12164
rect 9660 12114 9716 12126
rect 10108 12068 10164 13356
rect 10556 13300 10612 13694
rect 11564 13748 11620 13758
rect 11788 13748 11844 15092
rect 12348 14980 12404 18172
rect 12460 18004 12516 18014
rect 12460 16210 12516 17948
rect 12796 17668 12852 17678
rect 12796 17574 12852 17612
rect 13020 17668 13076 17678
rect 12908 16884 12964 16894
rect 12796 16882 12964 16884
rect 12796 16830 12910 16882
rect 12962 16830 12964 16882
rect 12796 16828 12964 16830
rect 12628 16660 12684 16670
rect 12628 16566 12684 16604
rect 12460 16158 12462 16210
rect 12514 16158 12516 16210
rect 12460 16146 12516 16158
rect 12572 16054 12628 16066
rect 12572 16002 12574 16054
rect 12626 16002 12628 16054
rect 12572 15316 12628 16002
rect 12572 15250 12628 15260
rect 12796 15988 12852 16828
rect 12908 16818 12964 16828
rect 13020 16882 13076 17612
rect 13020 16830 13022 16882
rect 13074 16830 13076 16882
rect 13020 16818 13076 16830
rect 12908 16100 12964 16110
rect 12908 16006 12964 16044
rect 12796 15148 12852 15932
rect 13132 15341 13188 18396
rect 13356 17108 13412 17118
rect 13356 16882 13412 17052
rect 13356 16830 13358 16882
rect 13410 16830 13412 16882
rect 13356 16818 13412 16830
rect 13580 16660 13636 20524
rect 13692 20514 13748 20524
rect 13972 20580 14028 20590
rect 14588 20580 14644 21420
rect 14812 21410 14868 21422
rect 14924 21420 15428 21476
rect 15484 21586 15540 21598
rect 15484 21534 15486 21586
rect 15538 21534 15540 21586
rect 14756 20804 14812 20814
rect 14756 20710 14812 20748
rect 14924 20802 14980 21420
rect 15484 21364 15540 21534
rect 15484 21298 15540 21308
rect 15148 21028 15204 21038
rect 14924 20750 14926 20802
rect 14978 20750 14980 20802
rect 14924 20692 14980 20750
rect 14924 20626 14980 20636
rect 15036 20802 15092 20814
rect 15036 20750 15038 20802
rect 15090 20750 15092 20802
rect 15036 20580 15092 20750
rect 14588 20524 14756 20580
rect 13692 20132 13748 20142
rect 13692 20018 13748 20076
rect 13972 20074 14028 20524
rect 13692 19966 13694 20018
rect 13746 19966 13748 20018
rect 13692 19954 13748 19966
rect 13804 20020 13860 20030
rect 13972 20022 13974 20074
rect 14026 20022 14028 20074
rect 14364 20132 14420 20142
rect 13972 20010 14028 20022
rect 14140 20018 14196 20030
rect 13692 19460 13748 19470
rect 13804 19460 13860 19964
rect 13692 19458 13860 19460
rect 13692 19406 13694 19458
rect 13746 19406 13860 19458
rect 13692 19404 13860 19406
rect 14140 19966 14142 20018
rect 14194 19966 14196 20018
rect 13692 19394 13748 19404
rect 14140 19348 14196 19966
rect 14364 19572 14420 20076
rect 14532 19908 14588 19918
rect 14532 19814 14588 19852
rect 14700 19796 14756 20524
rect 15036 20244 15092 20524
rect 15036 20178 15092 20188
rect 14812 20132 14868 20142
rect 14812 20018 14868 20076
rect 15148 20030 15204 20972
rect 15540 21028 15596 21038
rect 15540 20914 15596 20972
rect 15540 20862 15542 20914
rect 15594 20862 15596 20914
rect 15540 20850 15596 20862
rect 15708 20132 15764 20142
rect 14812 19966 14814 20018
rect 14866 19966 14868 20018
rect 14812 19954 14868 19966
rect 14924 20020 14980 20030
rect 14924 19908 14980 19964
rect 15092 20018 15204 20030
rect 15092 19966 15094 20018
rect 15146 19966 15204 20018
rect 15092 19964 15204 19966
rect 15260 20018 15316 20030
rect 15260 19966 15262 20018
rect 15314 19966 15316 20018
rect 15092 19944 15148 19964
rect 14924 19852 15036 19908
rect 14980 19796 15036 19852
rect 14700 19740 14924 19796
rect 14980 19740 15092 19796
rect 14700 19572 14756 19582
rect 14364 19516 14644 19572
rect 14140 19282 14196 19292
rect 14028 19236 14084 19246
rect 14028 19142 14084 19180
rect 14588 19234 14644 19516
rect 14588 19182 14590 19234
rect 14642 19182 14644 19234
rect 14308 19124 14364 19134
rect 14308 19030 14364 19068
rect 14588 19012 14644 19182
rect 14700 19234 14756 19516
rect 14700 19182 14702 19234
rect 14754 19182 14756 19234
rect 14868 19290 14924 19740
rect 15036 19572 15092 19740
rect 15036 19506 15092 19516
rect 15260 19460 15316 19966
rect 15708 20018 15764 20076
rect 15708 19966 15710 20018
rect 15762 19966 15764 20018
rect 15708 19954 15764 19966
rect 15596 19850 15652 19862
rect 15596 19798 15598 19850
rect 15650 19798 15652 19850
rect 14868 19238 14870 19290
rect 14922 19238 14924 19290
rect 14868 19226 14924 19238
rect 15036 19348 15092 19358
rect 15036 19234 15092 19292
rect 14700 19170 14756 19182
rect 15036 19182 15038 19234
rect 15090 19182 15092 19234
rect 15036 19170 15092 19182
rect 15148 19124 15204 19134
rect 14588 18956 14868 19012
rect 14812 18674 14868 18956
rect 14812 18622 14814 18674
rect 14866 18622 14868 18674
rect 14812 18610 14868 18622
rect 14308 18508 14532 18564
rect 14308 18479 14364 18508
rect 13916 18450 13972 18462
rect 13916 18398 13918 18450
rect 13970 18398 13972 18450
rect 14308 18427 14310 18479
rect 14362 18427 14364 18479
rect 14308 18415 14364 18427
rect 13916 18340 13972 18398
rect 14364 18340 14420 18350
rect 13916 18274 13972 18284
rect 14028 18338 14420 18340
rect 14028 18286 14366 18338
rect 14418 18286 14420 18338
rect 14028 18284 14420 18286
rect 13804 17780 13860 17790
rect 13804 17778 13972 17780
rect 13804 17726 13806 17778
rect 13858 17726 13972 17778
rect 13804 17724 13972 17726
rect 13804 17714 13860 17724
rect 13412 16604 13636 16660
rect 13412 16042 13468 16604
rect 13412 15990 13414 16042
rect 13466 15990 13468 16042
rect 13580 16100 13636 16110
rect 13580 16006 13636 16044
rect 13804 16098 13860 16110
rect 13804 16046 13806 16098
rect 13858 16046 13860 16098
rect 13412 15876 13468 15990
rect 13412 15810 13468 15820
rect 13580 15540 13636 15550
rect 13580 15446 13636 15484
rect 13132 15289 13134 15341
rect 13186 15289 13188 15341
rect 13132 15148 13188 15289
rect 12348 14914 12404 14924
rect 12684 15092 12852 15148
rect 13020 15092 13188 15148
rect 13468 15204 13524 15214
rect 13804 15148 13860 16046
rect 13916 15314 13972 17724
rect 14028 16772 14084 18284
rect 14364 18274 14420 18284
rect 14476 18116 14532 18508
rect 15148 18450 15204 19068
rect 15260 18676 15316 19404
rect 15428 19684 15484 19694
rect 15428 19458 15484 19628
rect 15428 19406 15430 19458
rect 15482 19406 15484 19458
rect 15428 19394 15484 19406
rect 15596 19012 15652 19798
rect 15820 19796 15876 21644
rect 15988 21474 16044 21486
rect 15988 21422 15990 21474
rect 16042 21422 16044 21474
rect 15988 21364 16044 21422
rect 15988 21298 16044 21308
rect 16156 21028 16212 21756
rect 15988 20972 16212 21028
rect 15988 20914 16044 20972
rect 15988 20862 15990 20914
rect 16042 20862 16044 20914
rect 15988 20850 16044 20862
rect 16156 20802 16212 20814
rect 16156 20750 16158 20802
rect 16210 20750 16212 20802
rect 16044 20468 16100 20478
rect 15932 20020 15988 20030
rect 15932 19926 15988 19964
rect 15820 19730 15876 19740
rect 16044 19302 16100 20412
rect 16156 20020 16212 20750
rect 16268 20356 16324 22540
rect 16380 22594 16492 22606
rect 16380 22542 16382 22594
rect 16434 22542 16492 22594
rect 16380 22540 16492 22542
rect 16380 22530 16436 22540
rect 16436 21476 16492 21486
rect 16436 20916 16492 21420
rect 16268 20290 16324 20300
rect 16380 20860 16492 20916
rect 16380 20244 16436 20860
rect 16604 20804 16660 23102
rect 16604 20738 16660 20748
rect 16716 23154 16772 23166
rect 16716 23102 16718 23154
rect 16770 23102 16772 23154
rect 16716 21140 16772 23102
rect 17388 23044 17444 25116
rect 17500 24948 17556 24958
rect 17500 24854 17556 24892
rect 17836 24722 17892 24734
rect 17836 24670 17838 24722
rect 17890 24670 17892 24722
rect 17836 24612 17892 24670
rect 18172 24612 18228 24622
rect 17836 24610 18228 24612
rect 17836 24558 18174 24610
rect 18226 24558 18228 24610
rect 17836 24556 18228 24558
rect 18172 24546 18228 24556
rect 17836 23940 17892 23950
rect 17948 23940 18004 23950
rect 17556 23938 18228 23940
rect 17556 23886 17838 23938
rect 17890 23886 17950 23938
rect 18002 23886 18228 23938
rect 17556 23884 18228 23886
rect 17556 23378 17612 23884
rect 17836 23874 17892 23884
rect 17948 23874 18004 23884
rect 17556 23326 17558 23378
rect 17610 23326 17612 23378
rect 17556 23314 17612 23326
rect 17948 23604 18004 23614
rect 17948 23378 18004 23548
rect 17948 23326 17950 23378
rect 18002 23326 18004 23378
rect 17948 23314 18004 23326
rect 17500 23044 17556 23054
rect 17388 22988 17500 23044
rect 16996 22596 17052 22606
rect 16996 22372 17052 22540
rect 16996 22278 17052 22316
rect 17388 22148 17444 22158
rect 17276 21812 17332 21822
rect 16884 21588 16940 21598
rect 17164 21588 17220 21598
rect 16940 21532 16996 21588
rect 16884 21494 16996 21532
rect 16492 20580 16548 20590
rect 16716 20580 16772 21084
rect 16492 20486 16548 20524
rect 16604 20524 16772 20580
rect 16828 20802 16884 20814
rect 16828 20750 16830 20802
rect 16882 20750 16884 20802
rect 16604 20468 16660 20524
rect 16604 20402 16660 20412
rect 16716 20356 16772 20366
rect 16380 20188 16548 20244
rect 16380 20020 16436 20030
rect 16156 19964 16380 20020
rect 16268 19796 16324 19806
rect 15988 19290 16100 19302
rect 15708 19234 15764 19246
rect 15708 19182 15710 19234
rect 15762 19182 15764 19234
rect 15708 19124 15764 19182
rect 15708 19058 15764 19068
rect 15820 19236 15876 19246
rect 15988 19238 15990 19290
rect 16042 19238 16100 19290
rect 15988 19236 16100 19238
rect 16156 19460 16212 19470
rect 15988 19226 16044 19236
rect 16156 19234 16212 19404
rect 15820 19124 15876 19180
rect 16156 19182 16158 19234
rect 16210 19182 16212 19234
rect 16156 19170 16212 19182
rect 15820 19122 15988 19124
rect 15820 19070 15822 19122
rect 15874 19070 15988 19122
rect 15820 19068 15988 19070
rect 15820 19058 15876 19068
rect 15596 18946 15652 18956
rect 15932 19012 15988 19068
rect 15932 18946 15988 18956
rect 15820 18900 15876 18910
rect 15484 18676 15540 18686
rect 15260 18674 15540 18676
rect 15260 18622 15486 18674
rect 15538 18622 15540 18674
rect 15260 18620 15540 18622
rect 15484 18610 15540 18620
rect 15148 18398 15150 18450
rect 15202 18398 15204 18450
rect 15148 18386 15204 18398
rect 15260 18452 15316 18462
rect 14364 18060 14532 18116
rect 14198 17892 14254 17902
rect 14198 17666 14254 17836
rect 14198 17614 14200 17666
rect 14252 17614 14254 17666
rect 14198 17602 14254 17614
rect 14364 17666 14420 18060
rect 15260 17780 15316 18396
rect 15820 18450 15876 18844
rect 15820 18398 15822 18450
rect 15874 18398 15876 18450
rect 15820 18386 15876 18398
rect 15932 18452 15988 18462
rect 15932 18358 15988 18396
rect 15092 17724 15316 17780
rect 14364 17614 14366 17666
rect 14418 17614 14420 17666
rect 14140 16772 14196 16782
rect 14028 16770 14196 16772
rect 14028 16718 14142 16770
rect 14194 16718 14196 16770
rect 14028 16716 14196 16718
rect 14140 16706 14196 16716
rect 14364 16436 14420 17614
rect 14476 17668 14532 17678
rect 14476 17574 14532 17612
rect 15092 17442 15148 17724
rect 15260 17666 15316 17724
rect 16044 18228 16100 18238
rect 16044 17778 16100 18172
rect 16044 17726 16046 17778
rect 16098 17726 16100 17778
rect 16044 17714 16100 17726
rect 15260 17614 15262 17666
rect 15314 17614 15316 17666
rect 15260 17602 15316 17614
rect 15092 17390 15094 17442
rect 15146 17390 15148 17442
rect 15092 17108 15148 17390
rect 15148 17052 15316 17108
rect 15092 17042 15148 17052
rect 15260 16548 15316 17052
rect 16268 16996 16324 19740
rect 16380 18900 16436 19964
rect 16380 18834 16436 18844
rect 16492 18116 16548 20188
rect 16716 20132 16772 20300
rect 16604 20130 16772 20132
rect 16604 20078 16718 20130
rect 16770 20078 16772 20130
rect 16604 20076 16772 20078
rect 16604 18900 16660 20076
rect 16716 20066 16772 20076
rect 16828 20020 16884 20750
rect 16828 19954 16884 19964
rect 16940 19908 16996 21494
rect 17164 20804 17220 21532
rect 17164 20710 17220 20748
rect 16772 19460 16828 19470
rect 16772 19346 16828 19404
rect 16772 19294 16774 19346
rect 16826 19294 16828 19346
rect 16772 19282 16828 19294
rect 16604 18834 16660 18844
rect 16940 18564 16996 19852
rect 17164 19348 17220 19358
rect 17164 19254 17220 19292
rect 16940 18498 16996 18508
rect 17052 19236 17108 19246
rect 16492 18050 16548 18060
rect 17052 18004 17108 19180
rect 17276 18452 17332 21756
rect 17388 19796 17444 22092
rect 17500 20580 17556 22988
rect 17780 22484 17836 22494
rect 17780 22426 17836 22428
rect 17612 22370 17668 22382
rect 17612 22318 17614 22370
rect 17666 22318 17668 22370
rect 17780 22374 17782 22426
rect 17834 22374 17836 22426
rect 17780 22362 17836 22374
rect 18060 22372 18116 22382
rect 17612 21700 17668 22318
rect 18060 22278 18116 22316
rect 17948 22258 18004 22270
rect 17948 22206 17950 22258
rect 18002 22206 18004 22258
rect 17612 21634 17668 21644
rect 17836 21924 17892 21934
rect 17948 21924 18004 22206
rect 17892 21868 18004 21924
rect 17668 21474 17724 21486
rect 17668 21422 17670 21474
rect 17722 21422 17724 21474
rect 17668 21028 17724 21422
rect 17836 21364 17892 21868
rect 18172 21812 18228 23884
rect 18284 23380 18340 25788
rect 18396 25620 18452 25630
rect 18396 25526 18452 25564
rect 18508 25508 18564 26238
rect 18620 26290 18676 26852
rect 18620 26238 18622 26290
rect 18674 26238 18676 26290
rect 18620 26226 18676 26238
rect 18732 26852 18788 27356
rect 18956 27188 19012 27198
rect 19012 27132 19124 27188
rect 18956 27094 19012 27132
rect 18732 26068 18788 26796
rect 18620 26012 18788 26068
rect 18844 26964 18900 26974
rect 18620 25732 18676 26012
rect 18620 25666 18676 25676
rect 18732 25844 18788 25854
rect 18564 25452 18676 25508
rect 18508 25442 18564 25452
rect 18620 24948 18676 25452
rect 18732 25284 18788 25788
rect 18844 25506 18900 26908
rect 18956 26628 19012 26638
rect 18956 26290 19012 26572
rect 18956 26238 18958 26290
rect 19010 26238 19012 26290
rect 18956 26226 19012 26238
rect 19068 25844 19124 27132
rect 19292 26908 19348 28700
rect 19404 28642 19460 29148
rect 19516 28868 19572 28878
rect 19516 28810 19572 28812
rect 19516 28758 19518 28810
rect 19570 28758 19572 28810
rect 19516 28746 19572 28758
rect 19404 28590 19406 28642
rect 19458 28590 19460 28642
rect 19404 27076 19460 28590
rect 19628 28644 19684 29708
rect 19740 29652 19796 29662
rect 20188 29652 20244 29932
rect 19740 29426 19796 29596
rect 19740 29374 19742 29426
rect 19794 29374 19796 29426
rect 19740 29362 19796 29374
rect 19852 29596 20244 29652
rect 19852 29426 19908 29596
rect 19852 29374 19854 29426
rect 19906 29374 19908 29426
rect 19852 28868 19908 29374
rect 20020 29428 20076 29438
rect 20020 29334 20076 29372
rect 20300 28868 20356 30044
rect 20412 30034 20468 30044
rect 20524 29428 20580 29438
rect 20412 29316 20468 29326
rect 20412 29222 20468 29260
rect 19852 28802 19908 28812
rect 20188 28812 20356 28868
rect 19740 28644 19796 28654
rect 19628 28588 19740 28644
rect 19740 28550 19796 28588
rect 19516 28532 19572 28542
rect 19516 28082 19572 28476
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19516 28030 19518 28082
rect 19570 28030 19572 28082
rect 19516 28018 19572 28030
rect 19740 28084 19796 28094
rect 20188 28084 20244 28812
rect 20412 28810 20468 28822
rect 20412 28758 20414 28810
rect 20466 28758 20468 28810
rect 20412 28756 20468 28758
rect 20412 28690 20468 28700
rect 20300 28644 20356 28654
rect 20300 28550 20356 28588
rect 20524 28642 20580 29372
rect 20524 28590 20526 28642
rect 20578 28590 20580 28642
rect 20524 28532 20580 28590
rect 20524 28466 20580 28476
rect 20188 28028 20580 28084
rect 19740 27188 19796 28028
rect 20244 27914 20300 27926
rect 20244 27862 20246 27914
rect 20298 27862 20300 27914
rect 20244 27860 20300 27862
rect 19404 27010 19460 27020
rect 19516 27036 19616 27076
rect 19516 26984 19562 27036
rect 19614 26984 19616 27036
rect 19516 26972 19616 26984
rect 19516 26908 19572 26972
rect 19740 26908 19796 27132
rect 19292 26852 19572 26908
rect 19628 26852 19796 26908
rect 19964 27802 20020 27814
rect 20244 27804 20356 27860
rect 19964 27750 19966 27802
rect 20018 27750 20020 27802
rect 19964 26852 20020 27750
rect 20300 27524 20356 27804
rect 20524 27748 20580 28028
rect 20636 27970 20692 30044
rect 20748 30098 20804 30110
rect 20748 30046 20750 30098
rect 20802 30046 20804 30098
rect 20748 29988 20804 30046
rect 20748 29922 20804 29932
rect 20860 29428 20916 30268
rect 21084 29988 21140 30828
rect 21644 30772 21700 30782
rect 21420 30660 21476 30670
rect 21420 30212 21476 30604
rect 21420 30210 21588 30212
rect 21084 29922 21140 29932
rect 21252 30154 21308 30166
rect 21252 30102 21254 30154
rect 21306 30102 21308 30154
rect 21420 30158 21422 30210
rect 21474 30158 21588 30210
rect 21420 30156 21588 30158
rect 21420 30146 21476 30156
rect 21252 29550 21308 30102
rect 21196 29540 21308 29550
rect 21252 29484 21308 29540
rect 20860 29362 20916 29372
rect 21084 29426 21140 29438
rect 21084 29374 21086 29426
rect 21138 29374 21140 29426
rect 20916 29202 20972 29214
rect 20916 29150 20918 29202
rect 20970 29150 20972 29202
rect 20916 28644 20972 29150
rect 21084 29204 21140 29374
rect 21084 29138 21140 29148
rect 21196 28644 21252 29484
rect 20916 28578 20972 28588
rect 21084 28642 21252 28644
rect 21084 28590 21198 28642
rect 21250 28590 21252 28642
rect 21084 28588 21252 28590
rect 20636 27918 20638 27970
rect 20690 27918 20692 27970
rect 20636 27906 20692 27918
rect 20804 27802 20860 27814
rect 20636 27748 20692 27758
rect 20524 27692 20636 27748
rect 20804 27750 20806 27802
rect 20858 27750 20860 27802
rect 20804 27748 20860 27750
rect 20804 27692 21028 27748
rect 20524 27524 20580 27534
rect 20300 27468 20468 27524
rect 20300 27300 20356 27310
rect 20300 27242 20356 27244
rect 20300 27190 20302 27242
rect 20354 27190 20356 27242
rect 20300 27178 20356 27190
rect 20300 27076 20356 27086
rect 20300 26982 20356 27020
rect 19068 25778 19124 25788
rect 18844 25454 18846 25506
rect 18898 25454 18900 25506
rect 18844 25442 18900 25454
rect 18956 25508 19012 25518
rect 18956 25414 19012 25452
rect 19122 25450 19178 25462
rect 19122 25398 19124 25450
rect 19176 25398 19178 25450
rect 18732 25228 18900 25284
rect 18620 24892 18788 24948
rect 18546 24759 18602 24771
rect 18546 24707 18548 24759
rect 18600 24707 18602 24759
rect 18546 24276 18602 24707
rect 18284 23314 18340 23324
rect 18396 24220 18602 24276
rect 18732 24722 18788 24892
rect 18732 24670 18734 24722
rect 18786 24670 18788 24722
rect 18284 23156 18340 23166
rect 18284 23062 18340 23100
rect 18396 22606 18452 24220
rect 18732 24164 18788 24670
rect 18844 24722 18900 25228
rect 19122 24836 19178 25398
rect 18844 24670 18846 24722
rect 18898 24670 18900 24722
rect 18844 24658 18900 24670
rect 18956 24780 19178 24836
rect 19292 25396 19348 25406
rect 18732 24108 18900 24164
rect 18732 23938 18788 23950
rect 18732 23886 18734 23938
rect 18786 23886 18788 23938
rect 18732 23604 18788 23886
rect 18844 23716 18900 24108
rect 18844 23650 18900 23660
rect 18732 23538 18788 23548
rect 18956 23380 19012 24780
rect 19292 24722 19348 25340
rect 19292 24670 19294 24722
rect 19346 24670 19348 24722
rect 19292 24658 19348 24670
rect 19404 24276 19460 26852
rect 19628 26290 19684 26852
rect 19964 26786 20020 26796
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19740 26458 19796 26470
rect 19740 26406 19742 26458
rect 19794 26406 19796 26458
rect 19740 26404 19796 26406
rect 19740 26338 19796 26348
rect 20412 26404 20468 27468
rect 19628 26238 19630 26290
rect 19682 26238 19684 26290
rect 19628 26226 19684 26238
rect 20300 26292 20356 26302
rect 20412 26292 20468 26348
rect 20300 26290 20468 26292
rect 20300 26238 20302 26290
rect 20354 26238 20468 26290
rect 20300 26236 20468 26238
rect 20300 26226 20356 26236
rect 19516 25620 19572 25630
rect 19516 25618 19908 25620
rect 19516 25566 19518 25618
rect 19570 25566 19908 25618
rect 19516 25564 19908 25566
rect 19516 25554 19572 25564
rect 19852 25506 19908 25564
rect 19852 25454 19854 25506
rect 19906 25454 19908 25506
rect 19852 25442 19908 25454
rect 20188 25282 20244 25294
rect 20188 25230 20190 25282
rect 20242 25230 20244 25282
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20188 24948 20244 25230
rect 20524 24948 20580 27468
rect 20636 26514 20692 27692
rect 20636 26462 20638 26514
rect 20690 26462 20692 26514
rect 20636 26450 20692 26462
rect 20972 27300 21028 27692
rect 20972 26292 21028 27244
rect 21084 26516 21140 28588
rect 21196 28578 21252 28588
rect 21420 29426 21476 29438
rect 21420 29374 21422 29426
rect 21474 29374 21476 29426
rect 21420 28980 21476 29374
rect 21532 29426 21588 30156
rect 21532 29374 21534 29426
rect 21586 29374 21588 29426
rect 21532 29362 21588 29374
rect 21644 30210 21700 30716
rect 21644 30158 21646 30210
rect 21698 30158 21700 30210
rect 21420 28756 21476 28924
rect 21420 28642 21476 28700
rect 21420 28590 21422 28642
rect 21474 28590 21476 28642
rect 21420 28578 21476 28590
rect 21532 29204 21588 29214
rect 21644 29204 21700 30158
rect 21756 29876 21812 30942
rect 21980 30994 22036 31006
rect 21980 30942 21982 30994
rect 22034 30942 22036 30994
rect 21980 30548 22036 30942
rect 22092 30826 22148 31612
rect 22204 31602 22260 31612
rect 22428 31780 22484 32386
rect 22540 32116 22596 32126
rect 22540 32002 22596 32060
rect 22540 31950 22542 32002
rect 22594 31950 22596 32002
rect 22540 31938 22596 31950
rect 22988 32004 23044 32510
rect 22988 31938 23044 31948
rect 22092 30774 22094 30826
rect 22146 30774 22148 30826
rect 22092 30762 22148 30774
rect 22316 30994 22372 31006
rect 22316 30942 22318 30994
rect 22370 30942 22372 30994
rect 21980 30482 22036 30492
rect 21868 30154 21924 30166
rect 21868 30102 21870 30154
rect 21922 30102 21924 30154
rect 21868 30100 21924 30102
rect 21868 30034 21924 30044
rect 21756 29810 21812 29820
rect 22316 29540 22372 30942
rect 22428 30548 22484 31724
rect 22876 31778 22932 31790
rect 22876 31726 22878 31778
rect 22930 31726 22932 31778
rect 22540 30996 22596 31006
rect 22876 30996 22932 31726
rect 23100 31444 23156 32956
rect 23212 32676 23268 32686
rect 23212 32562 23268 32620
rect 23548 32676 23604 32686
rect 23548 32582 23604 32620
rect 23212 32510 23214 32562
rect 23266 32510 23268 32562
rect 23212 32498 23268 32510
rect 23660 31780 23716 33740
rect 23772 33684 23828 33694
rect 23772 33460 23828 33628
rect 23772 33012 23828 33404
rect 23772 32946 23828 32956
rect 23791 32593 23847 32605
rect 23791 32541 23793 32593
rect 23845 32564 23847 32593
rect 23845 32541 23940 32564
rect 23791 32508 23940 32541
rect 23100 31378 23156 31388
rect 23436 31724 23716 31780
rect 23772 32004 23828 32014
rect 22540 30994 22932 30996
rect 22540 30942 22542 30994
rect 22594 30942 22932 30994
rect 22540 30940 22932 30942
rect 23212 30996 23268 31006
rect 22540 30930 22596 30940
rect 23212 30902 23268 30940
rect 22876 30772 22932 30782
rect 23436 30772 23492 31724
rect 23604 31554 23660 31566
rect 23604 31502 23606 31554
rect 23658 31502 23660 31554
rect 23604 31444 23660 31502
rect 23660 31388 23716 31444
rect 23604 31378 23716 31388
rect 23548 31108 23604 31118
rect 23548 30994 23604 31052
rect 23548 30942 23550 30994
rect 23602 30942 23604 30994
rect 23548 30930 23604 30942
rect 22876 30770 23156 30772
rect 22876 30718 22878 30770
rect 22930 30718 23156 30770
rect 22876 30716 23156 30718
rect 23436 30716 23604 30772
rect 22876 30706 22932 30716
rect 22428 30492 22932 30548
rect 22540 30212 22596 30222
rect 22540 29652 22596 30156
rect 22540 29586 22596 29596
rect 22764 29652 22820 29662
rect 22316 29474 22372 29484
rect 21812 29428 21868 29438
rect 21812 29334 21868 29372
rect 22204 29428 22260 29438
rect 22540 29426 22596 29438
rect 22204 29334 22260 29372
rect 22372 29370 22428 29382
rect 21588 29148 21700 29204
rect 22372 29318 22374 29370
rect 22426 29318 22428 29370
rect 21308 27858 21364 27870
rect 21308 27806 21310 27858
rect 21362 27806 21364 27858
rect 21196 27074 21252 27086
rect 21196 27022 21198 27074
rect 21250 27022 21252 27074
rect 21196 26852 21252 27022
rect 21308 26964 21364 27806
rect 21308 26898 21364 26908
rect 21420 27074 21476 27086
rect 21420 27022 21422 27074
rect 21474 27022 21476 27074
rect 21196 26786 21252 26796
rect 21308 26516 21364 26526
rect 21084 26514 21364 26516
rect 21084 26462 21310 26514
rect 21362 26462 21364 26514
rect 21084 26460 21364 26462
rect 21308 26450 21364 26460
rect 21420 26292 21476 27022
rect 21532 26908 21588 29148
rect 22372 29092 22428 29318
rect 22316 29036 22428 29092
rect 22540 29374 22542 29426
rect 22594 29374 22596 29426
rect 21700 28868 21756 28878
rect 21700 28774 21756 28812
rect 22316 28654 22372 29036
rect 22260 28644 22372 28654
rect 22092 28588 22148 28598
rect 21868 28586 22148 28588
rect 21868 28534 22094 28586
rect 22146 28534 22148 28586
rect 22316 28588 22372 28644
rect 22428 28868 22484 28878
rect 22540 28868 22596 29374
rect 22484 28812 22596 28868
rect 22652 29426 22708 29438
rect 22652 29374 22654 29426
rect 22706 29374 22708 29426
rect 22652 29316 22708 29374
rect 22428 28642 22484 28812
rect 22428 28590 22430 28642
rect 22482 28590 22484 28642
rect 22260 28550 22316 28588
rect 22428 28578 22484 28590
rect 22540 28644 22596 28654
rect 22652 28644 22708 29260
rect 22540 28642 22708 28644
rect 22540 28590 22542 28642
rect 22594 28590 22708 28642
rect 22540 28588 22708 28590
rect 22540 28578 22596 28588
rect 21868 28532 22148 28534
rect 21644 27887 21756 27972
rect 21644 27835 21702 27887
rect 21754 27835 21756 27887
rect 21644 27823 21756 27835
rect 21644 27198 21700 27823
rect 21756 27748 21812 27758
rect 21868 27748 21924 28532
rect 22092 28522 22148 28532
rect 22764 28420 22820 29596
rect 21756 27746 21924 27748
rect 21756 27694 21758 27746
rect 21810 27694 21924 27746
rect 21756 27692 21924 27694
rect 22428 28364 22820 28420
rect 21756 27682 21812 27692
rect 21644 27188 21756 27198
rect 21644 27132 21700 27188
rect 21700 27094 21756 27132
rect 22260 27076 22316 27114
rect 22260 27010 22316 27020
rect 21980 26964 22036 26974
rect 21532 26852 21700 26908
rect 20972 26290 21476 26292
rect 20972 26238 20974 26290
rect 21026 26238 21476 26290
rect 20972 26236 21476 26238
rect 21644 26292 21700 26852
rect 21980 26514 22036 26908
rect 21980 26462 21982 26514
rect 22034 26462 22036 26514
rect 21980 26450 22036 26462
rect 21644 26290 21924 26292
rect 21644 26238 21646 26290
rect 21698 26238 21924 26290
rect 21644 26236 21924 26238
rect 20972 26226 21028 26236
rect 21644 26226 21700 26236
rect 21196 25508 21252 25518
rect 20804 25396 20860 25406
rect 20804 25302 20860 25340
rect 20076 24892 20244 24948
rect 20300 24892 20580 24948
rect 20076 24722 20132 24892
rect 20076 24670 20078 24722
rect 20130 24670 20132 24722
rect 20076 24658 20132 24670
rect 19404 24210 19460 24220
rect 20188 24388 20244 24398
rect 20188 23940 20244 24332
rect 18844 23324 19012 23380
rect 19180 23716 19236 23726
rect 18620 23156 18676 23166
rect 18620 23042 18676 23100
rect 18620 22990 18622 23042
rect 18674 22990 18676 23042
rect 18620 22978 18676 22990
rect 18844 22708 18900 23324
rect 19034 23191 19090 23203
rect 19034 23139 19036 23191
rect 19088 23139 19090 23191
rect 19034 22820 19090 23139
rect 18340 22594 18452 22606
rect 18340 22542 18342 22594
rect 18394 22542 18452 22594
rect 18340 22540 18452 22542
rect 18620 22652 18900 22708
rect 18956 22764 19090 22820
rect 19180 23154 19236 23660
rect 19180 23102 19182 23154
rect 19234 23102 19236 23154
rect 18340 22530 18396 22540
rect 18396 22372 18452 22382
rect 18172 21746 18228 21756
rect 18284 21924 18340 21934
rect 18284 21698 18340 21868
rect 18284 21646 18286 21698
rect 18338 21646 18340 21698
rect 18284 21634 18340 21646
rect 17948 21588 18004 21598
rect 18396 21588 18452 22316
rect 18620 21710 18676 22652
rect 18844 22372 18900 22382
rect 18844 22278 18900 22316
rect 18620 21698 18732 21710
rect 18620 21646 18678 21698
rect 18730 21646 18732 21698
rect 18620 21644 18732 21646
rect 18676 21634 18732 21644
rect 18396 21586 18564 21588
rect 17948 21494 18004 21532
rect 18116 21530 18172 21542
rect 18116 21478 18118 21530
rect 18170 21478 18172 21530
rect 18396 21534 18398 21586
rect 18450 21534 18564 21586
rect 18396 21532 18564 21534
rect 18396 21522 18452 21532
rect 17836 21308 18004 21364
rect 17668 20962 17724 20972
rect 17612 20804 17668 20814
rect 17948 20802 18004 21308
rect 18116 21028 18172 21478
rect 18116 20962 18172 20972
rect 18340 21364 18396 21374
rect 18340 21026 18396 21308
rect 18340 20974 18342 21026
rect 18394 20974 18396 21026
rect 18340 20962 18396 20974
rect 17612 20710 17668 20748
rect 17780 20746 17836 20758
rect 17500 20514 17556 20524
rect 17780 20694 17782 20746
rect 17834 20694 17836 20746
rect 17948 20750 17950 20802
rect 18002 20750 18004 20802
rect 17948 20738 18004 20750
rect 18060 20802 18116 20814
rect 18060 20750 18062 20802
rect 18114 20750 18116 20802
rect 17780 20580 17836 20694
rect 17780 20244 17836 20524
rect 18060 20244 18116 20750
rect 18508 20244 18564 21532
rect 18956 21476 19012 22764
rect 19180 22596 19236 23102
rect 19292 23604 19348 23614
rect 19292 23154 19348 23548
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 20188 23380 20244 23884
rect 19292 23102 19294 23154
rect 19346 23102 19348 23154
rect 19292 23090 19348 23102
rect 19964 23324 20244 23380
rect 19068 22540 19236 22596
rect 19068 22538 19124 22540
rect 19068 22486 19070 22538
rect 19122 22486 19124 22538
rect 19964 22494 20020 23324
rect 20076 22932 20132 22942
rect 20076 22838 20132 22876
rect 19068 22474 19124 22486
rect 19908 22482 20020 22494
rect 19908 22430 19910 22482
rect 19962 22430 20020 22482
rect 19908 22428 20020 22430
rect 19908 22418 19964 22428
rect 19068 22370 19124 22382
rect 19068 22318 19070 22370
rect 19122 22318 19124 22370
rect 19068 21924 19124 22318
rect 20076 22370 20132 22382
rect 20076 22318 20078 22370
rect 20130 22318 20132 22370
rect 19068 21812 19124 21868
rect 19628 22260 19684 22270
rect 19180 21812 19236 21822
rect 19068 21810 19236 21812
rect 19068 21758 19182 21810
rect 19234 21758 19236 21810
rect 19068 21756 19236 21758
rect 19628 21812 19684 22204
rect 20076 22148 20132 22318
rect 20076 22082 20132 22092
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20300 21822 20356 24892
rect 21196 24276 21252 25452
rect 21532 25506 21588 25518
rect 21532 25454 21534 25506
rect 21586 25454 21588 25506
rect 21532 25396 21588 25454
rect 21532 25330 21588 25340
rect 21868 24836 21924 26236
rect 22428 26180 22484 28364
rect 22876 28196 22932 30492
rect 23100 30324 23156 30716
rect 23324 30324 23380 30334
rect 23100 30322 23380 30324
rect 23100 30270 23326 30322
rect 23378 30270 23380 30322
rect 23100 30268 23380 30270
rect 23324 30258 23380 30268
rect 23436 29540 23492 29550
rect 22876 28130 22932 28140
rect 22988 29428 23044 29438
rect 22764 27972 22820 27982
rect 22988 27972 23044 29372
rect 23212 29202 23268 29214
rect 23212 29150 23214 29202
rect 23266 29150 23268 29202
rect 23212 29092 23268 29150
rect 23212 29026 23268 29036
rect 23100 28868 23156 28878
rect 23100 28774 23156 28812
rect 23436 28644 23492 29484
rect 23548 29428 23604 30716
rect 23660 30548 23716 31378
rect 23772 30826 23828 31948
rect 23884 31892 23940 32508
rect 23996 32116 24052 33740
rect 25004 33458 25060 34076
rect 25116 33684 25172 34412
rect 25228 33796 25284 38098
rect 25340 36260 25396 38220
rect 25452 36428 25508 38332
rect 25900 38164 25956 39788
rect 26012 39396 26068 39900
rect 26236 39620 26292 39630
rect 26292 39564 26404 39620
rect 26236 39526 26292 39564
rect 26012 39340 26292 39396
rect 26124 39172 26180 39182
rect 26124 38877 26180 39116
rect 26236 38948 26292 39340
rect 26348 39284 26404 39564
rect 26348 39228 26852 39284
rect 26348 38948 26404 38958
rect 26236 38946 26404 38948
rect 26236 38894 26350 38946
rect 26402 38894 26404 38946
rect 26236 38892 26404 38894
rect 26348 38882 26404 38892
rect 26104 38865 26180 38877
rect 26104 38813 26106 38865
rect 26158 38813 26180 38865
rect 26104 38801 26180 38813
rect 26124 38276 26180 38801
rect 26796 38834 26852 39228
rect 26796 38782 26798 38834
rect 26850 38782 26852 38834
rect 26796 38770 26852 38782
rect 26124 38210 26180 38220
rect 25788 38108 25956 38164
rect 25620 37826 25676 37838
rect 25620 37774 25622 37826
rect 25674 37774 25676 37826
rect 25620 37604 25676 37774
rect 25620 37538 25676 37548
rect 25564 37380 25620 37390
rect 25564 37156 25620 37324
rect 25676 37380 25732 37390
rect 25788 37380 25844 38108
rect 26236 38052 26292 38062
rect 26124 38050 26292 38052
rect 26124 37998 26238 38050
rect 26290 37998 26292 38050
rect 26124 37996 26292 37998
rect 25956 37938 26012 37950
rect 25956 37886 25958 37938
rect 26010 37886 26012 37938
rect 25956 37716 26012 37886
rect 25956 37650 26012 37660
rect 25676 37378 25844 37380
rect 25676 37326 25678 37378
rect 25730 37326 25844 37378
rect 25676 37324 25844 37326
rect 25676 37314 25732 37324
rect 26124 37296 26180 37996
rect 26236 37986 26292 37996
rect 26348 38050 26404 38062
rect 26348 37998 26350 38050
rect 26402 37998 26404 38050
rect 26124 37244 26126 37296
rect 26178 37244 26180 37296
rect 25956 37210 26012 37222
rect 25956 37158 25958 37210
rect 26010 37158 26012 37210
rect 25564 37100 25732 37156
rect 25564 36596 25620 36634
rect 25564 36530 25620 36540
rect 25452 36372 25620 36428
rect 25340 36204 25508 36260
rect 25340 35728 25396 35740
rect 25340 35676 25342 35728
rect 25394 35676 25396 35728
rect 25340 35364 25396 35676
rect 25340 34972 25396 35308
rect 25452 35140 25508 36204
rect 25452 35074 25508 35084
rect 25340 34916 25488 34972
rect 25432 34886 25488 34916
rect 25432 34883 25508 34886
rect 25432 34831 25434 34883
rect 25486 34831 25508 34883
rect 25432 34819 25508 34831
rect 25452 34244 25508 34819
rect 25452 34178 25508 34188
rect 25396 34020 25452 34030
rect 25396 33926 25452 33964
rect 25228 33730 25284 33740
rect 25116 33618 25172 33628
rect 25004 33406 25006 33458
rect 25058 33406 25060 33458
rect 25004 33394 25060 33406
rect 25340 33460 25396 33470
rect 25116 33348 25172 33358
rect 24836 33290 24892 33302
rect 24444 33236 24500 33246
rect 24836 33238 24838 33290
rect 24890 33238 24892 33290
rect 24444 33234 24724 33236
rect 24444 33182 24446 33234
rect 24498 33182 24724 33234
rect 24444 33180 24724 33182
rect 24444 33170 24500 33180
rect 24668 32564 24724 33180
rect 24836 32900 24892 33238
rect 24836 32844 25060 32900
rect 24668 32562 24948 32564
rect 24668 32510 24670 32562
rect 24722 32510 24948 32562
rect 24668 32508 24948 32510
rect 24668 32498 24724 32508
rect 24892 32228 24948 32508
rect 24668 32172 24948 32228
rect 25004 32228 25060 32844
rect 23996 32060 24164 32116
rect 23884 31332 23940 31836
rect 23996 31666 24052 31678
rect 23996 31614 23998 31666
rect 24050 31614 24052 31666
rect 23996 31556 24052 31614
rect 23996 31490 24052 31500
rect 24108 31332 24164 32060
rect 24556 32004 24612 32014
rect 24556 31739 24612 31948
rect 24276 31722 24332 31734
rect 24276 31670 24278 31722
rect 24330 31670 24332 31722
rect 24556 31687 24558 31739
rect 24610 31687 24612 31739
rect 24556 31675 24612 31687
rect 24276 31556 24332 31670
rect 24668 31556 24724 32172
rect 24276 31500 24724 31556
rect 24780 31722 24836 31734
rect 24780 31670 24782 31722
rect 24834 31670 24836 31722
rect 24780 31556 24836 31670
rect 24780 31490 24836 31500
rect 24892 31444 24948 31454
rect 24108 31276 24836 31332
rect 23884 31266 23940 31276
rect 24668 31108 24724 31118
rect 23772 30774 23774 30826
rect 23826 30774 23828 30826
rect 23772 30762 23828 30774
rect 23884 30994 23940 31006
rect 23884 30942 23886 30994
rect 23938 30942 23940 30994
rect 23884 30548 23940 30942
rect 24276 30996 24332 31006
rect 24276 30902 24332 30940
rect 24556 30994 24612 31006
rect 24556 30942 24558 30994
rect 24610 30942 24612 30994
rect 23884 30492 24500 30548
rect 23660 30482 23716 30492
rect 23996 29988 24052 29998
rect 23828 29652 23884 29662
rect 23828 29558 23884 29596
rect 23548 29372 23828 29428
rect 23660 28754 23716 28766
rect 23660 28702 23662 28754
rect 23714 28702 23716 28754
rect 23548 28644 23604 28654
rect 23436 28642 23604 28644
rect 23436 28590 23550 28642
rect 23602 28590 23604 28642
rect 23436 28588 23604 28590
rect 23548 28578 23604 28588
rect 22764 27970 23044 27972
rect 22540 27914 22596 27926
rect 22540 27862 22542 27914
rect 22594 27862 22596 27914
rect 22764 27918 22766 27970
rect 22818 27918 23044 27970
rect 22764 27916 23044 27918
rect 23436 28420 23492 28430
rect 22764 27906 22820 27916
rect 22540 27018 22596 27862
rect 23100 27858 23156 27870
rect 23100 27806 23102 27858
rect 23154 27806 23156 27858
rect 22540 26966 22542 27018
rect 22594 26966 22596 27018
rect 22652 27748 22708 27758
rect 22652 27046 22708 27692
rect 23100 27748 23156 27806
rect 23100 27682 23156 27692
rect 23436 27310 23492 28364
rect 23380 27298 23492 27310
rect 23380 27246 23382 27298
rect 23434 27246 23492 27298
rect 23380 27244 23492 27246
rect 23660 27914 23716 28702
rect 23660 27862 23662 27914
rect 23714 27862 23716 27914
rect 23380 27234 23436 27244
rect 23100 27188 23156 27198
rect 22652 26994 22654 27046
rect 22706 26994 22708 27046
rect 22652 26982 22708 26994
rect 22876 27076 22932 27086
rect 22876 26994 22878 27020
rect 22930 26994 22932 27020
rect 22876 26982 22932 26994
rect 23100 27046 23156 27132
rect 23100 26994 23102 27046
rect 23154 26994 23156 27046
rect 23660 27076 23716 27862
rect 23660 27010 23716 27020
rect 23100 26982 23156 26994
rect 22540 26964 22596 26966
rect 22540 26898 22596 26908
rect 23212 26964 23268 26974
rect 22596 26180 22652 26190
rect 22428 26178 22652 26180
rect 22428 26126 22598 26178
rect 22650 26126 22652 26178
rect 22428 26124 22652 26126
rect 22316 25506 22372 25518
rect 22316 25454 22318 25506
rect 22370 25454 22372 25506
rect 22316 24948 22372 25454
rect 22316 24882 22372 24892
rect 22428 25396 22484 26124
rect 22596 26114 22652 26124
rect 23212 25844 23268 26908
rect 23772 26516 23828 29372
rect 23884 28756 23940 28766
rect 23884 28615 23940 28700
rect 23884 28563 23886 28615
rect 23938 28563 23940 28615
rect 23884 28551 23940 28563
rect 23996 26908 24052 29932
rect 24220 29652 24276 29662
rect 24220 28980 24276 29596
rect 24332 29426 24388 29438
rect 24332 29374 24334 29426
rect 24386 29374 24388 29426
rect 24332 29316 24388 29374
rect 24332 29250 24388 29260
rect 24444 29258 24500 30492
rect 24556 29540 24612 30942
rect 24668 30994 24724 31052
rect 24668 30942 24670 30994
rect 24722 30942 24724 30994
rect 24668 30930 24724 30942
rect 24556 29474 24612 29484
rect 24668 30100 24724 30110
rect 24668 29426 24724 30044
rect 24668 29374 24670 29426
rect 24722 29374 24724 29426
rect 24668 29362 24724 29374
rect 24444 29206 24446 29258
rect 24498 29206 24500 29258
rect 24444 29194 24500 29206
rect 24220 28924 24612 28980
rect 24220 28644 24276 28654
rect 24220 28550 24276 28588
rect 24444 28308 24500 28318
rect 24108 27914 24164 27926
rect 24108 27862 24110 27914
rect 24162 27862 24164 27914
rect 24108 27188 24164 27862
rect 24108 27122 24164 27132
rect 23660 26460 23828 26516
rect 23884 26852 24052 26908
rect 23492 26404 23548 26414
rect 23492 26310 23548 26348
rect 23212 25788 23492 25844
rect 21980 24836 22036 24846
rect 21868 24834 22036 24836
rect 21868 24782 21982 24834
rect 22034 24782 22036 24834
rect 21868 24780 22036 24782
rect 21980 24770 22036 24780
rect 22204 24836 22260 24846
rect 20972 24220 21252 24276
rect 22092 24724 22148 24734
rect 20636 24052 20692 24062
rect 20636 23958 20692 23996
rect 20412 23156 20468 23166
rect 20412 22594 20468 23100
rect 20748 22932 20804 22942
rect 20972 22932 21028 24220
rect 21532 23940 21588 23950
rect 21924 23940 21980 23950
rect 21532 23846 21588 23884
rect 21868 23884 21924 23940
rect 21868 23846 21980 23884
rect 21364 23716 21420 23726
rect 21308 23714 21420 23716
rect 21308 23662 21366 23714
rect 21418 23662 21420 23714
rect 21308 23650 21420 23662
rect 21084 23156 21140 23166
rect 21196 23156 21252 23166
rect 21140 23154 21252 23156
rect 21140 23102 21198 23154
rect 21250 23102 21252 23154
rect 21140 23100 21252 23102
rect 21084 23062 21140 23100
rect 20748 22930 21028 22932
rect 20748 22878 20750 22930
rect 20802 22878 21028 22930
rect 20748 22876 21028 22878
rect 20748 22866 20804 22876
rect 20412 22542 20414 22594
rect 20466 22542 20468 22594
rect 20412 22530 20468 22542
rect 20244 21812 20356 21822
rect 20692 21812 20748 21822
rect 19628 21756 19796 21812
rect 19180 21746 19236 21756
rect 19516 21588 19572 21598
rect 19516 21586 19684 21588
rect 19516 21534 19518 21586
rect 19570 21534 19684 21586
rect 19516 21532 19684 21534
rect 19516 21522 19572 21532
rect 18956 21420 19460 21476
rect 18900 21140 18956 21150
rect 18900 20858 18956 21084
rect 19404 21038 19460 21420
rect 19404 21026 19516 21038
rect 19404 20974 19462 21026
rect 19514 20974 19516 21026
rect 19404 20972 19516 20974
rect 19460 20962 19516 20972
rect 18732 20804 18788 20814
rect 18900 20806 18902 20858
rect 18954 20806 18956 20858
rect 18900 20794 18956 20806
rect 19180 20802 19236 20814
rect 18732 20710 18788 20748
rect 19180 20750 19182 20802
rect 19234 20750 19236 20802
rect 19068 20690 19124 20702
rect 19068 20638 19070 20690
rect 19122 20638 19124 20690
rect 19068 20468 19124 20638
rect 19068 20402 19124 20412
rect 19180 20244 19236 20750
rect 19628 20356 19684 21532
rect 19740 21028 19796 21756
rect 20244 21810 20580 21812
rect 20244 21758 20246 21810
rect 20298 21758 20580 21810
rect 20244 21756 20580 21758
rect 20244 21746 20300 21756
rect 19908 21028 19964 21038
rect 19740 21026 19964 21028
rect 19740 20974 19910 21026
rect 19962 20974 19964 21026
rect 19740 20972 19964 20974
rect 19908 20962 19964 20972
rect 20524 20916 20580 21756
rect 20692 21718 20748 21756
rect 20300 20860 20804 20916
rect 20188 20804 20244 20814
rect 20188 20722 20190 20748
rect 20242 20722 20244 20748
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19628 20300 19740 20356
rect 19836 20346 20100 20356
rect 18060 20242 18564 20244
rect 18060 20190 18510 20242
rect 18562 20190 18564 20242
rect 18060 20188 18564 20190
rect 17780 20178 17836 20188
rect 18508 20178 18564 20188
rect 18956 20188 19236 20244
rect 19684 20244 19740 20300
rect 19684 20188 19796 20244
rect 17500 20020 17556 20030
rect 17500 19926 17556 19964
rect 17836 20018 17892 20030
rect 17836 19966 17838 20018
rect 17890 19966 17892 20018
rect 17836 19796 17892 19966
rect 17388 19740 17892 19796
rect 18844 20020 18900 20030
rect 18956 20020 19012 20188
rect 19572 20132 19628 20142
rect 19572 20038 19628 20076
rect 18844 20018 19012 20020
rect 18844 19966 18846 20018
rect 18898 19966 19012 20018
rect 18844 19964 19012 19966
rect 19068 20018 19124 20030
rect 19068 19966 19070 20018
rect 19122 19966 19124 20018
rect 17388 18788 17444 19740
rect 18340 19684 18396 19694
rect 18340 19290 18396 19628
rect 17500 19234 17556 19246
rect 17500 19182 17502 19234
rect 17554 19182 17556 19234
rect 17500 18900 17556 19182
rect 18060 19236 18116 19246
rect 18340 19238 18342 19290
rect 18394 19238 18396 19290
rect 18340 19226 18396 19238
rect 18508 19234 18564 19246
rect 18060 19142 18116 19180
rect 18508 19182 18510 19234
rect 18562 19182 18564 19234
rect 17780 19124 17836 19134
rect 17780 19030 17836 19068
rect 18172 19122 18228 19134
rect 18508 19124 18564 19182
rect 18172 19070 18174 19122
rect 18226 19070 18228 19122
rect 18172 18900 18228 19070
rect 17500 18844 18228 18900
rect 17388 18732 17556 18788
rect 17276 18386 17332 18396
rect 17388 18477 17444 18489
rect 17388 18425 17390 18477
rect 17442 18425 17444 18477
rect 17388 18340 17444 18425
rect 17052 17948 17220 18004
rect 16604 17444 16660 17454
rect 17164 17444 17220 17948
rect 16604 17106 16660 17388
rect 16604 17054 16606 17106
rect 16658 17054 16660 17106
rect 16604 17042 16660 17054
rect 16940 17388 17220 17444
rect 16268 16930 16324 16940
rect 16156 16884 16212 16894
rect 16044 16772 16100 16782
rect 14364 16370 14420 16380
rect 14980 16492 15316 16548
rect 15596 16770 16100 16772
rect 15596 16718 16046 16770
rect 16098 16718 16100 16770
rect 15596 16716 16100 16718
rect 14980 16210 15036 16492
rect 14980 16158 14982 16210
rect 15034 16158 15036 16210
rect 14980 16146 15036 16158
rect 14140 16042 14196 16054
rect 14140 15990 14142 16042
rect 14194 15990 14196 16042
rect 14140 15540 14196 15990
rect 14924 15988 14980 15998
rect 14756 15876 14812 15886
rect 14140 15484 14532 15540
rect 13916 15262 13918 15314
rect 13970 15262 13972 15314
rect 13916 15250 13972 15262
rect 14196 15316 14252 15326
rect 14196 15222 14252 15260
rect 14476 15314 14532 15484
rect 14756 15370 14812 15820
rect 14476 15262 14478 15314
rect 14530 15262 14532 15314
rect 12460 14532 12516 14542
rect 12460 14438 12516 14476
rect 12684 14530 12740 15092
rect 12852 14980 12908 14990
rect 12852 14754 12908 14924
rect 12852 14702 12854 14754
rect 12906 14702 12908 14754
rect 12852 14690 12908 14702
rect 12684 14478 12686 14530
rect 12738 14478 12740 14530
rect 12684 14466 12740 14478
rect 12348 14420 12404 14430
rect 11564 13746 11844 13748
rect 11564 13694 11566 13746
rect 11618 13694 11844 13746
rect 11564 13692 11844 13694
rect 11900 14196 11956 14206
rect 10892 13524 10948 13534
rect 10892 13522 11396 13524
rect 10892 13470 10894 13522
rect 10946 13470 11396 13522
rect 10892 13468 11396 13470
rect 10892 13458 10948 13468
rect 9996 12012 10164 12068
rect 10220 13244 10612 13300
rect 10220 12066 10276 13244
rect 11340 13074 11396 13468
rect 11340 13022 11342 13074
rect 11394 13022 11396 13074
rect 11340 13010 11396 13022
rect 10220 12014 10222 12066
rect 10274 12014 10276 12066
rect 9324 11900 9772 11956
rect 9716 11506 9772 11900
rect 9716 11454 9718 11506
rect 9770 11454 9772 11506
rect 9716 11442 9772 11454
rect 9100 11396 9156 11406
rect 8932 11338 9044 11363
rect 8932 11286 8934 11338
rect 8986 11286 9044 11338
rect 9100 11302 9156 11340
rect 8932 11274 9044 11286
rect 8988 10948 9044 11274
rect 8988 10892 9716 10948
rect 9660 10778 9716 10892
rect 9660 10726 9662 10778
rect 9714 10726 9716 10778
rect 9660 10714 9716 10726
rect 9996 10651 10052 12012
rect 10220 12002 10276 12014
rect 10780 12740 10836 12750
rect 10780 12178 10836 12684
rect 11564 12740 11620 13692
rect 11900 13300 11956 14140
rect 12348 13746 12404 14364
rect 13020 13972 13076 15092
rect 12348 13694 12350 13746
rect 12402 13694 12404 13746
rect 12348 13682 12404 13694
rect 12572 13916 13076 13972
rect 11900 13234 11956 13244
rect 11564 12674 11620 12684
rect 12124 12962 12180 12974
rect 12124 12910 12126 12962
rect 12178 12910 12180 12962
rect 12124 12740 12180 12910
rect 12572 12964 12628 13916
rect 12964 13412 13020 13422
rect 12964 13074 13020 13356
rect 13468 13188 13524 15148
rect 12964 13022 12966 13074
rect 13018 13022 13020 13074
rect 12964 13010 13020 13022
rect 13356 13132 13524 13188
rect 13692 15092 13860 15148
rect 12572 12908 12740 12964
rect 12124 12674 12180 12684
rect 12516 12740 12572 12750
rect 12516 12646 12572 12684
rect 10780 12126 10782 12178
rect 10834 12126 10836 12178
rect 10108 11844 10164 11854
rect 10108 11394 10164 11788
rect 10108 11342 10110 11394
rect 10162 11342 10164 11394
rect 10108 11330 10164 11342
rect 10780 11844 10836 12126
rect 11564 12068 11620 12078
rect 11564 11974 11620 12012
rect 10780 10846 10836 11788
rect 10892 11394 10948 11406
rect 10892 11342 10894 11394
rect 10946 11342 10948 11394
rect 10892 11284 10948 11342
rect 10892 11218 10948 11228
rect 12684 10846 12740 12908
rect 13356 12740 13412 13132
rect 13356 12674 13412 12684
rect 13468 12962 13524 12974
rect 13468 12910 13470 12962
rect 13522 12910 13524 12962
rect 13468 12066 13524 12910
rect 13692 12964 13748 15092
rect 14476 14756 14532 15262
rect 14588 15314 14644 15326
rect 14588 15262 14590 15314
rect 14642 15262 14644 15314
rect 14756 15318 14758 15370
rect 14810 15318 14812 15370
rect 14756 15306 14812 15318
rect 14924 15314 14980 15932
rect 14588 15148 14644 15262
rect 14924 15262 14926 15314
rect 14978 15262 14980 15314
rect 14924 15204 14980 15262
rect 14588 15092 14756 15148
rect 14924 15138 14980 15148
rect 15148 15148 15204 16492
rect 15596 16098 15652 16716
rect 16044 16706 16100 16716
rect 16044 16212 16100 16222
rect 16156 16212 16212 16828
rect 16940 16882 16996 17388
rect 16940 16830 16942 16882
rect 16994 16830 16996 16882
rect 16492 16772 16548 16782
rect 16044 16210 16212 16212
rect 16044 16158 16046 16210
rect 16098 16158 16212 16210
rect 16044 16156 16212 16158
rect 16268 16324 16324 16334
rect 16044 16146 16100 16156
rect 15596 16046 15598 16098
rect 15650 16046 15652 16098
rect 15596 16034 15652 16046
rect 15820 16100 15876 16110
rect 16268 16100 16324 16268
rect 15820 16006 15876 16044
rect 16156 16083 16324 16100
rect 16156 16031 16158 16083
rect 16210 16044 16324 16083
rect 16492 16098 16548 16716
rect 16828 16212 16884 16222
rect 16940 16212 16996 16830
rect 16828 16210 16996 16212
rect 16828 16158 16830 16210
rect 16882 16158 16996 16210
rect 16828 16156 16996 16158
rect 17052 16324 17108 16334
rect 16828 16146 16884 16156
rect 16492 16046 16494 16098
rect 16546 16046 16548 16098
rect 16210 16031 16212 16044
rect 16492 16034 16548 16046
rect 16604 16100 16660 16110
rect 17052 16100 17108 16268
rect 15316 15988 15372 15998
rect 15316 15986 15540 15988
rect 15316 15934 15318 15986
rect 15370 15934 15540 15986
rect 15316 15932 15540 15934
rect 15316 15922 15372 15932
rect 15148 15092 15316 15148
rect 14476 14700 14644 14756
rect 14028 14532 14084 14542
rect 14476 14532 14532 14542
rect 14028 14438 14084 14476
rect 14252 14474 14308 14486
rect 14252 14422 14254 14474
rect 14306 14422 14308 14474
rect 13860 14308 13916 14318
rect 14252 14308 14308 14422
rect 13860 14306 14308 14308
rect 13860 14254 13862 14306
rect 13914 14254 14308 14306
rect 13860 14252 14308 14254
rect 14364 14474 14420 14486
rect 14364 14422 14366 14474
rect 14418 14422 14420 14474
rect 13860 14242 13916 14252
rect 13804 14084 13860 14094
rect 13804 12964 13860 14028
rect 14364 14084 14420 14422
rect 14364 14018 14420 14028
rect 14252 13748 14308 13758
rect 14252 13654 14308 13692
rect 14476 13748 14532 14476
rect 14588 13776 14644 14700
rect 14700 13972 14756 15092
rect 15260 14530 15316 15092
rect 15484 15092 15540 15932
rect 16156 15876 16212 16031
rect 15764 15820 16212 15876
rect 15764 15538 15820 15820
rect 15764 15486 15766 15538
rect 15818 15486 15820 15538
rect 15764 15148 15820 15486
rect 16604 15538 16660 16044
rect 16940 16083 17108 16100
rect 16940 16031 16942 16083
rect 16994 16044 17108 16083
rect 17276 16098 17332 16110
rect 17276 16046 17278 16098
rect 17330 16046 17332 16098
rect 16994 16031 16996 16044
rect 16940 16019 16996 16031
rect 17276 15988 17332 16046
rect 17388 16100 17444 18284
rect 17388 16034 17444 16044
rect 17276 15922 17332 15932
rect 17500 15764 17556 18732
rect 17612 18564 17668 18574
rect 17612 16882 17668 18508
rect 17948 17668 18004 17678
rect 17948 17574 18004 17612
rect 18172 17668 18228 18844
rect 18396 19068 18564 19124
rect 18396 18452 18452 19068
rect 18844 19012 18900 19964
rect 19068 19908 19124 19966
rect 19068 19842 19124 19852
rect 19292 20018 19348 20030
rect 19292 19966 19294 20018
rect 19346 19966 19348 20018
rect 19180 19796 19236 19806
rect 19068 19460 19124 19470
rect 19068 19234 19124 19404
rect 19068 19182 19070 19234
rect 19122 19182 19124 19234
rect 19068 19170 19124 19182
rect 18172 17602 18228 17612
rect 18284 18396 18452 18452
rect 18508 18956 18900 19012
rect 17612 16830 17614 16882
rect 17666 16830 17668 16882
rect 17948 17444 18004 17454
rect 18284 17444 18340 18396
rect 18508 17902 18564 18956
rect 19180 18788 19236 19740
rect 19292 19572 19348 19966
rect 19740 20020 19796 20188
rect 20188 20132 20244 20722
rect 20188 20074 20244 20076
rect 20188 20022 20190 20074
rect 20242 20022 20244 20074
rect 20188 20010 20244 20022
rect 19740 19954 19796 19964
rect 20300 19908 20356 20860
rect 20748 20767 20804 20860
rect 20412 20746 20468 20758
rect 20412 20694 20414 20746
rect 20466 20694 20468 20746
rect 20412 20132 20468 20694
rect 20636 20746 20692 20758
rect 20636 20694 20638 20746
rect 20690 20694 20692 20746
rect 20748 20715 20750 20767
rect 20802 20715 20804 20767
rect 20748 20703 20804 20715
rect 20636 20244 20692 20694
rect 20636 20188 20804 20244
rect 20412 20076 20692 20132
rect 20188 19852 20356 19908
rect 20636 20074 20692 20076
rect 20636 20022 20638 20074
rect 20690 20022 20692 20074
rect 19292 19506 19348 19516
rect 19628 19684 19684 19694
rect 19516 19460 19572 19470
rect 19292 19348 19348 19358
rect 19292 19195 19348 19292
rect 19292 19143 19294 19195
rect 19346 19143 19348 19195
rect 19292 19131 19348 19143
rect 19180 18722 19236 18732
rect 19404 19066 19460 19078
rect 19404 19014 19406 19066
rect 19458 19014 19460 19066
rect 18732 18452 18788 18462
rect 18452 17890 18564 17902
rect 18452 17838 18454 17890
rect 18506 17838 18564 17890
rect 18452 17836 18564 17838
rect 18620 18396 18732 18452
rect 18452 17826 18508 17836
rect 17948 16926 18004 17388
rect 17948 16874 17950 16926
rect 18002 16874 18004 16926
rect 17948 16862 18004 16874
rect 18060 17388 18340 17444
rect 18060 16996 18116 17388
rect 17612 16324 17668 16830
rect 18060 16770 18116 16940
rect 18060 16718 18062 16770
rect 18114 16718 18116 16770
rect 18060 16706 18116 16718
rect 17612 16258 17668 16268
rect 18508 16658 18564 16670
rect 18508 16606 18510 16658
rect 18562 16606 18564 16658
rect 16604 15486 16606 15538
rect 16658 15486 16660 15538
rect 15484 15026 15540 15036
rect 15596 15092 15820 15148
rect 16212 15428 16268 15438
rect 16212 15204 16268 15372
rect 16212 15138 16268 15148
rect 16604 15204 16660 15486
rect 17276 15708 17556 15764
rect 17836 16098 17892 16110
rect 17836 16046 17838 16098
rect 17890 16046 17892 16098
rect 16940 15316 16996 15326
rect 17276 15316 17332 15708
rect 16940 15314 17332 15316
rect 16940 15262 16942 15314
rect 16994 15262 17332 15314
rect 16940 15260 17332 15262
rect 17388 15316 17444 15326
rect 16940 15250 16996 15260
rect 16604 15138 16660 15148
rect 15092 14474 15148 14486
rect 14924 14420 14980 14430
rect 14924 14326 14980 14364
rect 15092 14422 15094 14474
rect 15146 14422 15148 14474
rect 15260 14478 15262 14530
rect 15314 14478 15316 14530
rect 15260 14466 15316 14478
rect 15092 14420 15148 14422
rect 15092 14354 15148 14364
rect 14700 13906 14756 13916
rect 15596 13860 15652 15092
rect 16044 14644 16100 14654
rect 16044 14550 16100 14588
rect 15484 13804 15652 13860
rect 16268 13916 16660 13972
rect 14588 13748 15092 13776
rect 15148 13774 15204 13786
rect 15148 13748 15150 13774
rect 14588 13722 15150 13748
rect 15202 13722 15204 13774
rect 14588 13720 15204 13722
rect 14476 13682 14532 13692
rect 15036 13692 15204 13720
rect 15372 13748 15428 13758
rect 14924 13636 14980 13646
rect 14812 13188 14868 13198
rect 14700 13132 14812 13188
rect 14028 12964 14084 12974
rect 13804 12908 13972 12964
rect 13692 12898 13748 12908
rect 13636 12794 13692 12806
rect 13636 12742 13638 12794
rect 13690 12742 13692 12794
rect 13636 12292 13692 12742
rect 13636 12226 13692 12236
rect 13804 12740 13860 12750
rect 13916 12740 13972 12908
rect 14028 12962 14196 12964
rect 14028 12910 14030 12962
rect 14082 12910 14196 12962
rect 14028 12908 14196 12910
rect 14028 12898 14084 12908
rect 13916 12684 14028 12740
rect 13468 12014 13470 12066
rect 13522 12014 13524 12066
rect 10780 10836 10892 10846
rect 11284 10836 11340 10846
rect 11732 10836 11788 10846
rect 12180 10836 12236 10846
rect 9940 10639 10052 10651
rect 8876 10612 8932 10622
rect 9548 10612 9604 10622
rect 8876 10610 9604 10612
rect 8876 10558 8878 10610
rect 8930 10558 9550 10610
rect 9602 10558 9604 10610
rect 8876 10556 9604 10558
rect 9940 10587 9942 10639
rect 9994 10612 10052 10639
rect 10556 10834 12236 10836
rect 10556 10782 10838 10834
rect 10890 10782 11286 10834
rect 11338 10782 11734 10834
rect 11786 10782 12182 10834
rect 12234 10782 12236 10834
rect 10556 10780 12236 10782
rect 9994 10587 10164 10612
rect 9940 10556 10164 10587
rect 8876 10546 8932 10556
rect 8876 9940 8932 9950
rect 8652 9650 8708 9660
rect 8764 9938 8932 9940
rect 8764 9886 8878 9938
rect 8930 9886 8932 9938
rect 8764 9884 8932 9886
rect 8428 9548 8596 9604
rect 8204 9042 8372 9044
rect 8204 8990 8206 9042
rect 8258 8990 8372 9042
rect 8204 8988 8372 8990
rect 8204 8978 8260 8988
rect 7756 8194 7812 8204
rect 8204 8260 8260 8270
rect 8204 8166 8260 8204
rect 7532 7700 7588 7710
rect 7532 7642 7588 7644
rect 7532 7590 7534 7642
rect 7586 7590 7588 7642
rect 7532 7578 7588 7590
rect 8316 7588 8372 8988
rect 8428 9069 8484 9081
rect 8428 9017 8430 9069
rect 8482 9017 8484 9069
rect 8428 8932 8484 9017
rect 8428 8866 8484 8876
rect 8540 8214 8596 9548
rect 8764 9042 8820 9884
rect 8876 9874 8932 9884
rect 9212 9826 9268 10556
rect 9548 10546 9604 10556
rect 8988 9782 9044 9794
rect 8988 9730 8990 9782
rect 9042 9730 9044 9782
rect 9212 9774 9214 9826
rect 9266 9774 9268 9826
rect 9212 9762 9268 9774
rect 10108 9826 10164 10556
rect 10556 9950 10612 10780
rect 10836 10770 10892 10780
rect 11284 10770 11340 10780
rect 11452 9950 11508 10780
rect 11732 10770 11788 10780
rect 12180 10770 12236 10780
rect 12628 10834 12740 10846
rect 12628 10782 12630 10834
rect 12682 10782 12740 10834
rect 12628 10780 12740 10782
rect 12796 11282 12852 11294
rect 12796 11230 12798 11282
rect 12850 11230 12852 11282
rect 12628 10770 12684 10780
rect 12796 10724 12852 11230
rect 12796 10658 12852 10668
rect 13356 10948 13412 10958
rect 13020 10610 13076 10622
rect 13020 10558 13022 10610
rect 13074 10558 13076 10610
rect 10108 9774 10110 9826
rect 10162 9774 10164 9826
rect 10108 9762 10164 9774
rect 10500 9938 10612 9950
rect 10500 9886 10502 9938
rect 10554 9886 10612 9938
rect 10500 9884 10612 9886
rect 11396 9940 11508 9950
rect 12124 10052 12180 10062
rect 11396 9938 11620 9940
rect 11396 9886 11398 9938
rect 11450 9886 11620 9938
rect 11396 9884 11620 9886
rect 8988 9716 9044 9730
rect 8988 9650 9044 9660
rect 9772 9604 9828 9614
rect 9772 9602 9940 9604
rect 9772 9550 9774 9602
rect 9826 9550 9940 9602
rect 9772 9548 9940 9550
rect 9772 9538 9828 9548
rect 8764 8990 8766 9042
rect 8818 8990 8820 9042
rect 8764 8978 8820 8990
rect 8876 9210 8932 9222
rect 8876 9158 8878 9210
rect 8930 9158 8932 9210
rect 8876 9044 8932 9158
rect 9436 9044 9492 9054
rect 8876 9042 9492 9044
rect 8876 8990 9438 9042
rect 9490 8990 9492 9042
rect 8876 8988 9492 8990
rect 9436 8978 9492 8988
rect 9772 8818 9828 8830
rect 9772 8766 9774 8818
rect 9826 8766 9828 8818
rect 8540 8162 8542 8214
rect 8594 8162 8596 8214
rect 8540 7812 8596 8162
rect 8652 8370 8708 8382
rect 8652 8318 8654 8370
rect 8706 8318 8708 8370
rect 8652 7924 8708 8318
rect 9772 8372 9828 8766
rect 9772 8306 9828 8316
rect 9100 8260 9156 8270
rect 9100 8166 9156 8204
rect 9884 8260 9940 9548
rect 10500 9268 10556 9884
rect 11396 9874 11452 9884
rect 10500 9266 10724 9268
rect 10500 9214 10502 9266
rect 10554 9214 10724 9266
rect 10500 9212 10724 9214
rect 10500 9202 10556 9212
rect 10668 9042 10724 9212
rect 10668 8990 10670 9042
rect 10722 8990 10724 9042
rect 10668 8978 10724 8990
rect 11452 9044 11508 9054
rect 11452 8950 11508 8988
rect 11564 8708 11620 9884
rect 12124 9793 12180 9996
rect 13020 10052 13076 10558
rect 13244 10612 13300 10622
rect 13244 10518 13300 10556
rect 13356 10442 13412 10892
rect 13468 10612 13524 12014
rect 13804 11528 13860 12684
rect 13972 12628 14028 12684
rect 13972 12572 14084 12628
rect 13916 12292 13972 12302
rect 13916 12234 13972 12236
rect 13916 12182 13918 12234
rect 13970 12182 13972 12234
rect 13916 12170 13972 12182
rect 14028 12234 14084 12572
rect 14028 12182 14030 12234
rect 14082 12182 14084 12234
rect 14028 12170 14084 12182
rect 13748 11506 13860 11528
rect 13748 11454 13750 11506
rect 13802 11454 13860 11506
rect 13748 11442 13860 11454
rect 13804 11363 13860 11442
rect 14140 11396 14196 12908
rect 14700 12852 14756 13132
rect 14812 13122 14868 13132
rect 14924 12974 14980 13580
rect 14904 12962 14980 12974
rect 14904 12910 14906 12962
rect 14958 12910 14980 12962
rect 14904 12908 14980 12910
rect 14904 12898 14960 12908
rect 14700 12796 14812 12852
rect 14028 11363 14084 11373
rect 13804 11361 14084 11363
rect 13804 11309 14030 11361
rect 14082 11309 14084 11361
rect 14476 12628 14532 12638
rect 14140 11330 14196 11340
rect 14364 11338 14420 11350
rect 13804 11307 14084 11309
rect 14028 11172 14084 11307
rect 14028 11106 14084 11116
rect 14364 11286 14366 11338
rect 14418 11286 14420 11338
rect 14364 10948 14420 11286
rect 14364 10882 14420 10892
rect 13962 10724 14018 10734
rect 13962 10660 14018 10668
rect 13692 10612 13748 10622
rect 13468 10610 13748 10612
rect 13468 10558 13694 10610
rect 13746 10558 13748 10610
rect 13468 10556 13748 10558
rect 13692 10546 13748 10556
rect 13804 10610 13860 10622
rect 13804 10558 13806 10610
rect 13858 10558 13860 10610
rect 13962 10608 13964 10660
rect 14016 10608 14018 10660
rect 13962 10596 14018 10608
rect 14364 10612 14420 10622
rect 13356 10390 13358 10442
rect 13410 10390 13412 10442
rect 13356 10378 13412 10390
rect 13804 10388 13860 10558
rect 14364 10498 14420 10556
rect 14364 10446 14366 10498
rect 14418 10446 14420 10498
rect 14364 10434 14420 10446
rect 13804 10322 13860 10332
rect 14476 10164 14532 12572
rect 14756 12234 14812 12796
rect 14756 12182 14758 12234
rect 14810 12182 14812 12234
rect 14756 12170 14812 12182
rect 14588 12068 14644 12078
rect 14588 11974 14644 12012
rect 15036 11844 15092 13692
rect 15372 13654 15428 13692
rect 15148 13524 15204 13534
rect 15148 13186 15204 13468
rect 15484 13412 15540 13804
rect 16156 13784 16212 13796
rect 15764 13748 15820 13758
rect 15764 13654 15820 13692
rect 16156 13732 16158 13784
rect 16210 13732 16212 13784
rect 15596 13636 15652 13646
rect 15596 13542 15652 13580
rect 16156 13524 16212 13732
rect 16156 13458 16212 13468
rect 15148 13134 15150 13186
rect 15202 13134 15204 13186
rect 15148 13122 15204 13134
rect 15372 13356 15540 13412
rect 15372 12414 15428 13356
rect 15316 12402 15428 12414
rect 15316 12350 15318 12402
rect 15370 12350 15428 12402
rect 15316 12338 15428 12350
rect 14588 11788 15092 11844
rect 14588 10388 14644 11788
rect 14812 11396 14868 11406
rect 14812 11309 14814 11340
rect 14866 11309 14868 11340
rect 14812 11060 14868 11309
rect 15122 11396 15178 11406
rect 15122 11309 15124 11340
rect 15176 11309 15178 11340
rect 15122 11297 15178 11309
rect 15260 11284 15316 11294
rect 15260 11190 15316 11228
rect 14812 11004 15260 11060
rect 15204 10722 15260 11004
rect 15372 10836 15428 12338
rect 15372 10770 15428 10780
rect 15484 13076 15540 13086
rect 15484 12962 15540 13020
rect 16268 13074 16324 13916
rect 16604 13860 16660 13916
rect 16716 13860 16772 13870
rect 16604 13858 16772 13860
rect 16604 13806 16718 13858
rect 16770 13806 16772 13858
rect 16604 13804 16772 13806
rect 16716 13794 16772 13804
rect 16268 13022 16270 13074
rect 16322 13022 16324 13074
rect 16268 13010 16324 13022
rect 16380 13748 16436 13758
rect 15484 12910 15486 12962
rect 15538 12910 15540 12962
rect 15204 10670 15206 10722
rect 15258 10670 15260 10722
rect 15204 10658 15260 10670
rect 14588 10322 14644 10332
rect 14700 10610 14756 10622
rect 14700 10558 14702 10610
rect 14754 10558 14756 10610
rect 14476 10108 14644 10164
rect 13020 9986 13076 9996
rect 13524 10052 13580 10062
rect 14364 10052 14420 10062
rect 13524 9958 13580 9996
rect 13804 10050 14420 10052
rect 13804 9998 14366 10050
rect 14418 9998 14420 10050
rect 13804 9996 14420 9998
rect 11844 9770 11900 9782
rect 11676 9714 11732 9726
rect 11676 9662 11678 9714
rect 11730 9662 11732 9714
rect 11676 9044 11732 9662
rect 11844 9718 11846 9770
rect 11898 9718 11900 9770
rect 12124 9741 12126 9793
rect 12178 9741 12180 9793
rect 13804 9826 13860 9996
rect 14364 9986 14420 9996
rect 12124 9729 12180 9741
rect 12572 9770 12628 9782
rect 11844 9492 11900 9718
rect 11844 9426 11900 9436
rect 12572 9718 12574 9770
rect 12626 9718 12628 9770
rect 11676 8978 11732 8988
rect 12572 8820 12628 9718
rect 12908 9770 12964 9782
rect 12908 9718 12910 9770
rect 12962 9718 12964 9770
rect 12908 9268 12964 9718
rect 13804 9774 13806 9826
rect 13858 9774 13860 9826
rect 13468 9492 13524 9502
rect 12908 9202 12964 9212
rect 13356 9380 13412 9390
rect 13356 9156 13412 9324
rect 12572 8754 12628 8764
rect 13020 9154 13412 9156
rect 13020 9102 13358 9154
rect 13410 9102 13412 9154
rect 13020 9100 13412 9102
rect 11564 8652 11844 8708
rect 11004 8372 11060 8382
rect 11004 8278 11060 8316
rect 9884 8194 9940 8204
rect 10892 8260 10948 8270
rect 8652 7868 9940 7924
rect 8540 7756 9156 7812
rect 7980 7501 8036 7513
rect 7084 7474 7252 7476
rect 7084 7422 7086 7474
rect 7138 7422 7252 7474
rect 7084 7420 7252 7422
rect 7084 7410 7140 7420
rect 6636 7196 6804 7252
rect 6524 6804 6580 6814
rect 6300 6802 6580 6804
rect 6300 6750 6526 6802
rect 6578 6750 6580 6802
rect 6300 6748 6580 6750
rect 6524 6738 6580 6748
rect 6076 6692 6132 6702
rect 5964 6690 6132 6692
rect 5964 6638 6078 6690
rect 6130 6638 6132 6690
rect 5964 6636 6132 6638
rect 5796 6598 5852 6636
rect 6076 6626 6132 6636
rect 6412 6646 6468 6658
rect 6412 6594 6414 6646
rect 6466 6594 6468 6646
rect 6412 6580 6468 6594
rect 6636 6580 6692 7196
rect 7084 6692 7140 6702
rect 7084 6598 7140 6636
rect 6412 6524 6692 6580
rect 4844 5906 5012 5908
rect 4844 5854 4846 5906
rect 4898 5854 5012 5906
rect 4844 5852 5012 5854
rect 5628 6468 5684 6478
rect 5628 5906 5684 6412
rect 7196 6020 7252 7420
rect 7644 7476 7700 7486
rect 7644 7382 7700 7420
rect 7980 7449 7982 7501
rect 8034 7449 8036 7501
rect 7868 6690 7924 6702
rect 7868 6638 7870 6690
rect 7922 6638 7924 6690
rect 7868 6132 7924 6638
rect 7868 6066 7924 6076
rect 7532 6020 7588 6030
rect 7196 6018 7588 6020
rect 7196 5966 7534 6018
rect 7586 5966 7588 6018
rect 7196 5964 7588 5966
rect 7532 5954 7588 5964
rect 5628 5854 5630 5906
rect 5682 5854 5684 5906
rect 4844 5842 4900 5852
rect 5628 5842 5684 5854
rect 7980 5796 8036 7449
rect 8316 7474 8372 7532
rect 8316 7422 8318 7474
rect 8370 7422 8372 7474
rect 8316 7410 8372 7422
rect 8988 6804 9044 6814
rect 8148 6692 8204 6702
rect 8148 6130 8204 6636
rect 8148 6078 8150 6130
rect 8202 6078 8204 6130
rect 8148 6066 8204 6078
rect 8708 5935 8764 5947
rect 8708 5883 8710 5935
rect 8762 5908 8764 5935
rect 8762 5883 8932 5908
rect 8708 5852 8932 5883
rect 7980 5730 8036 5740
rect 8540 5796 8596 5806
rect 8540 5702 8596 5740
rect 8876 5684 8932 5852
rect 8988 5906 9044 6748
rect 8988 5854 8990 5906
rect 9042 5854 9044 5906
rect 8988 5842 9044 5854
rect 9100 5684 9156 7756
rect 9772 7642 9828 7654
rect 9548 7588 9604 7598
rect 9548 7474 9604 7532
rect 9772 7590 9774 7642
rect 9826 7590 9828 7642
rect 9548 7422 9550 7474
rect 9602 7422 9604 7474
rect 9548 7410 9604 7422
rect 9660 7476 9716 7486
rect 9660 6804 9716 7420
rect 9772 6804 9828 7590
rect 9884 7530 9940 7868
rect 9884 7478 9886 7530
rect 9938 7478 9940 7530
rect 10892 7518 10948 8204
rect 11788 8258 11844 8652
rect 12180 8372 12236 8382
rect 12180 8278 12236 8316
rect 11788 8206 11790 8258
rect 11842 8206 11844 8258
rect 11788 8194 11844 8206
rect 12516 8260 12572 8270
rect 12516 8166 12572 8204
rect 12796 8258 12852 8270
rect 12796 8206 12798 8258
rect 12850 8206 12852 8258
rect 12068 8148 12124 8158
rect 12068 7698 12124 8092
rect 12068 7646 12070 7698
rect 12122 7646 12124 7698
rect 12068 7634 12124 7646
rect 12796 7700 12852 8206
rect 13020 8258 13076 9100
rect 13356 9090 13412 9100
rect 13468 8426 13524 9436
rect 13804 9044 13860 9774
rect 14028 9826 14084 9838
rect 14028 9774 14030 9826
rect 14082 9774 14084 9826
rect 13916 9044 13972 9054
rect 13804 9042 13972 9044
rect 13804 8990 13918 9042
rect 13970 8990 13972 9042
rect 13804 8988 13972 8990
rect 14028 9044 14084 9774
rect 14476 9380 14532 9390
rect 14252 9044 14308 9054
rect 14028 9042 14420 9044
rect 14028 8990 14254 9042
rect 14306 8990 14420 9042
rect 14028 8988 14420 8990
rect 13916 8978 13972 8988
rect 14252 8978 14308 8988
rect 13804 8874 13860 8886
rect 13804 8822 13806 8874
rect 13858 8822 13860 8874
rect 13804 8820 13860 8822
rect 13804 8754 13860 8764
rect 13468 8374 13470 8426
rect 13522 8374 13524 8426
rect 13468 8362 13524 8374
rect 13020 8206 13022 8258
rect 13074 8206 13076 8258
rect 13020 8194 13076 8206
rect 13580 8260 13636 8270
rect 13580 8166 13636 8204
rect 13804 8258 13860 8270
rect 13804 8206 13806 8258
rect 13858 8206 13860 8258
rect 13804 8148 13860 8206
rect 13804 8082 13860 8092
rect 14252 8148 14308 8158
rect 12796 7634 12852 7644
rect 13860 7700 13916 7710
rect 9884 7466 9940 7478
rect 10220 7474 10276 7486
rect 10220 7422 10222 7474
rect 10274 7422 10276 7474
rect 10892 7466 10894 7518
rect 10946 7466 10948 7518
rect 13468 7588 13524 7598
rect 10892 7454 10948 7466
rect 11116 7476 11172 7486
rect 10220 7364 10276 7422
rect 11116 7382 11172 7420
rect 12684 7474 12740 7486
rect 12684 7422 12686 7474
rect 12738 7422 12740 7474
rect 10780 7364 10836 7374
rect 10220 7362 10836 7364
rect 10220 7310 10782 7362
rect 10834 7310 10836 7362
rect 10220 7308 10836 7310
rect 10780 7298 10836 7308
rect 12684 7364 12740 7422
rect 12684 7298 12740 7308
rect 12796 7476 12852 7486
rect 12404 7250 12460 7262
rect 12404 7198 12406 7250
rect 12458 7198 12460 7250
rect 9772 6748 10052 6804
rect 9660 6580 9716 6748
rect 9772 6580 9828 6590
rect 9660 6578 9828 6580
rect 9660 6526 9774 6578
rect 9826 6526 9828 6578
rect 9660 6524 9828 6526
rect 9772 6514 9828 6524
rect 9660 6132 9716 6142
rect 9660 6038 9716 6076
rect 9996 5906 10052 6748
rect 10892 6802 10948 6814
rect 10892 6750 10894 6802
rect 10946 6750 10948 6802
rect 10108 6692 10164 6702
rect 10108 6598 10164 6636
rect 10388 6692 10444 6702
rect 10388 6132 10444 6636
rect 10388 6038 10444 6076
rect 10892 6020 10948 6750
rect 12404 6692 12460 7198
rect 12404 6626 12460 6636
rect 12796 6690 12852 7420
rect 12908 7476 12964 7486
rect 12908 7474 13412 7476
rect 12908 7422 12910 7474
rect 12962 7422 13412 7474
rect 12908 7420 13412 7422
rect 12908 7410 12964 7420
rect 13188 7252 13244 7262
rect 12796 6638 12798 6690
rect 12850 6638 12852 6690
rect 12796 6626 12852 6638
rect 12908 7250 13244 7252
rect 12908 7198 13190 7250
rect 13242 7198 13244 7250
rect 12908 7196 13244 7198
rect 10892 5954 10948 5964
rect 11900 6132 11956 6142
rect 9996 5854 9998 5906
rect 10050 5854 10052 5906
rect 9996 5842 10052 5854
rect 8876 5628 9156 5684
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 11732 4564 11788 4574
rect 11900 4564 11956 6076
rect 12068 6132 12124 6142
rect 12068 6038 12124 6076
rect 12348 6020 12404 6030
rect 12348 5926 12404 5964
rect 12796 6020 12852 6030
rect 12796 5962 12852 5964
rect 12507 5939 12563 5951
rect 12507 5887 12509 5939
rect 12561 5908 12563 5939
rect 12796 5910 12798 5962
rect 12850 5910 12852 5962
rect 12561 5887 12572 5908
rect 12796 5898 12852 5910
rect 12507 5852 12572 5887
rect 12516 5684 12572 5852
rect 12516 5628 12628 5684
rect 12572 5290 12628 5628
rect 12572 5238 12574 5290
rect 12626 5238 12628 5290
rect 12572 5226 12628 5238
rect 11732 4562 11956 4564
rect 11732 4510 11734 4562
rect 11786 4510 11956 4562
rect 11732 4508 11956 4510
rect 11732 4498 11788 4508
rect 11900 4338 11956 4508
rect 11900 4286 11902 4338
rect 11954 4286 11956 4338
rect 11900 4274 11956 4286
rect 12572 5122 12628 5134
rect 12572 5070 12574 5122
rect 12626 5070 12628 5122
rect 12572 4004 12628 5070
rect 12796 5124 12852 5134
rect 12908 5124 12964 7196
rect 13188 7186 13244 7196
rect 13132 6692 13188 6702
rect 13132 5962 13188 6636
rect 13132 5910 13134 5962
rect 13186 5910 13188 5962
rect 13132 5898 13188 5910
rect 13356 5908 13412 7420
rect 13468 7474 13524 7532
rect 13468 7422 13470 7474
rect 13522 7422 13524 7474
rect 13468 7410 13524 7422
rect 13580 7588 13636 7598
rect 13580 6916 13636 7532
rect 13860 7530 13916 7644
rect 13692 7476 13748 7486
rect 13860 7478 13862 7530
rect 13914 7478 13916 7530
rect 13860 7476 13916 7478
rect 13748 7420 13916 7476
rect 14140 7476 14196 7486
rect 13692 7382 13748 7420
rect 14028 7364 14084 7374
rect 13804 7308 14028 7364
rect 13580 6860 13662 6916
rect 13606 6804 13662 6860
rect 13606 6748 13748 6804
rect 13580 6634 13636 6646
rect 13356 5842 13412 5852
rect 13468 6580 13524 6590
rect 13468 5962 13524 6524
rect 13468 5910 13470 5962
rect 13522 5910 13524 5962
rect 13468 5236 13524 5910
rect 13580 6582 13582 6634
rect 13634 6582 13636 6634
rect 13580 5908 13636 6582
rect 13580 5842 13636 5852
rect 13692 5460 13748 6748
rect 13804 6692 13860 7308
rect 14028 7270 14084 7308
rect 14140 6916 14196 7420
rect 14252 7474 14308 8092
rect 14252 7422 14254 7474
rect 14306 7422 14308 7474
rect 14252 7410 14308 7422
rect 13804 6598 13860 6636
rect 13916 6860 14196 6916
rect 14252 6916 14308 6926
rect 14364 6916 14420 8988
rect 14476 8258 14532 9324
rect 14588 9044 14644 10108
rect 14700 10052 14756 10558
rect 14924 10612 14980 10622
rect 14924 10518 14980 10556
rect 14700 9986 14756 9996
rect 15036 10500 15092 10510
rect 14924 9826 14980 9838
rect 14756 9770 14812 9782
rect 14756 9718 14758 9770
rect 14810 9718 14812 9770
rect 14756 9380 14812 9718
rect 14756 9314 14812 9324
rect 14924 9774 14926 9826
rect 14978 9774 14980 9826
rect 14700 9044 14756 9054
rect 14588 9042 14756 9044
rect 14588 8990 14702 9042
rect 14754 8990 14756 9042
rect 14588 8988 14756 8990
rect 14476 8206 14478 8258
rect 14530 8206 14532 8258
rect 14476 8194 14532 8206
rect 14588 8484 14644 8494
rect 14588 7530 14644 8428
rect 14700 8372 14756 8988
rect 14924 8596 14980 9774
rect 15036 9826 15092 10444
rect 15036 9774 15038 9826
rect 15090 9774 15092 9826
rect 15036 9762 15092 9774
rect 15372 10388 15428 10398
rect 15260 9604 15316 9614
rect 15372 9604 15428 10332
rect 15484 9828 15540 12910
rect 16156 12516 16212 12526
rect 15708 12180 15764 12190
rect 16044 12180 16100 12190
rect 16156 12180 16212 12460
rect 15708 12178 15876 12180
rect 15708 12126 15710 12178
rect 15762 12126 15876 12178
rect 15708 12124 15876 12126
rect 15708 12114 15764 12124
rect 15596 12010 15652 12022
rect 15596 11958 15598 12010
rect 15650 11958 15652 12010
rect 15596 11396 15652 11958
rect 15820 11732 15876 12124
rect 16044 12178 16212 12180
rect 16044 12126 16046 12178
rect 16098 12126 16212 12178
rect 16044 12124 16212 12126
rect 16044 12114 16100 12124
rect 15820 11676 16044 11732
rect 15988 11618 16044 11676
rect 15988 11566 15990 11618
rect 16042 11566 16044 11618
rect 15988 11554 16044 11566
rect 16156 11396 16212 12124
rect 16380 11732 16436 13692
rect 16380 11666 16436 11676
rect 16492 13746 16548 13758
rect 16492 13694 16494 13746
rect 16546 13694 16548 13746
rect 16492 13412 16548 13694
rect 16884 13690 16940 13702
rect 16884 13638 16886 13690
rect 16938 13638 16940 13690
rect 16884 13636 16940 13638
rect 16884 13570 16940 13580
rect 15596 11330 15652 11340
rect 16044 11340 16212 11396
rect 16268 11394 16324 11406
rect 16268 11342 16270 11394
rect 16322 11342 16324 11394
rect 15596 11172 15652 11182
rect 15596 10052 15652 11116
rect 15764 10836 15820 10846
rect 15764 10742 15820 10780
rect 15596 9996 15764 10052
rect 15596 9828 15652 9838
rect 15484 9826 15652 9828
rect 15484 9774 15598 9826
rect 15650 9774 15652 9826
rect 15484 9772 15652 9774
rect 15596 9762 15652 9772
rect 15372 9548 15652 9604
rect 15036 9268 15092 9278
rect 15036 9174 15092 9212
rect 14924 8530 14980 8540
rect 14700 8306 14756 8316
rect 14924 8370 14980 8382
rect 14924 8318 14926 8370
rect 14978 8318 14980 8370
rect 14812 8214 14868 8226
rect 14812 8162 14814 8214
rect 14866 8162 14868 8214
rect 14812 7700 14868 8162
rect 14812 7634 14868 7644
rect 14588 7478 14590 7530
rect 14642 7478 14644 7530
rect 14588 7466 14644 7478
rect 14924 7476 14980 8318
rect 15260 8260 15316 9548
rect 15596 9266 15652 9548
rect 15596 9214 15598 9266
rect 15650 9214 15652 9266
rect 15596 9202 15652 9214
rect 15708 8932 15764 9996
rect 16044 9604 16100 11340
rect 16044 9538 16100 9548
rect 16156 10648 16212 10660
rect 16156 10596 16158 10648
rect 16210 10596 16212 10648
rect 15540 8876 15764 8932
rect 15932 9042 15988 9054
rect 15932 8990 15934 9042
rect 15986 8990 15988 9042
rect 15540 8370 15596 8876
rect 15932 8484 15988 8990
rect 15932 8418 15988 8428
rect 16156 8372 16212 10596
rect 16268 9156 16324 11342
rect 16380 11396 16436 11406
rect 16380 10724 16436 11340
rect 16380 10658 16436 10668
rect 16492 10612 16548 13356
rect 17388 12740 17444 15260
rect 17500 15316 17556 15326
rect 17836 15316 17892 16046
rect 17500 15314 17892 15316
rect 17500 15262 17502 15314
rect 17554 15262 17892 15314
rect 17500 15260 17892 15262
rect 17948 15988 18004 15998
rect 17500 13076 17556 15260
rect 17948 14642 18004 15932
rect 17948 14590 17950 14642
rect 18002 14590 18004 14642
rect 17948 14578 18004 14590
rect 18396 14644 18452 14654
rect 18396 14550 18452 14588
rect 18508 14515 18564 16606
rect 18620 15316 18676 18396
rect 18732 18358 18788 18396
rect 18844 18340 18900 18350
rect 18844 17892 18900 18284
rect 18732 17836 18900 17892
rect 18732 17666 18788 17836
rect 19292 17780 19348 17790
rect 18732 17614 18734 17666
rect 18786 17614 18788 17666
rect 18732 16884 18788 17614
rect 18844 17668 18900 17678
rect 18844 17574 18900 17612
rect 19012 17668 19068 17678
rect 19012 17574 19068 17612
rect 19180 17666 19236 17678
rect 19180 17614 19182 17666
rect 19234 17614 19236 17666
rect 19180 17556 19236 17614
rect 19180 17490 19236 17500
rect 18732 16818 18788 16828
rect 18922 16919 18978 16931
rect 18922 16867 18924 16919
rect 18976 16867 18978 16919
rect 18922 16436 18978 16867
rect 19068 16884 19124 16894
rect 19068 16790 19124 16828
rect 19180 16882 19236 16894
rect 19180 16830 19182 16882
rect 19234 16830 19236 16882
rect 19180 16772 19236 16830
rect 19068 16660 19124 16670
rect 18922 16380 19012 16436
rect 18956 15428 19012 16380
rect 18956 15362 19012 15372
rect 18732 15316 18788 15326
rect 18676 15314 18788 15316
rect 18676 15262 18734 15314
rect 18786 15262 18788 15314
rect 18676 15260 18788 15262
rect 18620 15222 18676 15260
rect 18732 15250 18788 15260
rect 18508 14463 18510 14515
rect 18562 14463 18564 14515
rect 18508 14451 18564 14463
rect 18732 14530 18788 14542
rect 18732 14478 18734 14530
rect 18786 14478 18788 14530
rect 17612 13748 17668 13758
rect 17612 13654 17668 13692
rect 17836 13746 17892 13758
rect 17836 13694 17838 13746
rect 17890 13694 17892 13746
rect 17556 13020 17668 13076
rect 17500 13010 17556 13020
rect 16884 12684 17444 12740
rect 16884 12402 16940 12684
rect 16884 12350 16886 12402
rect 16938 12350 16940 12402
rect 16884 12338 16940 12350
rect 17500 12180 17556 12190
rect 17500 12086 17556 12124
rect 17388 12010 17444 12022
rect 17388 11958 17390 12010
rect 17442 11958 17444 12010
rect 16716 11732 16772 11742
rect 16716 11394 16772 11676
rect 17164 11508 17220 11518
rect 17164 11414 17220 11452
rect 16716 11342 16718 11394
rect 16770 11342 16772 11394
rect 16716 11330 16772 11342
rect 17052 11396 17108 11406
rect 17052 11327 17054 11340
rect 17106 11327 17108 11340
rect 17052 11302 17108 11327
rect 17388 10948 17444 11958
rect 17612 11844 17668 13020
rect 17836 12628 17892 13694
rect 17948 13748 18004 13758
rect 17948 13188 18004 13692
rect 18116 13748 18172 13758
rect 18116 13654 18172 13692
rect 18620 13748 18676 13758
rect 18620 13654 18676 13692
rect 18508 13636 18564 13646
rect 18508 13578 18564 13580
rect 18508 13526 18510 13578
rect 18562 13526 18564 13578
rect 18508 13514 18564 13526
rect 18732 13300 18788 14478
rect 18620 13244 18788 13300
rect 18956 13748 19012 13758
rect 19068 13748 19124 16604
rect 19180 15876 19236 16716
rect 19180 15810 19236 15820
rect 19292 15316 19348 17724
rect 19404 15540 19460 19014
rect 19516 16884 19572 19404
rect 19628 19234 19684 19628
rect 19628 19182 19630 19234
rect 19682 19182 19684 19234
rect 19628 17668 19684 19182
rect 20188 19460 20244 19852
rect 20524 19684 20580 19694
rect 20188 19236 20244 19404
rect 20412 19572 20468 19582
rect 20188 19142 20244 19180
rect 20300 19348 20356 19358
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 20076 18452 20132 18462
rect 19628 17108 19684 17612
rect 19964 18396 20076 18452
rect 19964 17444 20020 18396
rect 20076 18358 20132 18396
rect 20076 17780 20132 17790
rect 20076 17666 20132 17724
rect 20076 17614 20078 17666
rect 20130 17614 20132 17666
rect 20076 17602 20132 17614
rect 20300 17668 20356 19292
rect 20412 18564 20468 19516
rect 20524 19458 20580 19628
rect 20524 19406 20526 19458
rect 20578 19406 20580 19458
rect 20524 19394 20580 19406
rect 20636 18788 20692 20022
rect 20748 19908 20804 20188
rect 20748 19842 20804 19852
rect 20412 18450 20468 18508
rect 20412 18398 20414 18450
rect 20466 18398 20468 18450
rect 20412 18386 20468 18398
rect 20524 18732 20692 18788
rect 20524 17778 20580 18732
rect 20860 18676 20916 22876
rect 21196 22370 21252 23100
rect 21196 22318 21198 22370
rect 21250 22318 21252 22370
rect 21196 22306 21252 22318
rect 21308 22148 21364 23650
rect 21532 23156 21588 23166
rect 21532 23062 21588 23100
rect 21308 22082 21364 22092
rect 21532 22596 21588 22606
rect 21532 22036 21588 22540
rect 21532 21970 21588 21980
rect 21700 22148 21756 22158
rect 21700 21698 21756 22092
rect 21868 21812 21924 23846
rect 22092 23042 22148 24668
rect 22092 22990 22094 23042
rect 22146 22990 22148 23042
rect 22092 22978 22148 22990
rect 22204 22820 22260 24780
rect 22316 24724 22372 24734
rect 22316 24630 22372 24668
rect 22428 24062 22484 25340
rect 22652 24948 22708 24958
rect 22652 24854 22708 24892
rect 23324 24500 23380 24510
rect 23436 24500 23492 25788
rect 23660 24948 23716 26460
rect 23324 24498 23492 24500
rect 23324 24446 23326 24498
rect 23378 24446 23492 24498
rect 23324 24444 23492 24446
rect 23548 24892 23716 24948
rect 23772 26290 23828 26302
rect 23772 26238 23774 26290
rect 23826 26238 23828 26290
rect 23772 24948 23828 26238
rect 23884 25508 23940 26852
rect 23996 26292 24052 26302
rect 24332 26292 24388 26302
rect 23996 26290 24388 26292
rect 23996 26238 23998 26290
rect 24050 26238 24334 26290
rect 24386 26238 24388 26290
rect 23996 26236 24388 26238
rect 23996 26226 24052 26236
rect 23884 25442 23940 25452
rect 24108 26068 24164 26078
rect 23324 24388 23380 24444
rect 22372 24050 22484 24062
rect 22372 23998 22374 24050
rect 22426 23998 22484 24050
rect 22372 23996 22484 23998
rect 22988 24332 23380 24388
rect 22372 23986 22428 23996
rect 22876 23940 22932 23950
rect 22876 23846 22932 23884
rect 22876 23604 22932 23614
rect 22466 23191 22522 23203
rect 22466 23156 22468 23191
rect 22204 22754 22260 22764
rect 22428 23139 22468 23156
rect 22520 23139 22522 23191
rect 22428 23100 22522 23139
rect 22652 23154 22708 23166
rect 22652 23102 22654 23154
rect 22706 23102 22708 23154
rect 22092 22596 22148 22606
rect 22428 22596 22484 23100
rect 22092 22594 22484 22596
rect 22092 22542 22094 22594
rect 22146 22542 22484 22594
rect 22092 22540 22484 22542
rect 22540 22932 22596 22942
rect 22092 22530 22148 22540
rect 22540 22382 22596 22876
rect 22652 22708 22708 23102
rect 22764 23154 22820 23166
rect 22764 23102 22766 23154
rect 22818 23102 22820 23154
rect 22764 22820 22820 23102
rect 22764 22754 22820 22764
rect 22652 22642 22708 22652
rect 22486 22370 22596 22382
rect 22486 22318 22488 22370
rect 22540 22318 22596 22370
rect 22486 22316 22596 22318
rect 22652 22370 22708 22382
rect 22652 22318 22654 22370
rect 22706 22318 22708 22370
rect 22486 22306 22542 22316
rect 22652 22148 22708 22318
rect 22764 22370 22820 22382
rect 22764 22318 22766 22370
rect 22818 22318 22820 22370
rect 22764 22260 22820 22318
rect 22764 22194 22820 22204
rect 22652 22082 22708 22092
rect 21868 21746 21924 21756
rect 21700 21646 21702 21698
rect 21754 21646 21756 21698
rect 21700 21634 21756 21646
rect 21980 21614 22036 21626
rect 21420 21588 21476 21598
rect 21084 21362 21140 21374
rect 21084 21310 21086 21362
rect 21138 21310 21140 21362
rect 21084 20580 21140 21310
rect 21420 20804 21476 21532
rect 21980 21588 21982 21614
rect 22034 21588 22036 21614
rect 22148 21621 22204 21633
rect 22148 21588 22150 21621
rect 21980 21522 22036 21532
rect 22092 21569 22150 21588
rect 22202 21569 22204 21621
rect 22092 21532 22204 21569
rect 22428 21614 22484 21626
rect 22428 21562 22430 21614
rect 22482 21562 22484 21614
rect 21420 20738 21476 20748
rect 21756 20746 21812 20758
rect 21756 20694 21758 20746
rect 21810 20694 21812 20746
rect 22092 20746 22148 21532
rect 22428 20916 22484 21562
rect 22428 20850 22484 20860
rect 22540 21621 22596 21633
rect 22540 21569 22542 21621
rect 22594 21569 22596 21621
rect 21756 20580 21812 20694
rect 21084 20524 21812 20580
rect 21644 20018 21700 20030
rect 21644 19966 21646 20018
rect 21698 19966 21700 20018
rect 21644 19908 21700 19966
rect 21644 19842 21700 19852
rect 21364 19460 21420 19470
rect 21196 19458 21420 19460
rect 21196 19406 21366 19458
rect 21418 19406 21420 19458
rect 21196 19404 21420 19406
rect 20524 17726 20526 17778
rect 20578 17726 20580 17778
rect 20524 17714 20580 17726
rect 20636 18620 20916 18676
rect 21028 19236 21084 19246
rect 21028 18674 21084 19180
rect 21028 18622 21030 18674
rect 21082 18622 21084 18674
rect 20300 17575 20302 17612
rect 20354 17575 20356 17612
rect 19964 17378 20020 17388
rect 20188 17556 20244 17566
rect 20300 17563 20356 17575
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20188 17220 20244 17500
rect 20636 17444 20692 18620
rect 21028 18610 21084 18622
rect 21196 18452 21252 19404
rect 21364 19394 21420 19404
rect 21532 19236 21588 19246
rect 21532 19142 21588 19180
rect 21532 18506 21644 18564
rect 21196 18386 21252 18396
rect 21308 18450 21364 18462
rect 21308 18398 21310 18450
rect 21362 18398 21364 18450
rect 21308 17892 21364 18398
rect 21420 18452 21476 18462
rect 21420 18338 21476 18396
rect 21420 18286 21422 18338
rect 21474 18286 21476 18338
rect 21420 18274 21476 18286
rect 21532 18454 21590 18506
rect 21642 18454 21644 18506
rect 21532 18442 21644 18454
rect 21084 17836 21364 17892
rect 20748 17668 20804 17678
rect 21084 17668 21140 17836
rect 21532 17780 21588 18442
rect 21756 18116 21812 20524
rect 21868 20692 21924 20702
rect 21868 20130 21924 20636
rect 21868 20078 21870 20130
rect 21922 20078 21924 20130
rect 21868 20066 21924 20078
rect 22092 20694 22094 20746
rect 22146 20694 22148 20746
rect 22092 19908 22148 20694
rect 21868 19852 22148 19908
rect 22540 20244 22596 21569
rect 22540 20074 22596 20188
rect 22540 20022 22542 20074
rect 22594 20022 22596 20074
rect 21868 18452 21924 19852
rect 22092 19684 22148 19694
rect 22092 18788 22148 19628
rect 22540 19684 22596 20022
rect 22540 19618 22596 19628
rect 22764 20018 22820 20030
rect 22764 19966 22766 20018
rect 22818 19966 22820 20018
rect 22260 19572 22316 19582
rect 22260 19346 22316 19516
rect 22764 19358 22820 19966
rect 22260 19294 22262 19346
rect 22314 19294 22316 19346
rect 22260 19282 22316 19294
rect 22708 19348 22820 19358
rect 22764 19292 22820 19348
rect 22708 19254 22764 19292
rect 22764 19012 22820 19022
rect 22092 18732 22260 18788
rect 21868 18386 21924 18396
rect 21980 18450 22036 18462
rect 21980 18398 21982 18450
rect 22034 18398 22036 18450
rect 21980 18340 22036 18398
rect 21980 18274 22036 18284
rect 22092 18452 22148 18462
rect 21868 18116 21924 18126
rect 21756 18060 21868 18116
rect 20748 17666 21140 17668
rect 20748 17614 20750 17666
rect 20802 17614 21140 17666
rect 20748 17612 21140 17614
rect 21196 17724 21588 17780
rect 21196 17668 21252 17724
rect 20748 17602 20804 17612
rect 19628 17042 19684 17052
rect 20188 16938 20244 17164
rect 19684 16884 19740 16894
rect 19516 16882 19740 16884
rect 19516 16830 19686 16882
rect 19738 16830 19740 16882
rect 20188 16886 20190 16938
rect 20242 16886 20244 16938
rect 20188 16874 20244 16886
rect 20300 17388 20692 17444
rect 19516 16828 19740 16830
rect 19684 16818 19740 16828
rect 19404 15474 19460 15484
rect 19516 16548 19572 16558
rect 19292 15260 19460 15316
rect 19404 15148 19460 15260
rect 19516 15314 19572 16492
rect 20300 16324 20356 17388
rect 20412 16884 20468 16894
rect 20412 16882 20580 16884
rect 20412 16830 20414 16882
rect 20466 16830 20580 16882
rect 20412 16828 20580 16830
rect 20412 16818 20468 16828
rect 20524 16324 20580 16828
rect 20804 16826 20860 16838
rect 20636 16770 20692 16782
rect 20636 16718 20638 16770
rect 20690 16718 20692 16770
rect 20636 16548 20692 16718
rect 20636 16482 20692 16492
rect 20804 16774 20806 16826
rect 20858 16774 20860 16826
rect 20524 16268 20692 16324
rect 20300 16258 20356 16268
rect 19740 16100 19796 16110
rect 19740 16018 19742 16044
rect 19794 16018 19796 16044
rect 19740 15988 19796 16018
rect 19516 15262 19518 15314
rect 19570 15262 19572 15314
rect 19516 15250 19572 15262
rect 19628 15932 19796 15988
rect 20300 16098 20356 16110
rect 20300 16046 20302 16098
rect 20354 16046 20356 16098
rect 20300 15988 20356 16046
rect 19404 15092 19572 15148
rect 19348 14532 19404 14542
rect 19348 14308 19404 14476
rect 19516 14530 19572 15092
rect 19516 14478 19518 14530
rect 19570 14478 19572 14530
rect 19516 14466 19572 14478
rect 19628 14532 19684 15932
rect 20300 15922 20356 15932
rect 20468 15876 20524 15886
rect 20468 15782 20524 15820
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19740 15540 19796 15550
rect 19740 14980 19796 15484
rect 20636 14980 20692 16268
rect 20804 16212 20860 16774
rect 20972 16772 21028 17612
rect 21196 17574 21252 17612
rect 21756 17666 21812 17678
rect 21756 17614 21758 17666
rect 21810 17614 21812 17666
rect 21364 17556 21420 17566
rect 21364 17498 21420 17500
rect 21364 17446 21366 17498
rect 21418 17446 21420 17498
rect 21364 17434 21420 17446
rect 21196 17108 21252 17118
rect 21196 17014 21252 17052
rect 21756 17108 21812 17614
rect 21756 17042 21812 17052
rect 21532 16884 21588 16894
rect 20972 16706 21028 16716
rect 21308 16882 21588 16884
rect 21308 16830 21534 16882
rect 21586 16830 21588 16882
rect 21308 16828 21588 16830
rect 20804 16156 21028 16212
rect 20972 15428 21028 16156
rect 21196 16100 21252 16110
rect 21308 16100 21364 16828
rect 21532 16818 21588 16828
rect 21756 16882 21812 16894
rect 21756 16830 21758 16882
rect 21810 16830 21812 16882
rect 21196 16098 21364 16100
rect 21196 16046 21198 16098
rect 21250 16046 21364 16098
rect 21196 16044 21364 16046
rect 21756 16772 21812 16830
rect 21196 15428 21252 16044
rect 21532 15988 21588 15998
rect 21364 15874 21420 15886
rect 21364 15822 21366 15874
rect 21418 15822 21420 15874
rect 21364 15652 21420 15822
rect 21364 15586 21420 15596
rect 21420 15428 21476 15438
rect 21196 15426 21476 15428
rect 21196 15374 21422 15426
rect 21474 15374 21476 15426
rect 21196 15372 21476 15374
rect 20972 15362 21028 15372
rect 21420 15362 21476 15372
rect 19740 14924 20244 14980
rect 19628 14466 19684 14476
rect 20188 14530 20244 14924
rect 20636 14914 20692 14924
rect 21196 14980 21252 14990
rect 20188 14478 20190 14530
rect 20242 14478 20244 14530
rect 19852 14308 19908 14318
rect 19348 14242 19404 14252
rect 19516 14306 19908 14308
rect 19516 14254 19854 14306
rect 19906 14254 19908 14306
rect 19516 14252 19908 14254
rect 18956 13746 19124 13748
rect 18956 13694 18958 13746
rect 19010 13694 19124 13746
rect 18956 13692 19124 13694
rect 19404 14084 19460 14094
rect 17948 13132 18228 13188
rect 18172 13074 18228 13132
rect 18172 13022 18174 13074
rect 18226 13022 18228 13074
rect 18172 13010 18228 13022
rect 18620 12628 18676 13244
rect 18788 13076 18844 13086
rect 18788 12982 18844 13020
rect 17836 12572 18228 12628
rect 18620 12572 18788 12628
rect 18060 12404 18116 12414
rect 17724 12348 18060 12404
rect 17724 12178 17780 12348
rect 17724 12126 17726 12178
rect 17778 12126 17780 12178
rect 17724 12114 17780 12126
rect 17836 12180 17892 12190
rect 17612 11508 17668 11788
rect 16884 10892 17444 10948
rect 17500 11452 17668 11508
rect 17724 11508 17780 11518
rect 16884 10666 16940 10892
rect 17500 10846 17556 11452
rect 17612 11282 17668 11294
rect 17612 11230 17614 11282
rect 17666 11230 17668 11282
rect 17612 11172 17668 11230
rect 17612 11106 17668 11116
rect 17500 10834 17612 10846
rect 17500 10782 17558 10834
rect 17610 10782 17612 10834
rect 17500 10780 17612 10782
rect 17556 10770 17612 10780
rect 16884 10614 16886 10666
rect 16938 10614 16940 10666
rect 16884 10602 16940 10614
rect 17500 10612 17556 10622
rect 16492 10518 16548 10556
rect 16716 10500 16772 10510
rect 16604 10498 16772 10500
rect 16604 10446 16718 10498
rect 16770 10446 16772 10498
rect 16604 10444 16772 10446
rect 16604 10164 16660 10444
rect 16716 10434 16772 10444
rect 16380 10108 16660 10164
rect 16380 9938 16436 10108
rect 16380 9886 16382 9938
rect 16434 9886 16436 9938
rect 16380 9874 16436 9886
rect 16268 9090 16324 9100
rect 16380 9604 16436 9614
rect 16380 8942 16436 9548
rect 16772 9156 16828 9166
rect 16772 9062 16828 9100
rect 16324 8930 16436 8942
rect 16324 8878 16326 8930
rect 16378 8878 16436 8930
rect 16324 8876 16436 8878
rect 16324 8866 16380 8876
rect 17500 8596 17556 10556
rect 17724 10500 17780 11452
rect 17836 10734 17892 12124
rect 17836 10722 17948 10734
rect 17836 10670 17894 10722
rect 17946 10670 17948 10722
rect 17836 10668 17948 10670
rect 17892 10658 17948 10668
rect 17724 10444 17892 10500
rect 17668 9492 17724 9502
rect 17668 9266 17724 9436
rect 17668 9214 17670 9266
rect 17722 9214 17724 9266
rect 17668 9202 17724 9214
rect 17836 8708 17892 10444
rect 18060 9278 18116 12348
rect 18172 12068 18228 12572
rect 18564 12404 18620 12414
rect 18564 12310 18620 12348
rect 18172 10610 18228 12012
rect 18732 11732 18788 12572
rect 18956 12404 19012 13692
rect 19404 13578 19460 14028
rect 19516 13748 19572 14252
rect 19852 14242 19908 14252
rect 19836 14140 20100 14150
rect 19516 13654 19572 13692
rect 19628 14084 19684 14094
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19404 13526 19406 13578
rect 19458 13526 19460 13578
rect 19404 13524 19460 13526
rect 19292 13468 19460 13524
rect 19292 12404 19348 13468
rect 19460 13076 19516 13086
rect 19628 13076 19684 14028
rect 19852 13860 19908 13870
rect 19852 13746 19908 13804
rect 19852 13694 19854 13746
rect 19906 13694 19908 13746
rect 19852 13186 19908 13694
rect 19852 13134 19854 13186
rect 19906 13134 19908 13186
rect 19852 13122 19908 13134
rect 19460 13074 19684 13076
rect 19460 13022 19462 13074
rect 19514 13022 19684 13074
rect 19460 13020 19684 13022
rect 19460 13010 19516 13020
rect 20188 12962 20244 14478
rect 20412 14420 20468 14430
rect 20188 12910 20190 12962
rect 20242 12910 20244 12962
rect 20188 12898 20244 12910
rect 20300 13748 20356 13758
rect 20300 12962 20356 13692
rect 20412 13524 20468 14364
rect 20524 14308 20580 14318
rect 20524 14306 20804 14308
rect 20524 14254 20526 14306
rect 20578 14254 20804 14306
rect 20524 14252 20804 14254
rect 20524 14242 20580 14252
rect 20580 13524 20636 13534
rect 20412 13522 20636 13524
rect 20412 13470 20582 13522
rect 20634 13470 20636 13522
rect 20412 13468 20636 13470
rect 20580 13458 20636 13468
rect 20748 13076 20804 14252
rect 20972 14196 21028 14206
rect 21196 14196 21252 14924
rect 20860 13748 20916 13758
rect 20860 13654 20916 13692
rect 20972 13746 21028 14140
rect 20972 13694 20974 13746
rect 21026 13694 21028 13746
rect 21140 14140 21252 14196
rect 21420 14306 21476 14318
rect 21420 14254 21422 14306
rect 21474 14254 21476 14306
rect 21420 14196 21476 14254
rect 21140 13802 21196 14140
rect 21420 14130 21476 14140
rect 21140 13750 21142 13802
rect 21194 13750 21196 13802
rect 21140 13738 21196 13750
rect 21308 13746 21364 13758
rect 20972 13412 21028 13694
rect 20972 13346 21028 13356
rect 21308 13694 21310 13746
rect 21362 13694 21364 13746
rect 21308 13636 21364 13694
rect 21532 13636 21588 15932
rect 21756 15652 21812 16716
rect 21868 16884 21924 18060
rect 21868 16100 21924 16828
rect 21980 17778 22036 17790
rect 21980 17726 21982 17778
rect 22034 17726 22036 17778
rect 21980 16436 22036 17726
rect 22092 17610 22148 18396
rect 22092 17558 22094 17610
rect 22146 17558 22148 17610
rect 22092 17556 22148 17558
rect 22092 17490 22148 17500
rect 22204 16938 22260 18732
rect 22428 18564 22484 18574
rect 22204 16886 22206 16938
rect 22258 16886 22260 16938
rect 22204 16874 22260 16886
rect 22316 18340 22372 18350
rect 22316 16884 22372 18284
rect 22428 17666 22484 18508
rect 22652 18488 22708 18500
rect 22652 18436 22654 18488
rect 22706 18436 22708 18488
rect 22652 18116 22708 18436
rect 22652 18050 22708 18060
rect 22764 18004 22820 18956
rect 22764 17938 22820 17948
rect 22428 17614 22430 17666
rect 22482 17614 22484 17666
rect 22428 17602 22484 17614
rect 22764 17780 22820 17790
rect 22764 17666 22820 17724
rect 22764 17614 22766 17666
rect 22818 17614 22820 17666
rect 22764 17602 22820 17614
rect 22316 16818 22372 16828
rect 22428 17332 22484 17342
rect 22428 16882 22484 17276
rect 22428 16830 22430 16882
rect 22482 16830 22484 16882
rect 22428 16818 22484 16830
rect 22540 17050 22596 17062
rect 22540 16998 22542 17050
rect 22594 16998 22596 17050
rect 22540 16772 22596 16998
rect 22540 16706 22596 16716
rect 21980 16380 22820 16436
rect 22204 16268 22652 16324
rect 22036 16212 22092 16222
rect 22036 16118 22092 16156
rect 21868 16044 21980 16100
rect 21924 15988 21980 16044
rect 21924 15932 22036 15988
rect 21868 15652 21924 15662
rect 21756 15596 21868 15652
rect 21868 15314 21924 15596
rect 21868 15262 21870 15314
rect 21922 15262 21924 15314
rect 21868 15250 21924 15262
rect 21980 15314 22036 15932
rect 22204 15540 22260 16268
rect 22316 16098 22372 16110
rect 22316 16046 22318 16098
rect 22370 16046 22372 16098
rect 22316 15652 22372 16046
rect 22428 16100 22484 16110
rect 22428 16006 22484 16044
rect 22596 16042 22652 16268
rect 22764 16100 22820 16380
rect 22876 16324 22932 23548
rect 22988 22260 23044 24332
rect 23548 23604 23604 24892
rect 23772 24882 23828 24892
rect 24108 24750 24164 26012
rect 23660 24722 23716 24734
rect 23660 24670 23662 24722
rect 23714 24670 23716 24722
rect 23660 24164 23716 24670
rect 24108 24698 24110 24750
rect 24162 24698 24164 24750
rect 24108 24500 24164 24698
rect 24108 24434 24164 24444
rect 24220 25394 24276 25406
rect 24220 25342 24222 25394
rect 24274 25342 24276 25394
rect 24220 24276 24276 25342
rect 24332 25396 24388 26236
rect 24444 26122 24500 28252
rect 24556 27198 24612 28924
rect 24780 28420 24836 31276
rect 24892 29988 24948 31388
rect 24892 29922 24948 29932
rect 25004 29876 25060 32172
rect 25116 32004 25172 33292
rect 25228 33346 25284 33358
rect 25228 33294 25230 33346
rect 25282 33294 25284 33346
rect 25228 32676 25284 33294
rect 25228 32610 25284 32620
rect 25340 32562 25396 33404
rect 25452 33348 25508 33358
rect 25452 33266 25454 33292
rect 25506 33266 25508 33292
rect 25452 33254 25508 33266
rect 25340 32510 25342 32562
rect 25394 32510 25396 32562
rect 25340 32498 25396 32510
rect 25116 31938 25172 31948
rect 25116 31778 25172 31790
rect 25116 31726 25118 31778
rect 25170 31726 25172 31778
rect 25116 31332 25172 31726
rect 25284 31556 25340 31566
rect 25284 31462 25340 31500
rect 25116 31266 25172 31276
rect 25564 31220 25620 36372
rect 25676 36260 25732 37100
rect 25956 36820 26012 37158
rect 26124 36932 26180 37244
rect 26124 36866 26180 36876
rect 26348 36932 26404 37998
rect 26572 38050 26628 38062
rect 26796 38052 26852 38062
rect 26572 37998 26574 38050
rect 26626 37998 26628 38050
rect 26572 37716 26628 37998
rect 26572 37650 26628 37660
rect 26684 38050 26852 38052
rect 26684 37998 26798 38050
rect 26850 37998 26852 38050
rect 26684 37996 26852 37998
rect 26460 37296 26516 37308
rect 26460 37244 26462 37296
rect 26514 37244 26516 37296
rect 26460 37156 26516 37244
rect 26460 37090 26516 37100
rect 26348 36866 26404 36876
rect 25788 36764 26012 36820
rect 25788 36596 25844 36764
rect 25788 36484 25844 36540
rect 26012 36484 26068 36494
rect 25788 36482 26068 36484
rect 25788 36430 26014 36482
rect 26066 36430 26068 36482
rect 25788 36428 26068 36430
rect 26012 36418 26068 36428
rect 26124 36484 26180 36494
rect 25676 36204 26068 36260
rect 25676 35728 25732 35740
rect 25676 35676 25678 35728
rect 25730 35676 25732 35728
rect 25676 35252 25732 35676
rect 25844 35642 25900 35654
rect 25844 35590 25846 35642
rect 25898 35590 25900 35642
rect 25844 35588 25900 35590
rect 25844 35522 25900 35532
rect 25676 35186 25732 35196
rect 26012 35140 26068 36204
rect 26124 35700 26180 36428
rect 26124 35606 26180 35644
rect 26236 35924 26292 35934
rect 26236 35364 26292 35868
rect 26684 35810 26740 37996
rect 26796 37986 26852 37996
rect 26908 37044 26964 40012
rect 27112 39562 27168 39574
rect 27112 39510 27114 39562
rect 27166 39510 27168 39562
rect 27112 39172 27168 39510
rect 27112 39106 27168 39116
rect 27132 38834 27188 38846
rect 27132 38782 27134 38834
rect 27186 38782 27188 38834
rect 27132 38724 27188 38782
rect 27244 38836 27300 41692
rect 27448 41692 27524 41748
rect 27448 41130 27504 41692
rect 27636 41524 27692 41974
rect 27804 42000 27860 42012
rect 27804 41948 27806 42000
rect 27858 41948 27860 42000
rect 27804 41860 27860 41948
rect 27804 41794 27860 41804
rect 28140 42000 28196 42012
rect 28140 41948 28142 42000
rect 28194 41948 28196 42000
rect 27636 41458 27692 41468
rect 27448 41078 27450 41130
rect 27502 41078 27504 41130
rect 27448 40740 27504 41078
rect 27448 40674 27504 40684
rect 27692 41074 27748 41086
rect 27692 41022 27694 41074
rect 27746 41022 27748 41074
rect 27524 40404 27580 40414
rect 27692 40404 27748 41022
rect 28140 40964 28196 41948
rect 28140 40740 28196 40908
rect 28364 40740 28420 44044
rect 28476 43577 28532 43589
rect 28476 43525 28478 43577
rect 28530 43525 28532 43577
rect 28476 43316 28532 43525
rect 29260 43540 29316 44044
rect 30156 43876 30212 46956
rect 30268 46116 30324 49200
rect 30268 46050 30324 46060
rect 30380 46060 30660 46116
rect 30268 45892 30324 45902
rect 30268 45798 30324 45836
rect 29260 43474 29316 43484
rect 29820 43820 30212 43876
rect 29652 43428 29708 43438
rect 29652 43334 29708 43372
rect 28476 43250 28532 43260
rect 29036 43314 29092 43326
rect 29036 43262 29038 43314
rect 29090 43262 29092 43314
rect 28476 42980 28532 42990
rect 28476 42886 28532 42924
rect 29036 42644 29092 43262
rect 29820 43204 29876 43820
rect 29932 43652 29988 43662
rect 29932 43538 29988 43596
rect 29932 43486 29934 43538
rect 29986 43486 29988 43538
rect 29932 43474 29988 43486
rect 30156 43540 30212 43550
rect 30156 43446 30212 43484
rect 30380 43316 30436 46060
rect 30492 45890 30548 45902
rect 30492 45838 30494 45890
rect 30546 45838 30548 45890
rect 30492 45220 30548 45838
rect 30604 45890 30660 46060
rect 30604 45838 30606 45890
rect 30658 45838 30660 45890
rect 30604 45826 30660 45838
rect 30940 45892 30996 45902
rect 30940 45798 30996 45836
rect 31444 45780 31500 45790
rect 31444 45722 31500 45724
rect 31444 45670 31446 45722
rect 31498 45670 31500 45722
rect 31444 45658 31500 45670
rect 31836 45332 31892 49200
rect 33180 46116 33236 46126
rect 33180 46022 33236 46060
rect 33404 46116 33460 49200
rect 34972 46340 35028 49200
rect 33404 46050 33460 46060
rect 34860 46284 35028 46340
rect 35196 46284 35460 46294
rect 32172 45892 32228 45902
rect 32172 45810 32174 45836
rect 32226 45810 32228 45836
rect 32172 45798 32228 45810
rect 33628 45780 33684 45790
rect 31836 45276 32340 45332
rect 30492 45164 30660 45220
rect 30492 44994 30548 45006
rect 30492 44942 30494 44994
rect 30546 44942 30548 44994
rect 30492 44548 30548 44942
rect 30492 44482 30548 44492
rect 30492 44210 30548 44222
rect 30492 44158 30494 44210
rect 30546 44158 30548 44210
rect 30492 43764 30548 44158
rect 30492 43698 30548 43708
rect 30380 43250 30436 43260
rect 30492 43568 30548 43580
rect 30492 43516 30494 43568
rect 30546 43516 30548 43568
rect 29036 42578 29092 42588
rect 29708 43148 29876 43204
rect 30492 43204 30548 43516
rect 29708 42754 29764 43148
rect 30492 43138 30548 43148
rect 29708 42702 29710 42754
rect 29762 42702 29764 42754
rect 29372 42532 29428 42542
rect 29372 42438 29428 42476
rect 28588 42308 28644 42318
rect 28588 42082 28644 42252
rect 28588 42030 28590 42082
rect 28642 42030 28644 42082
rect 28588 42018 28644 42030
rect 28700 42196 28756 42206
rect 28700 41310 28756 42140
rect 28644 41298 28756 41310
rect 28644 41246 28646 41298
rect 28698 41246 28756 41298
rect 28644 41244 28756 41246
rect 28812 41972 28868 41982
rect 28644 41234 28700 41244
rect 28680 40740 28736 40750
rect 28364 40684 28532 40740
rect 28140 40674 28196 40684
rect 27804 40404 27860 40414
rect 27692 40402 27860 40404
rect 27692 40350 27806 40402
rect 27858 40350 27860 40402
rect 27692 40348 27860 40350
rect 27524 40310 27580 40348
rect 27804 40338 27860 40348
rect 27468 40068 27524 40078
rect 27356 39620 27412 39630
rect 27356 39526 27412 39564
rect 27244 38770 27300 38780
rect 27132 38658 27188 38668
rect 27244 38668 27300 38678
rect 27468 38668 27524 40012
rect 28476 39956 28532 40684
rect 28680 40458 28736 40684
rect 28680 40406 28682 40458
rect 28734 40406 28736 40458
rect 28680 40394 28736 40406
rect 28812 40628 28868 41916
rect 29148 41970 29204 41982
rect 29148 41918 29150 41970
rect 29202 41918 29204 41970
rect 27804 39900 28532 39956
rect 27804 39070 27860 39900
rect 28532 39732 28588 39742
rect 28812 39732 28868 40572
rect 29036 41186 29092 41198
rect 29036 41134 29038 41186
rect 29090 41134 29092 41186
rect 28924 40516 28980 40526
rect 28924 40422 28980 40460
rect 29036 40404 29092 41134
rect 29036 39844 29092 40348
rect 29148 40068 29204 41918
rect 29484 41972 29540 41982
rect 29484 41878 29540 41916
rect 29596 41802 29652 41814
rect 29484 41748 29540 41758
rect 29372 40964 29428 40974
rect 29372 40870 29428 40908
rect 29148 40002 29204 40012
rect 29036 39788 29428 39844
rect 28532 39730 28868 39732
rect 28532 39678 28534 39730
rect 28586 39678 28868 39730
rect 28532 39676 28868 39678
rect 28532 39666 28588 39676
rect 28140 39618 28196 39630
rect 28140 39566 28142 39618
rect 28194 39566 28196 39618
rect 28140 39508 28196 39566
rect 27748 39058 27860 39070
rect 27748 39006 27750 39058
rect 27802 39006 27860 39058
rect 27748 39004 27860 39006
rect 28028 39452 28140 39508
rect 27748 38994 27804 39004
rect 28028 38834 28084 39452
rect 28140 39442 28196 39452
rect 28252 39618 28308 39630
rect 28252 39566 28254 39618
rect 28306 39566 28308 39618
rect 28252 39396 28308 39566
rect 29036 39620 29092 39630
rect 29036 39526 29092 39564
rect 29204 39508 29260 39518
rect 29204 39450 29260 39452
rect 28252 39330 28308 39340
rect 28904 39396 28960 39406
rect 29204 39398 29206 39450
rect 29258 39398 29260 39450
rect 29204 39386 29260 39398
rect 29372 39396 29428 39788
rect 28028 38782 28030 38834
rect 28082 38782 28084 38834
rect 28904 38890 28960 39340
rect 29372 39330 29428 39340
rect 28904 38838 28906 38890
rect 28958 38838 28960 38890
rect 28904 38826 28960 38838
rect 29148 38836 29204 38846
rect 28028 38770 28084 38782
rect 29148 38742 29204 38780
rect 27244 38666 27524 38668
rect 27244 38614 27246 38666
rect 27298 38614 27524 38666
rect 27244 38612 27524 38614
rect 28700 38724 28756 38734
rect 27244 38602 27300 38612
rect 28700 38388 28756 38668
rect 29484 38668 29540 41692
rect 29596 41750 29598 41802
rect 29650 41750 29652 41802
rect 29596 41188 29652 41750
rect 29708 41524 29764 42702
rect 29932 42756 29988 42766
rect 29932 42662 29988 42700
rect 30156 42196 30212 42206
rect 30156 41970 30212 42140
rect 30156 41918 30158 41970
rect 30210 41918 30212 41970
rect 30156 41906 30212 41918
rect 30492 41748 30548 41758
rect 30492 41654 30548 41692
rect 30604 41524 30660 45164
rect 31612 44324 31668 44334
rect 31612 44322 31780 44324
rect 30735 44266 30791 44278
rect 30735 44214 30737 44266
rect 30789 44214 30791 44266
rect 31612 44270 31614 44322
rect 31666 44270 31780 44322
rect 31612 44268 31780 44270
rect 31612 44258 31668 44268
rect 30735 44212 30791 44214
rect 30735 44146 30791 44156
rect 30716 43652 30772 43662
rect 30716 43092 30772 43596
rect 30716 43026 30772 43036
rect 30828 43568 30884 43580
rect 30828 43516 30830 43568
rect 30882 43516 30884 43568
rect 30828 42980 30884 43516
rect 31276 43540 31332 43550
rect 30828 42914 30884 42924
rect 30996 43482 31052 43494
rect 30996 43430 30998 43482
rect 31050 43430 31052 43482
rect 31276 43446 31332 43484
rect 31612 43540 31668 43550
rect 30996 42868 31052 43430
rect 30940 42812 31052 42868
rect 30808 42698 30864 42710
rect 30808 42646 30810 42698
rect 30862 42646 30864 42698
rect 30808 42308 30864 42646
rect 30808 42242 30864 42252
rect 30940 42084 30996 42812
rect 31612 42754 31668 43484
rect 31612 42702 31614 42754
rect 31666 42702 31668 42754
rect 31612 42690 31668 42702
rect 31724 43538 31780 44268
rect 32284 44322 32340 45276
rect 32396 45276 33012 45332
rect 32396 45218 32452 45276
rect 32396 45166 32398 45218
rect 32450 45166 32452 45218
rect 32396 45154 32452 45166
rect 32284 44270 32286 44322
rect 32338 44270 32340 44322
rect 32284 44258 32340 44270
rect 32732 45108 32788 45118
rect 31724 43486 31726 43538
rect 31778 43486 31780 43538
rect 31052 42642 31108 42654
rect 31052 42590 31054 42642
rect 31106 42590 31108 42642
rect 31052 42308 31108 42590
rect 31724 42644 31780 43486
rect 31836 44212 31892 44222
rect 31836 43538 31892 44156
rect 31836 43486 31838 43538
rect 31890 43486 31892 43538
rect 31836 43474 31892 43486
rect 31982 43575 32038 43587
rect 31982 43540 31984 43575
rect 32036 43540 32038 43575
rect 31982 43316 32038 43484
rect 32396 43316 32452 43326
rect 31982 43260 32116 43316
rect 31948 43092 32004 43102
rect 31948 42739 32004 43036
rect 32060 42866 32116 43260
rect 32396 43222 32452 43260
rect 32452 42980 32508 42990
rect 32452 42886 32508 42924
rect 32060 42814 32062 42866
rect 32114 42814 32116 42866
rect 32060 42802 32116 42814
rect 31948 42687 31950 42739
rect 32002 42687 32004 42739
rect 31948 42675 32004 42687
rect 32172 42756 32228 42766
rect 31724 42578 31780 42588
rect 31052 42252 31872 42308
rect 29708 41458 29764 41468
rect 30492 41468 30660 41524
rect 30716 42028 30996 42084
rect 29596 41122 29652 41132
rect 29820 41188 29876 41198
rect 29820 41186 29988 41188
rect 29820 41134 29822 41186
rect 29874 41134 29988 41186
rect 29820 41132 29988 41134
rect 29820 41122 29876 41132
rect 29932 40516 29988 41132
rect 30492 40852 30548 41468
rect 30716 41412 30772 42028
rect 30940 41970 30996 42028
rect 30940 41918 30942 41970
rect 30994 41918 30996 41970
rect 31816 42026 31872 42252
rect 31816 41974 31818 42026
rect 31870 41974 31872 42026
rect 31816 41962 31872 41974
rect 32060 41972 32116 41982
rect 32172 41972 32228 42700
rect 32284 42754 32340 42766
rect 32284 42702 32286 42754
rect 32338 42702 32340 42754
rect 32284 42308 32340 42702
rect 32284 42242 32340 42252
rect 32620 42756 32676 42766
rect 32060 41970 32228 41972
rect 30940 41906 30996 41918
rect 32060 41918 32062 41970
rect 32114 41918 32228 41970
rect 32060 41916 32228 41918
rect 32060 41906 32116 41916
rect 30716 41356 30884 41412
rect 30696 41188 30752 41198
rect 30696 41094 30752 41132
rect 30380 40796 30548 40852
rect 29932 40450 29988 40460
rect 30156 40516 30212 40526
rect 30156 40458 30212 40460
rect 29764 40404 29820 40414
rect 30156 40406 30158 40458
rect 30210 40406 30212 40458
rect 30156 40394 30212 40406
rect 29764 40310 29820 40348
rect 29708 39618 29764 39630
rect 29708 39566 29710 39618
rect 29762 39566 29764 39618
rect 29708 38836 29764 39566
rect 29708 38770 29764 38780
rect 29932 39284 29988 39294
rect 29932 38834 29988 39228
rect 30380 38948 30436 40796
rect 30660 40516 30716 40526
rect 30828 40516 30884 41356
rect 30940 41188 30996 41198
rect 30940 41094 30996 41132
rect 31388 41186 31444 41198
rect 31388 41134 31390 41186
rect 31442 41134 31444 41186
rect 31052 40964 31108 40974
rect 30940 40516 30996 40526
rect 30828 40514 30996 40516
rect 30828 40462 30942 40514
rect 30994 40462 30996 40514
rect 30828 40460 30996 40462
rect 30660 40458 30716 40460
rect 30492 40432 30548 40444
rect 30492 40404 30494 40432
rect 30546 40404 30548 40432
rect 30660 40406 30662 40458
rect 30714 40406 30716 40458
rect 30940 40450 30996 40460
rect 30660 40394 30716 40406
rect 30492 40338 30548 40348
rect 30828 39620 30884 39630
rect 30584 39562 30640 39574
rect 30584 39510 30586 39562
rect 30638 39510 30640 39562
rect 30828 39526 30884 39564
rect 30584 39284 30640 39510
rect 30584 39218 30640 39228
rect 30716 39060 30772 39070
rect 30716 39002 30772 39004
rect 30716 38950 30718 39002
rect 30770 38950 30772 39002
rect 30716 38938 30772 38950
rect 30380 38882 30436 38892
rect 29932 38782 29934 38834
rect 29986 38782 29988 38834
rect 29932 38724 29988 38782
rect 30492 38836 30548 38874
rect 30492 38770 30548 38780
rect 28476 38332 28756 38388
rect 28812 38612 28868 38622
rect 29484 38612 29876 38668
rect 29932 38658 29988 38668
rect 30380 38724 30436 38734
rect 30380 38612 30548 38668
rect 28476 38274 28532 38332
rect 28476 38222 28478 38274
rect 28530 38222 28532 38274
rect 28476 38210 28532 38222
rect 28028 38052 28084 38062
rect 27524 37994 27580 38006
rect 27076 37940 27132 37950
rect 27076 37846 27132 37884
rect 27524 37942 27526 37994
rect 27578 37942 27580 37994
rect 27524 37604 27580 37942
rect 27244 37548 27580 37604
rect 27804 37994 27860 38006
rect 27804 37942 27806 37994
rect 27858 37942 27860 37994
rect 28028 37968 28030 37996
rect 28082 37968 28084 37996
rect 28028 37956 28084 37968
rect 27804 37604 27860 37942
rect 28476 37940 28532 37950
rect 27804 37548 27972 37604
rect 27244 37492 27300 37548
rect 27244 37266 27300 37436
rect 27244 37214 27246 37266
rect 27298 37214 27300 37266
rect 27244 37202 27300 37214
rect 27916 37156 27972 37548
rect 28364 37380 28420 37390
rect 28364 37286 28420 37324
rect 26908 36988 27076 37044
rect 27020 36932 27076 36988
rect 27020 36876 27300 36932
rect 26888 36820 26944 36830
rect 26888 36484 26944 36764
rect 27020 36708 27076 36718
rect 26888 36482 26964 36484
rect 26888 36430 26890 36482
rect 26942 36430 26964 36482
rect 26888 36418 26964 36430
rect 26908 35924 26964 36418
rect 26684 35758 26686 35810
rect 26738 35758 26740 35810
rect 26684 35746 26740 35758
rect 26796 35868 26964 35924
rect 27020 36372 27076 36652
rect 27132 36372 27188 36382
rect 27020 36370 27188 36372
rect 27020 36318 27134 36370
rect 27186 36318 27188 36370
rect 27020 36316 27188 36318
rect 26236 35298 26292 35308
rect 26516 35642 26572 35654
rect 26516 35590 26518 35642
rect 26570 35590 26572 35642
rect 26516 35252 26572 35590
rect 26796 35476 26852 35868
rect 26908 35700 26964 35710
rect 27020 35700 27076 36316
rect 27132 36306 27188 36316
rect 26908 35698 27076 35700
rect 26908 35646 26910 35698
rect 26962 35646 27076 35698
rect 26908 35644 27076 35646
rect 27132 35726 27188 35738
rect 27132 35700 27134 35726
rect 27186 35700 27188 35726
rect 26908 35634 26964 35644
rect 27132 35634 27188 35644
rect 26796 35420 27076 35476
rect 26908 35252 26964 35262
rect 26516 35196 26740 35252
rect 26516 35140 26572 35196
rect 26012 35084 26572 35140
rect 26068 34860 26124 34870
rect 25900 34858 26124 34860
rect 25676 34802 25732 34814
rect 25676 34750 25678 34802
rect 25730 34750 25732 34802
rect 25676 34692 25732 34750
rect 25676 34626 25732 34636
rect 25900 34806 26070 34858
rect 26122 34806 26124 34858
rect 25900 34804 26124 34806
rect 25676 34130 25732 34142
rect 25676 34078 25678 34130
rect 25730 34078 25732 34130
rect 25676 34020 25732 34078
rect 25676 33954 25732 33964
rect 25900 33962 25956 34804
rect 26068 34794 26124 34804
rect 26236 34804 26292 34814
rect 26236 34710 26292 34748
rect 26012 34132 26068 34142
rect 26516 34132 26572 34142
rect 26012 34130 26572 34132
rect 26012 34078 26014 34130
rect 26066 34078 26518 34130
rect 26570 34078 26572 34130
rect 26012 34076 26572 34078
rect 26012 34066 26068 34076
rect 26516 34066 26572 34076
rect 25900 33910 25902 33962
rect 25954 33910 25956 33962
rect 25900 33898 25956 33910
rect 26012 33796 26068 33806
rect 26012 32116 26068 33740
rect 26292 33124 26348 33134
rect 26684 33124 26740 35196
rect 26908 34970 26964 35196
rect 26908 34918 26910 34970
rect 26962 34918 26964 34970
rect 26796 34858 26852 34870
rect 26796 34806 26798 34858
rect 26850 34806 26852 34858
rect 26796 34692 26852 34806
rect 26796 34130 26852 34636
rect 26796 34078 26798 34130
rect 26850 34078 26852 34130
rect 26796 34066 26852 34078
rect 26908 34130 26964 34918
rect 26908 34078 26910 34130
rect 26962 34078 26964 34130
rect 26908 33908 26964 34078
rect 26908 33842 26964 33852
rect 27020 33796 27076 35420
rect 27244 35140 27300 36876
rect 27916 36820 27972 37100
rect 27804 36764 27972 36820
rect 28120 37266 28176 37278
rect 28120 37214 28122 37266
rect 28174 37214 28176 37266
rect 28120 36820 28176 37214
rect 27804 36596 27860 36764
rect 28120 36754 28176 36764
rect 28476 36706 28532 37884
rect 28476 36654 28478 36706
rect 28530 36654 28532 36706
rect 28476 36642 28532 36654
rect 27580 36540 27860 36596
rect 27916 36596 27972 36606
rect 27580 35364 27636 36540
rect 27692 36426 27748 36438
rect 27692 36374 27694 36426
rect 27746 36374 27748 36426
rect 27692 35476 27748 36374
rect 27916 36426 27972 36540
rect 27916 36374 27918 36426
rect 27970 36374 27972 36426
rect 27916 36260 27972 36374
rect 27804 36204 27972 36260
rect 28196 36426 28252 36438
rect 28196 36374 28198 36426
rect 28250 36374 28252 36426
rect 27804 35812 27860 36204
rect 28196 36036 28252 36374
rect 27804 35746 27860 35756
rect 27916 35980 28252 36036
rect 27916 35924 27972 35980
rect 28812 35924 28868 38556
rect 29148 38050 29204 38062
rect 29148 37998 29150 38050
rect 29202 37998 29204 38050
rect 29148 37380 29204 37998
rect 29820 37940 29876 38612
rect 30380 38500 30436 38510
rect 30024 38052 30080 38062
rect 30024 37958 30080 37996
rect 30268 38052 30324 38062
rect 30268 37958 30324 37996
rect 29820 37884 29932 37940
rect 29876 37828 29932 37884
rect 29876 37772 29988 37828
rect 29148 37314 29204 37324
rect 29764 37716 29820 37726
rect 28980 37156 29036 37166
rect 27916 35698 27972 35868
rect 27916 35646 27918 35698
rect 27970 35646 27972 35698
rect 27916 35634 27972 35646
rect 28588 35868 28868 35924
rect 28924 37154 29036 37156
rect 28924 37102 28982 37154
rect 29034 37102 29036 37154
rect 28924 37090 29036 37102
rect 29764 37156 29820 37660
rect 27692 35410 27748 35420
rect 28588 35364 28644 35868
rect 28792 35698 28848 35710
rect 28792 35646 28794 35698
rect 28846 35646 28848 35698
rect 28792 35476 28848 35646
rect 28792 35410 28848 35420
rect 28924 35588 28980 37090
rect 29764 37062 29820 37100
rect 29260 36484 29316 36494
rect 29036 36482 29316 36484
rect 29036 36430 29262 36482
rect 29314 36430 29316 36482
rect 29036 36428 29316 36430
rect 29036 35810 29092 36428
rect 29260 36418 29316 36428
rect 29932 36260 29988 37772
rect 30380 37492 30436 38444
rect 30212 37268 30268 37278
rect 30212 37174 30268 37212
rect 30380 37044 30436 37436
rect 30492 37268 30548 38612
rect 31052 38500 31108 40908
rect 31388 40516 31444 41134
rect 32264 41188 32320 41198
rect 32264 41094 32320 41132
rect 32508 41074 32564 41086
rect 32508 41022 32510 41074
rect 32562 41022 32564 41074
rect 32284 40964 32340 40974
rect 31276 40402 31332 40414
rect 31276 40350 31278 40402
rect 31330 40350 31332 40402
rect 31276 40068 31332 40350
rect 31276 40002 31332 40012
rect 31388 39730 31444 40460
rect 31500 40628 31556 40638
rect 31500 40402 31556 40572
rect 32284 40626 32340 40908
rect 32284 40574 32286 40626
rect 32338 40574 32340 40626
rect 32284 40562 32340 40574
rect 31500 40350 31502 40402
rect 31554 40350 31556 40402
rect 31500 40338 31556 40350
rect 31780 40404 31836 40414
rect 31780 40310 31836 40348
rect 32508 39844 32564 41022
rect 32620 40402 32676 42700
rect 32732 42756 32788 45052
rect 32732 42754 32900 42756
rect 32732 42702 32734 42754
rect 32786 42702 32900 42754
rect 32732 42700 32900 42702
rect 32732 42690 32788 42700
rect 32620 40350 32622 40402
rect 32674 40350 32676 40402
rect 32620 40338 32676 40350
rect 32844 40404 32900 42700
rect 32956 41970 33012 45276
rect 33068 45108 33124 45118
rect 33068 45014 33124 45052
rect 33628 44996 33684 45724
rect 34860 45668 34916 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 35028 45892 35084 45902
rect 35028 45798 35084 45836
rect 35308 45890 35364 45902
rect 35308 45838 35310 45890
rect 35362 45838 35364 45890
rect 35308 45668 35364 45838
rect 34860 45612 35028 45668
rect 33404 44940 33684 44996
rect 33852 44994 33908 45006
rect 33852 44942 33854 44994
rect 33906 44942 33908 44994
rect 33068 43540 33124 43550
rect 33068 43446 33124 43484
rect 32956 41918 32958 41970
rect 33010 41918 33012 41970
rect 32956 41906 33012 41918
rect 33068 43204 33124 43214
rect 33068 41410 33124 43148
rect 33292 43092 33348 43102
rect 33292 41970 33348 43036
rect 33292 41918 33294 41970
rect 33346 41918 33348 41970
rect 33292 41906 33348 41918
rect 33068 41358 33070 41410
rect 33122 41358 33124 41410
rect 33068 41346 33124 41358
rect 33404 41186 33460 44940
rect 33740 43538 33796 43550
rect 33740 43486 33742 43538
rect 33794 43486 33796 43538
rect 33740 43428 33796 43486
rect 33740 43362 33796 43372
rect 33852 43204 33908 44942
rect 34188 44294 34244 44306
rect 34188 44242 34190 44294
rect 34242 44242 34244 44294
rect 34076 43428 34132 43438
rect 34076 43334 34132 43372
rect 33852 43138 33908 43148
rect 34188 43092 34244 44242
rect 34972 43652 35028 45612
rect 35308 45602 35364 45612
rect 35532 45890 35588 45902
rect 35532 45838 35534 45890
rect 35586 45838 35588 45890
rect 34972 43586 35028 43596
rect 35084 45444 35140 45454
rect 34412 43538 34468 43550
rect 34412 43486 34414 43538
rect 34466 43486 34468 43538
rect 34412 43316 34468 43486
rect 34412 43250 34468 43260
rect 34748 43314 34804 43326
rect 34748 43262 34750 43314
rect 34802 43262 34804 43314
rect 34188 43026 34244 43036
rect 33740 42980 33796 42990
rect 33516 42754 33572 42766
rect 33516 42702 33518 42754
rect 33570 42702 33572 42754
rect 33516 41972 33572 42702
rect 33740 42420 33796 42924
rect 34748 42980 34804 43262
rect 34748 42914 34804 42924
rect 35084 42532 35140 45388
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 35532 44548 35588 45838
rect 35980 45862 36036 45874
rect 35980 45810 35982 45862
rect 36034 45810 36036 45862
rect 35980 45444 36036 45810
rect 35980 45378 36036 45388
rect 36428 45556 36484 45566
rect 36260 45162 36316 45174
rect 36260 45110 36262 45162
rect 36314 45110 36316 45162
rect 35756 44996 35812 45006
rect 36260 44996 36316 45110
rect 36428 45162 36484 45500
rect 36540 45332 36596 49200
rect 36988 46116 37044 46126
rect 36988 46022 37044 46060
rect 38108 46116 38164 49200
rect 38108 46050 38164 46060
rect 38668 45892 38724 45902
rect 38668 45798 38724 45836
rect 38892 45890 38948 45902
rect 38892 45838 38894 45890
rect 38946 45838 38948 45890
rect 36540 45266 36596 45276
rect 36652 45668 36708 45678
rect 36428 45110 36430 45162
rect 36482 45110 36484 45162
rect 36428 45098 36484 45110
rect 36652 45162 36708 45612
rect 36652 45110 36654 45162
rect 36706 45110 36708 45162
rect 37660 45444 37716 45454
rect 35756 44994 36316 44996
rect 35756 44942 35758 44994
rect 35810 44942 36316 44994
rect 35756 44940 36316 44942
rect 35756 44930 35812 44940
rect 36260 44772 36316 44940
rect 36652 44996 36708 45110
rect 36652 44930 36708 44940
rect 37548 45106 37604 45118
rect 37548 45054 37550 45106
rect 37602 45054 37604 45106
rect 37212 44884 37268 44894
rect 37212 44790 37268 44828
rect 36260 44716 36484 44772
rect 36428 44660 36484 44716
rect 36428 44604 36708 44660
rect 35420 44492 35588 44548
rect 35756 44548 35812 44558
rect 35308 44212 35364 44222
rect 35420 44212 35476 44492
rect 35551 44324 35607 44362
rect 35551 44258 35607 44268
rect 35364 44156 35476 44212
rect 35308 44118 35364 44156
rect 35756 43988 35812 44492
rect 36428 44322 36484 44334
rect 36428 44270 36430 44322
rect 36482 44270 36484 44322
rect 35756 43932 35924 43988
rect 35532 43565 35588 43577
rect 35532 43513 35534 43565
rect 35586 43513 35588 43565
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 35420 42868 35476 42878
rect 35420 42774 35476 42812
rect 33740 42354 33796 42364
rect 34188 42476 35140 42532
rect 33964 41972 34020 41982
rect 33516 41970 34020 41972
rect 33516 41918 33966 41970
rect 34018 41918 34020 41970
rect 33516 41916 34020 41918
rect 33964 41906 34020 41916
rect 34076 41188 34132 41198
rect 33404 41134 33406 41186
rect 33458 41134 33460 41186
rect 33404 41122 33460 41134
rect 33964 41186 34132 41188
rect 33964 41134 34078 41186
rect 34130 41134 34132 41186
rect 33964 41132 34132 41134
rect 33740 40962 33796 40974
rect 33740 40910 33742 40962
rect 33794 40910 33796 40962
rect 32956 40404 33012 40414
rect 32844 40402 33012 40404
rect 32844 40350 32958 40402
rect 33010 40350 33012 40402
rect 32844 40348 33012 40350
rect 32508 39778 32564 39788
rect 32620 39786 32676 39798
rect 31388 39678 31390 39730
rect 31442 39678 31444 39730
rect 31388 39666 31444 39678
rect 32620 39734 32622 39786
rect 32674 39734 32676 39786
rect 32620 39732 32676 39734
rect 32620 39666 32676 39676
rect 31612 39620 31668 39630
rect 31220 39562 31276 39574
rect 31220 39510 31222 39562
rect 31274 39510 31276 39562
rect 32396 39620 32452 39630
rect 31612 39526 31668 39564
rect 31780 39562 31836 39574
rect 31780 39518 31782 39562
rect 31220 39060 31276 39510
rect 31724 39510 31782 39518
rect 31834 39510 31836 39562
rect 32396 39526 32452 39564
rect 32732 39618 32788 39630
rect 32732 39566 32734 39618
rect 32786 39566 32788 39618
rect 31724 39508 31836 39510
rect 31780 39452 31836 39508
rect 32732 39508 32788 39566
rect 31724 39396 31780 39452
rect 32732 39442 32788 39452
rect 31220 38994 31276 39004
rect 31612 39340 31780 39396
rect 31388 38948 31444 38958
rect 31612 38948 31668 39340
rect 31388 38946 31668 38948
rect 31388 38894 31390 38946
rect 31442 38894 31668 38946
rect 31388 38892 31668 38894
rect 31388 38882 31444 38892
rect 31780 38890 31836 38902
rect 31780 38838 31782 38890
rect 31834 38838 31836 38890
rect 32340 38890 32396 38902
rect 31780 38836 31836 38838
rect 31052 38434 31108 38444
rect 31724 38780 31836 38836
rect 32172 38864 32228 38876
rect 32172 38812 32174 38864
rect 32226 38812 32228 38864
rect 30716 38052 30772 38062
rect 31724 38052 31780 38780
rect 31948 38724 32004 38734
rect 31836 38668 31948 38724
rect 31836 38274 31892 38668
rect 31948 38658 32004 38668
rect 31836 38222 31838 38274
rect 31890 38222 31892 38274
rect 31836 38210 31892 38222
rect 32060 38612 32116 38622
rect 30716 37958 30772 37996
rect 31592 37996 31780 38052
rect 31592 37994 31648 37996
rect 31592 37942 31594 37994
rect 31646 37942 31648 37994
rect 31592 37940 31648 37942
rect 31592 37874 31648 37884
rect 30660 37492 30716 37502
rect 30660 37398 30716 37436
rect 30604 37268 30660 37278
rect 31052 37268 31108 37278
rect 30492 37212 30604 37268
rect 30268 36988 30436 37044
rect 30136 36596 30192 36606
rect 30136 36482 30192 36540
rect 30136 36430 30138 36482
rect 30190 36430 30192 36482
rect 30136 36418 30192 36430
rect 30268 36484 30324 36988
rect 30380 36708 30436 36718
rect 30380 36614 30436 36652
rect 30268 36428 30492 36484
rect 29932 36204 30212 36260
rect 29036 35758 29038 35810
rect 29090 35758 29092 35810
rect 29036 35746 29092 35758
rect 29148 36148 29204 36158
rect 28588 35308 28756 35364
rect 27580 35298 27636 35308
rect 28364 35252 28420 35262
rect 27244 35084 28308 35140
rect 28028 34916 28084 34926
rect 27524 34860 27580 34870
rect 27244 34858 27580 34860
rect 27244 34806 27526 34858
rect 27578 34806 27580 34858
rect 27244 34804 27580 34806
rect 27244 34468 27300 34804
rect 27524 34794 27580 34804
rect 27804 34860 27860 34870
rect 27804 34858 27972 34860
rect 27804 34806 27806 34858
rect 27858 34806 27972 34858
rect 28028 34832 28030 34860
rect 28082 34832 28084 34860
rect 28028 34820 28084 34832
rect 27804 34804 27972 34806
rect 27804 34794 27860 34804
rect 27244 34130 27300 34412
rect 27244 34078 27246 34130
rect 27298 34078 27300 34130
rect 27244 34066 27300 34078
rect 27916 33796 27972 34804
rect 28120 34130 28176 34142
rect 28120 34078 28122 34130
rect 28174 34078 28176 34130
rect 28120 34020 28176 34078
rect 27020 33740 27300 33796
rect 26852 33684 26908 33694
rect 26908 33628 27020 33684
rect 26852 33618 26908 33628
rect 26964 33458 27020 33628
rect 26964 33406 26966 33458
rect 27018 33406 27020 33458
rect 26964 33394 27020 33406
rect 26292 33122 26740 33124
rect 26292 33070 26294 33122
rect 26346 33070 26740 33122
rect 26292 33068 26740 33070
rect 26292 32564 26348 33068
rect 26292 32498 26348 32508
rect 26124 32450 26180 32462
rect 26124 32398 26126 32450
rect 26178 32398 26180 32450
rect 26124 32228 26180 32398
rect 27244 32228 27300 33740
rect 27916 33730 27972 33740
rect 28028 33964 28176 34020
rect 27356 33684 27412 33694
rect 27356 33570 27412 33628
rect 27356 33518 27358 33570
rect 27410 33518 27412 33570
rect 27356 33506 27412 33518
rect 27636 33290 27692 33302
rect 27636 33238 27638 33290
rect 27690 33238 27692 33290
rect 27636 32788 27692 33238
rect 27916 33290 27972 33302
rect 27916 33238 27918 33290
rect 27970 33238 27972 33290
rect 27636 32732 27748 32788
rect 27692 32452 27748 32732
rect 27916 32676 27972 33238
rect 28028 32788 28084 33964
rect 28140 33796 28196 33806
rect 28140 33290 28196 33740
rect 28140 33238 28142 33290
rect 28194 33238 28196 33290
rect 28140 32900 28196 33238
rect 28252 33012 28308 35084
rect 28364 34916 28420 35196
rect 28476 35140 28532 35150
rect 28476 35046 28532 35084
rect 28364 34860 28532 34916
rect 28364 34244 28420 34254
rect 28364 34150 28420 34188
rect 28476 33684 28532 34860
rect 28476 33618 28532 33628
rect 28252 32956 28420 33012
rect 28140 32844 28308 32900
rect 28028 32732 28196 32788
rect 27916 32610 27972 32620
rect 28028 32452 28084 32462
rect 27692 32450 28084 32452
rect 27692 32398 28030 32450
rect 28082 32398 28084 32450
rect 27692 32396 28084 32398
rect 26124 32172 26740 32228
rect 26012 32060 26348 32116
rect 26292 31890 26348 32060
rect 26292 31838 26294 31890
rect 26346 31838 26348 31890
rect 25844 31780 25900 31790
rect 25844 31554 25900 31724
rect 25844 31502 25846 31554
rect 25898 31502 25900 31554
rect 25844 31444 25900 31502
rect 25844 31378 25900 31388
rect 26292 31220 26348 31838
rect 26572 32004 26628 32014
rect 25564 31164 25844 31220
rect 25228 31108 25284 31118
rect 25228 31006 25284 31052
rect 25228 30994 25340 31006
rect 25564 30996 25620 31006
rect 25228 30942 25286 30994
rect 25338 30942 25340 30994
rect 25228 30940 25340 30942
rect 25284 30930 25340 30940
rect 25452 30994 25620 30996
rect 25452 30942 25566 30994
rect 25618 30942 25620 30994
rect 25452 30940 25620 30942
rect 25452 30212 25508 30940
rect 25564 30930 25620 30940
rect 25676 30996 25732 31006
rect 25676 30902 25732 30940
rect 25788 30660 25844 31164
rect 26292 31218 26404 31220
rect 26292 31166 26294 31218
rect 26346 31166 26404 31218
rect 26292 31154 26404 31166
rect 25788 30594 25844 30604
rect 25228 30100 25284 30110
rect 25228 30006 25284 30044
rect 25004 29820 25228 29876
rect 25172 29482 25228 29820
rect 25172 29430 25174 29482
rect 25226 29430 25228 29482
rect 25340 29540 25396 29550
rect 25340 29446 25396 29484
rect 25172 29418 25228 29430
rect 25228 29204 25284 29214
rect 25452 29204 25508 30156
rect 25676 30210 25732 30222
rect 25676 30158 25678 30210
rect 25730 30158 25732 30210
rect 25676 30100 25732 30158
rect 25676 30034 25732 30044
rect 26124 29876 26180 29886
rect 26012 29652 26068 29662
rect 25732 29482 25788 29494
rect 25564 29428 25620 29438
rect 25732 29430 25734 29482
rect 25786 29430 25788 29482
rect 25732 29428 25788 29430
rect 25564 29334 25620 29372
rect 25676 29372 25788 29428
rect 26012 29428 26068 29596
rect 25676 29204 25732 29372
rect 26012 29362 26068 29372
rect 25452 29148 25732 29204
rect 25228 28644 25284 29148
rect 25228 28588 25396 28644
rect 25172 28420 25228 28430
rect 24780 28418 25228 28420
rect 24780 28366 25174 28418
rect 25226 28366 25228 28418
rect 24780 28364 25228 28366
rect 24556 27186 24668 27198
rect 24556 27134 24614 27186
rect 24666 27134 24668 27186
rect 24556 27132 24668 27134
rect 24612 27122 24668 27132
rect 24892 27188 24948 27198
rect 24892 27074 24948 27132
rect 24892 27022 24894 27074
rect 24946 27022 24948 27074
rect 24892 26964 24948 27022
rect 24892 26898 24948 26908
rect 24668 26628 24724 26638
rect 24444 26070 24446 26122
rect 24498 26070 24500 26122
rect 24556 26290 24612 26302
rect 24556 26238 24558 26290
rect 24610 26238 24612 26290
rect 24556 26180 24612 26238
rect 24556 26114 24612 26124
rect 24444 26058 24500 26070
rect 24668 25956 24724 26572
rect 24556 25900 24724 25956
rect 24332 25340 24500 25396
rect 24332 24722 24388 24734
rect 24332 24670 24334 24722
rect 24386 24670 24388 24722
rect 24332 24276 24388 24670
rect 24444 24612 24500 25340
rect 24556 24834 24612 25900
rect 24836 25284 24892 25294
rect 24836 25190 24892 25228
rect 24556 24782 24558 24834
rect 24610 24782 24612 24834
rect 24556 24770 24612 24782
rect 24724 24724 24780 24734
rect 24724 24630 24780 24668
rect 24444 24546 24500 24556
rect 24892 24500 24948 24510
rect 24332 24220 24836 24276
rect 24220 24210 24276 24220
rect 23660 24098 23716 24108
rect 23660 23940 23716 23950
rect 23660 23938 23940 23940
rect 23660 23886 23662 23938
rect 23714 23886 23940 23938
rect 23660 23884 23940 23886
rect 23660 23874 23716 23884
rect 23548 23538 23604 23548
rect 23884 23492 23940 23884
rect 24780 23492 24836 24220
rect 23884 23436 24500 23492
rect 24444 23378 24500 23436
rect 24444 23326 24446 23378
rect 24498 23326 24500 23378
rect 24444 23314 24500 23326
rect 23884 23268 23940 23278
rect 23626 23191 23682 23203
rect 23626 23156 23628 23191
rect 23680 23156 23682 23191
rect 23772 23156 23828 23166
rect 23682 23100 23716 23156
rect 23626 23062 23716 23100
rect 23772 23062 23828 23100
rect 23884 23154 23940 23212
rect 23884 23102 23886 23154
rect 23938 23102 23940 23154
rect 23884 23090 23940 23102
rect 24108 23154 24164 23166
rect 24108 23102 24110 23154
rect 24162 23102 24164 23154
rect 23212 22932 23268 22942
rect 23212 22930 23434 22932
rect 23212 22878 23214 22930
rect 23266 22878 23434 22930
rect 23212 22876 23434 22878
rect 23212 22866 23268 22876
rect 23212 22708 23268 22718
rect 23100 22372 23156 22382
rect 23100 22278 23156 22316
rect 23212 22370 23268 22652
rect 23212 22318 23214 22370
rect 23266 22318 23268 22370
rect 22988 22194 23044 22204
rect 23044 21924 23100 21934
rect 23044 21810 23100 21868
rect 23044 21758 23046 21810
rect 23098 21758 23100 21810
rect 23044 21746 23100 21758
rect 23100 20916 23156 20926
rect 23100 20802 23156 20860
rect 23100 20750 23102 20802
rect 23154 20750 23156 20802
rect 23100 20738 23156 20750
rect 23212 20804 23268 22318
rect 23378 22370 23434 22876
rect 23378 22318 23380 22370
rect 23432 22318 23434 22370
rect 23378 22306 23434 22318
rect 23548 22820 23604 22830
rect 23548 22148 23604 22764
rect 23436 22092 23604 22148
rect 23436 21140 23492 22092
rect 23660 21924 23716 23062
rect 23772 22596 23828 22606
rect 24108 22596 24164 23102
rect 23772 22594 24164 22596
rect 23772 22542 23774 22594
rect 23826 22542 24164 22594
rect 23772 22540 24164 22542
rect 23772 22530 23828 22540
rect 24780 22370 24836 23436
rect 24892 22820 24948 24444
rect 25004 24388 25060 28364
rect 25172 28354 25228 28364
rect 25116 28196 25172 28206
rect 25116 26068 25172 28140
rect 25340 28094 25396 28588
rect 25452 28642 25508 28654
rect 25452 28590 25454 28642
rect 25506 28590 25508 28642
rect 25452 28308 25508 28590
rect 25452 28242 25508 28252
rect 25564 28644 25620 28654
rect 25340 28082 25452 28094
rect 25340 28030 25398 28082
rect 25450 28030 25452 28082
rect 25340 28028 25452 28030
rect 25396 28018 25452 28028
rect 25564 27186 25620 28588
rect 26012 27873 26068 27898
rect 25788 27860 25844 27870
rect 26012 27860 26014 27873
rect 26066 27860 26068 27873
rect 25788 27858 25956 27860
rect 25788 27806 25790 27858
rect 25842 27806 25956 27858
rect 25788 27804 25956 27806
rect 25788 27794 25844 27804
rect 25564 27134 25566 27186
rect 25618 27134 25620 27186
rect 25564 27122 25620 27134
rect 25676 27188 25732 27198
rect 25340 27074 25396 27086
rect 25340 27022 25342 27074
rect 25394 27022 25396 27074
rect 25340 26908 25396 27022
rect 25676 26908 25732 27132
rect 25788 27076 25844 27114
rect 25788 27010 25844 27020
rect 25340 26852 25620 26908
rect 25676 26852 25844 26908
rect 25340 26628 25396 26638
rect 25340 26346 25396 26572
rect 25228 26325 25284 26337
rect 25228 26292 25230 26325
rect 25282 26292 25284 26325
rect 25340 26294 25342 26346
rect 25394 26294 25396 26346
rect 25340 26282 25396 26294
rect 25564 26404 25620 26852
rect 25564 26346 25620 26348
rect 25564 26294 25566 26346
rect 25618 26294 25620 26346
rect 25564 26282 25620 26294
rect 25788 26346 25844 26852
rect 25788 26294 25790 26346
rect 25842 26294 25844 26346
rect 25788 26282 25844 26294
rect 25228 26226 25284 26236
rect 25116 26002 25172 26012
rect 25116 25478 25172 25490
rect 25116 25426 25118 25478
rect 25170 25426 25172 25478
rect 25116 25284 25172 25426
rect 25116 25218 25172 25228
rect 25788 25172 25844 25182
rect 25676 25060 25732 25070
rect 25452 24722 25508 24734
rect 25452 24670 25454 24722
rect 25506 24670 25508 24722
rect 25284 24612 25340 24622
rect 25284 24554 25340 24556
rect 25284 24502 25286 24554
rect 25338 24502 25340 24554
rect 25284 24490 25340 24502
rect 25452 24612 25508 24670
rect 25676 24666 25732 25004
rect 25788 24948 25844 25116
rect 25788 24778 25844 24892
rect 25788 24726 25790 24778
rect 25842 24726 25844 24778
rect 25900 24836 25956 27804
rect 26012 27794 26068 27804
rect 26124 27746 26180 29820
rect 26348 29876 26404 31154
rect 26572 30436 26628 31948
rect 26684 32002 26740 32172
rect 26684 31950 26686 32002
rect 26738 31950 26740 32002
rect 26684 31938 26740 31950
rect 26908 32172 27300 32228
rect 26908 31556 26964 32172
rect 27020 31892 27076 31902
rect 27020 31778 27076 31836
rect 27020 31726 27022 31778
rect 27074 31726 27076 31778
rect 27020 31714 27076 31726
rect 27244 31780 27300 31790
rect 27244 31686 27300 31724
rect 27916 31780 27972 32396
rect 28028 32386 28084 32396
rect 28140 31790 28196 32732
rect 27916 31714 27972 31724
rect 28120 31780 28196 31790
rect 28176 31724 28196 31780
rect 28120 31686 28176 31724
rect 28252 31556 28308 32844
rect 28364 32004 28420 32956
rect 28364 31938 28420 31948
rect 28532 32338 28588 32350
rect 28532 32286 28534 32338
rect 28586 32286 28588 32338
rect 28532 31892 28588 32286
rect 28532 31826 28588 31836
rect 26908 31500 27076 31556
rect 26740 31220 26796 31230
rect 26796 31164 26964 31220
rect 26740 31126 26796 31164
rect 26908 30994 26964 31164
rect 26908 30942 26910 30994
rect 26962 30942 26964 30994
rect 26908 30930 26964 30942
rect 26572 30380 26740 30436
rect 26552 30156 26608 30166
rect 26552 30154 26628 30156
rect 26552 30102 26554 30154
rect 26606 30102 26628 30154
rect 26552 30090 26628 30102
rect 26572 29988 26628 30090
rect 26348 29810 26404 29820
rect 26460 29932 26628 29988
rect 26460 29316 26516 29932
rect 26684 29876 26740 30380
rect 26796 30212 26852 30222
rect 26796 30118 26852 30156
rect 26460 29250 26516 29260
rect 26572 29820 26740 29876
rect 26572 28756 26628 29820
rect 27020 29764 27076 31500
rect 27916 31500 28308 31556
rect 28364 31780 28420 31790
rect 27804 31444 27860 31454
rect 27804 31106 27860 31388
rect 27804 31054 27806 31106
rect 27858 31054 27860 31106
rect 27804 31042 27860 31054
rect 27636 30938 27692 30950
rect 27636 30886 27638 30938
rect 27690 30886 27692 30938
rect 27244 30770 27300 30782
rect 27244 30718 27246 30770
rect 27298 30718 27300 30770
rect 27244 29988 27300 30718
rect 27636 30436 27692 30886
rect 27580 30380 27692 30436
rect 27412 29988 27468 29998
rect 27244 29986 27468 29988
rect 27244 29934 27414 29986
rect 27466 29934 27468 29986
rect 27244 29932 27468 29934
rect 27412 29876 27468 29932
rect 27580 29876 27636 30380
rect 27916 30378 27972 31500
rect 28364 31220 28420 31724
rect 28028 31164 28420 31220
rect 28476 31668 28532 31678
rect 28028 30994 28084 31164
rect 28476 31108 28532 31612
rect 28700 31220 28756 35308
rect 28812 35252 28868 35262
rect 28812 33236 28868 35196
rect 28924 34030 28980 35532
rect 29148 35252 29204 36092
rect 29148 35186 29204 35196
rect 29820 36036 29876 36046
rect 29148 34914 29204 34926
rect 29148 34862 29150 34914
rect 29202 34862 29204 34914
rect 29148 34244 29204 34862
rect 29820 34356 29876 35980
rect 29988 36036 30044 36046
rect 29988 35588 30044 35980
rect 29988 35494 30044 35532
rect 30024 34916 30080 34926
rect 30024 34822 30080 34860
rect 29148 34178 29204 34188
rect 29484 34300 29876 34356
rect 28924 34018 29036 34030
rect 28924 33966 28982 34018
rect 29034 33966 29036 34018
rect 28924 33964 29036 33966
rect 28980 33460 29036 33964
rect 28980 33394 29036 33404
rect 29260 33346 29316 33358
rect 29260 33294 29262 33346
rect 29314 33294 29316 33346
rect 28812 33180 28980 33236
rect 28812 32562 28868 32574
rect 28812 32510 28814 32562
rect 28866 32510 28868 32562
rect 28812 31444 28868 32510
rect 28812 31378 28868 31388
rect 28700 31154 28756 31164
rect 28028 30942 28030 30994
rect 28082 30942 28084 30994
rect 28364 31052 28532 31108
rect 28364 31032 28420 31052
rect 28364 30980 28366 31032
rect 28418 30980 28420 31032
rect 28924 30996 28980 33180
rect 29036 32562 29092 32574
rect 29036 32510 29038 32562
rect 29090 32510 29092 32562
rect 29036 32004 29092 32510
rect 29260 32564 29316 33294
rect 29372 33346 29428 33358
rect 29372 33294 29374 33346
rect 29426 33294 29428 33346
rect 29372 32788 29428 33294
rect 29484 33348 29540 34300
rect 29596 34132 29652 34142
rect 29764 34132 29820 34142
rect 29596 34130 29708 34132
rect 29596 34078 29598 34130
rect 29650 34078 29708 34130
rect 29596 34066 29708 34078
rect 29652 33570 29708 34066
rect 29764 34038 29820 34076
rect 29932 34130 29988 34142
rect 29932 34078 29934 34130
rect 29986 34078 29988 34130
rect 29932 33684 29988 34078
rect 29652 33518 29654 33570
rect 29706 33518 29708 33570
rect 29652 33506 29708 33518
rect 29820 33628 29988 33684
rect 30044 34130 30100 34142
rect 30044 34078 30046 34130
rect 30098 34078 30100 34130
rect 30044 33684 30100 34078
rect 30156 33796 30212 36204
rect 30436 35922 30492 36428
rect 30436 35870 30438 35922
rect 30490 35870 30492 35922
rect 30436 35858 30492 35870
rect 30268 35812 30324 35822
rect 30268 35138 30324 35756
rect 30604 35700 30660 37212
rect 30828 37266 31108 37268
rect 30828 37214 31054 37266
rect 31106 37214 31108 37266
rect 30828 37212 31108 37214
rect 30828 36708 30884 37212
rect 31052 37202 31108 37212
rect 31928 37266 31984 37278
rect 31928 37214 31930 37266
rect 31982 37214 31984 37266
rect 31928 36820 31984 37214
rect 32060 37044 32116 38556
rect 32172 38276 32228 38812
rect 32340 38838 32342 38890
rect 32394 38838 32396 38890
rect 32340 38668 32396 38838
rect 32732 38836 32788 38846
rect 32340 38612 32564 38668
rect 32340 38276 32396 38286
rect 32172 38274 32396 38276
rect 32172 38222 32342 38274
rect 32394 38222 32396 38274
rect 32172 38220 32396 38222
rect 32340 38210 32396 38220
rect 32172 38052 32228 38062
rect 32172 37958 32228 37996
rect 32508 37828 32564 38612
rect 32620 38050 32676 38062
rect 32620 37998 32622 38050
rect 32674 37998 32676 38050
rect 32620 37828 32676 37998
rect 32732 37940 32788 38780
rect 32844 38052 32900 40348
rect 32956 40338 33012 40348
rect 33740 40402 33796 40910
rect 33740 40350 33742 40402
rect 33794 40350 33796 40402
rect 33740 40338 33796 40350
rect 33852 40740 33908 40750
rect 33852 39732 33908 40684
rect 33740 39676 33908 39732
rect 33068 39620 33124 39630
rect 33068 39526 33124 39564
rect 33292 39618 33348 39630
rect 33292 39566 33294 39618
rect 33346 39566 33348 39618
rect 33292 39508 33348 39566
rect 33572 39620 33628 39630
rect 33572 39526 33628 39564
rect 33292 39442 33348 39452
rect 33068 38836 33124 38874
rect 33068 38770 33124 38780
rect 33740 38052 33796 39676
rect 33964 39060 34020 41132
rect 34076 41122 34132 41132
rect 34188 40964 34244 42476
rect 34412 42308 34468 42318
rect 35532 42308 35588 43513
rect 35868 42922 35924 43932
rect 36204 43652 36260 43662
rect 36204 43426 36260 43596
rect 36428 43652 36484 44270
rect 36428 43586 36484 43596
rect 36652 43540 36708 44604
rect 36652 43474 36708 43484
rect 36988 44294 37044 44306
rect 36988 44242 36990 44294
rect 37042 44242 37044 44294
rect 36204 43374 36206 43426
rect 36258 43374 36260 43426
rect 36204 43362 36260 43374
rect 35868 42870 35870 42922
rect 35922 42870 35924 42922
rect 35868 42858 35924 42870
rect 35980 42754 36036 42766
rect 35980 42702 35982 42754
rect 36034 42702 36036 42754
rect 35532 42252 35700 42308
rect 34300 42196 34356 42206
rect 34300 41970 34356 42140
rect 34300 41918 34302 41970
rect 34354 41918 34356 41970
rect 34300 41906 34356 41918
rect 34412 41188 34468 42252
rect 34580 42196 34636 42206
rect 34580 42194 34916 42196
rect 34580 42142 34582 42194
rect 34634 42142 34916 42194
rect 34580 42140 34916 42142
rect 34580 42130 34636 42140
rect 34748 41970 34804 41982
rect 34748 41918 34750 41970
rect 34802 41918 34804 41970
rect 34748 41748 34804 41918
rect 34860 41972 34916 42140
rect 34972 41972 35028 41982
rect 34860 41970 35028 41972
rect 34860 41918 34974 41970
rect 35026 41918 35028 41970
rect 34860 41916 35028 41918
rect 34972 41906 35028 41916
rect 34748 41682 34804 41692
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35532 41300 35588 41310
rect 34748 41188 34804 41198
rect 34412 41186 34804 41188
rect 34412 41134 34750 41186
rect 34802 41134 34804 41186
rect 34412 41132 34804 41134
rect 34748 41122 34804 41132
rect 35084 41186 35140 41198
rect 35084 41134 35086 41186
rect 35138 41134 35140 41186
rect 34412 40964 34468 40974
rect 34188 40962 34468 40964
rect 34188 40910 34414 40962
rect 34466 40910 34468 40962
rect 34188 40908 34468 40910
rect 34412 40898 34468 40908
rect 35084 40628 35140 41134
rect 35084 40562 35140 40572
rect 35420 40962 35476 40974
rect 35420 40910 35422 40962
rect 35474 40910 35476 40962
rect 34860 40404 34916 40414
rect 34860 40068 34916 40348
rect 35420 40180 35476 40910
rect 35420 40114 35476 40124
rect 34300 40012 34916 40068
rect 35196 40012 35460 40022
rect 34300 39618 34356 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35532 39844 35588 41244
rect 35644 40740 35700 42252
rect 35980 42084 36036 42702
rect 35980 42018 36036 42028
rect 36204 42754 36260 42766
rect 36876 42756 36932 42766
rect 36204 42702 36206 42754
rect 36258 42702 36260 42754
rect 35848 41972 35904 41982
rect 35848 41878 35904 41916
rect 36092 41860 36148 41870
rect 36092 41766 36148 41804
rect 36204 41524 36260 42702
rect 36764 42754 36932 42756
rect 36764 42702 36878 42754
rect 36930 42702 36932 42754
rect 36764 42700 36932 42702
rect 36652 42084 36708 42094
rect 36652 42026 36708 42028
rect 36652 41974 36654 42026
rect 36706 41974 36708 42026
rect 36652 41962 36708 41974
rect 36204 41458 36260 41468
rect 36316 41860 36372 41870
rect 35924 41412 35980 41422
rect 35924 41318 35980 41356
rect 36204 41188 36260 41198
rect 36204 41094 36260 41132
rect 36316 41186 36372 41804
rect 36764 41412 36820 42700
rect 36876 42690 36932 42700
rect 36988 42196 37044 44242
rect 36876 42140 37044 42196
rect 37100 42754 37156 42766
rect 37100 42702 37102 42754
rect 37154 42702 37156 42754
rect 36876 42084 36932 42140
rect 36876 42018 36932 42028
rect 37100 42084 37156 42702
rect 37380 42642 37436 42654
rect 37380 42590 37382 42642
rect 37434 42590 37436 42642
rect 37380 42196 37436 42590
rect 37380 42130 37436 42140
rect 37100 42018 37156 42028
rect 36764 41346 36820 41356
rect 36988 42000 37044 42012
rect 36988 41948 36990 42000
rect 37042 41948 37044 42000
rect 36988 41748 37044 41948
rect 37324 41972 37380 41982
rect 37548 41972 37604 45054
rect 37156 41916 37212 41926
rect 36316 41134 36318 41186
rect 36370 41134 36372 41186
rect 36316 41122 36372 41134
rect 36988 41188 37044 41692
rect 37100 41914 37212 41916
rect 37100 41862 37158 41914
rect 37210 41862 37212 41914
rect 37380 41916 37492 41972
rect 37324 41906 37380 41916
rect 37100 41850 37212 41862
rect 37436 41858 37492 41916
rect 37100 41636 37156 41850
rect 37436 41806 37438 41858
rect 37490 41806 37492 41858
rect 37436 41794 37492 41806
rect 37436 41636 37492 41646
rect 37100 41580 37436 41636
rect 37436 41570 37492 41580
rect 35644 40684 36260 40740
rect 35644 40404 35700 40414
rect 35644 40310 35700 40348
rect 35196 39788 35588 39844
rect 34300 39566 34302 39618
rect 34354 39566 34356 39618
rect 34300 39554 34356 39566
rect 34524 39618 34580 39630
rect 34524 39566 34526 39618
rect 34578 39566 34580 39618
rect 34132 39396 34188 39406
rect 34524 39396 34580 39566
rect 34132 39394 34580 39396
rect 34132 39342 34134 39394
rect 34186 39342 34580 39394
rect 34132 39340 34580 39342
rect 34636 39396 34692 39406
rect 34132 39330 34188 39340
rect 34636 39060 34692 39340
rect 33964 38994 34020 39004
rect 34524 39004 34692 39060
rect 35084 39060 35140 39070
rect 33944 38834 34000 38846
rect 33944 38782 33946 38834
rect 33998 38782 34000 38834
rect 33944 38724 34000 38782
rect 33944 38658 34000 38668
rect 34188 38610 34244 38622
rect 34188 38558 34190 38610
rect 34242 38558 34244 38610
rect 34188 38276 34244 38558
rect 34188 38210 34244 38220
rect 34524 38274 34580 39004
rect 34804 38836 34860 38846
rect 34804 38742 34860 38780
rect 35084 38834 35140 39004
rect 35084 38782 35086 38834
rect 35138 38782 35140 38834
rect 35084 38770 35140 38782
rect 35196 38668 35252 39788
rect 35756 39732 35812 40684
rect 36204 40458 36260 40684
rect 36204 40406 36206 40458
rect 36258 40406 36260 40458
rect 36708 40516 36764 40526
rect 36708 40458 36764 40460
rect 36204 40394 36260 40406
rect 36428 40441 36484 40453
rect 36428 40389 36430 40441
rect 36482 40389 36484 40441
rect 36204 40292 36260 40302
rect 36204 39842 36260 40236
rect 36204 39790 36206 39842
rect 36258 39790 36260 39842
rect 36204 39778 36260 39790
rect 35400 39676 35812 39732
rect 35400 39618 35456 39676
rect 35400 39566 35402 39618
rect 35454 39566 35456 39618
rect 35400 39554 35456 39566
rect 35644 39506 35700 39518
rect 35644 39454 35646 39506
rect 35698 39454 35700 39506
rect 35644 39396 35700 39454
rect 35308 39340 35700 39396
rect 35308 38948 35364 39340
rect 35756 39060 35812 39676
rect 36204 39172 36260 39182
rect 35644 39004 35812 39060
rect 35868 39060 35924 39070
rect 35308 38892 35588 38948
rect 35308 38834 35364 38892
rect 35308 38782 35310 38834
rect 35362 38782 35364 38834
rect 35532 38890 35588 38892
rect 35532 38838 35534 38890
rect 35586 38838 35588 38890
rect 35532 38826 35588 38838
rect 35308 38770 35364 38782
rect 35644 38724 35700 39004
rect 35868 38948 35924 39004
rect 35812 38892 35924 38948
rect 36204 38948 36260 39116
rect 36428 39060 36484 40389
rect 36540 40404 36596 40414
rect 36708 40406 36710 40458
rect 36762 40406 36764 40458
rect 36988 40514 37044 41132
rect 37212 41188 37268 41198
rect 37212 41106 37214 41132
rect 37266 41106 37268 41132
rect 37212 41094 37268 41106
rect 37436 41186 37492 41198
rect 37436 41134 37438 41186
rect 37490 41134 37492 41186
rect 37436 41076 37492 41134
rect 37548 41188 37604 41916
rect 37660 41298 37716 45388
rect 38892 45444 38948 45838
rect 39172 45780 39228 45790
rect 39172 45686 39228 45724
rect 38892 45378 38948 45388
rect 37996 45332 38052 45342
rect 37996 44546 38052 45276
rect 38332 44996 38388 45006
rect 38332 44994 38612 44996
rect 38332 44942 38334 44994
rect 38386 44942 38612 44994
rect 38332 44940 38612 44942
rect 38332 44930 38388 44940
rect 37996 44494 37998 44546
rect 38050 44494 38052 44546
rect 37996 44482 38052 44494
rect 38052 43706 38108 43718
rect 38052 43654 38054 43706
rect 38106 43654 38108 43706
rect 38052 43652 38108 43654
rect 38556 43708 38612 44940
rect 39004 44772 39060 44782
rect 38799 44100 38855 44110
rect 38556 43652 38724 43708
rect 38052 43586 38108 43596
rect 37884 43540 37940 43550
rect 37884 43446 37940 43484
rect 38556 43540 38612 43550
rect 38108 42642 38164 42654
rect 38108 42590 38110 42642
rect 38162 42590 38164 42642
rect 38108 42308 38164 42590
rect 38108 42242 38164 42252
rect 37996 42084 38052 42094
rect 37996 41990 38052 42028
rect 38556 42084 38612 43484
rect 38556 42018 38612 42028
rect 38444 41998 38500 42010
rect 38220 41970 38276 41982
rect 37828 41914 37884 41926
rect 37828 41862 37830 41914
rect 37882 41862 37884 41914
rect 37828 41860 37884 41862
rect 38220 41918 38222 41970
rect 38274 41918 38276 41970
rect 38220 41860 38276 41918
rect 37828 41804 38164 41860
rect 37660 41246 37662 41298
rect 37714 41246 37716 41298
rect 37660 41234 37716 41246
rect 37828 41636 37884 41646
rect 37828 41242 37884 41580
rect 38108 41524 38164 41804
rect 38220 41794 38276 41804
rect 38444 41946 38446 41998
rect 38498 41946 38500 41998
rect 38444 41748 38500 41946
rect 38444 41682 38500 41692
rect 38332 41524 38388 41534
rect 38108 41468 38276 41524
rect 37828 41190 37830 41242
rect 37882 41190 37884 41242
rect 37828 41178 37884 41190
rect 38108 41188 38164 41198
rect 37548 41122 37604 41132
rect 37996 41132 38108 41188
rect 37436 41010 37492 41020
rect 36988 40462 36990 40514
rect 37042 40462 37044 40514
rect 36988 40450 37044 40462
rect 37660 40516 37716 40526
rect 36708 40394 36764 40406
rect 37324 40404 37380 40414
rect 37212 40402 37380 40404
rect 36540 39618 36596 40348
rect 37212 40350 37326 40402
rect 37378 40350 37380 40402
rect 37212 40348 37380 40350
rect 36540 39566 36542 39618
rect 36594 39566 36596 39618
rect 36540 39554 36596 39566
rect 36652 40180 36708 40190
rect 36652 39172 36708 40124
rect 37212 39742 37268 40348
rect 37324 40338 37380 40348
rect 37548 40402 37604 40414
rect 37548 40350 37550 40402
rect 37602 40350 37604 40402
rect 37548 39844 37604 40350
rect 37156 39732 37268 39742
rect 37212 39676 37268 39732
rect 37324 39788 37604 39844
rect 37660 39854 37716 40460
rect 37828 40404 37884 40414
rect 37828 40310 37884 40348
rect 37884 40068 37940 40078
rect 37660 39842 37772 39854
rect 37660 39790 37718 39842
rect 37770 39790 37772 39842
rect 37660 39788 37772 39790
rect 37156 39674 37212 39676
rect 36988 39618 37044 39630
rect 36988 39566 36990 39618
rect 37042 39566 37044 39618
rect 37156 39622 37158 39674
rect 37210 39622 37212 39674
rect 37156 39610 37212 39622
rect 37324 39620 37380 39788
rect 37716 39778 37772 39788
rect 36988 39172 37044 39566
rect 37324 39526 37380 39564
rect 37436 39620 37492 39630
rect 37884 39620 37940 40012
rect 37436 39618 37940 39620
rect 37436 39566 37438 39618
rect 37490 39566 37940 39618
rect 37436 39564 37940 39566
rect 36988 39116 37268 39172
rect 36652 39106 36708 39116
rect 36428 38994 36484 39004
rect 36988 38948 37044 38958
rect 36204 38892 36372 38948
rect 35812 38890 35868 38892
rect 35812 38838 35814 38890
rect 35866 38838 35868 38890
rect 35812 38724 35868 38838
rect 36316 38846 36372 38892
rect 36316 38834 36428 38846
rect 36316 38782 36374 38834
rect 36426 38782 36428 38834
rect 36316 38780 36428 38782
rect 36372 38770 36428 38780
rect 36540 38836 36596 38874
rect 36540 38770 36596 38780
rect 36764 38834 36820 38846
rect 36764 38782 36766 38834
rect 36818 38782 36820 38834
rect 34524 38222 34526 38274
rect 34578 38222 34580 38274
rect 34524 38210 34580 38222
rect 35084 38612 35252 38668
rect 35420 38668 35700 38724
rect 35756 38668 35868 38724
rect 36204 38722 36260 38734
rect 36204 38670 36206 38722
rect 36258 38670 36260 38722
rect 36204 38668 36260 38670
rect 36764 38668 36820 38782
rect 35420 38612 35588 38668
rect 34860 38164 34916 38174
rect 34188 38052 34244 38062
rect 32844 37996 33012 38052
rect 33740 38050 34244 38052
rect 33740 37998 34190 38050
rect 34242 37998 34244 38050
rect 33740 37996 34244 37998
rect 32732 37884 32844 37940
rect 32284 37772 32676 37828
rect 32788 37882 32844 37884
rect 32788 37830 32790 37882
rect 32842 37830 32844 37882
rect 32788 37818 32844 37830
rect 32172 37268 32228 37278
rect 32172 37174 32228 37212
rect 32060 36988 32228 37044
rect 31724 36764 31984 36820
rect 30828 36642 30884 36652
rect 31500 36708 31556 36718
rect 31500 36452 31556 36652
rect 31500 36400 31502 36452
rect 31554 36400 31556 36452
rect 31500 36388 31556 36400
rect 31724 36426 31780 36764
rect 32004 36596 32060 36606
rect 32004 36538 32060 36540
rect 31724 36374 31726 36426
rect 31778 36374 31780 36426
rect 31108 36258 31164 36270
rect 31108 36206 31110 36258
rect 31162 36206 31164 36258
rect 31108 36036 31164 36206
rect 31108 35970 31164 35980
rect 30492 35644 30660 35700
rect 30716 35812 30772 35822
rect 30716 35698 30772 35756
rect 30716 35646 30718 35698
rect 30770 35646 30772 35698
rect 30492 35364 30548 35644
rect 30716 35634 30772 35646
rect 31592 35698 31648 35710
rect 31592 35646 31594 35698
rect 31646 35646 31648 35698
rect 31592 35364 31648 35646
rect 31724 35476 31780 36374
rect 31836 36484 31892 36494
rect 32004 36486 32006 36538
rect 32058 36486 32060 36538
rect 32004 36474 32060 36486
rect 31836 35810 31892 36428
rect 31836 35758 31838 35810
rect 31890 35758 31892 35810
rect 31836 35746 31892 35758
rect 31724 35410 31780 35420
rect 30492 35308 30660 35364
rect 30268 35086 30270 35138
rect 30322 35086 30324 35138
rect 30268 35074 30324 35086
rect 30492 35140 30548 35150
rect 30324 34244 30380 34254
rect 30492 34244 30548 35084
rect 30324 34242 30548 34244
rect 30324 34190 30326 34242
rect 30378 34190 30548 34242
rect 30324 34188 30548 34190
rect 30324 34178 30380 34188
rect 30604 34132 30660 35308
rect 31592 35298 31648 35308
rect 31780 34860 31836 34870
rect 31780 34858 31892 34860
rect 31556 34804 31612 34814
rect 31780 34806 31782 34858
rect 31834 34806 31892 34858
rect 31780 34794 31892 34806
rect 31108 34692 31164 34702
rect 31108 34598 31164 34636
rect 31556 34468 31612 34748
rect 31556 34402 31612 34412
rect 30492 34076 30660 34132
rect 30716 34132 30772 34170
rect 31592 34132 31648 34142
rect 30492 33796 30548 34076
rect 30716 34066 30772 34076
rect 31388 34130 31648 34132
rect 31388 34078 31594 34130
rect 31646 34078 31648 34130
rect 31388 34076 31648 34078
rect 30492 33740 30772 33796
rect 30156 33730 30212 33740
rect 29484 33282 29540 33292
rect 29820 33124 29876 33628
rect 30044 33618 30100 33628
rect 30044 33348 30100 33358
rect 30044 33254 30100 33292
rect 29820 33058 29876 33068
rect 29372 32722 29428 32732
rect 30136 32788 30192 32798
rect 30136 32618 30192 32732
rect 30136 32566 30138 32618
rect 30190 32566 30192 32618
rect 30380 32676 30436 32686
rect 30380 32582 30436 32620
rect 30136 32554 30192 32566
rect 29260 32498 29316 32508
rect 29036 31938 29092 31948
rect 29148 32228 29204 32238
rect 29036 31780 29092 31790
rect 29036 31686 29092 31724
rect 29148 31108 29204 32172
rect 29540 32004 29596 32014
rect 29540 31910 29596 31948
rect 29260 31778 29316 31790
rect 29260 31726 29262 31778
rect 29314 31726 29316 31778
rect 29260 31668 29316 31726
rect 29260 31602 29316 31612
rect 30212 31722 30268 31734
rect 30212 31670 30214 31722
rect 30266 31670 30268 31722
rect 30212 31556 30268 31670
rect 30436 31724 30492 31734
rect 30436 31722 30548 31724
rect 30436 31670 30438 31722
rect 30490 31670 30548 31722
rect 30436 31658 30548 31670
rect 30212 31490 30268 31500
rect 28364 30968 28420 30980
rect 28028 30930 28084 30942
rect 28700 30940 28980 30996
rect 29036 31052 29204 31108
rect 29596 31332 29652 31342
rect 27916 30326 27918 30378
rect 27970 30326 27972 30378
rect 27916 30314 27972 30326
rect 28028 30772 28084 30782
rect 27916 30210 27972 30222
rect 27916 30158 27918 30210
rect 27970 30158 27972 30210
rect 27916 30100 27972 30158
rect 27916 30034 27972 30044
rect 27412 29820 27636 29876
rect 27020 29708 27412 29764
rect 27188 29428 27244 29438
rect 27188 29334 27244 29372
rect 26740 29314 26796 29326
rect 26740 29262 26742 29314
rect 26794 29262 26796 29314
rect 26740 29204 26796 29262
rect 27356 29314 27412 29708
rect 27580 29652 27636 29820
rect 27580 29586 27636 29596
rect 27356 29262 27358 29314
rect 27410 29262 27412 29314
rect 27356 29250 27412 29262
rect 27580 29426 27636 29438
rect 27580 29374 27582 29426
rect 27634 29374 27636 29426
rect 26740 29138 26796 29148
rect 26572 28700 26740 28756
rect 26328 28586 26384 28598
rect 26328 28534 26330 28586
rect 26382 28534 26384 28586
rect 26328 28084 26384 28534
rect 26572 28532 26628 28570
rect 26572 28466 26628 28476
rect 26572 28308 26628 28318
rect 26328 28028 26516 28084
rect 26348 27860 26404 27870
rect 26348 27766 26404 27804
rect 26124 27694 26126 27746
rect 26178 27694 26180 27746
rect 26124 27682 26180 27694
rect 26460 27310 26516 28028
rect 26572 27858 26628 28252
rect 26572 27806 26574 27858
rect 26626 27806 26628 27858
rect 26572 27794 26628 27806
rect 26012 27244 26292 27300
rect 26460 27298 26572 27310
rect 26460 27246 26518 27298
rect 26570 27246 26572 27298
rect 26460 27244 26572 27246
rect 26012 26414 26068 27244
rect 26124 27074 26180 27086
rect 26124 27022 26126 27074
rect 26178 27022 26180 27074
rect 26124 26908 26180 27022
rect 26236 27076 26292 27244
rect 26516 27234 26572 27244
rect 26684 27076 26740 28700
rect 27300 28644 27356 28654
rect 27300 28550 27356 28588
rect 27580 28420 27636 29374
rect 27916 29428 27972 29438
rect 27748 29204 27804 29214
rect 27748 28754 27804 29148
rect 27748 28702 27750 28754
rect 27802 28702 27804 28754
rect 27748 28690 27804 28702
rect 27580 28354 27636 28364
rect 26852 27972 26908 27982
rect 26852 27878 26908 27916
rect 27020 27860 27076 27870
rect 26236 27020 26740 27076
rect 26796 27074 26852 27086
rect 26796 27022 26798 27074
rect 26850 27022 26852 27074
rect 26796 26908 26852 27022
rect 27020 27074 27076 27804
rect 27468 27860 27524 27870
rect 27636 27860 27692 27870
rect 27468 27858 27580 27860
rect 27468 27806 27470 27858
rect 27522 27806 27580 27858
rect 27468 27794 27580 27806
rect 27524 27298 27580 27794
rect 27524 27246 27526 27298
rect 27578 27246 27580 27298
rect 27524 27234 27580 27246
rect 27636 27076 27692 27804
rect 27804 27860 27860 27870
rect 27804 27766 27860 27804
rect 27916 27860 27972 29372
rect 28028 28878 28084 30716
rect 28252 30212 28308 30222
rect 28252 30118 28308 30156
rect 28252 29426 28308 29438
rect 28252 29374 28254 29426
rect 28306 29374 28308 29426
rect 28028 28866 28140 28878
rect 28028 28814 28086 28866
rect 28138 28814 28140 28866
rect 28028 28812 28140 28814
rect 28084 28802 28140 28812
rect 28252 27972 28308 29374
rect 28588 29426 28644 29438
rect 28588 29374 28590 29426
rect 28642 29374 28644 29426
rect 28252 27906 28308 27916
rect 28364 28642 28420 28654
rect 28364 28590 28366 28642
rect 28418 28590 28420 28642
rect 27916 27858 28084 27860
rect 27916 27806 27918 27858
rect 27970 27806 28084 27858
rect 27916 27804 28084 27806
rect 27916 27794 27972 27804
rect 27020 27022 27022 27074
rect 27074 27022 27076 27074
rect 27020 27010 27076 27022
rect 27580 27020 27692 27076
rect 27804 27300 27860 27310
rect 27804 27076 27860 27244
rect 26124 26852 26516 26908
rect 26012 26402 26124 26414
rect 26012 26350 26070 26402
rect 26122 26350 26124 26402
rect 26012 26348 26124 26350
rect 26068 26338 26124 26348
rect 26460 26292 26516 26852
rect 26460 26122 26516 26236
rect 26572 26852 26852 26908
rect 26572 26404 26628 26852
rect 27468 26516 27524 26526
rect 27580 26516 27636 27020
rect 27804 26982 27860 27020
rect 27916 27074 27972 27086
rect 27916 27022 27918 27074
rect 27970 27022 27972 27074
rect 27468 26514 27636 26516
rect 27468 26462 27470 26514
rect 27522 26462 27636 26514
rect 27468 26460 27636 26462
rect 27468 26450 27524 26460
rect 26572 26290 26628 26348
rect 26572 26238 26574 26290
rect 26626 26238 26628 26290
rect 26572 26226 26628 26238
rect 26908 26292 26964 26302
rect 26908 26198 26964 26236
rect 27132 26290 27188 26302
rect 27132 26238 27134 26290
rect 27186 26238 27188 26290
rect 26460 26070 26462 26122
rect 26514 26070 26516 26122
rect 26460 26058 26516 26070
rect 26796 26068 26852 26078
rect 26348 25956 26404 25966
rect 25900 24770 25956 24780
rect 26236 25172 26292 25182
rect 25788 24714 25844 24726
rect 25676 24614 25678 24666
rect 25730 24614 25732 24666
rect 25676 24612 25732 24614
rect 25452 24556 25732 24612
rect 25004 24322 25060 24332
rect 25452 23268 25508 24556
rect 26124 24500 26180 24510
rect 26236 24500 26292 25116
rect 26348 24834 26404 25900
rect 26796 25730 26852 26012
rect 26796 25678 26798 25730
rect 26850 25678 26852 25730
rect 26796 25666 26852 25678
rect 26348 24782 26350 24834
rect 26402 24782 26404 24834
rect 26348 24770 26404 24782
rect 26516 24948 26572 24958
rect 26516 24724 26572 24892
rect 27132 24948 27188 26238
rect 27916 25844 27972 27022
rect 28028 26908 28084 27804
rect 28196 27748 28252 27758
rect 28196 27654 28252 27692
rect 28364 27524 28420 28590
rect 28364 27458 28420 27468
rect 28476 28642 28532 28654
rect 28476 28590 28478 28642
rect 28530 28590 28532 28642
rect 28476 28420 28532 28590
rect 28364 27300 28420 27310
rect 28476 27300 28532 28364
rect 28364 27298 28532 27300
rect 28364 27246 28366 27298
rect 28418 27246 28532 27298
rect 28364 27244 28532 27246
rect 28588 28532 28644 29374
rect 28364 27234 28420 27244
rect 28588 26908 28644 28476
rect 28700 27636 28756 30940
rect 29036 30324 29092 31052
rect 29372 30996 29428 31006
rect 29372 30902 29428 30940
rect 29596 30994 29652 31276
rect 29596 30942 29598 30994
rect 29650 30942 29652 30994
rect 29596 30930 29652 30942
rect 30268 31332 30324 31342
rect 29204 30884 29260 30894
rect 29204 30826 29260 30828
rect 29204 30774 29206 30826
rect 29258 30774 29260 30826
rect 29204 30762 29260 30774
rect 29540 30660 29596 30670
rect 29540 30434 29596 30604
rect 29540 30382 29542 30434
rect 29594 30382 29596 30434
rect 29540 30370 29596 30382
rect 29708 30436 29764 30446
rect 28812 30268 29092 30324
rect 28812 28308 28868 30268
rect 29148 30212 29204 30222
rect 28812 28242 28868 28252
rect 28924 30100 28980 30110
rect 28812 27972 28868 27982
rect 28812 27858 28868 27916
rect 28812 27806 28814 27858
rect 28866 27806 28868 27858
rect 28812 27794 28868 27806
rect 28924 27636 28980 30044
rect 29148 29652 29204 30156
rect 29260 30210 29316 30222
rect 29260 30158 29262 30210
rect 29314 30158 29316 30210
rect 29260 30100 29316 30158
rect 29260 30034 29316 30044
rect 29148 29596 29316 29652
rect 29036 29461 29092 29473
rect 29036 29409 29038 29461
rect 29090 29409 29092 29461
rect 29036 28420 29092 29409
rect 29148 29454 29204 29466
rect 29148 29428 29150 29454
rect 29202 29428 29204 29454
rect 29148 29362 29204 29372
rect 29148 28868 29204 28878
rect 29148 28810 29204 28812
rect 29148 28758 29150 28810
rect 29202 28758 29204 28810
rect 29148 28746 29204 28758
rect 29260 28642 29316 29596
rect 29708 29540 29764 30380
rect 30156 30212 30212 30222
rect 30268 30212 30324 31276
rect 30492 31062 30548 31658
rect 30472 31050 30548 31062
rect 30472 30998 30474 31050
rect 30526 30998 30548 31050
rect 30604 31722 30660 31734
rect 30604 31670 30606 31722
rect 30658 31670 30660 31722
rect 30604 31108 30660 31670
rect 30716 31556 30772 33740
rect 31052 33684 31108 33694
rect 31388 33684 31444 34076
rect 31592 34066 31648 34076
rect 31836 34132 31892 34794
rect 31836 34038 31892 34076
rect 31948 34858 32004 34870
rect 31948 34806 31950 34858
rect 32002 34806 32004 34858
rect 31948 34244 32004 34806
rect 31948 33908 32004 34188
rect 31724 33852 32004 33908
rect 32060 34692 32116 34702
rect 31724 33796 31780 33852
rect 30920 33460 30976 33470
rect 30920 33348 30976 33404
rect 30920 33346 30996 33348
rect 30920 33294 30922 33346
rect 30974 33294 30996 33346
rect 30920 33282 30996 33294
rect 30828 33124 30884 33134
rect 30828 32394 30884 33068
rect 30940 32562 30996 33282
rect 30940 32510 30942 32562
rect 30994 32510 30996 32562
rect 30940 32498 30996 32510
rect 30828 32342 30830 32394
rect 30882 32342 30884 32394
rect 30828 32330 30884 32342
rect 31052 32228 31108 33628
rect 31164 33628 31444 33684
rect 31612 33740 31780 33796
rect 31164 33570 31220 33628
rect 31164 33518 31166 33570
rect 31218 33518 31220 33570
rect 31164 33506 31220 33518
rect 31164 33348 31220 33358
rect 31164 32562 31220 33292
rect 31500 33348 31556 33358
rect 31500 33254 31556 33292
rect 31164 32510 31166 32562
rect 31218 32510 31220 32562
rect 31164 32498 31220 32510
rect 30716 31490 30772 31500
rect 30828 32172 31108 32228
rect 30604 31042 30660 31052
rect 30472 30986 30548 30998
rect 30492 30772 30548 30986
rect 30716 30996 30772 31006
rect 30716 30902 30772 30940
rect 30828 30772 30884 32172
rect 31164 32004 31220 32014
rect 31612 32004 31668 33740
rect 31836 33684 31892 33694
rect 31724 33460 31780 33470
rect 31724 33346 31780 33404
rect 31724 33294 31726 33346
rect 31778 33294 31780 33346
rect 31724 33282 31780 33294
rect 31836 33012 31892 33628
rect 31948 33572 32004 33582
rect 31948 33246 32004 33516
rect 32060 33460 32116 34636
rect 32172 33796 32228 36988
rect 32284 36706 32340 37772
rect 32956 37716 33012 37996
rect 34188 37986 34244 37996
rect 34860 38050 34916 38108
rect 34860 37998 34862 38050
rect 34914 37998 34916 38050
rect 34860 37986 34916 37998
rect 34972 38050 35028 38062
rect 34972 37998 34974 38050
rect 35026 37998 35028 38050
rect 32844 37660 33012 37716
rect 33460 37826 33516 37838
rect 33460 37774 33462 37826
rect 33514 37774 33516 37826
rect 32284 36654 32286 36706
rect 32338 36654 32340 36706
rect 32284 36642 32340 36654
rect 32396 37604 32452 37614
rect 32396 37156 32452 37548
rect 32396 36372 32452 37100
rect 32732 37380 32788 37390
rect 32732 36596 32788 37324
rect 32844 37156 32900 37660
rect 33460 37604 33516 37774
rect 33852 37828 33908 37838
rect 33852 37734 33908 37772
rect 33460 37538 33516 37548
rect 34972 37390 35028 37998
rect 35084 37604 35140 38612
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35308 38276 35364 38286
rect 35532 38276 35588 38612
rect 35308 38274 35588 38276
rect 35308 38222 35310 38274
rect 35362 38222 35588 38274
rect 35308 38220 35588 38222
rect 35644 38276 35700 38286
rect 35308 38210 35364 38220
rect 35644 38050 35700 38220
rect 35644 37998 35646 38050
rect 35698 37998 35700 38050
rect 35644 37986 35700 37998
rect 35084 37548 35252 37604
rect 33068 37380 33124 37390
rect 34972 37378 35084 37390
rect 34972 37326 35030 37378
rect 35082 37326 35084 37378
rect 34972 37324 35084 37326
rect 33068 37266 33124 37324
rect 35028 37314 35084 37324
rect 33068 37214 33070 37266
rect 33122 37214 33124 37266
rect 33068 37202 33124 37214
rect 33944 37268 34000 37278
rect 33944 37174 34000 37212
rect 34188 37268 34244 37278
rect 34188 37174 34244 37212
rect 34636 37266 34692 37278
rect 34636 37214 34638 37266
rect 34690 37214 34692 37266
rect 32844 36932 32900 37100
rect 32844 36876 33124 36932
rect 32844 36596 32900 36606
rect 32732 36540 32844 36596
rect 32844 36502 32900 36540
rect 32284 34858 32340 34870
rect 32284 34806 32286 34858
rect 32338 34806 32340 34858
rect 32284 34804 32340 34806
rect 32284 34738 32340 34748
rect 32284 34020 32340 34030
rect 32396 34020 32452 36316
rect 32564 36148 32620 36158
rect 32564 35922 32620 36092
rect 32564 35870 32566 35922
rect 32618 35870 32620 35922
rect 32564 35858 32620 35870
rect 33068 35924 33124 36876
rect 34300 36650 34356 36662
rect 34300 36598 34302 36650
rect 34354 36598 34356 36650
rect 34300 36596 34356 36598
rect 34300 36530 34356 36540
rect 34636 36596 34692 37214
rect 34636 36530 34692 36540
rect 34748 37266 34804 37278
rect 34748 37214 34750 37266
rect 34802 37214 34804 37266
rect 33404 36484 33460 36494
rect 33238 36426 33294 36438
rect 33238 36374 33240 36426
rect 33292 36374 33294 36426
rect 33404 36390 33460 36428
rect 33516 36484 33572 36494
rect 33852 36484 33908 36494
rect 33516 36482 33908 36484
rect 33516 36430 33518 36482
rect 33570 36430 33854 36482
rect 33906 36430 33908 36482
rect 33516 36428 33908 36430
rect 33238 36036 33294 36374
rect 33238 35980 33460 36036
rect 32732 35700 32788 35710
rect 32732 35138 32788 35644
rect 32732 35086 32734 35138
rect 32786 35086 32788 35138
rect 32732 35074 32788 35086
rect 33068 34916 33124 35868
rect 33404 35866 33460 35980
rect 33180 35812 33236 35822
rect 33404 35814 33406 35866
rect 33458 35814 33460 35866
rect 33404 35802 33460 35814
rect 33180 35698 33236 35756
rect 33180 35646 33182 35698
rect 33234 35646 33236 35698
rect 33180 35634 33236 35646
rect 33516 35700 33572 36428
rect 33852 36418 33908 36428
rect 34188 36484 34244 36494
rect 33516 35634 33572 35644
rect 33852 35698 33908 35710
rect 33852 35646 33854 35698
rect 33906 35646 33908 35698
rect 33852 35364 33908 35646
rect 34076 35700 34132 35710
rect 34188 35700 34244 36428
rect 34580 36260 34636 36270
rect 34580 35810 34636 36204
rect 34748 36260 34804 37214
rect 35196 37044 35252 37548
rect 35644 37492 35700 37502
rect 35644 37398 35700 37436
rect 35308 37268 35364 37278
rect 35308 37174 35364 37212
rect 35084 36988 35252 37044
rect 34916 36372 34972 36382
rect 34916 36278 34972 36316
rect 34748 36194 34804 36204
rect 34580 35758 34582 35810
rect 34634 35758 34636 35810
rect 34580 35746 34636 35758
rect 34300 35700 34356 35710
rect 34188 35698 34356 35700
rect 34188 35646 34302 35698
rect 34354 35646 34356 35698
rect 34188 35644 34356 35646
rect 34076 35606 34132 35644
rect 34300 35634 34356 35644
rect 33852 35298 33908 35308
rect 32844 34914 33124 34916
rect 32844 34862 33070 34914
rect 33122 34862 33124 34914
rect 32844 34860 33124 34862
rect 32732 34804 32788 34814
rect 32564 34020 32620 34030
rect 32396 34018 32620 34020
rect 32396 33966 32566 34018
rect 32618 33966 32620 34018
rect 32396 33964 32620 33966
rect 32284 33908 32340 33964
rect 32284 33852 32508 33908
rect 32172 33730 32228 33740
rect 32452 33514 32508 33852
rect 32564 33684 32620 33964
rect 32564 33618 32620 33628
rect 32452 33462 32454 33514
rect 32506 33462 32508 33514
rect 32060 33404 32172 33460
rect 32452 33450 32508 33462
rect 31948 33234 32060 33246
rect 31948 33182 32006 33234
rect 32058 33182 32060 33234
rect 31948 33180 32060 33182
rect 32004 33170 32060 33180
rect 31164 32002 31668 32004
rect 31164 31950 31166 32002
rect 31218 31950 31668 32002
rect 31164 31948 31668 31950
rect 31724 32956 31892 33012
rect 31164 31938 31220 31948
rect 30492 30706 30548 30716
rect 30716 30716 30884 30772
rect 30940 31780 30996 31790
rect 30604 30378 30660 30390
rect 30156 30210 30324 30212
rect 30156 30158 30158 30210
rect 30210 30158 30324 30210
rect 30156 30156 30324 30158
rect 30492 30324 30548 30334
rect 30492 30210 30548 30268
rect 30492 30158 30494 30210
rect 30546 30158 30548 30210
rect 29876 29540 29932 29550
rect 29708 29538 29932 29540
rect 29708 29486 29878 29538
rect 29930 29486 29932 29538
rect 29708 29484 29932 29486
rect 29876 29474 29932 29484
rect 29260 28590 29262 28642
rect 29314 28590 29316 28642
rect 29092 28364 29204 28420
rect 29036 28354 29092 28364
rect 28700 27580 28868 27636
rect 28028 26852 28196 26908
rect 28028 26292 28084 26302
rect 28028 26198 28084 26236
rect 27132 24882 27188 24892
rect 27580 25788 27972 25844
rect 26908 24836 26964 24846
rect 26684 24780 26908 24836
rect 26572 24668 26628 24724
rect 26516 24630 26628 24668
rect 26236 24444 26516 24500
rect 26124 24388 26180 24444
rect 26124 24332 26292 24388
rect 26120 24164 26176 24174
rect 26120 23900 26176 24108
rect 26120 23848 26122 23900
rect 26174 23848 26176 23900
rect 25452 23202 25508 23212
rect 25564 23826 25620 23838
rect 26120 23836 26176 23848
rect 25564 23774 25566 23826
rect 25618 23774 25620 23826
rect 24892 22754 24948 22764
rect 25004 23156 25060 23166
rect 25004 22596 25060 23100
rect 25564 23156 25620 23774
rect 25788 23268 25844 23278
rect 25788 23174 25844 23212
rect 25564 23090 25620 23100
rect 26124 23156 26180 23166
rect 26124 23062 26180 23100
rect 26236 22932 26292 24332
rect 26460 23378 26516 24444
rect 26572 24106 26628 24630
rect 26572 24054 26574 24106
rect 26626 24054 26628 24106
rect 26684 24164 26740 24780
rect 26908 24770 26964 24780
rect 26684 24098 26740 24108
rect 27020 24724 27076 24734
rect 26572 24042 26628 24054
rect 26796 23940 26852 23950
rect 26796 23846 26852 23884
rect 26460 23326 26462 23378
rect 26514 23326 26516 23378
rect 26460 23314 26516 23326
rect 27020 23268 27076 24668
rect 27468 24724 27524 24734
rect 27468 24630 27524 24668
rect 27580 24612 27636 25788
rect 27580 24546 27636 24556
rect 27692 25676 28084 25732
rect 27692 24276 27748 25676
rect 28028 25674 28084 25676
rect 28028 25622 28030 25674
rect 28082 25622 28084 25674
rect 28028 25610 28084 25622
rect 27916 25506 27972 25518
rect 28140 25508 28196 26852
rect 28476 26852 28644 26908
rect 28700 27074 28756 27086
rect 28700 27022 28702 27074
rect 28754 27022 28756 27074
rect 28364 26290 28420 26302
rect 28364 26238 28366 26290
rect 28418 26238 28420 26290
rect 27916 25454 27918 25506
rect 27970 25454 27972 25506
rect 27804 25172 27860 25182
rect 27804 24722 27860 25116
rect 27916 25060 27972 25454
rect 27916 24994 27972 25004
rect 28028 25452 28196 25508
rect 28252 25506 28308 25518
rect 28252 25454 28254 25506
rect 28306 25454 28308 25506
rect 27804 24670 27806 24722
rect 27858 24670 27860 24722
rect 27804 24658 27860 24670
rect 28028 24610 28084 25452
rect 28252 25172 28308 25454
rect 28364 25508 28420 26238
rect 28476 26122 28532 26852
rect 28476 26070 28478 26122
rect 28530 26070 28532 26122
rect 28476 26058 28532 26070
rect 28700 25956 28756 27022
rect 28700 25890 28756 25900
rect 28812 25732 28868 27580
rect 28924 27570 28980 27580
rect 29036 27897 29092 27909
rect 29036 27860 29038 27897
rect 29090 27860 29092 27897
rect 29036 26852 29092 27804
rect 29148 27039 29204 28364
rect 29260 27746 29316 28590
rect 29372 29454 29428 29466
rect 29372 29402 29374 29454
rect 29426 29402 29428 29454
rect 29372 28084 29428 29402
rect 29596 29454 29652 29466
rect 29596 29402 29598 29454
rect 29650 29402 29652 29454
rect 29596 28868 29652 29402
rect 30044 29092 30100 29102
rect 30156 29092 30212 30156
rect 30492 30146 30548 30158
rect 30604 30326 30606 30378
rect 30658 30326 30660 30378
rect 30604 30212 30660 30326
rect 30604 30146 30660 30156
rect 30548 29764 30604 29774
rect 30548 29650 30604 29708
rect 30548 29598 30550 29650
rect 30602 29598 30604 29650
rect 30548 29586 30604 29598
rect 30716 29428 30772 30716
rect 30940 30378 30996 31724
rect 31612 31778 31668 31790
rect 31612 31726 31614 31778
rect 31666 31726 31668 31778
rect 31612 31332 31668 31726
rect 31724 31556 31780 32956
rect 32116 32452 32172 33404
rect 32732 33348 32788 34748
rect 32284 33290 32340 33302
rect 32284 33238 32286 33290
rect 32338 33238 32340 33290
rect 32732 33282 32788 33292
rect 32284 32676 32340 33238
rect 32844 33124 32900 34860
rect 33068 34850 33124 34860
rect 33852 34914 33908 34926
rect 33852 34862 33854 34914
rect 33906 34862 33908 34914
rect 33852 34356 33908 34862
rect 35084 34356 35140 36988
rect 35644 36932 35700 36942
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 36708 35252 36718
rect 35196 36482 35252 36652
rect 35196 36430 35198 36482
rect 35250 36430 35252 36482
rect 35364 36596 35420 36606
rect 35364 36538 35420 36540
rect 35364 36486 35366 36538
rect 35418 36486 35420 36538
rect 35364 36474 35420 36486
rect 35644 36482 35700 36876
rect 35196 36418 35252 36430
rect 35644 36430 35646 36482
rect 35698 36430 35700 36482
rect 35644 36418 35700 36430
rect 35532 36370 35588 36382
rect 35532 36318 35534 36370
rect 35586 36318 35588 36370
rect 35532 36260 35588 36318
rect 35532 36194 35588 36204
rect 35420 35812 35476 35822
rect 35756 35812 35812 38668
rect 36204 38612 36820 38668
rect 36988 38668 37044 38892
rect 36988 38612 37100 38668
rect 37044 38610 37100 38612
rect 37044 38558 37046 38610
rect 37098 38558 37100 38610
rect 37044 38546 37100 38558
rect 35980 38388 36036 38398
rect 35980 38274 36036 38332
rect 35980 38222 35982 38274
rect 36034 38222 36036 38274
rect 35980 38210 36036 38222
rect 36988 38276 37044 38286
rect 36988 37828 37044 38220
rect 37212 37940 37268 39116
rect 37436 38668 37492 39564
rect 37996 39284 38052 41132
rect 38108 41094 38164 41132
rect 37772 39228 38052 39284
rect 38108 40628 38164 40638
rect 37604 39060 37660 39070
rect 37604 38966 37660 39004
rect 37772 38668 37828 39228
rect 38108 39060 38164 40572
rect 38220 40180 38276 41468
rect 38332 40628 38388 41468
rect 38668 40964 38724 43652
rect 38799 43540 38855 44044
rect 38780 43538 38855 43540
rect 38780 43486 38801 43538
rect 38853 43486 38855 43538
rect 38780 43474 38855 43486
rect 38780 41188 38836 43474
rect 39004 43428 39060 44716
rect 39676 44548 39732 49200
rect 40796 46116 40852 46126
rect 40796 46022 40852 46060
rect 41132 45892 41188 45902
rect 39788 45862 39844 45874
rect 39788 45810 39790 45862
rect 39842 45810 39844 45862
rect 39788 45556 39844 45810
rect 39788 45490 39844 45500
rect 40460 45780 40516 45790
rect 40236 44996 40292 45006
rect 40348 44996 40404 45006
rect 40236 44994 40348 44996
rect 40236 44942 40238 44994
rect 40290 44942 40348 44994
rect 40236 44940 40348 44942
rect 40236 44930 40292 44940
rect 39676 44482 39732 44492
rect 39900 44294 39956 44306
rect 39900 44242 39902 44294
rect 39954 44242 39956 44294
rect 39900 44100 39956 44242
rect 39900 44034 39956 44044
rect 39676 43652 40180 43708
rect 39676 43538 39732 43652
rect 39676 43486 39678 43538
rect 39730 43486 39732 43538
rect 39676 43474 39732 43486
rect 39900 43538 39956 43550
rect 39900 43486 39902 43538
rect 39954 43486 39956 43538
rect 38892 43372 39060 43428
rect 38892 42532 38948 43372
rect 38892 42476 39172 42532
rect 39116 42026 39172 42476
rect 39116 41974 39118 42026
rect 39170 41974 39172 42026
rect 39116 41962 39172 41974
rect 39228 42420 39284 42430
rect 39228 41860 39284 42364
rect 39900 42308 39956 43486
rect 39564 42252 39956 42308
rect 40012 42754 40068 42766
rect 40012 42702 40014 42754
rect 40066 42702 40068 42754
rect 39452 42084 39508 42094
rect 39452 41970 39508 42028
rect 39452 41918 39454 41970
rect 39506 41918 39508 41970
rect 39452 41906 39508 41918
rect 39228 41636 39284 41804
rect 39228 41570 39284 41580
rect 39564 41524 39620 42252
rect 40012 42084 40068 42702
rect 40124 42206 40180 43652
rect 40236 43314 40292 43326
rect 40236 43262 40238 43314
rect 40290 43262 40292 43314
rect 40236 43204 40292 43262
rect 40236 42420 40292 43148
rect 40236 42354 40292 42364
rect 40124 42194 40236 42206
rect 40124 42142 40182 42194
rect 40234 42142 40236 42194
rect 40124 42140 40236 42142
rect 40180 42130 40236 42140
rect 40012 42018 40068 42028
rect 40348 41970 40404 44940
rect 39844 41914 39900 41926
rect 39676 41858 39732 41870
rect 39676 41806 39678 41858
rect 39730 41806 39732 41858
rect 39676 41524 39732 41806
rect 39844 41862 39846 41914
rect 39898 41862 39900 41914
rect 40348 41918 40350 41970
rect 40402 41918 40404 41970
rect 40348 41906 40404 41918
rect 39844 41860 39900 41862
rect 39844 41794 39900 41804
rect 39676 41468 40292 41524
rect 39564 41458 39620 41468
rect 38780 41122 38836 41132
rect 38892 41188 38948 41198
rect 38892 41186 39172 41188
rect 38892 41134 38894 41186
rect 38946 41134 39172 41186
rect 38892 41132 39172 41134
rect 38892 41122 38948 41132
rect 38668 40908 39060 40964
rect 38332 40562 38388 40572
rect 38332 40404 38388 40414
rect 38332 40310 38388 40348
rect 38444 40404 38500 40414
rect 38444 40402 38612 40404
rect 38444 40350 38446 40402
rect 38498 40350 38612 40402
rect 38444 40348 38612 40350
rect 38444 40338 38500 40348
rect 38220 40114 38276 40124
rect 38220 39620 38276 39630
rect 38220 39526 38276 39564
rect 38108 38994 38164 39004
rect 38444 39508 38500 39518
rect 37212 37874 37268 37884
rect 37324 38612 37492 38668
rect 37548 38612 37828 38668
rect 37884 38948 37940 38958
rect 37884 38834 37940 38892
rect 38332 38948 38388 38958
rect 38142 38871 38198 38883
rect 37884 38782 37886 38834
rect 37938 38782 37940 38834
rect 36988 37762 37044 37772
rect 37100 37826 37156 37838
rect 37100 37774 37102 37826
rect 37154 37774 37156 37826
rect 37100 37492 37156 37774
rect 37324 37828 37380 38612
rect 37436 38052 37492 38062
rect 37548 38052 37604 38612
rect 37884 38388 37940 38782
rect 37996 38834 38052 38846
rect 37996 38782 37998 38834
rect 38050 38782 38052 38834
rect 37996 38724 38052 38782
rect 38142 38819 38144 38871
rect 38196 38819 38198 38871
rect 38142 38668 38198 38819
rect 37996 38658 38052 38668
rect 38108 38612 38198 38668
rect 38108 38500 38164 38612
rect 38332 38500 38388 38892
rect 38108 38434 38164 38444
rect 38220 38444 38388 38500
rect 37884 38322 37940 38332
rect 38220 38276 38276 38444
rect 38108 38220 38276 38276
rect 38444 38276 38500 39452
rect 38556 38722 38612 40348
rect 38724 40180 38780 40190
rect 38724 40178 38948 40180
rect 38724 40126 38726 40178
rect 38778 40126 38948 40178
rect 38724 40124 38948 40126
rect 38724 40114 38780 40124
rect 38892 39172 38948 40124
rect 39004 39956 39060 40908
rect 39116 40404 39172 41132
rect 39452 40516 39508 40526
rect 39116 40348 39396 40404
rect 39172 40180 39228 40190
rect 39004 39890 39060 39900
rect 39116 40178 39228 40180
rect 39116 40126 39174 40178
rect 39226 40126 39228 40178
rect 39116 40114 39228 40126
rect 38892 39106 38948 39116
rect 39004 39618 39060 39630
rect 39004 39566 39006 39618
rect 39058 39566 39060 39618
rect 39004 39060 39060 39566
rect 39004 38994 39060 39004
rect 38556 38670 38558 38722
rect 38610 38670 38612 38722
rect 38556 38658 38612 38670
rect 38892 38834 38948 38846
rect 38892 38782 38894 38834
rect 38946 38782 38948 38834
rect 37548 37996 37610 38052
rect 37436 37958 37492 37996
rect 37554 37828 37610 37996
rect 37996 38050 38052 38062
rect 37996 37998 37998 38050
rect 38050 37998 38052 38050
rect 37324 37772 37492 37828
rect 36876 37436 37156 37492
rect 37324 37492 37380 37502
rect 36260 37156 36316 37166
rect 36260 37062 36316 37100
rect 36652 37156 36708 37166
rect 36652 37062 36708 37100
rect 36876 37044 36932 37436
rect 37046 37268 37102 37278
rect 37046 37174 37102 37212
rect 37212 37266 37268 37278
rect 37212 37214 37214 37266
rect 37266 37214 37268 37266
rect 37212 37044 37268 37214
rect 37324 37266 37380 37436
rect 37324 37214 37326 37266
rect 37378 37214 37380 37266
rect 37324 37202 37380 37214
rect 36876 36988 37044 37044
rect 36876 36482 36932 36494
rect 36876 36430 36878 36482
rect 36930 36430 36932 36482
rect 35924 36370 35980 36382
rect 35924 36318 35926 36370
rect 35978 36318 35980 36370
rect 35924 35924 35980 36318
rect 36876 36372 36932 36430
rect 36876 36306 36932 36316
rect 36484 36260 36540 36270
rect 36484 36258 36596 36260
rect 36484 36206 36486 36258
rect 36538 36206 36596 36258
rect 36484 36194 36596 36206
rect 35924 35858 35980 35868
rect 35420 35810 35812 35812
rect 35420 35758 35422 35810
rect 35474 35758 35812 35810
rect 35420 35756 35812 35758
rect 35420 35746 35476 35756
rect 36372 35754 36428 35766
rect 35868 35728 35924 35740
rect 35868 35676 35870 35728
rect 35922 35676 35924 35728
rect 35644 35588 35700 35598
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 33852 34290 33908 34300
rect 34412 34300 35140 34356
rect 33964 34244 34020 34254
rect 33944 34188 33964 34244
rect 33944 34186 34020 34188
rect 33068 34132 33124 34170
rect 33944 34134 33946 34186
rect 33998 34178 34020 34186
rect 33998 34134 34000 34178
rect 33944 34122 34000 34134
rect 33068 34066 33124 34076
rect 34300 34020 34356 34030
rect 34188 33908 34244 33918
rect 33944 33906 34244 33908
rect 33944 33854 34190 33906
rect 34242 33854 34244 33906
rect 33944 33852 34244 33854
rect 32564 33068 32900 33124
rect 32564 32786 32620 33068
rect 32564 32734 32566 32786
rect 32618 32734 32620 32786
rect 32564 32722 32620 32734
rect 32844 32788 32900 33068
rect 32844 32722 32900 32732
rect 33068 33348 33124 33358
rect 32284 32610 32340 32620
rect 33068 32564 33124 33292
rect 33944 33346 34000 33852
rect 34188 33842 34244 33852
rect 34188 33572 34244 33582
rect 34300 33572 34356 33964
rect 34188 33570 34356 33572
rect 34188 33518 34190 33570
rect 34242 33518 34356 33570
rect 34188 33516 34356 33518
rect 34188 33506 34244 33516
rect 33944 33294 33946 33346
rect 33998 33294 34000 33346
rect 33944 33282 34000 33294
rect 33740 33236 33796 33246
rect 33404 33012 33460 33022
rect 32732 32508 33124 32564
rect 33180 32900 33236 32910
rect 33180 32674 33236 32844
rect 33180 32622 33182 32674
rect 33234 32622 33236 32674
rect 32116 32450 32452 32452
rect 32116 32398 32118 32450
rect 32170 32398 32452 32450
rect 32116 32396 32452 32398
rect 32116 32386 32172 32396
rect 31836 31780 31892 31790
rect 31836 31686 31892 31724
rect 32116 31666 32172 31678
rect 32116 31614 32118 31666
rect 32170 31614 32172 31666
rect 31724 31500 31892 31556
rect 31612 31266 31668 31276
rect 31164 31108 31220 31118
rect 31164 30994 31220 31052
rect 31164 30942 31166 30994
rect 31218 30942 31220 30994
rect 31164 30930 31220 30942
rect 30940 30326 30942 30378
rect 30994 30326 30996 30378
rect 30940 30324 30996 30326
rect 30940 30248 30996 30268
rect 31052 30210 31108 30222
rect 31052 30158 31054 30210
rect 31106 30158 31108 30210
rect 30100 29036 30212 29092
rect 30604 29372 30772 29428
rect 30828 30100 30884 30110
rect 30828 29764 30884 30044
rect 31052 29764 31108 30158
rect 31276 30210 31332 30222
rect 31276 30158 31278 30210
rect 31330 30158 31332 30210
rect 31276 30100 31332 30158
rect 31276 30034 31332 30044
rect 31052 29708 31760 29764
rect 30828 29426 30884 29708
rect 30828 29374 30830 29426
rect 30882 29374 30884 29426
rect 30044 29026 30100 29036
rect 30604 28980 30660 29372
rect 30828 29362 30884 29374
rect 31500 28980 31556 29708
rect 31704 29482 31760 29708
rect 31704 29430 31706 29482
rect 31758 29430 31760 29482
rect 31704 29418 31760 29430
rect 30604 28924 30996 28980
rect 29484 28812 29652 28868
rect 29484 28532 29540 28812
rect 29708 28756 29764 28766
rect 29484 28466 29540 28476
rect 29596 28642 29652 28654
rect 29596 28590 29598 28642
rect 29650 28590 29652 28642
rect 29596 28196 29652 28590
rect 29708 28644 29764 28700
rect 29932 28644 29988 28654
rect 29708 28642 29988 28644
rect 29708 28590 29934 28642
rect 29986 28590 29988 28642
rect 29708 28588 29988 28590
rect 29932 28578 29988 28588
rect 30604 28644 30660 28654
rect 30940 28644 30996 28924
rect 31052 28924 31556 28980
rect 31612 29316 31668 29326
rect 31836 29316 31892 31500
rect 32116 31220 32172 31614
rect 32116 31154 32172 31164
rect 32040 30994 32096 31006
rect 32284 30996 32340 31006
rect 32040 30942 32042 30994
rect 32094 30942 32096 30994
rect 32040 30884 32096 30942
rect 32040 30818 32096 30828
rect 32172 30940 32284 30996
rect 32172 30660 32228 30940
rect 32284 30902 32340 30940
rect 32396 30772 32452 32396
rect 32004 30604 32228 30660
rect 32284 30716 32452 30772
rect 32508 31668 32564 31678
rect 32004 30154 32060 30604
rect 32004 30102 32006 30154
rect 32058 30102 32060 30154
rect 32172 30212 32228 30222
rect 32172 30128 32174 30156
rect 32226 30128 32228 30156
rect 32172 30116 32228 30128
rect 32004 30090 32060 30102
rect 31948 29428 32004 29438
rect 31948 29334 32004 29372
rect 31052 28866 31108 28924
rect 31052 28814 31054 28866
rect 31106 28814 31108 28866
rect 31052 28802 31108 28814
rect 30044 28308 30100 28318
rect 29596 28140 29876 28196
rect 29372 28018 29428 28028
rect 29260 27694 29262 27746
rect 29314 27694 29316 27746
rect 29260 27682 29316 27694
rect 29372 27858 29428 27870
rect 29372 27806 29374 27858
rect 29426 27806 29428 27858
rect 29148 26987 29150 27039
rect 29202 26987 29204 27039
rect 29148 26975 29204 26987
rect 29260 27076 29316 27086
rect 29260 26994 29262 27020
rect 29314 26994 29316 27020
rect 29260 26982 29316 26994
rect 29036 26404 29092 26796
rect 28980 26348 29092 26404
rect 29148 26628 29204 26638
rect 29148 26458 29204 26572
rect 29148 26406 29150 26458
rect 29202 26406 29204 26458
rect 29148 26394 29204 26406
rect 28980 26346 29036 26348
rect 28980 26294 28982 26346
rect 29034 26294 29036 26346
rect 28980 26282 29036 26294
rect 29260 26292 29316 26302
rect 29372 26292 29428 27806
rect 29820 27690 29876 28140
rect 29596 27636 29652 27646
rect 29820 27638 29822 27690
rect 29874 27638 29876 27690
rect 29820 27626 29876 27638
rect 29932 27858 29988 27870
rect 29932 27806 29934 27858
rect 29986 27806 29988 27858
rect 29484 27018 29540 27030
rect 29484 26966 29486 27018
rect 29538 26966 29540 27018
rect 29484 26628 29540 26966
rect 29484 26562 29540 26572
rect 29260 26290 29428 26292
rect 29260 26238 29262 26290
rect 29314 26238 29428 26290
rect 29260 26236 29428 26238
rect 29260 26226 29316 26236
rect 28812 25666 28868 25676
rect 28364 25442 28420 25452
rect 29036 25506 29092 25518
rect 29036 25454 29038 25506
rect 29090 25454 29092 25506
rect 28252 25106 28308 25116
rect 29036 24836 29092 25454
rect 29036 24770 29092 24780
rect 29260 25508 29316 25518
rect 28028 24558 28030 24610
rect 28082 24558 28084 24610
rect 28028 24546 28084 24558
rect 28252 24722 28308 24734
rect 28252 24670 28254 24722
rect 28306 24670 28308 24722
rect 27692 24210 27748 24220
rect 27692 23938 27748 23950
rect 27692 23886 27694 23938
rect 27746 23886 27748 23938
rect 27692 23828 27748 23886
rect 27692 23762 27748 23772
rect 28252 23492 28308 24670
rect 28476 24724 28532 24734
rect 28476 24106 28532 24668
rect 29148 24722 29204 24734
rect 29148 24670 29150 24722
rect 29202 24670 29204 24722
rect 28868 24610 28924 24622
rect 28868 24558 28870 24610
rect 28922 24558 28924 24610
rect 28868 24388 28924 24558
rect 29148 24612 29204 24670
rect 29148 24546 29204 24556
rect 29260 24554 29316 25452
rect 29260 24502 29262 24554
rect 29314 24502 29316 24554
rect 29260 24490 29316 24502
rect 29372 24500 29428 26236
rect 29484 26292 29540 26302
rect 29484 26198 29540 26236
rect 29596 25742 29652 27580
rect 29820 27524 29876 27534
rect 29708 27188 29764 27198
rect 29708 27046 29764 27132
rect 29708 26994 29710 27046
rect 29762 26994 29764 27046
rect 29708 26982 29764 26994
rect 29540 25730 29652 25742
rect 29540 25678 29542 25730
rect 29594 25678 29652 25730
rect 29540 25676 29652 25678
rect 29708 26290 29764 26302
rect 29708 26238 29710 26290
rect 29762 26238 29764 26290
rect 29540 25666 29596 25676
rect 29708 25508 29764 26238
rect 29708 25442 29764 25452
rect 29820 26292 29876 27468
rect 29932 27300 29988 27806
rect 29932 27234 29988 27244
rect 30044 27086 30100 28252
rect 30604 28196 30660 28588
rect 30808 28586 30864 28598
rect 30940 28588 31108 28644
rect 30808 28534 30810 28586
rect 30862 28534 30864 28586
rect 30808 28308 30864 28534
rect 30808 28252 30996 28308
rect 30604 28140 30828 28196
rect 30772 28082 30828 28140
rect 30772 28030 30774 28082
rect 30826 28030 30828 28082
rect 30772 28018 30828 28030
rect 29988 27074 30100 27086
rect 29988 27022 29990 27074
rect 30042 27022 30100 27074
rect 29988 27020 30100 27022
rect 30156 27858 30212 27870
rect 30156 27806 30158 27858
rect 30210 27806 30212 27858
rect 29988 27010 30044 27020
rect 30156 26852 30212 27806
rect 30940 27858 30996 28252
rect 30940 27806 30942 27858
rect 30994 27806 30996 27858
rect 30940 27748 30996 27806
rect 30940 27682 30996 27692
rect 30492 27524 30548 27534
rect 30380 27242 30436 27254
rect 30380 27190 30382 27242
rect 30434 27190 30436 27242
rect 30380 27076 30436 27190
rect 30380 27010 30436 27020
rect 30492 27074 30548 27468
rect 30492 27022 30494 27074
rect 30546 27022 30548 27074
rect 30492 27010 30548 27022
rect 30716 27074 30772 27086
rect 30716 27022 30718 27074
rect 30770 27022 30772 27074
rect 29820 25284 29876 26236
rect 29988 26404 30044 26414
rect 29988 25508 30044 26348
rect 29988 25442 30044 25452
rect 30156 25396 30212 26796
rect 30716 26404 30772 27022
rect 31052 26628 31108 28588
rect 31612 28642 31668 29260
rect 31612 28590 31614 28642
rect 31666 28590 31668 28642
rect 31612 28578 31668 28590
rect 31724 29260 31892 29316
rect 31724 28644 31780 29260
rect 32284 29204 32340 30716
rect 32508 30436 32564 31612
rect 32732 30660 32788 32508
rect 32900 31780 32956 31790
rect 32900 31610 32956 31724
rect 33068 31780 33124 31790
rect 33180 31780 33236 32622
rect 33404 31902 33460 32956
rect 33740 32452 33796 33180
rect 34412 33012 34468 34300
rect 35644 34142 35700 35532
rect 35868 35252 35924 35676
rect 36092 35736 36148 35748
rect 36092 35684 36094 35736
rect 36146 35684 36148 35736
rect 36092 35588 36148 35684
rect 36092 35522 36148 35532
rect 36372 35702 36374 35754
rect 36426 35702 36428 35754
rect 36372 35252 36428 35702
rect 35868 35186 35924 35196
rect 36204 35196 36428 35252
rect 35756 34916 35812 34926
rect 36092 34916 36148 34926
rect 36204 34916 36260 35196
rect 36540 35028 36596 36194
rect 36540 34962 36596 34972
rect 36652 35698 36708 35710
rect 36652 35646 36654 35698
rect 36706 35646 36708 35698
rect 36652 34916 36708 35646
rect 36764 35698 36820 35710
rect 36988 35700 37044 36988
rect 36764 35646 36766 35698
rect 36818 35646 36820 35698
rect 36764 35028 36820 35646
rect 36876 35644 37044 35700
rect 37212 35700 37268 36988
rect 37436 36932 37492 37772
rect 37436 36866 37492 36876
rect 37548 37772 37610 37828
rect 37716 37938 37772 37950
rect 37716 37886 37718 37938
rect 37770 37886 37772 37938
rect 37716 37828 37772 37886
rect 37548 37266 37604 37772
rect 37716 37762 37772 37772
rect 37548 37214 37550 37266
rect 37602 37214 37604 37266
rect 37548 36596 37604 37214
rect 36876 35140 36932 35644
rect 37212 35634 37268 35644
rect 37324 36372 37380 36382
rect 37548 36372 37604 36540
rect 37884 37604 37940 37614
rect 37380 36316 37604 36372
rect 37660 36482 37716 36494
rect 37660 36430 37662 36482
rect 37714 36430 37716 36482
rect 37044 35476 37100 35486
rect 37044 35474 37268 35476
rect 37044 35422 37046 35474
rect 37098 35422 37268 35474
rect 37044 35420 37268 35422
rect 37044 35410 37100 35420
rect 36876 35074 36932 35084
rect 37100 35252 37156 35262
rect 36764 34962 36820 34972
rect 35756 34914 36260 34916
rect 35756 34862 35758 34914
rect 35810 34862 36094 34914
rect 36146 34862 36260 34914
rect 35756 34860 36260 34862
rect 35756 34850 35812 34860
rect 36092 34850 36148 34860
rect 36650 34804 36708 34916
rect 36988 34860 37044 34870
rect 36260 34692 36316 34702
rect 36260 34690 36596 34692
rect 36260 34638 36262 34690
rect 36314 34638 36596 34690
rect 36260 34636 36596 34638
rect 36260 34626 36316 34636
rect 33348 31890 33460 31902
rect 33348 31838 33350 31890
rect 33402 31838 33460 31890
rect 33348 31836 33460 31838
rect 33628 32396 33796 32452
rect 33852 32956 34468 33012
rect 34524 34130 34580 34142
rect 34524 34078 34526 34130
rect 34578 34078 34580 34130
rect 34524 33012 34580 34078
rect 34692 34132 34748 34142
rect 35644 34130 35719 34142
rect 35644 34078 35665 34130
rect 35717 34078 35719 34130
rect 35644 34076 35719 34078
rect 34692 33570 34748 34076
rect 35663 34020 35719 34076
rect 36540 34130 36596 34636
rect 36540 34078 36542 34130
rect 36594 34078 36596 34130
rect 36540 34066 36596 34078
rect 36652 34132 36708 34804
rect 36652 34066 36708 34076
rect 36876 34858 37044 34860
rect 36876 34806 36990 34858
rect 37042 34806 37044 34858
rect 36876 34804 37044 34806
rect 35663 33954 35719 33964
rect 34692 33518 34694 33570
rect 34746 33518 34748 33570
rect 34692 33506 34748 33518
rect 34860 33906 34916 33918
rect 34860 33854 34862 33906
rect 34914 33854 34916 33906
rect 34860 33124 34916 33854
rect 35420 33908 35476 33918
rect 35420 33906 35588 33908
rect 35420 33854 35422 33906
rect 35474 33854 35588 33906
rect 35420 33852 35588 33854
rect 35420 33842 35476 33852
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 33572 35252 33582
rect 34972 33348 35028 33358
rect 34972 33254 35028 33292
rect 35196 33346 35252 33516
rect 35532 33572 35588 33852
rect 35532 33506 35588 33516
rect 36316 33684 36372 33694
rect 35196 33294 35198 33346
rect 35250 33294 35252 33346
rect 36316 33348 36372 33628
rect 36876 33572 36932 34804
rect 36988 34794 37044 34804
rect 37100 34858 37156 35196
rect 37100 34806 37102 34858
rect 37154 34806 37156 34858
rect 36988 34356 37044 34366
rect 36988 34262 37044 34300
rect 36876 33506 36932 33516
rect 36988 34132 37044 34142
rect 36988 33358 37044 34076
rect 37100 33684 37156 34806
rect 37212 34132 37268 35420
rect 37324 34860 37380 36316
rect 37660 36036 37716 36430
rect 37660 35970 37716 35980
rect 37436 35700 37492 35710
rect 37436 35606 37492 35644
rect 37548 35698 37604 35710
rect 37548 35646 37550 35698
rect 37602 35646 37604 35698
rect 37548 35588 37604 35646
rect 37548 35522 37604 35532
rect 37716 35698 37772 35710
rect 37716 35646 37718 35698
rect 37770 35646 37772 35698
rect 37716 35252 37772 35646
rect 37884 35588 37940 37548
rect 37996 37156 38052 37998
rect 38108 38050 38164 38220
rect 38444 38210 38500 38220
rect 38556 38500 38612 38510
rect 38108 37998 38110 38050
rect 38162 37998 38164 38050
rect 38556 38052 38612 38444
rect 38108 37986 38164 37998
rect 38332 37994 38388 38006
rect 38332 37942 38334 37994
rect 38386 37942 38388 37994
rect 38556 37986 38612 37996
rect 38220 37828 38276 37838
rect 38332 37828 38388 37942
rect 38668 37828 38724 37838
rect 38276 37772 38388 37828
rect 38444 37826 38724 37828
rect 38444 37774 38670 37826
rect 38722 37774 38724 37826
rect 38444 37772 38724 37774
rect 38220 37762 38276 37772
rect 38332 37268 38388 37278
rect 38444 37268 38500 37772
rect 38668 37762 38724 37772
rect 38892 37492 38948 38782
rect 39116 38668 39172 40114
rect 39340 39956 39396 40348
rect 39452 40402 39508 40460
rect 39452 40350 39454 40402
rect 39506 40350 39508 40402
rect 39452 40338 39508 40350
rect 39676 40516 39732 40526
rect 39676 40402 39732 40460
rect 39676 40350 39678 40402
rect 39730 40350 39732 40402
rect 39676 40338 39732 40350
rect 40236 40402 40292 41468
rect 40236 40350 40238 40402
rect 40290 40350 40292 40402
rect 40236 40338 40292 40350
rect 40460 40402 40516 45724
rect 40852 45162 40908 45174
rect 40852 45110 40854 45162
rect 40906 45110 40908 45162
rect 40852 44996 40908 45110
rect 40852 44930 40908 44940
rect 41020 45136 41076 45148
rect 41020 45084 41022 45136
rect 41074 45084 41076 45136
rect 40908 44548 40964 44558
rect 40908 44454 40964 44492
rect 41020 44100 41076 45084
rect 41020 44034 41076 44044
rect 41020 43652 41076 43662
rect 41132 43652 41188 45836
rect 41244 45332 41300 49200
rect 42476 45890 42532 45902
rect 42476 45838 42478 45890
rect 42530 45838 42532 45890
rect 41244 45266 41300 45276
rect 41356 45444 41412 45454
rect 41244 45145 41300 45157
rect 41244 45093 41246 45145
rect 41298 45093 41300 45145
rect 41244 44884 41300 45093
rect 41244 44818 41300 44828
rect 41356 43708 41412 45388
rect 42252 45108 42308 45118
rect 42252 45014 42308 45052
rect 41804 44882 41860 44894
rect 41804 44830 41806 44882
rect 41858 44830 41860 44882
rect 41020 43650 41188 43652
rect 41020 43598 41022 43650
rect 41074 43598 41188 43650
rect 41020 43596 41188 43598
rect 41244 43652 41412 43708
rect 41468 44436 41524 44446
rect 41244 43596 41319 43652
rect 41020 43586 41076 43596
rect 41132 42868 41188 43596
rect 41263 43594 41319 43596
rect 41263 43542 41265 43594
rect 41317 43542 41319 43594
rect 41263 42980 41319 43542
rect 41468 43092 41524 44380
rect 41804 44436 41860 44830
rect 41804 44370 41860 44380
rect 42140 44100 42196 44110
rect 42140 43538 42196 44044
rect 42140 43486 42142 43538
rect 42194 43486 42196 43538
rect 42140 43474 42196 43486
rect 42476 43540 42532 45838
rect 42700 45890 42756 45902
rect 42700 45838 42702 45890
rect 42754 45838 42756 45890
rect 42476 43474 42532 43484
rect 42588 45108 42644 45118
rect 42420 43204 42476 43214
rect 42252 43092 42308 43102
rect 41468 43036 41748 43092
rect 41263 42924 41412 42980
rect 41132 42802 41188 42812
rect 40796 42756 40852 42766
rect 41020 42756 41076 42766
rect 40460 40350 40462 40402
rect 40514 40350 40516 40402
rect 40460 40338 40516 40350
rect 40684 42754 40852 42756
rect 40684 42702 40798 42754
rect 40850 42702 40852 42754
rect 40684 42700 40852 42702
rect 39956 40180 40012 40190
rect 39956 40178 40292 40180
rect 39956 40126 39958 40178
rect 40010 40126 40292 40178
rect 39956 40124 40292 40126
rect 39956 40114 40012 40124
rect 39228 39900 39396 39956
rect 40124 39956 40180 39966
rect 39228 39396 39284 39900
rect 39228 39340 39396 39396
rect 39228 38948 39284 38958
rect 39228 38854 39284 38892
rect 39004 38612 39172 38668
rect 39004 38050 39060 38612
rect 39340 38274 39396 39340
rect 39564 39172 39620 39182
rect 39564 38834 39620 39116
rect 39900 39060 39956 39070
rect 39900 38966 39956 39004
rect 39564 38782 39566 38834
rect 39618 38782 39620 38834
rect 39564 38770 39620 38782
rect 40124 38668 40180 39900
rect 39340 38222 39342 38274
rect 39394 38222 39396 38274
rect 39340 38210 39396 38222
rect 39452 38612 39508 38622
rect 39004 37998 39006 38050
rect 39058 37998 39060 38050
rect 39004 37986 39060 37998
rect 38892 37426 38948 37436
rect 38332 37266 38500 37268
rect 38332 37214 38334 37266
rect 38386 37214 38500 37266
rect 38332 37212 38500 37214
rect 38332 37202 38388 37212
rect 37996 37090 38052 37100
rect 39452 36148 39508 38556
rect 39900 38612 40180 38668
rect 39900 38274 39956 38612
rect 39900 38222 39902 38274
rect 39954 38222 39956 38274
rect 39900 38210 39956 38222
rect 40236 38050 40292 40124
rect 40684 39620 40740 42700
rect 40796 42690 40852 42700
rect 40908 42754 41076 42756
rect 40908 42702 41022 42754
rect 41074 42702 41076 42754
rect 40908 42700 41076 42702
rect 40908 42532 40964 42700
rect 41020 42690 41076 42700
rect 41188 42532 41244 42542
rect 40908 42466 40964 42476
rect 41020 42530 41244 42532
rect 41020 42478 41190 42530
rect 41242 42478 41244 42530
rect 41020 42476 41244 42478
rect 40796 41972 40852 41982
rect 40796 41878 40852 41916
rect 40684 39554 40740 39564
rect 40796 41074 40852 41086
rect 40796 41022 40798 41074
rect 40850 41022 40852 41074
rect 40796 39060 40852 41022
rect 40684 39004 40852 39060
rect 40908 39506 40964 39518
rect 40908 39454 40910 39506
rect 40962 39454 40964 39506
rect 40684 38724 40740 39004
rect 40796 38836 40852 38846
rect 40796 38742 40852 38780
rect 40684 38658 40740 38668
rect 40908 38276 40964 39454
rect 40908 38210 40964 38220
rect 40236 37998 40238 38050
rect 40290 37998 40292 38050
rect 40236 37986 40292 37998
rect 40852 37940 40908 37950
rect 40852 37846 40908 37884
rect 40012 37492 40068 37502
rect 39564 36484 39620 36494
rect 39564 36390 39620 36428
rect 39004 36092 39508 36148
rect 38612 35812 38668 35822
rect 38612 35718 38668 35756
rect 37716 35186 37772 35196
rect 37828 35532 37940 35588
rect 38108 35700 38164 35710
rect 38108 35586 38164 35644
rect 38892 35700 38948 35710
rect 38892 35606 38948 35644
rect 38108 35534 38110 35586
rect 38162 35534 38164 35586
rect 37660 35028 37716 35038
rect 37660 34934 37716 34972
rect 37828 34970 37884 35532
rect 38108 35522 38164 35534
rect 37828 34918 37830 34970
rect 37882 34918 37884 34970
rect 38276 35084 38612 35140
rect 38276 35026 38332 35084
rect 38276 34974 38278 35026
rect 38330 34974 38332 35026
rect 38276 34962 38332 34974
rect 37324 34804 37492 34860
rect 37324 34132 37380 34142
rect 37212 34130 37380 34132
rect 37212 34078 37326 34130
rect 37378 34078 37380 34130
rect 37212 34076 37380 34078
rect 37324 34066 37380 34076
rect 37436 34132 37492 34804
rect 37828 34356 37884 34918
rect 37828 34290 37884 34300
rect 38444 34914 38500 34926
rect 38444 34862 38446 34914
rect 38498 34862 38500 34914
rect 38444 34132 38500 34862
rect 37436 34130 38500 34132
rect 37436 34078 37438 34130
rect 37490 34078 38500 34130
rect 37436 34076 38500 34078
rect 37436 34066 37492 34076
rect 37100 33618 37156 33628
rect 35196 33282 35252 33294
rect 35364 33290 35420 33302
rect 35364 33238 35366 33290
rect 35418 33238 35420 33290
rect 34860 33068 35140 33124
rect 33348 31826 33404 31836
rect 33068 31778 33236 31780
rect 33068 31726 33070 31778
rect 33122 31726 33236 31778
rect 33068 31724 33236 31726
rect 33628 31778 33684 32396
rect 33628 31726 33630 31778
rect 33682 31726 33684 31778
rect 33068 31714 33124 31724
rect 33628 31714 33684 31726
rect 33740 31778 33796 31790
rect 33740 31726 33742 31778
rect 33794 31726 33796 31778
rect 32900 31558 32902 31610
rect 32954 31558 32956 31610
rect 32900 31546 32956 31558
rect 33068 30996 33124 31006
rect 33068 30902 33124 30940
rect 32732 30604 33012 30660
rect 32508 30370 32564 30380
rect 32396 30324 32452 30334
rect 32396 30171 32452 30268
rect 32396 30119 32398 30171
rect 32450 30119 32452 30171
rect 32396 30107 32452 30119
rect 32564 30100 32620 30110
rect 32564 29650 32620 30044
rect 32956 30098 33012 30604
rect 33516 30436 33572 30446
rect 33404 30378 33460 30390
rect 33180 30324 33236 30334
rect 33404 30326 33406 30378
rect 33458 30326 33460 30378
rect 33404 30324 33460 30326
rect 33236 30268 33460 30324
rect 33180 30258 33236 30268
rect 33516 30212 33572 30380
rect 32956 30046 32958 30098
rect 33010 30046 33012 30098
rect 32956 30034 33012 30046
rect 33292 30156 33572 30212
rect 33628 30212 33684 30222
rect 32564 29598 32566 29650
rect 32618 29598 32620 29650
rect 32564 29586 32620 29598
rect 33180 29988 33236 29998
rect 32284 29138 32340 29148
rect 31836 28980 31892 28990
rect 31836 28810 31892 28924
rect 31836 28758 31838 28810
rect 31890 28758 31892 28810
rect 31836 28746 31892 28758
rect 32844 28868 32900 28878
rect 31724 28578 31780 28588
rect 31836 28642 31892 28654
rect 31836 28590 31838 28642
rect 31890 28590 31892 28642
rect 31836 28196 31892 28590
rect 32564 28644 32620 28654
rect 32564 28550 32620 28588
rect 31052 26562 31108 26572
rect 31276 28140 31892 28196
rect 32732 28420 32788 28430
rect 31276 28082 31332 28140
rect 31276 28030 31278 28082
rect 31330 28030 31332 28082
rect 30492 26348 30772 26404
rect 30492 26180 30548 26348
rect 30828 26292 30884 26302
rect 30380 26124 30492 26180
rect 30156 25340 30324 25396
rect 29708 25228 29876 25284
rect 29484 24724 29540 24734
rect 29484 24630 29540 24668
rect 29372 24444 29540 24500
rect 28868 24322 28924 24332
rect 28476 24054 28478 24106
rect 28530 24054 28532 24106
rect 28476 24042 28532 24054
rect 29484 24106 29540 24444
rect 29484 24054 29486 24106
rect 29538 24054 29540 24106
rect 27020 23202 27076 23212
rect 27692 23268 27748 23278
rect 26796 23154 26852 23166
rect 26796 23102 26798 23154
rect 26850 23102 26852 23154
rect 24780 22318 24782 22370
rect 24834 22318 24836 22370
rect 24780 22306 24836 22318
rect 24892 22540 25060 22596
rect 26124 22876 26292 22932
rect 26572 22932 26628 22942
rect 24892 22370 24948 22540
rect 25452 22484 25508 22494
rect 25452 22482 25732 22484
rect 25452 22430 25454 22482
rect 25506 22430 25732 22482
rect 25452 22428 25732 22430
rect 25452 22418 25508 22428
rect 24892 22318 24894 22370
rect 24946 22318 24948 22370
rect 23660 21858 23716 21868
rect 24500 22146 24556 22158
rect 24500 22094 24502 22146
rect 24554 22094 24556 22146
rect 24500 21924 24556 22094
rect 24892 22148 24948 22318
rect 24892 22082 24948 22092
rect 25060 22314 25116 22326
rect 25060 22262 25062 22314
rect 25114 22262 25116 22314
rect 24500 21858 24556 21868
rect 25060 21924 25116 22262
rect 25676 22036 25732 22428
rect 25788 22372 25844 22382
rect 25788 22370 26068 22372
rect 25788 22318 25790 22370
rect 25842 22318 26068 22370
rect 25788 22316 26068 22318
rect 25788 22306 25844 22316
rect 25676 21980 25878 22036
rect 25060 21858 25116 21868
rect 24276 21700 24332 21710
rect 23324 20804 23380 20814
rect 23212 20748 23324 20804
rect 23324 20710 23380 20748
rect 23436 20356 23492 21084
rect 24220 21644 24276 21700
rect 24220 21606 24332 21644
rect 25116 21700 25172 21710
rect 23436 20290 23492 20300
rect 23548 20746 23604 20758
rect 23548 20694 23550 20746
rect 23602 20694 23604 20746
rect 23548 20244 23604 20694
rect 23548 20178 23604 20188
rect 24108 20132 24164 20142
rect 24108 20074 24164 20076
rect 23492 20020 23548 20030
rect 23100 19796 23156 19806
rect 23100 19702 23156 19740
rect 23156 19572 23212 19582
rect 23156 19346 23212 19516
rect 23492 19458 23548 19964
rect 23772 20018 23828 20030
rect 23772 19966 23774 20018
rect 23826 19966 23828 20018
rect 24108 20022 24110 20074
rect 24162 20022 24164 20074
rect 24108 20010 24164 20022
rect 23772 19796 23828 19966
rect 24108 19908 24164 19918
rect 24108 19814 24164 19852
rect 23492 19406 23494 19458
rect 23546 19406 23548 19458
rect 23492 19394 23548 19406
rect 23660 19572 23716 19582
rect 23156 19294 23158 19346
rect 23210 19294 23212 19346
rect 23156 19282 23212 19294
rect 23660 19292 23716 19516
rect 23548 19236 23716 19292
rect 22988 18452 23044 18462
rect 23548 18450 23604 19236
rect 23772 19234 23828 19740
rect 24220 19684 24276 21606
rect 24724 21588 24780 21598
rect 24724 21494 24780 21532
rect 24892 20916 24948 20926
rect 24892 20822 24948 20860
rect 24556 20804 24612 20814
rect 24332 20802 24612 20804
rect 24332 20750 24558 20802
rect 24610 20750 24612 20802
rect 25116 20802 25172 21644
rect 25822 21624 25878 21980
rect 24332 20748 24612 20750
rect 24332 19796 24388 20748
rect 24556 20738 24612 20748
rect 24948 20746 25004 20758
rect 24948 20694 24950 20746
rect 25002 20694 25004 20746
rect 25116 20750 25118 20802
rect 25170 20750 25172 20802
rect 25116 20738 25172 20750
rect 25452 21588 25508 21598
rect 25564 21588 25620 21598
rect 25508 21586 25620 21588
rect 25508 21534 25566 21586
rect 25618 21534 25620 21586
rect 25508 21532 25620 21534
rect 24948 20692 25004 20694
rect 24948 20636 25060 20692
rect 25004 20468 25060 20636
rect 25004 20412 25172 20468
rect 25116 20132 25172 20412
rect 25452 20356 25508 21532
rect 25564 21522 25620 21532
rect 25676 21586 25732 21598
rect 25676 21534 25678 21586
rect 25730 21534 25732 21586
rect 25822 21572 25824 21624
rect 25876 21572 25878 21624
rect 25822 21560 25878 21572
rect 26012 21588 26068 22316
rect 26124 21700 26180 22876
rect 26124 21634 26180 21644
rect 26236 22708 26292 22718
rect 25676 20804 25732 21534
rect 25452 20290 25508 20300
rect 25564 20580 25620 20590
rect 25676 20580 25732 20748
rect 25788 20804 25844 20814
rect 26012 20804 26068 21532
rect 26236 21474 26292 22652
rect 26572 22482 26628 22876
rect 26796 22820 26852 23102
rect 26796 22754 26852 22764
rect 26908 23154 26964 23166
rect 26908 23102 26910 23154
rect 26962 23102 26964 23154
rect 26908 22708 26964 23102
rect 27244 22932 27300 22942
rect 27244 22838 27300 22876
rect 26908 22642 26964 22652
rect 26572 22430 26574 22482
rect 26626 22430 26628 22482
rect 26572 22418 26628 22430
rect 27692 22372 27748 23212
rect 27960 23192 28016 23204
rect 27960 23156 27962 23192
rect 28014 23156 28016 23192
rect 27960 23090 28016 23100
rect 28252 23156 28308 23436
rect 28252 23090 28308 23100
rect 28364 23938 28420 23950
rect 28364 23886 28366 23938
rect 28418 23886 28420 23938
rect 28364 23716 28420 23886
rect 29260 23938 29316 23950
rect 29260 23886 29262 23938
rect 29314 23886 29316 23938
rect 28364 22484 28420 23660
rect 28700 23828 28756 23838
rect 28700 23154 28756 23772
rect 29260 23828 29316 23886
rect 29260 23762 29316 23772
rect 29372 23940 29428 23950
rect 29260 23156 29316 23166
rect 29372 23156 29428 23884
rect 28700 23102 28702 23154
rect 28754 23102 28756 23154
rect 28700 22932 28756 23102
rect 28812 23154 29428 23156
rect 28812 23102 29262 23154
rect 29314 23102 29428 23154
rect 28812 23100 29428 23102
rect 29484 23154 29540 24054
rect 29484 23102 29486 23154
rect 29538 23102 29540 23154
rect 28812 22986 28868 23100
rect 29260 23090 29316 23100
rect 29484 23090 29540 23102
rect 28812 22934 28814 22986
rect 28866 22934 28868 22986
rect 28812 22922 28868 22934
rect 29484 22986 29540 22998
rect 29484 22934 29486 22986
rect 29538 22934 29540 22986
rect 29484 22932 29540 22934
rect 29708 22932 29764 25228
rect 30156 25172 30212 25182
rect 30156 24622 30212 25116
rect 30268 24836 30324 25340
rect 30268 24770 30324 24780
rect 30380 24790 30436 26124
rect 30492 26086 30548 26124
rect 30604 26290 30884 26292
rect 30604 26238 30830 26290
rect 30882 26238 30884 26290
rect 30604 26236 30884 26238
rect 30604 25956 30660 26236
rect 30828 26226 30884 26236
rect 30940 26290 30996 26302
rect 30940 26238 30942 26290
rect 30994 26238 30996 26290
rect 30492 25900 30660 25956
rect 30716 26068 30772 26078
rect 30492 25450 30548 25900
rect 30492 25398 30494 25450
rect 30546 25398 30548 25450
rect 30492 25396 30548 25398
rect 30492 25330 30548 25340
rect 30604 25508 30660 25518
rect 30380 24778 30473 24790
rect 30380 24726 30419 24778
rect 30471 24726 30473 24778
rect 30380 24724 30473 24726
rect 30417 24714 30473 24724
rect 30604 24778 30660 25452
rect 30604 24726 30606 24778
rect 30658 24726 30660 24778
rect 30604 24714 30660 24726
rect 30156 24612 30268 24622
rect 29484 22876 29764 22932
rect 29820 24610 30268 24612
rect 29820 24558 30214 24610
rect 30266 24558 30268 24610
rect 29820 24556 30268 24558
rect 28700 22866 28756 22876
rect 28588 22820 28644 22830
rect 28476 22484 28532 22494
rect 28364 22482 28532 22484
rect 28364 22430 28478 22482
rect 28530 22430 28532 22482
rect 28364 22428 28532 22430
rect 28476 22418 28532 22428
rect 27356 22148 27412 22158
rect 26236 21422 26238 21474
rect 26290 21422 26292 21474
rect 26236 21410 26292 21422
rect 26460 22036 26516 22046
rect 25788 20802 26068 20804
rect 25788 20750 25790 20802
rect 25842 20750 26068 20802
rect 25788 20748 26068 20750
rect 26124 21252 26180 21262
rect 25788 20738 25844 20748
rect 26124 20580 26180 21196
rect 25676 20524 25956 20580
rect 24332 19730 24388 19740
rect 24444 20020 24500 20030
rect 24444 20018 24724 20020
rect 24444 19966 24446 20018
rect 24498 19966 24724 20018
rect 24444 19964 24724 19966
rect 24052 19628 24276 19684
rect 24052 19572 24108 19628
rect 24052 19290 24108 19516
rect 24444 19292 24500 19964
rect 24668 19348 24724 19964
rect 25116 19796 25172 20076
rect 25564 20244 25620 20524
rect 25452 20020 25508 20030
rect 25564 20020 25620 20188
rect 25788 20020 25844 20030
rect 25564 20018 25844 20020
rect 25564 19966 25790 20018
rect 25842 19966 25844 20018
rect 25564 19964 25844 19966
rect 25452 19926 25508 19964
rect 25788 19954 25844 19964
rect 25900 20018 25956 20524
rect 25900 19966 25902 20018
rect 25954 19966 25956 20018
rect 26086 20524 26180 20580
rect 26086 20056 26142 20524
rect 26460 20132 26516 21980
rect 27198 21812 27254 21822
rect 27198 21636 27254 21756
rect 27198 21584 27200 21636
rect 27252 21584 27254 21636
rect 27198 21572 27254 21584
rect 27356 21586 27412 22092
rect 27356 21534 27358 21586
rect 27410 21534 27412 21586
rect 27356 21522 27412 21534
rect 27468 21588 27524 21598
rect 27692 21588 27748 22316
rect 27972 21812 28028 21822
rect 27972 21718 28028 21756
rect 28588 21754 28644 22764
rect 29640 22372 29696 22382
rect 29640 22280 29642 22316
rect 29694 22280 29696 22316
rect 29640 21812 29696 22280
rect 28588 21702 28590 21754
rect 28642 21702 28644 21754
rect 28588 21690 28644 21702
rect 29484 21756 29696 21812
rect 29820 21812 29876 24556
rect 30212 24546 30268 24556
rect 30492 24612 30548 24622
rect 30156 24276 30212 24286
rect 30000 23900 30056 23912
rect 30000 23848 30002 23900
rect 30054 23848 30056 23900
rect 30000 23716 30056 23848
rect 30000 23650 30056 23660
rect 29932 23156 29988 23166
rect 29932 22820 29988 23100
rect 30044 23156 30100 23166
rect 30156 23156 30212 24220
rect 30380 24164 30436 24174
rect 30380 23278 30436 24108
rect 30324 23266 30436 23278
rect 30324 23214 30326 23266
rect 30378 23214 30436 23266
rect 30324 23212 30436 23214
rect 30324 23202 30380 23212
rect 30044 23154 30212 23156
rect 30044 23102 30046 23154
rect 30098 23102 30212 23154
rect 30044 23100 30212 23102
rect 30044 23090 30100 23100
rect 29932 22754 29988 22764
rect 30492 22538 30548 24556
rect 30604 24276 30660 24286
rect 30604 23910 30660 24220
rect 30604 23858 30606 23910
rect 30658 23858 30660 23910
rect 30604 23846 30660 23858
rect 30716 22596 30772 26012
rect 30940 25956 30996 26238
rect 31108 26068 31164 26078
rect 31108 26066 31220 26068
rect 31108 26014 31110 26066
rect 31162 26014 31220 26066
rect 31108 26002 31220 26014
rect 30940 25890 30996 25900
rect 30828 25844 30884 25854
rect 30828 25618 30884 25788
rect 30828 25566 30830 25618
rect 30882 25566 30884 25618
rect 30828 25554 30884 25566
rect 31052 25508 31108 25518
rect 31052 25414 31108 25452
rect 31164 25396 31220 26002
rect 31276 25620 31332 28030
rect 32564 28084 32620 28094
rect 32564 27990 32620 28028
rect 32116 27972 32172 27982
rect 32116 27878 32172 27916
rect 32732 27188 32788 28364
rect 31612 27076 31668 27114
rect 32732 27086 32788 27132
rect 31836 27076 31892 27086
rect 31612 27010 31668 27020
rect 31724 27074 31892 27076
rect 31724 27022 31838 27074
rect 31890 27022 31892 27074
rect 31724 27020 31892 27022
rect 31444 26908 31500 26918
rect 31724 26908 31780 27020
rect 31836 27010 31892 27020
rect 32712 27074 32788 27086
rect 32712 27022 32714 27074
rect 32766 27022 32788 27074
rect 32712 27020 32788 27022
rect 32712 27010 32768 27020
rect 31444 26906 31780 26908
rect 31444 26854 31446 26906
rect 31498 26854 31780 26906
rect 31444 26852 31780 26854
rect 31836 26852 31892 26862
rect 31444 26842 31500 26852
rect 31668 26628 31724 26638
rect 31668 26514 31724 26572
rect 31668 26462 31670 26514
rect 31722 26462 31724 26514
rect 31668 26450 31724 26462
rect 31836 26068 31892 26796
rect 32116 26628 32172 26638
rect 32116 26516 32172 26572
rect 32732 26628 32788 26638
rect 31836 26002 31892 26012
rect 32060 26514 32172 26516
rect 32060 26462 32118 26514
rect 32170 26462 32172 26514
rect 32060 26450 32172 26462
rect 32564 26516 32620 26526
rect 32732 26516 32788 26572
rect 32564 26514 32788 26516
rect 32564 26462 32566 26514
rect 32618 26462 32788 26514
rect 32564 26460 32788 26462
rect 32564 26450 32620 26460
rect 31276 25564 31780 25620
rect 31164 24836 31220 25340
rect 31612 25450 31668 25462
rect 31612 25398 31614 25450
rect 31666 25398 31668 25450
rect 31108 24780 31220 24836
rect 31332 25284 31388 25294
rect 31332 24834 31388 25228
rect 31332 24782 31334 24834
rect 31386 24782 31388 24834
rect 31108 24778 31164 24780
rect 30884 24757 30940 24769
rect 30884 24705 30886 24757
rect 30938 24724 30940 24757
rect 31108 24726 31110 24778
rect 31162 24726 31164 24778
rect 31332 24770 31388 24782
rect 30938 24705 30996 24724
rect 31108 24714 31164 24726
rect 30884 24668 30996 24705
rect 30940 24612 30996 24668
rect 31612 24612 31668 25398
rect 31724 24724 31780 25564
rect 32060 25172 32116 26450
rect 32172 25450 32228 25462
rect 32172 25398 32174 25450
rect 32226 25398 32228 25450
rect 32172 25396 32228 25398
rect 32172 25330 32228 25340
rect 32060 25116 32228 25172
rect 32060 24948 32116 24958
rect 31948 24836 32004 24846
rect 31724 24658 31780 24668
rect 31836 24722 31892 24734
rect 31836 24670 31838 24722
rect 31890 24670 31892 24722
rect 30940 24556 31668 24612
rect 30940 24164 30996 24556
rect 30940 24098 30996 24108
rect 31724 24276 31780 24286
rect 30828 23940 30884 23950
rect 30828 23938 30996 23940
rect 30828 23886 30830 23938
rect 30882 23886 30996 23938
rect 30828 23884 30996 23886
rect 30828 23874 30884 23884
rect 30492 22486 30494 22538
rect 30546 22486 30548 22538
rect 30492 22474 30548 22486
rect 30604 22540 30772 22596
rect 30828 23716 30884 23726
rect 27468 21586 27748 21588
rect 27468 21534 27470 21586
rect 27522 21534 27748 21586
rect 27468 21532 27748 21534
rect 28700 21586 28756 21598
rect 28700 21534 28702 21586
rect 28754 21534 28756 21586
rect 27468 21522 27524 21532
rect 26796 21362 26852 21374
rect 26796 21310 26798 21362
rect 26850 21310 26852 21362
rect 26796 21252 26852 21310
rect 26796 21186 26852 21196
rect 26796 21028 26852 21038
rect 26086 20004 26088 20056
rect 26140 20004 26142 20056
rect 26086 19992 26142 20004
rect 26348 20076 26516 20132
rect 26572 20802 26628 20814
rect 26572 20750 26574 20802
rect 26626 20750 26628 20802
rect 26572 20132 26628 20750
rect 26796 20580 26852 20972
rect 28476 20916 28532 20926
rect 28700 20916 28756 21534
rect 29148 21588 29204 21598
rect 28476 20914 29092 20916
rect 28476 20862 28478 20914
rect 28530 20862 29092 20914
rect 28476 20860 29092 20862
rect 28476 20850 28532 20860
rect 29036 20802 29092 20860
rect 29036 20750 29038 20802
rect 29090 20750 29092 20802
rect 29036 20738 29092 20750
rect 26796 20524 26964 20580
rect 25900 19954 25956 19966
rect 25284 19850 25340 19862
rect 25284 19798 25286 19850
rect 25338 19798 25340 19850
rect 25284 19796 25340 19798
rect 25116 19740 25340 19796
rect 25004 19348 25060 19358
rect 24668 19292 24780 19348
rect 23772 19182 23774 19234
rect 23826 19182 23828 19234
rect 23772 18900 23828 19182
rect 23884 19236 23940 19246
rect 24052 19238 24054 19290
rect 24106 19238 24108 19290
rect 24052 19226 24108 19238
rect 24220 19234 24276 19246
rect 23884 19142 23940 19180
rect 24220 19182 24222 19234
rect 24274 19182 24276 19234
rect 24220 19012 24276 19182
rect 24220 18946 24276 18956
rect 24332 19236 24500 19292
rect 24724 19290 24780 19292
rect 23772 18834 23828 18844
rect 24332 18788 24388 19236
rect 24108 18732 24388 18788
rect 24556 19234 24612 19246
rect 24556 19182 24558 19234
rect 24610 19182 24612 19234
rect 24724 19238 24726 19290
rect 24778 19238 24780 19290
rect 24724 19226 24780 19238
rect 24836 19236 24948 19246
rect 24556 19012 24612 19182
rect 24892 19234 24948 19236
rect 24892 19182 24894 19234
rect 24946 19182 24948 19234
rect 24892 19180 24948 19182
rect 24836 19170 24948 19180
rect 25004 19234 25060 19292
rect 25004 19182 25006 19234
rect 25058 19182 25060 19234
rect 25004 19170 25060 19182
rect 23716 18676 23772 18686
rect 24108 18676 24164 18732
rect 23716 18674 24164 18676
rect 23716 18622 23718 18674
rect 23770 18622 24164 18674
rect 23716 18620 24164 18622
rect 23716 18610 23772 18620
rect 22988 18358 23044 18396
rect 23380 18394 23436 18406
rect 23212 18338 23268 18350
rect 23212 18286 23214 18338
rect 23266 18286 23268 18338
rect 23212 18228 23268 18286
rect 23212 18162 23268 18172
rect 23380 18342 23382 18394
rect 23434 18342 23436 18394
rect 23380 18004 23436 18342
rect 22876 16258 22932 16268
rect 22988 17948 23436 18004
rect 23548 18398 23550 18450
rect 23602 18398 23604 18450
rect 22988 16322 23044 17948
rect 23324 17834 23380 17846
rect 23324 17782 23326 17834
rect 23378 17782 23380 17834
rect 23324 17332 23380 17782
rect 23436 17780 23492 17790
rect 23436 17666 23492 17724
rect 23436 17614 23438 17666
rect 23490 17614 23492 17666
rect 23436 17602 23492 17614
rect 23548 17668 23604 18398
rect 23548 17602 23604 17612
rect 23660 18452 23716 18462
rect 23660 17666 23716 18396
rect 24108 18450 24164 18620
rect 24556 18564 24612 18956
rect 24556 18498 24612 18508
rect 24780 19012 24836 19022
rect 25116 19012 25172 19740
rect 26348 19460 26404 20076
rect 26572 20066 26628 20076
rect 26796 20018 26852 20030
rect 26796 19966 26798 20018
rect 26850 19966 26852 20018
rect 26460 19908 26516 19918
rect 26796 19908 26852 19966
rect 26460 19906 26852 19908
rect 26460 19854 26462 19906
rect 26514 19854 26852 19906
rect 26460 19852 26852 19854
rect 26460 19842 26516 19852
rect 26348 19404 26516 19460
rect 25676 19348 25732 19358
rect 25564 19236 25620 19246
rect 25284 19124 25340 19162
rect 25284 19058 25340 19068
rect 24108 18398 24110 18450
rect 24162 18398 24164 18450
rect 24108 18386 24164 18398
rect 24220 18450 24276 18462
rect 24444 18452 24500 18462
rect 24220 18398 24222 18450
rect 24274 18398 24276 18450
rect 23660 17614 23662 17666
rect 23714 17614 23716 17666
rect 23660 17602 23716 17614
rect 23324 17266 23380 17276
rect 23716 17332 23772 17342
rect 22988 16270 22990 16322
rect 23042 16270 23044 16322
rect 22988 16258 23044 16270
rect 23212 17220 23268 17230
rect 23212 16100 23268 17164
rect 23380 17108 23436 17118
rect 23716 17108 23772 17276
rect 23380 17014 23436 17052
rect 23548 17106 23772 17108
rect 23548 17054 23718 17106
rect 23770 17054 23772 17106
rect 23548 17052 23772 17054
rect 23436 16772 23492 16782
rect 22764 16044 23156 16100
rect 22596 15990 22598 16042
rect 22650 15990 22652 16042
rect 22596 15988 22652 15990
rect 22596 15932 22820 15988
rect 22316 15596 22484 15652
rect 21980 15262 21982 15314
rect 22034 15262 22036 15314
rect 22166 15484 22260 15540
rect 22166 15352 22222 15484
rect 22166 15300 22168 15352
rect 22220 15300 22222 15352
rect 22166 15288 22222 15300
rect 21980 15250 22036 15262
rect 21756 15204 21812 15214
rect 21756 14980 21812 15148
rect 22316 15204 22372 15214
rect 22148 15092 22204 15102
rect 21756 14924 21924 14980
rect 21756 14530 21812 14542
rect 21756 14478 21758 14530
rect 21810 14478 21812 14530
rect 21756 13860 21812 14478
rect 21868 14420 21924 14924
rect 22148 14642 22204 15036
rect 22148 14590 22150 14642
rect 22202 14590 22204 14642
rect 22148 14578 22204 14590
rect 22316 14530 22372 15148
rect 22428 14980 22484 15596
rect 22540 15428 22596 15438
rect 22540 15202 22596 15372
rect 22540 15150 22542 15202
rect 22594 15150 22596 15202
rect 22540 15138 22596 15150
rect 22428 14924 22596 14980
rect 22316 14478 22318 14530
rect 22370 14478 22372 14530
rect 22316 14420 22372 14478
rect 21868 14364 22372 14420
rect 22428 14756 22484 14766
rect 21756 13794 21812 13804
rect 21980 13748 22036 13758
rect 21980 13654 22036 13692
rect 22092 13746 22148 13758
rect 22092 13694 22094 13746
rect 22146 13694 22148 13746
rect 22428 13746 22484 14700
rect 20748 13010 20804 13020
rect 20300 12910 20302 12962
rect 20354 12910 20356 12962
rect 20300 12898 20356 12910
rect 20636 12964 20692 12974
rect 20636 12870 20692 12908
rect 21308 12962 21364 13580
rect 21308 12910 21310 12962
rect 21362 12910 21364 12962
rect 21476 13580 21588 13636
rect 21476 13018 21532 13580
rect 21700 13522 21756 13534
rect 21700 13470 21702 13522
rect 21754 13470 21756 13522
rect 21700 13188 21756 13470
rect 22092 13412 22148 13694
rect 22260 13690 22316 13702
rect 22260 13638 22262 13690
rect 22314 13638 22316 13690
rect 22260 13534 22316 13638
rect 22428 13694 22430 13746
rect 22482 13694 22484 13746
rect 22428 13636 22484 13694
rect 22428 13570 22484 13580
rect 22260 13524 22372 13534
rect 22260 13468 22316 13524
rect 22316 13458 22372 13468
rect 22540 13524 22596 14924
rect 22652 14306 22708 14318
rect 22652 14254 22654 14306
rect 22706 14254 22708 14306
rect 22652 14196 22708 14254
rect 22652 14130 22708 14140
rect 22540 13458 22596 13468
rect 22148 13356 22260 13412
rect 22092 13318 22148 13356
rect 21700 13122 21756 13132
rect 21476 12966 21478 13018
rect 21530 12966 21532 13018
rect 21476 12954 21532 12966
rect 21756 12964 21812 12974
rect 21308 12898 21364 12910
rect 21644 12850 21700 12862
rect 21644 12798 21646 12850
rect 21698 12798 21700 12850
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19684 12404 19740 12414
rect 19292 12348 19460 12404
rect 18956 12338 19012 12348
rect 19068 12206 19124 12218
rect 19068 12154 19070 12206
rect 19122 12154 19124 12206
rect 19068 11956 19124 12154
rect 19068 11890 19124 11900
rect 19292 12178 19348 12190
rect 19292 12126 19294 12178
rect 19346 12126 19348 12178
rect 18732 11666 18788 11676
rect 18844 11172 18900 11182
rect 18172 10558 18174 10610
rect 18226 10558 18228 10610
rect 18172 9492 18228 10558
rect 18172 9426 18228 9436
rect 18284 10610 18340 10622
rect 18284 10558 18286 10610
rect 18338 10558 18340 10610
rect 18284 9714 18340 10558
rect 18844 10612 18900 11116
rect 19012 10836 19068 10846
rect 19292 10836 19348 12126
rect 19404 12180 19460 12348
rect 19684 12234 19740 12348
rect 19684 12182 19686 12234
rect 19738 12182 19740 12234
rect 21644 12292 21700 12798
rect 21644 12226 21700 12236
rect 19684 12170 19740 12182
rect 19852 12180 19908 12190
rect 19404 12114 19460 12124
rect 19852 12086 19908 12124
rect 21756 12180 21812 12908
rect 22036 12852 22092 12862
rect 21756 12114 21812 12124
rect 21868 12850 22092 12852
rect 21868 12798 22038 12850
rect 22090 12798 22092 12850
rect 21868 12796 22092 12798
rect 19516 12066 19572 12078
rect 19516 12014 19518 12066
rect 19570 12014 19572 12066
rect 19012 10834 19348 10836
rect 19012 10782 19014 10834
rect 19066 10782 19348 10834
rect 19012 10780 19348 10782
rect 19404 11732 19460 11742
rect 19012 10770 19068 10780
rect 18844 10610 19012 10612
rect 18844 10558 18846 10610
rect 18898 10558 19012 10610
rect 18844 10556 19012 10558
rect 18844 10546 18900 10556
rect 18844 9828 18900 9838
rect 18284 9662 18286 9714
rect 18338 9662 18340 9714
rect 18060 9266 18172 9278
rect 18060 9214 18118 9266
rect 18170 9214 18172 9266
rect 18060 9212 18172 9214
rect 18116 9202 18172 9212
rect 17836 8652 18228 8708
rect 17500 8540 17892 8596
rect 15540 8318 15542 8370
rect 15594 8318 15596 8370
rect 15540 8306 15596 8318
rect 16044 8316 16212 8372
rect 16380 8484 16436 8494
rect 15260 8194 15316 8204
rect 16044 7588 16100 8316
rect 16156 8146 16212 8158
rect 16156 8094 16158 8146
rect 16210 8094 16212 8146
rect 16156 8036 16212 8094
rect 16212 7980 16324 8036
rect 16156 7970 16212 7980
rect 16156 7588 16212 7598
rect 16044 7586 16212 7588
rect 16044 7534 16158 7586
rect 16210 7534 16212 7586
rect 16044 7532 16212 7534
rect 16156 7522 16212 7532
rect 14812 7420 14980 7476
rect 15036 7476 15092 7514
rect 14308 6860 14420 6916
rect 14700 7028 14756 7038
rect 13916 6858 13972 6860
rect 13916 6806 13918 6858
rect 13970 6806 13972 6858
rect 13916 6020 13972 6806
rect 14252 6804 14308 6860
rect 13916 5954 13972 5964
rect 14028 6748 14308 6804
rect 13692 5404 13860 5460
rect 13468 5170 13524 5180
rect 12796 5122 12964 5124
rect 12796 5070 12798 5122
rect 12850 5070 12964 5122
rect 12796 5068 12964 5070
rect 13648 5082 13704 5094
rect 12796 5058 12852 5068
rect 13648 5030 13650 5082
rect 13702 5030 13704 5082
rect 12684 5012 12740 5022
rect 12684 4338 12740 4956
rect 13468 5012 13524 5022
rect 13468 4918 13524 4956
rect 13648 4564 13704 5030
rect 13804 4788 13860 5404
rect 14028 5124 14084 6748
rect 14476 6690 14532 6702
rect 14476 6638 14478 6690
rect 14530 6638 14532 6690
rect 14476 6580 14532 6638
rect 14700 6692 14756 6972
rect 14812 6916 14868 7420
rect 15036 7410 15092 7420
rect 15912 7474 15968 7486
rect 15912 7422 15914 7474
rect 15966 7422 15968 7474
rect 15912 7028 15968 7422
rect 15912 6962 15968 6972
rect 15148 6916 15204 6926
rect 14812 6860 14980 6916
rect 14812 6692 14868 6702
rect 14700 6690 14868 6692
rect 14700 6638 14814 6690
rect 14866 6638 14868 6690
rect 14700 6636 14868 6638
rect 14476 6514 14532 6524
rect 14700 6356 14756 6366
rect 14196 5794 14252 5806
rect 14196 5742 14198 5794
rect 14250 5742 14252 5794
rect 14196 5348 14252 5742
rect 14532 5684 14588 5694
rect 14196 5282 14252 5292
rect 14476 5682 14588 5684
rect 14476 5630 14534 5682
rect 14586 5630 14588 5682
rect 14476 5618 14588 5630
rect 14476 5124 14532 5618
rect 13972 5068 14084 5124
rect 14420 5068 14532 5124
rect 13972 5066 14028 5068
rect 13972 5014 13974 5066
rect 14026 5014 14028 5066
rect 13972 5002 14028 5014
rect 14420 5066 14476 5068
rect 14420 5014 14422 5066
rect 14474 5014 14476 5066
rect 14420 5002 14476 5014
rect 14588 5066 14644 5078
rect 14588 5014 14590 5066
rect 14642 5014 14644 5066
rect 14588 5012 14644 5014
rect 14588 4946 14644 4956
rect 13804 4722 13860 4732
rect 14476 4788 14532 4798
rect 13648 4508 13860 4564
rect 12684 4286 12686 4338
rect 12738 4286 12740 4338
rect 12684 4274 12740 4286
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 12572 3938 12628 3948
rect 13356 4004 13412 4014
rect 4476 3882 4740 3892
rect 13356 3780 13412 3948
rect 13356 3554 13412 3724
rect 13804 3722 13860 4508
rect 13804 3670 13806 3722
rect 13858 3670 13860 3722
rect 13804 3658 13860 3670
rect 14476 3668 14532 4732
rect 14588 4452 14644 4462
rect 14700 4452 14756 6300
rect 14812 5906 14868 6636
rect 14924 6468 14980 6860
rect 15148 6802 15204 6860
rect 15148 6750 15150 6802
rect 15202 6750 15204 6802
rect 15148 6738 15204 6750
rect 14924 6402 14980 6412
rect 15036 6692 15092 6702
rect 15036 6599 15038 6636
rect 15090 6599 15092 6636
rect 14924 6020 14980 6030
rect 15036 6020 15092 6599
rect 15484 6690 15540 6702
rect 15484 6638 15486 6690
rect 15538 6638 15540 6690
rect 16156 6692 16212 6702
rect 16268 6692 16324 7980
rect 16156 6690 16324 6692
rect 14924 6018 15092 6020
rect 14924 5966 14926 6018
rect 14978 5966 15092 6018
rect 14924 5964 15092 5966
rect 15260 6580 15316 6590
rect 14924 5954 14980 5964
rect 15148 5908 15204 5918
rect 14812 5854 14814 5906
rect 14866 5854 14868 5906
rect 14812 5842 14868 5854
rect 15092 5852 15148 5908
rect 15092 5850 15204 5852
rect 15092 5798 15094 5850
rect 15146 5842 15204 5850
rect 15260 5906 15316 6524
rect 15260 5854 15262 5906
rect 15314 5854 15316 5906
rect 15260 5842 15316 5854
rect 15484 6132 15540 6638
rect 15764 6634 15820 6646
rect 15764 6582 15766 6634
rect 15818 6582 15820 6634
rect 16156 6638 16158 6690
rect 16210 6638 16324 6690
rect 16156 6636 16324 6638
rect 16380 6692 16436 8428
rect 17836 8036 17892 8540
rect 18060 8484 18116 8494
rect 18060 8370 18116 8428
rect 18060 8318 18062 8370
rect 18114 8318 18116 8370
rect 18060 8306 18116 8318
rect 17556 7980 17892 8036
rect 17556 7698 17612 7980
rect 17556 7646 17558 7698
rect 17610 7646 17612 7698
rect 17556 7634 17612 7646
rect 16940 7476 16996 7486
rect 16940 7382 16996 7420
rect 17948 7476 18004 7486
rect 17948 7362 18004 7420
rect 17948 7310 17950 7362
rect 18002 7310 18004 7362
rect 17948 7298 18004 7310
rect 18060 7364 18116 7374
rect 16772 7250 16828 7262
rect 16772 7198 16774 7250
rect 16826 7198 16828 7250
rect 16772 7028 16828 7198
rect 16772 6962 16828 6972
rect 16156 6626 16212 6636
rect 16380 6610 16382 6636
rect 16434 6610 16436 6636
rect 16380 6598 16436 6610
rect 17052 6692 17108 6702
rect 17052 6598 17108 6636
rect 17388 6692 17444 6702
rect 17388 6598 17444 6636
rect 17836 6690 17892 6702
rect 17836 6638 17838 6690
rect 17890 6638 17892 6690
rect 15764 6356 15820 6582
rect 15932 6580 15988 6590
rect 15932 6486 15988 6524
rect 17836 6468 17892 6638
rect 17836 6402 17892 6412
rect 15764 6290 15820 6300
rect 17612 6356 17668 6366
rect 15484 6076 16436 6132
rect 15146 5798 15148 5842
rect 15092 5236 15148 5798
rect 14588 4450 14756 4452
rect 14588 4398 14590 4450
rect 14642 4398 14756 4450
rect 14588 4396 14756 4398
rect 14588 4386 14644 4396
rect 13356 3502 13358 3554
rect 13410 3502 13412 3554
rect 13356 3490 13412 3502
rect 13692 3556 13748 3566
rect 14196 3556 14252 3566
rect 13692 3554 14252 3556
rect 13692 3502 13694 3554
rect 13746 3502 14198 3554
rect 14250 3502 14252 3554
rect 13692 3500 14252 3502
rect 13692 3490 13748 3500
rect 14196 3490 14252 3500
rect 14476 3554 14532 3612
rect 14476 3502 14478 3554
rect 14530 3502 14532 3554
rect 14476 3490 14532 3502
rect 14700 3554 14756 4396
rect 15036 5180 15148 5236
rect 15260 5236 15316 5246
rect 15036 4340 15092 5180
rect 15260 5122 15316 5180
rect 15260 5070 15262 5122
rect 15314 5070 15316 5122
rect 15260 5058 15316 5070
rect 15372 5012 15428 5022
rect 15372 4394 15428 4956
rect 15372 4342 15374 4394
rect 15426 4342 15428 4394
rect 15372 4330 15428 4342
rect 15036 3778 15092 4284
rect 15036 3726 15038 3778
rect 15090 3726 15092 3778
rect 15036 3714 15092 3726
rect 14700 3502 14702 3554
rect 14754 3502 14756 3554
rect 14700 3490 14756 3502
rect 15372 3556 15428 3566
rect 15484 3556 15540 6076
rect 15708 5908 15764 5918
rect 15708 5814 15764 5852
rect 16044 5906 16100 5918
rect 16044 5854 16046 5906
rect 16098 5854 16100 5906
rect 16044 5796 16100 5854
rect 15596 5738 15652 5750
rect 15596 5686 15598 5738
rect 15650 5686 15652 5738
rect 16044 5730 16100 5740
rect 16380 5794 16436 6076
rect 16492 5921 16548 5946
rect 16492 5908 16494 5921
rect 16546 5908 16548 5921
rect 16492 5842 16548 5852
rect 16828 5906 16884 5918
rect 16828 5854 16830 5906
rect 16882 5854 16884 5906
rect 16380 5742 16382 5794
rect 16434 5742 16436 5794
rect 16380 5730 16436 5742
rect 16828 5796 16884 5854
rect 17612 5906 17668 6300
rect 17612 5854 17614 5906
rect 17666 5854 17668 5906
rect 18060 5962 18116 7308
rect 18172 6690 18228 8652
rect 18284 8036 18340 9662
rect 18732 9770 18788 9782
rect 18732 9718 18734 9770
rect 18786 9718 18788 9770
rect 18844 9736 18846 9772
rect 18898 9736 18900 9772
rect 18844 9724 18900 9736
rect 18732 9278 18788 9718
rect 18676 9266 18788 9278
rect 18676 9214 18678 9266
rect 18730 9214 18788 9266
rect 18676 9212 18788 9214
rect 18676 9202 18732 9212
rect 18508 9042 18564 9054
rect 18956 9044 19012 10556
rect 19404 9940 19460 11676
rect 19516 11506 19572 12014
rect 20804 12068 20860 12078
rect 20804 11974 20860 12012
rect 21252 12066 21308 12078
rect 21252 12014 21254 12066
rect 21306 12014 21308 12066
rect 19516 11454 19518 11506
rect 19570 11454 19572 11506
rect 19516 11442 19572 11454
rect 20188 11956 20244 11966
rect 19628 11396 19684 11406
rect 19628 10500 19684 11340
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19404 9874 19460 9884
rect 19572 10444 19684 10500
rect 19852 10500 19908 10510
rect 19572 9882 19628 10444
rect 19852 10406 19908 10444
rect 20188 10052 20244 11900
rect 20300 11844 20356 11854
rect 20300 11394 20356 11788
rect 21252 11844 21308 12014
rect 21252 11778 21308 11788
rect 21420 11956 21476 11966
rect 20692 11564 20748 11574
rect 20692 11562 21364 11564
rect 20692 11510 20694 11562
rect 20746 11510 21364 11562
rect 20692 11508 21364 11510
rect 20692 11498 20748 11508
rect 21308 11450 21364 11508
rect 20300 11342 20302 11394
rect 20354 11342 20356 11394
rect 20300 11330 20356 11342
rect 20524 11394 20580 11406
rect 20524 11342 20526 11394
rect 20578 11342 20580 11394
rect 21308 11398 21310 11450
rect 21362 11398 21364 11450
rect 21308 11386 21364 11398
rect 20524 10500 20580 11342
rect 21420 11356 21476 11900
rect 21420 11304 21422 11356
rect 21474 11304 21476 11356
rect 21700 11954 21756 11966
rect 21700 11902 21702 11954
rect 21754 11902 21756 11954
rect 21700 11396 21756 11902
rect 21868 11956 21924 12796
rect 22036 12786 22092 12796
rect 22204 12628 22260 13356
rect 22092 12572 22260 12628
rect 22316 13188 22372 13198
rect 22764 13188 22820 15932
rect 22988 15204 23044 15214
rect 22988 14530 23044 15148
rect 22988 14478 22990 14530
rect 23042 14478 23044 14530
rect 22988 14466 23044 14478
rect 22932 13972 22988 13982
rect 22932 13878 22988 13916
rect 23100 13412 23156 16044
rect 23212 16034 23268 16044
rect 23324 16098 23380 16110
rect 23324 16046 23326 16098
rect 23378 16046 23380 16098
rect 23324 15764 23380 16046
rect 23212 15708 23380 15764
rect 23212 15204 23268 15708
rect 23324 15540 23380 15550
rect 23324 15204 23380 15484
rect 23436 15428 23492 16716
rect 23436 15362 23492 15372
rect 23436 15204 23492 15214
rect 23324 15202 23492 15204
rect 23324 15150 23438 15202
rect 23490 15150 23492 15202
rect 23324 15148 23492 15150
rect 23212 15138 23268 15148
rect 23436 15138 23492 15148
rect 23324 14868 23380 14878
rect 23324 14754 23380 14812
rect 23324 14702 23326 14754
rect 23378 14702 23380 14754
rect 23324 14690 23380 14702
rect 23548 13636 23604 17052
rect 23716 17042 23772 17052
rect 23996 16996 24052 17006
rect 24220 16996 24276 18398
rect 24388 18396 24444 18452
rect 24388 18386 24500 18396
rect 24388 18004 24444 18386
rect 24500 18228 24556 18238
rect 24500 18226 24724 18228
rect 24500 18174 24502 18226
rect 24554 18174 24724 18226
rect 24500 18172 24724 18174
rect 24500 18162 24556 18172
rect 24388 17778 24444 17948
rect 24388 17726 24390 17778
rect 24442 17726 24444 17778
rect 24388 17714 24444 17726
rect 24332 17220 24388 17230
rect 24332 17106 24388 17164
rect 24332 17054 24334 17106
rect 24386 17054 24388 17106
rect 24332 17042 24388 17054
rect 24052 16940 24276 16996
rect 23660 16884 23716 16894
rect 23884 16884 23940 16894
rect 23716 16828 23828 16884
rect 23660 16818 23716 16828
rect 23772 15988 23828 16828
rect 23884 16212 23940 16828
rect 23996 16882 24052 16940
rect 23996 16830 23998 16882
rect 24050 16830 24052 16882
rect 23996 16818 24052 16830
rect 23884 16146 23940 16156
rect 23772 15932 23940 15988
rect 23660 15874 23716 15886
rect 23660 15822 23662 15874
rect 23714 15822 23716 15874
rect 23660 15316 23716 15822
rect 23772 15316 23828 15326
rect 23660 15314 23828 15316
rect 23660 15262 23774 15314
rect 23826 15262 23828 15314
rect 23660 15260 23828 15262
rect 23772 15148 23828 15260
rect 23884 15314 23940 15932
rect 23884 15262 23886 15314
rect 23938 15262 23940 15314
rect 23884 15250 23940 15262
rect 24556 15874 24612 15886
rect 24556 15822 24558 15874
rect 24610 15822 24612 15874
rect 23660 15092 23828 15148
rect 24220 15092 24276 15102
rect 23660 14532 23716 15092
rect 24220 14998 24276 15036
rect 24556 14980 24612 15822
rect 24668 15148 24724 18172
rect 24780 17890 24836 18956
rect 24780 17838 24782 17890
rect 24834 17838 24836 17890
rect 24780 17826 24836 17838
rect 24892 18956 25172 19012
rect 24892 16098 24948 18956
rect 25340 18900 25396 18910
rect 25340 18494 25396 18844
rect 25340 18442 25342 18494
rect 25394 18442 25396 18494
rect 25340 18430 25396 18442
rect 25564 18450 25620 19180
rect 25676 19234 25732 19292
rect 25676 19182 25678 19234
rect 25730 19182 25732 19234
rect 25676 19170 25732 19182
rect 26124 19236 26180 19246
rect 26348 19236 26404 19246
rect 26124 19142 26180 19180
rect 26236 19234 26404 19236
rect 26236 19182 26350 19234
rect 26402 19182 26404 19234
rect 26236 19180 26404 19182
rect 25844 19012 25900 19022
rect 26236 19012 26292 19180
rect 26348 19170 26404 19180
rect 25844 19010 26292 19012
rect 25844 18958 25846 19010
rect 25898 18958 26292 19010
rect 25844 18956 26292 18958
rect 25844 18946 25900 18956
rect 25564 18398 25566 18450
rect 25618 18398 25620 18450
rect 25564 18386 25620 18398
rect 26236 18452 26292 18956
rect 26460 18788 26516 19404
rect 26460 18722 26516 18732
rect 26628 19122 26684 19134
rect 26628 19070 26630 19122
rect 26682 19070 26684 19122
rect 26628 18564 26684 19070
rect 26460 18508 26684 18564
rect 26796 18564 26852 18574
rect 26236 18386 26292 18396
rect 26348 18450 26404 18462
rect 26348 18398 26350 18450
rect 26402 18398 26404 18450
rect 25228 18338 25284 18350
rect 25228 18286 25230 18338
rect 25282 18286 25284 18338
rect 25228 18116 25284 18286
rect 25228 18050 25284 18060
rect 26068 18226 26124 18238
rect 26068 18174 26070 18226
rect 26122 18174 26124 18226
rect 26068 17892 26124 18174
rect 26068 17826 26124 17836
rect 26236 18228 26292 18238
rect 25116 17666 25172 17678
rect 25116 17614 25118 17666
rect 25170 17614 25172 17666
rect 25116 17108 25172 17614
rect 25116 17042 25172 17052
rect 25228 17668 25284 17678
rect 24892 16046 24894 16098
rect 24946 16046 24948 16098
rect 24892 16034 24948 16046
rect 25004 16324 25060 16334
rect 25004 16098 25060 16268
rect 25004 16046 25006 16098
rect 25058 16046 25060 16098
rect 25004 15988 25060 16046
rect 25004 15922 25060 15932
rect 25228 15316 25284 17612
rect 25452 17666 25508 17678
rect 25452 17614 25454 17666
rect 25506 17614 25508 17666
rect 25340 17444 25396 17454
rect 25340 17106 25396 17388
rect 25452 17220 25508 17614
rect 25452 17154 25508 17164
rect 25732 17554 25788 17566
rect 25732 17502 25734 17554
rect 25786 17502 25788 17554
rect 25732 17220 25788 17502
rect 25732 17154 25788 17164
rect 25900 17556 25956 17566
rect 25340 17054 25342 17106
rect 25394 17054 25396 17106
rect 25340 17042 25396 17054
rect 25900 16996 25956 17500
rect 25788 16940 25956 16996
rect 26124 17108 26180 17118
rect 25676 16884 25732 16894
rect 25564 16828 25676 16884
rect 25452 16548 25508 16558
rect 25228 15250 25284 15260
rect 25340 16324 25396 16334
rect 25452 16324 25508 16492
rect 25340 16322 25508 16324
rect 25340 16270 25342 16322
rect 25394 16270 25508 16322
rect 25340 16268 25508 16270
rect 25340 15148 25396 16268
rect 24668 15092 25060 15148
rect 23996 14756 24052 14766
rect 23996 14662 24052 14700
rect 24332 14532 24388 14542
rect 23660 14530 24388 14532
rect 23660 14478 23662 14530
rect 23714 14478 24334 14530
rect 24386 14478 24388 14530
rect 23660 14476 24388 14478
rect 23660 14466 23716 14476
rect 23436 13580 23604 13636
rect 24108 13972 24164 13982
rect 23436 13412 23492 13580
rect 23884 13524 23940 13534
rect 23100 13346 23156 13356
rect 23324 13356 23492 13412
rect 23548 13522 23940 13524
rect 23548 13470 23886 13522
rect 23938 13470 23940 13522
rect 23548 13468 23940 13470
rect 22092 12292 22148 12572
rect 22316 12516 22372 13132
rect 22652 13132 22820 13188
rect 22092 12198 22148 12236
rect 22260 12460 22372 12516
rect 22484 12850 22540 12862
rect 22484 12798 22486 12850
rect 22538 12798 22540 12850
rect 22260 12234 22316 12460
rect 22484 12404 22540 12798
rect 22484 12338 22540 12348
rect 21980 12180 22036 12190
rect 22260 12182 22262 12234
rect 22314 12182 22316 12234
rect 22260 12170 22316 12182
rect 22428 12178 22484 12190
rect 21980 12086 22036 12124
rect 22428 12126 22430 12178
rect 22482 12126 22484 12178
rect 22428 12068 22484 12126
rect 22652 12180 22708 13132
rect 22876 13076 22932 13086
rect 22764 12964 22820 12974
rect 22764 12870 22820 12908
rect 22876 12962 22932 13020
rect 22876 12910 22878 12962
rect 22930 12910 22932 12962
rect 23212 12962 23268 12974
rect 22876 12628 22932 12910
rect 23044 12906 23100 12918
rect 23044 12854 23046 12906
rect 23098 12854 23100 12906
rect 23044 12852 23100 12854
rect 23044 12786 23100 12796
rect 23212 12910 23214 12962
rect 23266 12910 23268 12962
rect 23212 12740 23268 12910
rect 23324 12964 23380 13356
rect 23324 12898 23380 12908
rect 23436 13188 23492 13198
rect 23436 12962 23492 13132
rect 23436 12910 23438 12962
rect 23490 12910 23492 12962
rect 23436 12898 23492 12910
rect 23548 12964 23604 13468
rect 23884 13458 23940 13468
rect 23548 12740 23604 12908
rect 23772 12740 23828 12750
rect 23212 12684 23604 12740
rect 22876 12572 23268 12628
rect 23212 12290 23268 12572
rect 23212 12238 23214 12290
rect 23266 12238 23268 12290
rect 23212 12226 23268 12238
rect 23380 12292 23436 12302
rect 23380 12234 23436 12236
rect 23100 12180 23156 12190
rect 22652 12124 23044 12180
rect 22428 12002 22484 12012
rect 22820 11956 22876 11966
rect 21868 11900 22204 11956
rect 21700 11330 21756 11340
rect 21868 11732 21924 11742
rect 21420 11292 21476 11304
rect 21756 10836 21812 10846
rect 21756 10610 21812 10780
rect 21756 10558 21758 10610
rect 21810 10558 21812 10610
rect 21756 10546 21812 10558
rect 21868 10612 21924 11676
rect 22148 11450 22204 11900
rect 22764 11954 22876 11956
rect 22764 11902 22822 11954
rect 22874 11902 22876 11954
rect 22764 11890 22876 11902
rect 22596 11844 22652 11854
rect 22148 11398 22150 11450
rect 22202 11398 22204 11450
rect 22148 11386 22204 11398
rect 22428 11732 22484 11742
rect 22428 11394 22484 11676
rect 22596 11618 22652 11788
rect 22596 11566 22598 11618
rect 22650 11566 22652 11618
rect 22596 11554 22652 11566
rect 22428 11342 22430 11394
rect 22482 11342 22484 11394
rect 22428 11330 22484 11342
rect 21980 11282 22036 11294
rect 21980 11230 21982 11282
rect 22034 11230 22036 11282
rect 21980 10836 22036 11230
rect 21980 10770 22036 10780
rect 22540 10612 22596 10622
rect 21868 10610 22596 10612
rect 21868 10558 22542 10610
rect 22594 10558 22596 10610
rect 21868 10556 22596 10558
rect 20524 10434 20580 10444
rect 19572 9830 19574 9882
rect 19626 9830 19628 9882
rect 19572 9818 19628 9830
rect 20076 9996 20244 10052
rect 20804 10164 20860 10174
rect 20076 9828 20132 9996
rect 20804 9882 20860 10108
rect 20412 9828 20468 9838
rect 20076 9736 20078 9772
rect 20130 9736 20132 9772
rect 18508 8990 18510 9042
rect 18562 8990 18564 9042
rect 18508 8036 18564 8990
rect 18284 7980 18378 8036
rect 18322 7511 18378 7980
rect 18508 7970 18564 7980
rect 18620 8988 19012 9044
rect 19404 9714 19460 9726
rect 20076 9724 20132 9736
rect 20188 9826 20468 9828
rect 20188 9774 20414 9826
rect 20466 9774 20468 9826
rect 20804 9830 20806 9882
rect 20858 9830 20860 9882
rect 20804 9818 20860 9830
rect 20188 9772 20468 9774
rect 19404 9662 19406 9714
rect 19458 9662 19460 9714
rect 18322 7459 18324 7511
rect 18376 7459 18378 7511
rect 18322 7364 18378 7459
rect 18322 7298 18378 7308
rect 18508 7474 18564 7486
rect 18508 7422 18510 7474
rect 18562 7422 18564 7474
rect 18508 7028 18564 7422
rect 18620 7474 18676 8988
rect 19292 8930 19348 8942
rect 19292 8878 19294 8930
rect 19346 8878 19348 8930
rect 19292 8820 19348 8878
rect 18732 8764 19348 8820
rect 18732 8148 18788 8764
rect 19404 8484 19460 9662
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 20188 9268 20244 9772
rect 20412 9762 20468 9772
rect 20636 9714 20692 9726
rect 20636 9662 20638 9714
rect 20690 9662 20692 9714
rect 20636 9380 20692 9662
rect 21476 9604 21532 9614
rect 21868 9604 21924 10556
rect 22540 10546 22596 10556
rect 22652 10164 22708 10174
rect 22764 10164 22820 11890
rect 22708 10108 22820 10164
rect 22988 10836 23044 12124
rect 23100 12086 23156 12124
rect 23380 12182 23382 12234
rect 23434 12182 23436 12234
rect 23380 11844 23436 12182
rect 23548 12178 23604 12684
rect 23548 12126 23550 12178
rect 23602 12126 23604 12178
rect 23548 12068 23604 12126
rect 23548 12002 23604 12012
rect 23660 12684 23772 12740
rect 23380 11778 23436 11788
rect 23156 11732 23212 11742
rect 23156 11506 23212 11676
rect 23156 11454 23158 11506
rect 23210 11454 23212 11506
rect 23156 11442 23212 11454
rect 23100 10836 23156 10846
rect 22988 10834 23156 10836
rect 22988 10782 23102 10834
rect 23154 10782 23156 10834
rect 22988 10780 23156 10782
rect 22652 10098 22708 10108
rect 22540 9940 22596 9950
rect 22428 9828 22484 9838
rect 22428 9734 22484 9772
rect 22540 9826 22596 9884
rect 22540 9774 22542 9826
rect 22594 9774 22596 9826
rect 22708 9940 22764 9950
rect 22708 9882 22764 9884
rect 22708 9830 22710 9882
rect 22762 9830 22764 9882
rect 22708 9818 22764 9830
rect 22876 9828 22932 9838
rect 22988 9828 23044 10780
rect 23100 10770 23156 10780
rect 23436 10610 23492 10622
rect 23436 10558 23438 10610
rect 23490 10558 23492 10610
rect 23436 10164 23492 10558
rect 23436 10098 23492 10108
rect 23660 10052 23716 12684
rect 23772 12646 23828 12684
rect 23996 12516 24052 12526
rect 23996 12404 24052 12460
rect 23884 12402 24052 12404
rect 23884 12350 23998 12402
rect 24050 12350 24052 12402
rect 23884 12348 24052 12350
rect 23772 11956 23828 11966
rect 23772 10948 23828 11900
rect 23772 10882 23828 10892
rect 23660 9986 23716 9996
rect 23380 9940 23436 9950
rect 23884 9940 23940 12348
rect 23996 12338 24052 12348
rect 24108 11564 24164 13916
rect 24220 13746 24276 14476
rect 24332 14466 24388 14476
rect 24220 13694 24222 13746
rect 24274 13694 24276 13746
rect 24220 13682 24276 13694
rect 24556 13636 24612 14924
rect 24668 14532 24724 14542
rect 24668 14438 24724 14476
rect 24780 13972 24836 13982
rect 24556 13580 24668 13636
rect 24444 12964 24500 12974
rect 24444 12870 24500 12908
rect 24612 12906 24668 13580
rect 24332 12852 24388 12862
rect 24332 12178 24388 12796
rect 24612 12854 24614 12906
rect 24666 12854 24668 12906
rect 24780 12962 24836 13916
rect 24780 12910 24782 12962
rect 24834 12910 24836 12962
rect 24780 12898 24836 12910
rect 24892 13076 24948 13086
rect 24892 12962 24948 13020
rect 24892 12910 24894 12962
rect 24946 12910 24948 12962
rect 24892 12898 24948 12910
rect 24612 12852 24668 12854
rect 24612 12786 24668 12796
rect 24332 12126 24334 12178
rect 24386 12126 24388 12178
rect 24332 12114 24388 12126
rect 24780 12180 24836 12190
rect 24108 11508 24276 11564
rect 24052 11396 24108 11406
rect 24052 11302 24108 11340
rect 24220 10388 24276 11508
rect 24500 11508 24556 11518
rect 24500 11450 24556 11452
rect 24332 11396 24388 11406
rect 24500 11398 24502 11450
rect 24554 11398 24556 11450
rect 24500 11386 24556 11398
rect 24780 11394 24836 12124
rect 25004 11732 25060 15092
rect 25228 15092 25396 15148
rect 25452 16100 25508 16110
rect 25228 14756 25284 15092
rect 25116 14700 25284 14756
rect 25116 13524 25172 14700
rect 25228 14532 25284 14542
rect 25228 13746 25284 14476
rect 25452 14084 25508 16044
rect 25564 14980 25620 16828
rect 25676 16790 25732 16828
rect 25788 15242 25844 16940
rect 26124 16882 26180 17052
rect 26124 16830 26126 16882
rect 26178 16830 26180 16882
rect 26124 16818 26180 16830
rect 26236 16884 26292 18172
rect 26348 17220 26404 18398
rect 26460 18450 26516 18508
rect 26460 18398 26462 18450
rect 26514 18398 26516 18450
rect 26796 18450 26852 18508
rect 26460 18228 26516 18398
rect 26628 18394 26684 18406
rect 26628 18342 26630 18394
rect 26682 18342 26684 18394
rect 26796 18398 26798 18450
rect 26850 18398 26852 18450
rect 26796 18386 26852 18398
rect 26628 18340 26684 18342
rect 26628 18274 26684 18284
rect 26460 18162 26516 18172
rect 26796 18116 26852 18126
rect 26460 18004 26516 18014
rect 26460 17666 26516 17948
rect 26460 17614 26462 17666
rect 26514 17614 26516 17666
rect 26460 17602 26516 17614
rect 26628 18004 26684 18014
rect 26628 17610 26684 17948
rect 26628 17558 26630 17610
rect 26682 17558 26684 17610
rect 26628 17556 26684 17558
rect 26628 17490 26684 17500
rect 26796 17666 26852 18060
rect 26908 18004 26964 20524
rect 27020 20244 27076 20254
rect 27020 19460 27076 20188
rect 28028 20244 28084 20254
rect 27132 20132 27188 20142
rect 27132 20038 27188 20076
rect 28028 20020 28084 20188
rect 28420 20244 28476 20254
rect 28420 20150 28476 20188
rect 28868 20244 28924 20254
rect 28868 20150 28924 20188
rect 28028 19926 28084 19964
rect 27692 19794 27748 19806
rect 27692 19742 27694 19794
rect 27746 19742 27748 19794
rect 27132 19460 27188 19470
rect 27020 19458 27188 19460
rect 27020 19406 27134 19458
rect 27186 19406 27188 19458
rect 27020 19404 27188 19406
rect 27132 19394 27188 19404
rect 27468 19234 27524 19246
rect 27468 19182 27470 19234
rect 27522 19182 27524 19234
rect 27020 18452 27076 18462
rect 27020 18358 27076 18396
rect 27468 18340 27524 19182
rect 27692 19236 27748 19742
rect 27692 19170 27748 19180
rect 27860 19348 27916 19358
rect 27860 19012 27916 19292
rect 27860 18918 27916 18956
rect 28140 19236 28196 19246
rect 28140 18450 28196 19180
rect 29036 19236 29092 19246
rect 29148 19236 29204 21532
rect 29372 21586 29428 21598
rect 29372 21534 29374 21586
rect 29426 21534 29428 21586
rect 29372 21476 29428 21534
rect 29372 21410 29428 21420
rect 29372 21028 29428 21038
rect 29484 21028 29540 21756
rect 29820 21746 29876 21756
rect 30380 22370 30436 22382
rect 30380 22318 30382 22370
rect 30434 22318 30436 22370
rect 29708 21588 29764 21598
rect 29708 21494 29764 21532
rect 29372 21026 29540 21028
rect 29372 20974 29374 21026
rect 29426 20974 29540 21026
rect 29372 20972 29540 20974
rect 29372 20962 29428 20972
rect 30268 20020 30324 20030
rect 29932 20018 30324 20020
rect 29932 19966 30270 20018
rect 30322 19966 30324 20018
rect 29932 19964 30324 19966
rect 29036 19234 29204 19236
rect 29036 19182 29038 19234
rect 29090 19182 29204 19234
rect 29036 19180 29204 19182
rect 29820 19236 29876 19246
rect 28308 19012 28364 19022
rect 28308 18918 28364 18956
rect 27972 18396 28028 18406
rect 26908 17938 26964 17948
rect 27356 18226 27412 18238
rect 27356 18174 27358 18226
rect 27410 18174 27412 18226
rect 26796 17614 26798 17666
rect 26850 17614 26852 17666
rect 26348 17154 26404 17164
rect 26684 17108 26740 17118
rect 26460 17052 26684 17108
rect 26348 16884 26404 16894
rect 26236 16828 26348 16884
rect 26348 16790 26404 16828
rect 25956 16658 26012 16670
rect 25956 16606 25958 16658
rect 26010 16606 26012 16658
rect 25956 16324 26012 16606
rect 25956 16258 26012 16268
rect 26348 16660 26404 16670
rect 26236 16100 26292 16110
rect 26068 15876 26124 15886
rect 26068 15782 26124 15820
rect 26236 15652 26292 16044
rect 25732 15204 25844 15242
rect 25788 15148 25844 15204
rect 26012 15596 26292 15652
rect 25732 15138 25788 15148
rect 25564 14914 25620 14924
rect 25900 15092 25956 15102
rect 25900 14530 25956 15036
rect 25900 14478 25902 14530
rect 25954 14478 25956 14530
rect 25452 14018 25508 14028
rect 25732 14306 25788 14318
rect 25732 14254 25734 14306
rect 25786 14254 25788 14306
rect 25732 14084 25788 14254
rect 25732 14018 25788 14028
rect 25340 13972 25396 13982
rect 25340 13860 25396 13916
rect 25900 13972 25956 14478
rect 25900 13906 25956 13916
rect 25340 13804 25582 13860
rect 25228 13694 25230 13746
rect 25282 13694 25284 13746
rect 25526 13758 25582 13804
rect 25526 13746 25620 13758
rect 25228 13682 25284 13694
rect 25396 13690 25452 13702
rect 25526 13694 25566 13746
rect 25618 13694 25620 13746
rect 25526 13692 25620 13694
rect 25396 13638 25398 13690
rect 25450 13638 25452 13690
rect 25564 13682 25620 13692
rect 25676 13746 25732 13758
rect 26012 13748 26068 15596
rect 26348 15540 26404 16604
rect 26180 15484 26404 15540
rect 26180 15426 26236 15484
rect 26180 15374 26182 15426
rect 26234 15374 26236 15426
rect 26180 15148 26236 15374
rect 26180 15092 26404 15148
rect 25676 13694 25678 13746
rect 25730 13694 25732 13746
rect 25396 13524 25452 13638
rect 25116 13468 25284 13524
rect 25228 13188 25284 13468
rect 25396 13458 25452 13468
rect 25564 13412 25620 13422
rect 25228 13132 25396 13188
rect 25172 12964 25228 12974
rect 25172 12870 25228 12908
rect 25004 11676 25172 11732
rect 25116 11508 25172 11676
rect 25116 11452 25284 11508
rect 24332 11302 24388 11340
rect 24780 11342 24782 11394
rect 24834 11342 24836 11394
rect 24780 11330 24836 11342
rect 24668 11282 24724 11294
rect 25060 11284 25116 11294
rect 24668 11230 24670 11282
rect 24722 11230 24724 11282
rect 24668 10836 24724 11230
rect 25004 11282 25116 11284
rect 25004 11230 25062 11282
rect 25114 11230 25116 11282
rect 25004 11218 25116 11230
rect 24780 10836 24836 10846
rect 24668 10780 24780 10836
rect 24780 10610 24836 10780
rect 24780 10558 24782 10610
rect 24834 10558 24836 10610
rect 24780 10546 24836 10558
rect 24220 10322 24276 10332
rect 24444 10386 24500 10398
rect 24444 10334 24446 10386
rect 24498 10334 24500 10386
rect 23380 9882 23436 9884
rect 23212 9828 23268 9838
rect 22876 9826 23268 9828
rect 22148 9716 22204 9726
rect 22540 9716 22596 9774
rect 22876 9774 22878 9826
rect 22930 9774 23214 9826
rect 23266 9774 23268 9826
rect 23380 9830 23382 9882
rect 23434 9830 23436 9882
rect 23772 9884 23884 9940
rect 23380 9818 23436 9830
rect 23660 9828 23716 9838
rect 22876 9772 23268 9774
rect 22876 9762 22932 9772
rect 23212 9762 23268 9772
rect 23660 9734 23716 9772
rect 22148 9714 22372 9716
rect 22148 9662 22150 9714
rect 22202 9662 22372 9714
rect 22148 9660 22372 9662
rect 22148 9650 22204 9660
rect 21476 9602 21924 9604
rect 21476 9550 21478 9602
rect 21530 9550 21924 9602
rect 21476 9548 21924 9550
rect 21476 9538 21532 9548
rect 20636 9324 21252 9380
rect 20076 9212 20244 9268
rect 20076 8708 20132 9212
rect 21196 9042 21252 9324
rect 21196 8990 21198 9042
rect 21250 8990 21252 9042
rect 21196 8978 21252 8990
rect 21868 9044 21924 9548
rect 22316 9268 22372 9660
rect 22540 9650 22596 9660
rect 23548 9716 23604 9726
rect 23548 9622 23604 9660
rect 22988 9604 23044 9614
rect 22316 9212 22596 9268
rect 21980 9044 22036 9054
rect 22372 9044 22428 9054
rect 21868 9042 22428 9044
rect 21868 8990 21982 9042
rect 22034 8990 22374 9042
rect 22426 8990 22428 9042
rect 21868 8988 22428 8990
rect 21980 8978 22036 8988
rect 22316 8978 22428 8988
rect 21252 8820 21308 8830
rect 20076 8652 20524 8708
rect 19404 8418 19460 8428
rect 20132 8484 20188 8494
rect 18844 8260 18900 8270
rect 19236 8260 19292 8270
rect 19684 8260 19740 8270
rect 20132 8260 20188 8428
rect 20468 8482 20524 8652
rect 20468 8430 20470 8482
rect 20522 8430 20524 8482
rect 20468 8418 20524 8430
rect 21252 8314 21308 8764
rect 18844 8258 20188 8260
rect 18844 8206 18846 8258
rect 18898 8206 19238 8258
rect 19290 8206 19686 8258
rect 19738 8206 20134 8258
rect 20186 8206 20188 8258
rect 18844 8204 20188 8206
rect 18844 8194 18900 8204
rect 19236 8194 19292 8204
rect 18732 8082 18788 8092
rect 18620 7422 18622 7474
rect 18674 7422 18676 7474
rect 18620 7410 18676 7422
rect 19180 7476 19236 7486
rect 18508 6972 18900 7028
rect 18508 6804 18564 6814
rect 18172 6638 18174 6690
rect 18226 6638 18228 6690
rect 18172 6626 18228 6638
rect 18284 6802 18564 6804
rect 18284 6750 18510 6802
rect 18562 6750 18564 6802
rect 18284 6748 18564 6750
rect 18060 5910 18062 5962
rect 18114 5910 18116 5962
rect 18060 5898 18116 5910
rect 18284 5906 18340 6748
rect 18508 6738 18564 6748
rect 18732 6692 18788 6702
rect 18620 6690 18788 6692
rect 18508 6634 18564 6646
rect 18396 6580 18452 6590
rect 18396 6074 18452 6524
rect 18508 6582 18510 6634
rect 18562 6582 18564 6634
rect 18508 6468 18564 6582
rect 18508 6402 18564 6412
rect 18620 6638 18734 6690
rect 18786 6638 18788 6690
rect 18620 6636 18788 6638
rect 18396 6022 18398 6074
rect 18450 6022 18452 6074
rect 18396 6010 18452 6022
rect 17612 5842 17668 5854
rect 18284 5854 18286 5906
rect 18338 5854 18340 5906
rect 18284 5842 18340 5854
rect 16828 5730 16884 5740
rect 18172 5796 18228 5806
rect 15596 4394 15652 5686
rect 17164 5236 17220 5246
rect 16044 5124 16100 5134
rect 16044 5122 16212 5124
rect 16044 5070 16046 5122
rect 16098 5070 16212 5122
rect 16044 5068 16212 5070
rect 16044 5058 16100 5068
rect 15596 4342 15598 4394
rect 15650 4342 15652 4394
rect 15596 4330 15652 4342
rect 16044 4452 16100 4462
rect 16044 4394 16100 4396
rect 16044 4342 16046 4394
rect 16098 4342 16100 4394
rect 16044 4330 16100 4342
rect 16156 4228 16212 5068
rect 16354 4396 16548 4452
rect 16354 4378 16410 4396
rect 16354 4326 16356 4378
rect 16408 4326 16410 4378
rect 16354 4314 16410 4326
rect 16380 4228 16436 4238
rect 16156 4226 16436 4228
rect 16156 4174 16382 4226
rect 16434 4174 16436 4226
rect 16156 4172 16436 4174
rect 16380 4162 16436 4172
rect 16492 4004 16548 4396
rect 16380 3948 16548 4004
rect 15372 3554 15540 3556
rect 15372 3502 15374 3554
rect 15426 3502 15540 3554
rect 15372 3500 15540 3502
rect 16044 3780 16100 3790
rect 16044 3554 16100 3724
rect 16380 3722 16436 3948
rect 16380 3670 16382 3722
rect 16434 3670 16436 3722
rect 16380 3658 16436 3670
rect 17164 3678 17220 5180
rect 17948 5124 18004 5134
rect 17444 4506 17500 4518
rect 17444 4454 17446 4506
rect 17498 4454 17500 4506
rect 17444 4452 17500 4454
rect 17444 4386 17500 4396
rect 17276 4340 17332 4350
rect 17276 4246 17332 4284
rect 17948 4338 18004 5068
rect 17948 4286 17950 4338
rect 18002 4286 18004 4338
rect 17164 3666 17276 3678
rect 17164 3614 17222 3666
rect 17274 3614 17276 3666
rect 17164 3612 17276 3614
rect 17220 3602 17276 3612
rect 17836 3668 17892 3678
rect 16044 3502 16046 3554
rect 16098 3502 16100 3554
rect 15372 3490 15428 3500
rect 16044 3490 16100 3502
rect 16268 3556 16324 3566
rect 12628 3444 12684 3482
rect 16268 3462 16324 3500
rect 17556 3556 17612 3566
rect 17556 3462 17612 3500
rect 17836 3554 17892 3612
rect 17836 3502 17838 3554
rect 17890 3502 17892 3554
rect 17836 3490 17892 3502
rect 17948 3554 18004 4286
rect 17948 3502 17950 3554
rect 18002 3502 18004 3554
rect 17948 3490 18004 3502
rect 12628 3378 12684 3388
rect 18172 3444 18228 5740
rect 18620 5460 18676 6636
rect 18732 6626 18788 6636
rect 18844 6692 18900 6972
rect 18844 6626 18900 6636
rect 18396 5404 18676 5460
rect 18732 5908 18788 5918
rect 18284 5012 18340 5022
rect 18284 4382 18340 4956
rect 18284 4330 18286 4382
rect 18338 4330 18340 4382
rect 18284 4318 18340 4330
rect 18396 4226 18452 5404
rect 18508 5236 18564 5246
rect 18732 5236 18788 5852
rect 18956 5794 19012 5806
rect 18956 5742 18958 5794
rect 19010 5742 19012 5794
rect 18956 5348 19012 5742
rect 18956 5282 19012 5292
rect 18508 5234 18788 5236
rect 18508 5182 18510 5234
rect 18562 5182 18788 5234
rect 18508 5180 18788 5182
rect 18508 5170 18564 5180
rect 18900 5124 18956 5134
rect 18900 5030 18956 5068
rect 19068 5124 19124 5134
rect 19068 5030 19124 5068
rect 19180 5122 19236 7420
rect 19684 7364 19740 8204
rect 20132 8194 20188 8204
rect 20300 8258 20356 8270
rect 20300 8206 20302 8258
rect 20354 8206 20356 8258
rect 21252 8262 21254 8314
rect 21306 8262 21308 8314
rect 21980 8484 22036 8494
rect 21252 8250 21308 8262
rect 21868 8260 21924 8270
rect 20300 8148 20356 8206
rect 21868 8178 21870 8204
rect 21922 8178 21924 8204
rect 21868 8166 21924 8178
rect 20300 8082 20356 8092
rect 21420 8146 21476 8158
rect 21420 8094 21422 8146
rect 21474 8094 21476 8146
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 21420 7812 21476 8094
rect 21980 8036 22036 8428
rect 22316 8484 22372 8978
rect 22316 8258 22372 8428
rect 19836 7802 20100 7812
rect 21084 7756 21476 7812
rect 21868 7980 22036 8036
rect 22092 8202 22148 8214
rect 22092 8150 22094 8202
rect 22146 8150 22148 8202
rect 22316 8206 22318 8258
rect 22370 8206 22372 8258
rect 22316 8194 22372 8206
rect 21084 7474 21140 7756
rect 21084 7422 21086 7474
rect 21138 7422 21140 7474
rect 21084 7410 21140 7422
rect 21868 7474 21924 7980
rect 22092 7710 22148 8150
rect 22092 7698 22204 7710
rect 22092 7646 22150 7698
rect 22202 7646 22204 7698
rect 22092 7644 22204 7646
rect 22148 7634 22204 7644
rect 21868 7422 21870 7474
rect 21922 7422 21924 7474
rect 19684 7308 20020 7364
rect 19964 6814 20020 7308
rect 19964 6802 20076 6814
rect 19964 6750 20022 6802
rect 20074 6750 20076 6802
rect 19964 6748 20076 6750
rect 19180 5070 19182 5122
rect 19234 5070 19236 5122
rect 19180 5058 19236 5070
rect 19292 6692 19348 6702
rect 19292 6466 19348 6636
rect 19628 6690 19684 6702
rect 19628 6638 19630 6690
rect 19682 6638 19684 6690
rect 19628 6580 19684 6638
rect 20020 6692 20076 6748
rect 20020 6626 20076 6636
rect 20468 6692 20524 6702
rect 21756 6692 21812 6702
rect 20468 6598 20524 6636
rect 21532 6634 21588 6646
rect 19628 6514 19684 6524
rect 21532 6582 21534 6634
rect 21586 6582 21588 6634
rect 21756 6610 21758 6636
rect 21810 6610 21812 6636
rect 21756 6598 21812 6610
rect 19292 6414 19294 6466
rect 19346 6414 19348 6466
rect 19292 5124 19348 6414
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 20860 5908 20916 5918
rect 20860 5814 20916 5852
rect 20300 5348 20356 5358
rect 19292 5058 19348 5068
rect 19516 5236 19572 5246
rect 18396 4174 18398 4226
rect 18450 4174 18452 4226
rect 18396 4162 18452 4174
rect 19068 4338 19124 4350
rect 19068 4286 19070 4338
rect 19122 4286 19124 4338
rect 19068 4228 19124 4286
rect 19292 4338 19348 4350
rect 19292 4286 19294 4338
rect 19346 4286 19348 4338
rect 19068 4162 19124 4172
rect 19180 4170 19236 4182
rect 19180 4118 19182 4170
rect 19234 4118 19236 4170
rect 18732 3892 18788 3902
rect 18396 3668 18452 3678
rect 18396 3574 18452 3612
rect 18732 3556 18788 3836
rect 18732 3462 18788 3500
rect 19180 3556 19236 4118
rect 19292 4116 19348 4286
rect 19516 4340 19572 5180
rect 19628 5234 19684 5246
rect 19628 5182 19630 5234
rect 19682 5182 19684 5234
rect 19628 4564 19684 5182
rect 20188 5124 20244 5134
rect 20020 5066 20076 5078
rect 20020 5014 20022 5066
rect 20074 5014 20076 5066
rect 20188 5030 20244 5068
rect 20300 5122 20356 5292
rect 21196 5348 21252 5358
rect 20804 5236 20860 5246
rect 20804 5142 20860 5180
rect 20300 5070 20302 5122
rect 20354 5070 20356 5122
rect 20300 5058 20356 5070
rect 21196 5122 21252 5292
rect 21364 5348 21420 5358
rect 21532 5348 21588 6582
rect 21364 5346 21588 5348
rect 21364 5294 21366 5346
rect 21418 5294 21588 5346
rect 21364 5292 21588 5294
rect 21644 5908 21700 5918
rect 21868 5908 21924 7422
rect 21980 7494 22036 7506
rect 21980 7476 21982 7494
rect 22034 7476 22036 7494
rect 21980 7402 22036 7420
rect 22540 7252 22596 9212
rect 22988 9266 23044 9548
rect 22988 9214 22990 9266
rect 23042 9214 23044 9266
rect 22988 9202 23044 9214
rect 22372 7196 22596 7252
rect 22652 9042 22708 9054
rect 22652 8990 22654 9042
rect 22706 8990 22708 9042
rect 22652 8932 22708 8990
rect 22372 6746 22428 7196
rect 22652 6916 22708 8876
rect 23772 8596 23828 9884
rect 23884 9874 23940 9884
rect 24220 10164 24276 10174
rect 24220 9826 24276 10108
rect 24220 9774 24222 9826
rect 24274 9774 24276 9826
rect 24220 9762 24276 9774
rect 23940 9716 23996 9726
rect 24444 9716 24500 10334
rect 23940 9714 24164 9716
rect 23940 9662 23942 9714
rect 23994 9662 24164 9714
rect 23940 9660 24164 9662
rect 23940 9650 23996 9660
rect 23940 8820 23996 8830
rect 23940 8726 23996 8764
rect 24108 8596 24164 9660
rect 24220 9604 24276 9614
rect 24444 9604 24500 9660
rect 24220 9042 24276 9548
rect 24388 9548 24500 9604
rect 24556 9604 24612 9614
rect 24556 9602 24724 9604
rect 24556 9550 24558 9602
rect 24610 9550 24724 9602
rect 24556 9548 24724 9550
rect 24388 9492 24444 9548
rect 24556 9538 24612 9548
rect 24332 9436 24444 9492
rect 24332 9154 24388 9436
rect 24332 9102 24334 9154
rect 24386 9102 24388 9154
rect 24332 9090 24388 9102
rect 24500 9268 24556 9278
rect 24500 9098 24556 9212
rect 24220 8990 24222 9042
rect 24274 8990 24276 9042
rect 24500 9046 24502 9098
rect 24554 9046 24556 9098
rect 24500 9034 24556 9046
rect 24668 9042 24724 9548
rect 24220 8978 24276 8990
rect 24668 8990 24670 9042
rect 24722 8990 24724 9042
rect 24108 8540 24276 8596
rect 23772 8530 23828 8540
rect 23100 8258 23156 8270
rect 23100 8206 23102 8258
rect 23154 8206 23156 8258
rect 23100 7700 23156 8206
rect 23100 7634 23156 7644
rect 23324 8260 23380 8270
rect 23324 7812 23380 8204
rect 22372 6694 22374 6746
rect 22426 6694 22428 6746
rect 22372 6682 22428 6694
rect 22540 6860 22708 6916
rect 21644 5906 21924 5908
rect 21644 5854 21646 5906
rect 21698 5854 21870 5906
rect 21922 5854 21924 5906
rect 21644 5852 21924 5854
rect 21364 5282 21420 5292
rect 21644 5236 21700 5852
rect 21868 5842 21924 5852
rect 22204 6578 22260 6590
rect 22204 6526 22206 6578
rect 22258 6526 22260 6578
rect 22204 5908 22260 6526
rect 22204 5842 22260 5852
rect 21644 5170 21700 5180
rect 21756 5290 21812 5302
rect 21756 5238 21758 5290
rect 21810 5238 21812 5290
rect 21196 5070 21198 5122
rect 21250 5070 21252 5122
rect 21196 5058 21252 5070
rect 20020 5012 20076 5014
rect 20020 4946 20076 4956
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19628 4508 19796 4564
rect 19628 4340 19684 4350
rect 19516 4338 19684 4340
rect 19516 4286 19630 4338
rect 19682 4286 19684 4338
rect 19516 4284 19684 4286
rect 19628 4274 19684 4284
rect 19740 4116 19796 4508
rect 20300 4228 20356 4238
rect 19292 4060 20020 4116
rect 19180 3490 19236 3500
rect 19516 3668 19572 3678
rect 19516 3388 19572 3612
rect 18172 3378 18228 3388
rect 19460 3332 19572 3388
rect 19796 3554 19852 3566
rect 19796 3502 19798 3554
rect 19850 3502 19852 3554
rect 19796 3332 19852 3502
rect 19964 3556 20020 4060
rect 20076 3556 20132 3566
rect 19964 3554 20132 3556
rect 19964 3502 20078 3554
rect 20130 3502 20132 3554
rect 19964 3500 20132 3502
rect 20076 3490 20132 3500
rect 20300 3554 20356 4172
rect 20300 3502 20302 3554
rect 20354 3502 20356 3554
rect 20300 3490 20356 3502
rect 20412 4226 20468 4238
rect 20412 4174 20414 4226
rect 20466 4174 20468 4226
rect 20412 3444 20468 4174
rect 21756 3780 21812 5238
rect 21868 5124 21924 5134
rect 21868 5122 22036 5124
rect 21868 5070 21870 5122
rect 21922 5070 22036 5122
rect 21868 5068 22036 5070
rect 21868 5058 21924 5068
rect 21868 4900 21924 4910
rect 21868 4340 21924 4844
rect 21980 4452 22036 5068
rect 21980 4386 22036 4396
rect 22204 5122 22260 5134
rect 22204 5070 22206 5122
rect 22258 5070 22260 5122
rect 21868 4274 21924 4284
rect 20928 3724 21812 3780
rect 21980 4116 22036 4126
rect 20928 3521 20984 3724
rect 20928 3469 20930 3521
rect 20982 3469 20984 3521
rect 21532 3556 21588 3566
rect 20928 3457 20984 3469
rect 21084 3498 21140 3510
rect 20748 3444 20804 3454
rect 20412 3442 20804 3444
rect 20412 3390 20750 3442
rect 20802 3390 20804 3442
rect 20412 3388 20804 3390
rect 20748 3378 20804 3388
rect 21084 3446 21086 3498
rect 21138 3446 21140 3498
rect 21532 3465 21534 3500
rect 21586 3465 21588 3500
rect 21532 3453 21588 3465
rect 21980 3521 22036 4060
rect 22204 4004 22260 5070
rect 22316 4340 22372 4350
rect 22316 4246 22372 4284
rect 22204 3948 22484 4004
rect 22428 3780 22484 3948
rect 22428 3686 22484 3724
rect 22540 3668 22596 6860
rect 23324 6692 23380 7756
rect 23772 7700 23828 7710
rect 23772 7606 23828 7644
rect 24108 7476 24164 7486
rect 24108 7382 24164 7420
rect 24220 7252 24276 8540
rect 24668 8484 24724 8990
rect 25004 8484 25060 11218
rect 25228 11060 25284 11452
rect 25116 11004 25284 11060
rect 25116 10610 25172 11004
rect 25116 10558 25118 10610
rect 25170 10558 25172 10610
rect 25116 9940 25172 10558
rect 25116 9874 25172 9884
rect 25228 9492 25284 9502
rect 25228 8932 25284 9436
rect 25340 9268 25396 13132
rect 25452 12628 25508 12638
rect 25452 11060 25508 12572
rect 25564 11528 25620 13356
rect 25676 13076 25732 13694
rect 25676 13010 25732 13020
rect 25788 13692 26068 13748
rect 26124 14980 26180 14990
rect 25676 12180 25732 12190
rect 25788 12180 25844 13692
rect 25956 13522 26012 13534
rect 25956 13470 25958 13522
rect 26010 13470 26012 13522
rect 25956 13076 26012 13470
rect 25956 13010 26012 13020
rect 26012 12628 26068 12638
rect 26012 12402 26068 12572
rect 26012 12350 26014 12402
rect 26066 12350 26068 12402
rect 26012 12338 26068 12350
rect 26124 12180 26180 14924
rect 26236 14420 26292 14430
rect 26236 14326 26292 14364
rect 26348 13972 26404 15092
rect 25732 12124 25844 12180
rect 25900 12124 26180 12180
rect 26236 13916 26404 13972
rect 25676 12086 25732 12124
rect 25564 11508 25676 11528
rect 25620 11506 25676 11508
rect 25620 11454 25622 11506
rect 25674 11454 25676 11506
rect 25620 11452 25676 11454
rect 25564 11442 25676 11452
rect 25452 11004 25620 11060
rect 25452 10836 25508 10846
rect 25452 10742 25508 10780
rect 25452 9940 25508 9950
rect 25452 9826 25508 9884
rect 25452 9774 25454 9826
rect 25506 9774 25508 9826
rect 25452 9762 25508 9774
rect 25564 9828 25620 11004
rect 25564 9762 25620 9772
rect 25676 10052 25732 10062
rect 25396 9212 25620 9268
rect 25340 9202 25396 9212
rect 25228 8866 25284 8876
rect 25396 8932 25452 8942
rect 25396 8838 25452 8876
rect 25452 8484 25508 8494
rect 25004 8428 25396 8484
rect 24668 8418 24724 8428
rect 25004 8146 25060 8158
rect 25004 8094 25006 8146
rect 25058 8094 25060 8146
rect 24724 7364 24780 7374
rect 23940 7196 24276 7252
rect 24332 7362 24780 7364
rect 24332 7310 24726 7362
rect 24778 7310 24780 7362
rect 24332 7308 24780 7310
rect 23940 6746 23996 7196
rect 24332 6916 24388 7308
rect 24724 7298 24780 7308
rect 25004 7140 25060 8094
rect 25340 8036 25396 8428
rect 25452 8258 25508 8428
rect 25452 8206 25454 8258
rect 25506 8206 25508 8258
rect 25452 8194 25508 8206
rect 25564 8214 25620 9212
rect 25676 9044 25732 9996
rect 25788 9604 25844 9614
rect 25788 9510 25844 9548
rect 25676 8978 25732 8988
rect 25788 9044 25844 9054
rect 25900 9044 25956 12124
rect 26124 11732 26180 11742
rect 26124 11618 26180 11676
rect 26124 11566 26126 11618
rect 26178 11566 26180 11618
rect 26124 11554 26180 11566
rect 26236 11396 26292 13916
rect 26348 13748 26404 13758
rect 26348 13654 26404 13692
rect 26460 12292 26516 17052
rect 26684 17014 26740 17052
rect 26684 16324 26740 16334
rect 26684 15932 26740 16268
rect 26796 16100 26852 17614
rect 26908 17666 26964 17678
rect 26908 17614 26910 17666
rect 26962 17614 26964 17666
rect 26908 17444 26964 17614
rect 27188 17668 27244 17678
rect 27188 17574 27244 17612
rect 26908 17378 26964 17388
rect 27244 17444 27300 17454
rect 27244 17106 27300 17388
rect 27244 17054 27246 17106
rect 27298 17054 27300 17106
rect 27244 17042 27300 17054
rect 26796 16034 26852 16044
rect 26908 16884 26964 16894
rect 27356 16884 27412 18174
rect 26908 16098 26964 16828
rect 26908 16046 26910 16098
rect 26962 16046 26964 16098
rect 26908 16034 26964 16046
rect 27132 16828 27412 16884
rect 27468 17444 27524 18284
rect 27916 18394 28028 18396
rect 27916 18342 27974 18394
rect 28026 18342 28028 18394
rect 28140 18398 28142 18450
rect 28194 18398 28196 18450
rect 28140 18386 28196 18398
rect 28588 18478 28644 18490
rect 28588 18426 28590 18478
rect 28642 18426 28644 18478
rect 27916 18330 28028 18342
rect 27748 17444 27804 17454
rect 27468 17442 27804 17444
rect 27468 17390 27750 17442
rect 27802 17390 27804 17442
rect 27468 17388 27804 17390
rect 26572 15874 26628 15886
rect 26684 15876 26852 15932
rect 26572 15822 26574 15874
rect 26626 15822 26628 15874
rect 26572 15652 26628 15822
rect 26572 15586 26628 15596
rect 26572 15316 26628 15326
rect 26572 15214 26628 15260
rect 26572 15202 26684 15214
rect 26572 15150 26630 15202
rect 26682 15150 26684 15202
rect 26572 15148 26684 15150
rect 26628 15138 26684 15148
rect 26796 14542 26852 15876
rect 27132 14980 27188 16828
rect 27244 15874 27300 15886
rect 27244 15822 27246 15874
rect 27298 15822 27300 15874
rect 27244 15540 27300 15822
rect 27468 15876 27524 17388
rect 27748 17378 27804 17388
rect 27580 17220 27636 17230
rect 27580 16882 27636 17164
rect 27580 16830 27582 16882
rect 27634 16830 27636 16882
rect 27580 16098 27636 16830
rect 27580 16046 27582 16098
rect 27634 16046 27636 16098
rect 27580 16034 27636 16046
rect 27916 16100 27972 18330
rect 28028 18228 28084 18238
rect 28028 17834 28084 18172
rect 28588 18228 28644 18426
rect 29036 18450 29092 19180
rect 29820 19142 29876 19180
rect 28588 18162 28644 18172
rect 28812 18394 28868 18406
rect 28812 18342 28814 18394
rect 28866 18342 28868 18394
rect 28812 18228 28868 18342
rect 28812 18162 28868 18172
rect 29036 18398 29038 18450
rect 29090 18398 29092 18450
rect 28028 17782 28030 17834
rect 28082 17782 28084 17834
rect 29036 17892 29092 18398
rect 29036 17826 29092 17836
rect 29260 18340 29316 18350
rect 28028 16436 28084 17782
rect 28140 17780 28196 17790
rect 28140 17666 28196 17724
rect 28588 17780 28644 17790
rect 28140 17614 28142 17666
rect 28194 17614 28196 17666
rect 28140 17444 28196 17614
rect 28140 17378 28196 17388
rect 28476 17666 28532 17678
rect 28476 17614 28478 17666
rect 28530 17614 28532 17666
rect 28308 17332 28364 17342
rect 28028 16370 28084 16380
rect 28140 17220 28196 17230
rect 28140 16882 28196 17164
rect 28140 16830 28142 16882
rect 28194 16830 28196 16882
rect 28308 16938 28364 17276
rect 28308 16886 28310 16938
rect 28362 16886 28364 16938
rect 28476 17108 28532 17614
rect 28476 16994 28532 17052
rect 28476 16942 28478 16994
rect 28530 16942 28532 16994
rect 28476 16930 28532 16942
rect 28308 16874 28364 16886
rect 28588 16882 28644 17724
rect 29260 17778 29316 18284
rect 29820 18340 29876 18350
rect 29820 18246 29876 18284
rect 29260 17726 29262 17778
rect 29314 17726 29316 17778
rect 29260 17714 29316 17726
rect 29484 18116 29540 18126
rect 29484 17666 29540 18060
rect 29092 17612 29148 17622
rect 28924 17610 29148 17612
rect 28924 17558 29094 17610
rect 29146 17558 29148 17610
rect 29484 17614 29486 17666
rect 29538 17614 29540 17666
rect 29484 17602 29540 17614
rect 29708 18004 29764 18014
rect 29708 17638 29764 17948
rect 29708 17586 29710 17638
rect 29762 17586 29764 17638
rect 29708 17574 29764 17586
rect 28924 17556 29148 17558
rect 27916 16044 28084 16100
rect 27916 15876 27972 15886
rect 27468 15810 27524 15820
rect 27692 15820 27916 15876
rect 27244 15484 27636 15540
rect 27132 14914 27188 14924
rect 27244 15314 27300 15326
rect 27244 15262 27246 15314
rect 27298 15262 27300 15314
rect 27580 15314 27636 15484
rect 27244 14756 27300 15262
rect 27412 15258 27468 15270
rect 27412 15206 27414 15258
rect 27466 15206 27468 15258
rect 27412 15148 27468 15206
rect 27580 15262 27582 15314
rect 27634 15262 27636 15314
rect 27412 15092 27524 15148
rect 27244 14690 27300 14700
rect 27468 14644 27524 15092
rect 27468 14578 27524 14588
rect 26684 14532 26740 14542
rect 26796 14530 26908 14542
rect 26796 14478 26854 14530
rect 26906 14478 26908 14530
rect 26796 14476 26908 14478
rect 26684 14438 26740 14476
rect 26852 14466 26908 14476
rect 27132 14530 27188 14542
rect 27132 14478 27134 14530
rect 27186 14504 27188 14530
rect 27186 14478 27202 14504
rect 27132 14448 27202 14478
rect 27020 14418 27076 14430
rect 27020 14366 27022 14418
rect 27074 14366 27076 14418
rect 27020 14196 27076 14366
rect 27146 14308 27202 14448
rect 27412 14418 27468 14430
rect 27412 14366 27414 14418
rect 27466 14366 27468 14418
rect 27146 14252 27300 14308
rect 27020 14130 27076 14140
rect 26684 14084 26740 14094
rect 26740 14028 26964 14084
rect 26684 14018 26740 14028
rect 26572 13972 26628 13982
rect 26572 13748 26628 13916
rect 26572 13682 26628 13692
rect 26684 13860 26740 13870
rect 26684 13746 26740 13804
rect 26684 13694 26686 13746
rect 26738 13694 26740 13746
rect 26684 13682 26740 13694
rect 26796 13636 26852 13646
rect 26796 13578 26852 13580
rect 26796 13526 26798 13578
rect 26850 13526 26852 13578
rect 26796 13514 26852 13526
rect 26908 12962 26964 14028
rect 27020 13860 27076 13870
rect 27020 13746 27076 13804
rect 27020 13694 27022 13746
rect 27074 13694 27076 13746
rect 27020 13682 27076 13694
rect 27244 13636 27300 14252
rect 27412 13860 27468 14366
rect 27412 13794 27468 13804
rect 27356 13636 27412 13646
rect 27244 13580 27356 13636
rect 27356 13542 27412 13580
rect 27580 13412 27636 15262
rect 27692 15314 27748 15820
rect 27916 15782 27972 15820
rect 28028 15438 28084 16044
rect 27972 15426 28084 15438
rect 27972 15374 27974 15426
rect 28026 15374 28084 15426
rect 27972 15372 28084 15374
rect 28140 15540 28196 16830
rect 28588 16830 28590 16882
rect 28642 16830 28644 16882
rect 28588 16818 28644 16830
rect 28700 17332 28756 17342
rect 28700 16436 28756 17276
rect 28924 17006 28980 17556
rect 29092 17546 29148 17556
rect 29428 17108 29484 17118
rect 29428 17014 29484 17052
rect 28868 16994 28980 17006
rect 29932 16996 29988 19964
rect 30268 19954 30324 19964
rect 30380 19908 30436 22318
rect 30492 21474 30548 21486
rect 30492 21422 30494 21474
rect 30546 21422 30548 21474
rect 30492 20580 30548 21422
rect 30604 20804 30660 22540
rect 30716 22372 30772 22382
rect 30828 22372 30884 23660
rect 30940 23380 30996 23884
rect 31220 23882 31276 23894
rect 31052 23828 31108 23838
rect 31052 23734 31108 23772
rect 31220 23830 31222 23882
rect 31274 23830 31276 23882
rect 31220 23492 31276 23830
rect 31612 23826 31668 23838
rect 31612 23774 31614 23826
rect 31666 23774 31668 23826
rect 31612 23604 31668 23774
rect 31612 23538 31668 23548
rect 31220 23436 31500 23492
rect 30940 23314 30996 23324
rect 30996 23156 31052 23166
rect 31276 23156 31332 23166
rect 30716 22370 30884 22372
rect 30716 22318 30718 22370
rect 30770 22318 30884 22370
rect 30716 22316 30884 22318
rect 30940 23154 31332 23156
rect 30940 23102 30998 23154
rect 31050 23102 31278 23154
rect 31330 23102 31332 23154
rect 30940 23100 31332 23102
rect 30940 23090 31052 23100
rect 31276 23090 31332 23100
rect 31444 23098 31500 23436
rect 30716 22306 30772 22316
rect 30940 21812 30996 23090
rect 31444 23046 31446 23098
rect 31498 23046 31500 23098
rect 31052 22820 31108 22830
rect 31052 22594 31108 22764
rect 31052 22542 31054 22594
rect 31106 22542 31108 22594
rect 31052 22530 31108 22542
rect 31444 22596 31500 23046
rect 31612 23380 31668 23390
rect 31612 23266 31668 23324
rect 31612 23214 31614 23266
rect 31666 23214 31668 23266
rect 31612 22606 31668 23214
rect 31724 23154 31780 24220
rect 31836 23940 31892 24670
rect 31948 24554 32004 24780
rect 32060 24722 32116 24892
rect 32060 24670 32062 24722
rect 32114 24670 32116 24722
rect 32060 24658 32116 24670
rect 31948 24502 31950 24554
rect 32002 24502 32004 24554
rect 31948 24490 32004 24502
rect 31836 23874 31892 23884
rect 31948 23604 32004 23614
rect 31948 23492 32116 23548
rect 32060 23380 32116 23492
rect 32060 23314 32116 23324
rect 32172 23268 32228 25116
rect 32844 24948 32900 28812
rect 33012 28644 33068 28654
rect 33012 28550 33068 28588
rect 32956 26964 33012 27002
rect 32956 26898 33012 26908
rect 33180 26628 33236 29932
rect 33292 27300 33348 30156
rect 33628 29428 33684 30156
rect 33740 29876 33796 31726
rect 33852 31556 33908 32956
rect 34524 32946 34580 32956
rect 33964 32788 34020 32798
rect 33964 31778 34020 32732
rect 35084 32562 35140 33068
rect 35364 32900 35420 33238
rect 35364 32834 35420 32844
rect 35532 33290 35588 33302
rect 35532 33238 35534 33290
rect 35586 33238 35588 33290
rect 35084 32510 35086 32562
rect 35138 32510 35140 32562
rect 35084 32498 35140 32510
rect 35532 32452 35588 33238
rect 35868 33290 35924 33302
rect 35868 33238 35870 33290
rect 35922 33238 35924 33290
rect 36316 33254 36372 33292
rect 36932 33346 37044 33358
rect 36932 33294 36934 33346
rect 36986 33294 37044 33346
rect 36932 33292 37044 33294
rect 37324 33346 37380 33358
rect 37324 33294 37326 33346
rect 37378 33294 37380 33346
rect 38108 33346 38164 34076
rect 36932 33282 36988 33292
rect 35868 33124 35924 33238
rect 37100 33236 37156 33246
rect 37100 33142 37156 33180
rect 35868 33058 35924 33068
rect 35868 32788 35924 32798
rect 35868 32562 35924 32732
rect 37100 32788 37156 32798
rect 35868 32510 35870 32562
rect 35922 32510 35924 32562
rect 35868 32498 35924 32510
rect 36204 32676 36260 32686
rect 35532 32386 35588 32396
rect 36092 32452 36148 32462
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 36092 31790 36148 32396
rect 33964 31726 33966 31778
rect 34018 31726 34020 31778
rect 33964 31714 34020 31726
rect 35196 31780 35252 31790
rect 36072 31780 36148 31790
rect 35196 31686 35252 31724
rect 35868 31778 36148 31780
rect 35868 31726 36074 31778
rect 36126 31726 36148 31778
rect 35868 31724 36148 31726
rect 33852 31500 34132 31556
rect 33944 31220 34000 31230
rect 33944 31050 34000 31164
rect 33944 30998 33946 31050
rect 33998 30998 34000 31050
rect 33944 30986 34000 30998
rect 33740 29810 33796 29820
rect 34076 29764 34132 31500
rect 35756 31108 35812 31118
rect 35868 31108 35924 31724
rect 36072 31714 36128 31724
rect 36204 31556 36260 32620
rect 36428 32589 36484 32601
rect 36428 32537 36430 32589
rect 36482 32537 36484 32589
rect 35756 31106 35924 31108
rect 35756 31054 35758 31106
rect 35810 31054 35924 31106
rect 35756 31052 35924 31054
rect 36092 31500 36260 31556
rect 36316 31892 36372 31902
rect 36316 31666 36372 31836
rect 36316 31614 36318 31666
rect 36370 31614 36372 31666
rect 35756 31042 35812 31052
rect 34188 30996 34244 31006
rect 34636 30996 34692 31006
rect 34188 30902 34244 30940
rect 34412 30994 34692 30996
rect 34412 30942 34638 30994
rect 34690 30942 34692 30994
rect 34412 30940 34692 30942
rect 34412 30660 34468 30940
rect 34636 30930 34692 30940
rect 35512 30996 35568 31006
rect 35512 30902 35568 30940
rect 34412 30604 34580 30660
rect 34524 30378 34580 30604
rect 35196 30604 35460 30614
rect 34524 30326 34526 30378
rect 34578 30326 34580 30378
rect 34524 30314 34580 30326
rect 34748 30548 34804 30558
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 34188 30212 34244 30222
rect 34636 30212 34692 30222
rect 34188 30210 34692 30212
rect 34188 30158 34190 30210
rect 34242 30158 34638 30210
rect 34690 30158 34692 30210
rect 34188 30156 34692 30158
rect 34188 30146 34244 30156
rect 34076 29698 34132 29708
rect 33740 29428 33796 29466
rect 34636 29438 34692 30156
rect 33628 29372 33740 29428
rect 33740 29362 33796 29372
rect 34616 29426 34692 29438
rect 34616 29374 34618 29426
rect 34670 29374 34692 29426
rect 34616 29372 34692 29374
rect 33460 29314 33516 29326
rect 33460 29262 33462 29314
rect 33514 29262 33516 29314
rect 33460 29204 33516 29262
rect 33460 29138 33516 29148
rect 34616 28980 34672 29372
rect 34300 28924 34672 28980
rect 33404 28868 33460 28878
rect 33404 28644 33460 28812
rect 33404 27914 33460 28588
rect 33628 28642 33684 28654
rect 33628 28590 33630 28642
rect 33682 28590 33684 28642
rect 33628 28532 33684 28590
rect 33628 28308 33684 28476
rect 33628 28252 33964 28308
rect 33404 27862 33406 27914
rect 33458 27862 33460 27914
rect 33404 27850 33460 27862
rect 33740 28084 33796 28094
rect 33740 27914 33796 28028
rect 33740 27862 33742 27914
rect 33794 27862 33796 27914
rect 33740 27748 33796 27862
rect 33628 27692 33796 27748
rect 33908 27914 33964 28252
rect 33908 27862 33910 27914
rect 33962 27862 33964 27914
rect 34188 27972 34244 27982
rect 34300 27972 34356 28924
rect 34748 28868 34804 30492
rect 35312 30212 35368 30222
rect 35312 30120 35314 30156
rect 35366 30120 35368 30156
rect 35312 30108 35368 30120
rect 35812 30212 35868 30222
rect 35812 30118 35868 30156
rect 36092 29988 36148 31500
rect 36204 30884 36260 30894
rect 36204 30210 36260 30828
rect 36316 30660 36372 31614
rect 36316 30594 36372 30604
rect 36428 31780 36484 32537
rect 37100 31902 37156 32732
rect 37324 32004 37380 33294
rect 37660 33290 37716 33302
rect 37660 33238 37662 33290
rect 37714 33238 37716 33290
rect 38108 33294 38110 33346
rect 38162 33294 38164 33346
rect 38108 33282 38164 33294
rect 37660 33236 37716 33238
rect 37660 33180 37828 33236
rect 37772 33124 37828 33180
rect 37660 33012 37716 33022
rect 37436 32788 37492 32798
rect 37436 32694 37492 32732
rect 37324 31938 37380 31948
rect 37100 31890 37212 31902
rect 37100 31838 37158 31890
rect 37210 31838 37212 31890
rect 37100 31836 37212 31838
rect 37156 31826 37212 31836
rect 36428 31724 37044 31780
rect 36204 30158 36206 30210
rect 36258 30158 36260 30210
rect 36204 30146 36260 30158
rect 36428 30212 36484 31724
rect 36988 31668 37044 31724
rect 37548 31750 37604 31762
rect 37548 31698 37550 31750
rect 37602 31698 37604 31750
rect 37548 31668 37604 31698
rect 36988 31612 37604 31668
rect 37660 31220 37716 32956
rect 37324 31164 37716 31220
rect 36838 31108 36894 31118
rect 36838 31032 36894 31052
rect 36540 30996 36596 31006
rect 36540 30902 36596 30940
rect 36652 30994 36708 31006
rect 36652 30942 36654 30994
rect 36706 30942 36708 30994
rect 36838 30980 36840 31032
rect 36892 30980 36894 31032
rect 36838 30968 36894 30980
rect 36428 30146 36484 30156
rect 36540 30210 36596 30222
rect 36540 30158 36542 30210
rect 36594 30158 36596 30210
rect 36540 30100 36596 30158
rect 36540 30034 36596 30044
rect 35756 29932 36148 29988
rect 34860 29540 34916 29550
rect 34860 29446 34916 29484
rect 35756 29428 35812 29932
rect 36652 29764 36708 30942
rect 37212 30884 37268 30894
rect 37324 30884 37380 31164
rect 37548 30996 37604 31006
rect 37548 30994 37716 30996
rect 37548 30942 37550 30994
rect 37602 30942 37716 30994
rect 37548 30940 37716 30942
rect 37548 30930 37604 30940
rect 37212 30882 37380 30884
rect 37212 30830 37214 30882
rect 37266 30830 37380 30882
rect 37212 30828 37380 30830
rect 37212 30818 37268 30828
rect 37380 30154 37436 30166
rect 37100 30098 37156 30110
rect 37100 30046 37102 30098
rect 37154 30046 37156 30098
rect 37100 29988 37156 30046
rect 37100 29922 37156 29932
rect 37380 30102 37382 30154
rect 37434 30102 37436 30154
rect 36652 29698 36708 29708
rect 35924 29652 35980 29662
rect 35924 29650 36372 29652
rect 35924 29598 35926 29650
rect 35978 29598 36372 29650
rect 35924 29596 36372 29598
rect 35924 29586 35980 29596
rect 36092 29428 36148 29438
rect 35756 29372 35924 29428
rect 34748 28802 34804 28812
rect 34972 29316 35028 29326
rect 34504 28644 34560 28654
rect 34504 28550 34560 28588
rect 34748 28644 34804 28654
rect 34748 28550 34804 28588
rect 34972 28644 35028 29260
rect 35476 29316 35532 29326
rect 35476 29222 35532 29260
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 28644 35252 28654
rect 34972 28642 35252 28644
rect 34972 28590 35198 28642
rect 35250 28590 35252 28642
rect 34972 28588 35252 28590
rect 34972 28084 35028 28588
rect 35196 28578 35252 28588
rect 35868 28420 35924 29372
rect 36092 29334 36148 29372
rect 36316 29426 36372 29596
rect 36316 29374 36318 29426
rect 36370 29374 36372 29426
rect 37192 29540 37248 29550
rect 37380 29540 37436 30102
rect 37192 29482 37248 29484
rect 37192 29430 37194 29482
rect 37246 29430 37248 29482
rect 37192 29418 37248 29430
rect 37324 29484 37436 29540
rect 37548 30154 37604 30166
rect 37548 30102 37550 30154
rect 37602 30102 37604 30154
rect 37548 29540 37604 30102
rect 37324 29428 37380 29484
rect 37548 29474 37604 29484
rect 36316 29362 36372 29374
rect 37156 29092 37212 29102
rect 36316 28868 36372 28878
rect 36316 28774 36372 28812
rect 37156 28756 37212 29036
rect 37156 28662 37212 28700
rect 36072 28644 36128 28654
rect 37324 28644 37380 29372
rect 37436 29202 37492 29214
rect 37436 29150 37438 29202
rect 37490 29150 37492 29202
rect 37436 28868 37492 29150
rect 37660 29204 37716 30940
rect 37772 29988 37828 33068
rect 38444 32004 38500 34076
rect 38556 32788 38612 35084
rect 38668 34468 38724 34478
rect 38668 32900 38724 34412
rect 39004 34356 39060 36092
rect 39452 35924 39508 35934
rect 39116 35700 39172 35710
rect 39340 35700 39396 35710
rect 39116 35698 39396 35700
rect 39116 35646 39118 35698
rect 39170 35646 39342 35698
rect 39394 35646 39396 35698
rect 39116 35644 39396 35646
rect 39116 35634 39172 35644
rect 39228 35476 39284 35486
rect 39228 35026 39284 35420
rect 39228 34974 39230 35026
rect 39282 34974 39284 35026
rect 39228 34962 39284 34974
rect 39004 34290 39060 34300
rect 38948 34132 39004 34142
rect 39228 34132 39284 34142
rect 38668 32834 38724 32844
rect 38780 34130 39004 34132
rect 38780 34078 38950 34130
rect 39002 34078 39004 34130
rect 38780 34076 39004 34078
rect 38556 32722 38612 32732
rect 38556 32228 38612 32238
rect 38780 32228 38836 34076
rect 38948 34066 39004 34076
rect 39116 34130 39284 34132
rect 39116 34078 39230 34130
rect 39282 34078 39284 34130
rect 39116 34076 39284 34078
rect 39340 34132 39396 35644
rect 39452 35698 39508 35868
rect 39452 35646 39454 35698
rect 39506 35646 39508 35698
rect 39452 35634 39508 35646
rect 39732 35700 39788 35710
rect 39732 35606 39788 35644
rect 40012 35252 40068 37436
rect 40236 37492 40292 37502
rect 40236 37378 40292 37436
rect 40236 37326 40238 37378
rect 40290 37326 40292 37378
rect 40236 37314 40292 37326
rect 40572 37492 40628 37502
rect 40348 37268 40404 37278
rect 40348 36718 40404 37212
rect 40292 36706 40404 36718
rect 40292 36654 40294 36706
rect 40346 36654 40404 36706
rect 40292 36652 40404 36654
rect 40292 36642 40348 36652
rect 40124 36596 40180 36606
rect 40124 35924 40180 36540
rect 40572 36454 40628 37436
rect 41020 36596 41076 42476
rect 41188 42466 41244 42476
rect 41356 42084 41412 42924
rect 41580 42868 41636 42878
rect 41580 42810 41636 42812
rect 41580 42758 41582 42810
rect 41634 42758 41636 42810
rect 41580 42746 41636 42758
rect 41692 42716 41748 43036
rect 42252 42866 42308 43036
rect 42252 42814 42254 42866
rect 42306 42814 42308 42866
rect 42252 42802 42308 42814
rect 42420 42810 42476 43148
rect 42420 42758 42422 42810
rect 42474 42758 42476 42810
rect 42420 42746 42476 42758
rect 41692 42664 41694 42716
rect 41746 42664 41748 42716
rect 41692 42652 41748 42664
rect 42588 42196 42644 45052
rect 42700 44884 42756 45838
rect 42700 44818 42756 44828
rect 42812 44548 42868 49200
rect 43596 45862 43652 45874
rect 43596 45810 43598 45862
rect 43650 45810 43652 45862
rect 42980 45780 43036 45790
rect 42980 45686 43036 45724
rect 43260 45444 43316 45454
rect 43260 45332 43316 45388
rect 43596 45332 43652 45810
rect 43260 45276 43652 45332
rect 42812 44482 42868 44492
rect 43036 44994 43092 45006
rect 43036 44942 43038 44994
rect 43090 44942 43092 44994
rect 42812 44212 42868 44222
rect 42812 44210 42980 44212
rect 42812 44158 42814 44210
rect 42866 44158 42980 44210
rect 42812 44156 42980 44158
rect 42812 44146 42868 44156
rect 42700 43568 42756 43580
rect 42700 43516 42702 43568
rect 42754 43516 42756 43568
rect 42700 43428 42756 43516
rect 42700 43362 42756 43372
rect 42924 42756 42980 44156
rect 43036 43876 43092 44942
rect 43260 44660 43316 45276
rect 44380 45108 44436 49200
rect 44604 46002 44660 46014
rect 44604 45950 44606 46002
rect 44658 45950 44660 46002
rect 44604 45332 44660 45950
rect 45948 45556 46004 49200
rect 48076 45948 48356 46004
rect 46284 45892 46340 45902
rect 46508 45892 46564 45902
rect 46284 45798 46340 45836
rect 46396 45890 46564 45892
rect 46396 45838 46510 45890
rect 46562 45838 46564 45890
rect 48076 45852 48132 45948
rect 46396 45836 46564 45838
rect 45948 45500 46116 45556
rect 44604 45266 44660 45276
rect 45388 45108 45444 45118
rect 44380 45052 44660 45108
rect 43260 44604 43540 44660
rect 43260 44436 43316 44446
rect 43260 44292 43316 44380
rect 43260 44240 43262 44292
rect 43314 44240 43316 44292
rect 43260 44228 43316 44240
rect 43484 44283 43540 44604
rect 43484 44231 43486 44283
rect 43538 44231 43540 44283
rect 43484 44219 43540 44231
rect 43764 44324 43820 44334
rect 43764 44266 43820 44268
rect 43764 44214 43766 44266
rect 43818 44214 43820 44266
rect 44268 44324 44324 44334
rect 44268 44230 44324 44268
rect 43764 44202 43820 44214
rect 44100 44100 44156 44110
rect 44100 44006 44156 44044
rect 43036 43810 43092 43820
rect 43036 43568 43092 43580
rect 43036 43516 43038 43568
rect 43090 43516 43092 43568
rect 43036 42978 43092 43516
rect 43484 43540 43540 43550
rect 43932 43540 43988 43550
rect 43036 42926 43038 42978
rect 43090 42926 43092 42978
rect 43036 42914 43092 42926
rect 43204 43482 43260 43494
rect 43204 43430 43206 43482
rect 43258 43430 43260 43482
rect 43484 43446 43540 43484
rect 43708 43538 43988 43540
rect 43708 43486 43934 43538
rect 43986 43486 43988 43538
rect 43708 43484 43988 43486
rect 43204 42868 43260 43430
rect 43708 42868 43764 43484
rect 43932 43474 43988 43484
rect 44604 42980 44660 45052
rect 44940 44994 44996 45006
rect 44940 44942 44942 44994
rect 44994 44942 44996 44994
rect 44940 44324 44996 44942
rect 44940 44258 44996 44268
rect 45388 43708 45444 45052
rect 45612 44548 45668 44558
rect 45612 44454 45668 44492
rect 45052 43652 45108 43662
rect 45052 43558 45108 43596
rect 45164 43652 45444 43708
rect 44808 43538 44864 43550
rect 44808 43486 44810 43538
rect 44862 43486 44864 43538
rect 44808 42980 44864 43486
rect 44604 42914 44660 42924
rect 44716 42924 44864 42980
rect 44940 43540 44996 43550
rect 44156 42868 44212 42878
rect 43204 42812 43652 42868
rect 43708 42812 43876 42868
rect 42924 42700 43484 42756
rect 42588 42140 42756 42196
rect 41244 42028 41412 42084
rect 41804 42084 41860 42094
rect 41244 40402 41300 42028
rect 41580 41858 41636 41870
rect 41580 41806 41582 41858
rect 41634 41806 41636 41858
rect 41580 41636 41636 41806
rect 41356 41580 41636 41636
rect 41804 41636 41860 42028
rect 42700 41972 42756 42140
rect 42700 41906 42756 41916
rect 43260 41636 43316 42700
rect 43428 42698 43484 42700
rect 43428 42646 43430 42698
rect 43482 42646 43484 42698
rect 43428 42634 43484 42646
rect 41804 41580 42084 41636
rect 41356 41298 41412 41580
rect 41356 41246 41358 41298
rect 41410 41246 41412 41298
rect 41356 41234 41412 41246
rect 41468 41188 41524 41198
rect 41468 41119 41470 41132
rect 41522 41119 41524 41132
rect 41468 41094 41524 41119
rect 41804 41186 41860 41198
rect 41804 41134 41806 41186
rect 41858 41134 41860 41186
rect 41804 41076 41860 41134
rect 41804 41010 41860 41020
rect 41244 40350 41246 40402
rect 41298 40350 41300 40402
rect 41132 39060 41188 39070
rect 41244 39060 41300 40350
rect 41356 40402 41412 40414
rect 41356 40350 41358 40402
rect 41410 40350 41412 40402
rect 41356 39844 41412 40350
rect 41524 40402 41580 40414
rect 41524 40350 41526 40402
rect 41578 40350 41580 40402
rect 41524 40068 41580 40350
rect 41916 40404 41972 40414
rect 41916 40290 41972 40348
rect 41916 40238 41918 40290
rect 41970 40238 41972 40290
rect 41916 40226 41972 40238
rect 41524 40002 41580 40012
rect 41356 39778 41412 39788
rect 41356 39620 41412 39630
rect 41356 39526 41412 39564
rect 41132 39058 41300 39060
rect 41132 39006 41134 39058
rect 41186 39006 41300 39058
rect 41132 39004 41300 39006
rect 41692 39396 41748 39406
rect 41132 38994 41188 39004
rect 41505 38890 41561 38902
rect 41505 38838 41507 38890
rect 41559 38838 41561 38890
rect 41505 38836 41561 38838
rect 41132 38780 41561 38836
rect 41692 38890 41748 39340
rect 41692 38838 41694 38890
rect 41746 38838 41748 38890
rect 41692 38836 41748 38838
rect 41132 38724 41188 38780
rect 41692 38760 41748 38780
rect 41916 38862 41972 38874
rect 41916 38810 41918 38862
rect 41970 38810 41972 38862
rect 41132 38022 41188 38668
rect 41916 38724 41972 38810
rect 41132 37970 41134 38022
rect 41186 37970 41188 38022
rect 41132 37958 41188 37970
rect 41244 38612 41300 38622
rect 41244 37490 41300 38556
rect 41692 38276 41748 38286
rect 41692 38015 41748 38220
rect 41244 37438 41246 37490
rect 41298 37438 41300 37490
rect 41244 37426 41300 37438
rect 41356 37994 41412 38006
rect 41356 37942 41358 37994
rect 41410 37942 41412 37994
rect 41356 37044 41412 37942
rect 41580 37994 41636 38006
rect 41580 37942 41582 37994
rect 41634 37942 41636 37994
rect 41692 37963 41694 38015
rect 41746 37963 41748 38015
rect 41692 37951 41748 37963
rect 41580 37716 41636 37942
rect 41580 37650 41636 37660
rect 41916 37490 41972 38668
rect 42028 38668 42084 41580
rect 43204 41580 43316 41636
rect 43484 42532 43540 42542
rect 43484 41972 43540 42476
rect 43484 41858 43540 41916
rect 43484 41806 43486 41858
rect 43538 41806 43540 41858
rect 43204 41412 43260 41580
rect 42756 41356 43260 41412
rect 42756 41242 42812 41356
rect 42196 41188 42252 41198
rect 42196 41094 42252 41132
rect 42476 41188 42532 41198
rect 42756 41190 42758 41242
rect 42810 41190 42812 41242
rect 43204 41242 43260 41356
rect 42756 41178 42812 41190
rect 42924 41186 42980 41198
rect 42476 41094 42532 41132
rect 42924 41134 42926 41186
rect 42978 41134 42980 41186
rect 42588 41074 42644 41086
rect 42588 41022 42590 41074
rect 42642 41022 42644 41074
rect 42588 40964 42644 41022
rect 42588 40740 42644 40908
rect 42924 40852 42980 41134
rect 42924 40786 42980 40796
rect 43204 41190 43206 41242
rect 43258 41190 43260 41242
rect 42140 40684 42644 40740
rect 42756 40740 42812 40750
rect 42140 40180 42196 40684
rect 42252 40516 42308 40526
rect 42252 40402 42308 40460
rect 42756 40514 42812 40684
rect 42756 40462 42758 40514
rect 42810 40462 42812 40514
rect 42756 40450 42812 40462
rect 43204 40516 43260 41190
rect 43372 41076 43428 41086
rect 43372 40982 43428 41020
rect 43484 40628 43540 41806
rect 43596 41412 43652 42812
rect 43708 42698 43764 42710
rect 43708 42646 43710 42698
rect 43762 42646 43764 42698
rect 43708 42644 43764 42646
rect 43708 42578 43764 42588
rect 43820 42532 43876 42812
rect 43988 42756 44044 42766
rect 43988 42698 44044 42700
rect 43988 42646 43990 42698
rect 44042 42646 44044 42698
rect 43988 42634 44044 42646
rect 43820 42476 44044 42532
rect 43988 42194 44044 42476
rect 43988 42142 43990 42194
rect 44042 42142 44044 42194
rect 43988 42130 44044 42142
rect 44156 42000 44212 42812
rect 44492 42308 44548 42318
rect 44716 42308 44772 42924
rect 44940 42420 44996 43484
rect 44548 42252 44772 42308
rect 44828 42364 44996 42420
rect 45052 43428 45108 43438
rect 45052 42726 45108 43372
rect 45052 42674 45054 42726
rect 45106 42674 45108 42726
rect 44324 42026 44380 42038
rect 44324 42000 44326 42026
rect 44156 41974 44326 42000
rect 44378 41974 44380 42026
rect 44156 41970 44380 41974
rect 44156 41918 44158 41970
rect 44210 41944 44380 41970
rect 44492 42026 44548 42252
rect 44492 41974 44494 42026
rect 44546 41974 44548 42026
rect 44210 41918 44212 41944
rect 44156 41906 44212 41918
rect 44492 41860 44548 41974
rect 44380 41804 44492 41860
rect 43596 41346 43652 41356
rect 43932 41636 43988 41646
rect 43596 41186 43652 41198
rect 43596 41134 43598 41186
rect 43650 41134 43652 41186
rect 43596 40964 43652 41134
rect 43596 40898 43652 40908
rect 43932 41188 43988 41580
rect 43932 41096 43934 41132
rect 43986 41096 43988 41132
rect 43820 40852 43876 40862
rect 43484 40562 43540 40572
rect 43652 40740 43708 40750
rect 43372 40516 43428 40526
rect 43204 40460 43316 40516
rect 42252 40350 42254 40402
rect 42306 40350 42308 40402
rect 42252 40338 42308 40350
rect 42476 40404 42532 40414
rect 42476 40310 42532 40348
rect 42140 40124 42308 40180
rect 42140 39618 42196 39630
rect 42140 39566 42142 39618
rect 42194 39566 42196 39618
rect 42140 39508 42196 39566
rect 42140 39442 42196 39452
rect 42140 39284 42196 39294
rect 42140 38890 42196 39228
rect 42140 38838 42142 38890
rect 42194 38838 42196 38890
rect 42252 38948 42308 40124
rect 42364 40068 42420 40078
rect 42364 38958 42420 40012
rect 42700 39396 42756 39406
rect 42364 38946 42476 38958
rect 42364 38894 42422 38946
rect 42474 38894 42476 38946
rect 42364 38892 42476 38894
rect 42252 38882 42308 38892
rect 42420 38882 42476 38892
rect 42140 38826 42196 38838
rect 42588 38724 42644 38734
rect 42028 38612 42532 38668
rect 42084 38388 42140 38398
rect 42084 38274 42140 38332
rect 42084 38222 42086 38274
rect 42138 38222 42140 38274
rect 42084 38210 42140 38222
rect 42364 38276 42420 38286
rect 42364 38022 42420 38220
rect 42364 37970 42366 38022
rect 42418 37970 42420 38022
rect 42364 37958 42420 37970
rect 41916 37438 41918 37490
rect 41970 37438 41972 37490
rect 41916 37426 41972 37438
rect 42140 37716 42196 37726
rect 41580 37268 41636 37278
rect 41580 37174 41636 37212
rect 41356 36978 41412 36988
rect 42028 37044 42084 37054
rect 41524 36708 41580 36718
rect 41524 36614 41580 36652
rect 40572 36402 40574 36454
rect 40626 36402 40628 36454
rect 40572 36390 40628 36402
rect 40684 36540 41076 36596
rect 40684 36260 40740 36540
rect 41132 36484 41188 36494
rect 40572 36204 40740 36260
rect 40796 36426 40852 36438
rect 40796 36374 40798 36426
rect 40850 36374 40852 36426
rect 40292 35924 40348 35934
rect 40124 35922 40348 35924
rect 40124 35870 40294 35922
rect 40346 35870 40348 35922
rect 40124 35868 40348 35870
rect 40292 35858 40348 35868
rect 40012 35196 40404 35252
rect 40348 34692 40404 35196
rect 40236 34636 40404 34692
rect 39676 34300 39956 34356
rect 39452 34132 39508 34142
rect 39676 34132 39732 34300
rect 39340 34130 39732 34132
rect 39340 34078 39454 34130
rect 39506 34078 39678 34130
rect 39730 34078 39732 34130
rect 39340 34076 39732 34078
rect 38892 33684 38948 33694
rect 38892 33458 38948 33628
rect 38892 33406 38894 33458
rect 38946 33406 38948 33458
rect 38892 33394 38948 33406
rect 39116 33012 39172 34076
rect 39228 34066 39284 34076
rect 39452 34066 39508 34076
rect 39676 34066 39732 34076
rect 39788 34130 39844 34142
rect 39788 34078 39790 34130
rect 39842 34078 39844 34130
rect 39788 33684 39844 34078
rect 39900 33908 39956 34300
rect 40068 34132 40124 34142
rect 40068 34038 40124 34076
rect 39900 33852 40180 33908
rect 39788 33628 40068 33684
rect 40012 33124 40068 33628
rect 39116 32946 39172 32956
rect 39564 33068 40068 33124
rect 38892 32564 38948 32574
rect 38892 32470 38948 32508
rect 39004 32562 39060 32574
rect 39004 32510 39006 32562
rect 39058 32510 39060 32562
rect 39004 32452 39060 32510
rect 39172 32564 39228 32574
rect 39172 32470 39228 32508
rect 39004 32386 39060 32396
rect 39564 32450 39620 33068
rect 40012 32900 40068 32910
rect 39900 32788 39956 32798
rect 39564 32398 39566 32450
rect 39618 32398 39620 32450
rect 39564 32386 39620 32398
rect 39788 32452 39844 32462
rect 38612 32172 38836 32228
rect 38556 32162 38612 32172
rect 38556 32004 38612 32014
rect 38444 32002 38612 32004
rect 38444 31950 38558 32002
rect 38610 31950 38612 32002
rect 38444 31948 38612 31950
rect 38556 31938 38612 31948
rect 39676 31892 39732 31902
rect 39452 31220 39508 31230
rect 38332 30884 38388 30894
rect 38332 30790 38388 30828
rect 38332 30660 38388 30670
rect 37772 29922 37828 29932
rect 37884 30154 37940 30166
rect 37884 30102 37886 30154
rect 37938 30102 37940 30154
rect 37660 29138 37716 29148
rect 37884 29426 37940 30102
rect 37884 29374 37886 29426
rect 37938 29374 37940 29426
rect 37660 28980 37716 28990
rect 37660 28868 37716 28924
rect 37436 28812 37716 28868
rect 37548 28644 37604 28654
rect 37324 28642 37604 28644
rect 37324 28590 37550 28642
rect 37602 28590 37604 28642
rect 37324 28588 37604 28590
rect 36072 28550 36128 28588
rect 37548 28578 37604 28588
rect 35868 28354 35924 28364
rect 37436 28420 37492 28430
rect 34972 28018 35028 28028
rect 34188 27970 34356 27972
rect 34188 27918 34190 27970
rect 34242 27918 34356 27970
rect 34188 27916 34356 27918
rect 34188 27906 34244 27916
rect 33908 27748 33964 27862
rect 33516 27300 33572 27310
rect 33292 27298 33572 27300
rect 33292 27246 33518 27298
rect 33570 27246 33572 27298
rect 33292 27244 33572 27246
rect 33516 27234 33572 27244
rect 33628 26908 33684 27692
rect 33908 27682 33964 27692
rect 34524 27858 34580 27870
rect 34524 27806 34526 27858
rect 34578 27806 34580 27858
rect 33796 27524 33852 27534
rect 33796 27076 33852 27468
rect 34524 27412 34580 27806
rect 34748 27860 34804 27870
rect 35868 27860 35924 27870
rect 37324 27860 37380 27870
rect 34748 27858 34916 27860
rect 34748 27806 34750 27858
rect 34802 27806 34916 27858
rect 34748 27804 34916 27806
rect 34748 27794 34804 27804
rect 34524 27346 34580 27356
rect 34188 27188 34244 27198
rect 33796 27018 33852 27020
rect 33796 26966 33798 27018
rect 33850 26966 33852 27018
rect 33796 26954 33852 26966
rect 33964 27044 34020 27056
rect 33964 26992 33966 27044
rect 34018 26992 34020 27044
rect 33180 26562 33236 26572
rect 33516 26852 33684 26908
rect 33964 26908 34020 26992
rect 34188 27035 34244 27132
rect 34188 26983 34190 27035
rect 34242 26983 34244 27035
rect 34188 26971 34244 26983
rect 34860 27036 34916 27804
rect 35868 27858 36316 27860
rect 35868 27806 35870 27858
rect 35922 27806 36316 27858
rect 35868 27804 36316 27806
rect 35868 27794 35924 27804
rect 34860 26984 34862 27036
rect 34914 26984 34916 27036
rect 35028 27634 35084 27646
rect 35028 27582 35030 27634
rect 35082 27582 35084 27634
rect 35028 27076 35084 27582
rect 35532 27636 35588 27646
rect 35532 27634 36148 27636
rect 35532 27582 35534 27634
rect 35586 27582 36148 27634
rect 35532 27580 36148 27582
rect 35532 27570 35588 27580
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35196 27300 35252 27310
rect 35252 27244 35364 27300
rect 35196 27234 35252 27244
rect 35028 27010 35084 27020
rect 35196 27074 35252 27086
rect 35196 27022 35198 27074
rect 35250 27022 35252 27074
rect 34860 26908 34916 26984
rect 33964 26852 34916 26908
rect 35196 26964 35252 27022
rect 35196 26898 35252 26908
rect 33516 26516 33572 26852
rect 33516 26450 33572 26460
rect 33740 26516 33796 26526
rect 33012 26346 33068 26358
rect 33012 26294 33014 26346
rect 33066 26294 33068 26346
rect 33012 26292 33068 26294
rect 33012 26226 33068 26236
rect 33180 26320 33236 26332
rect 33180 26268 33182 26320
rect 33234 26268 33236 26320
rect 33180 25956 33236 26268
rect 33180 25890 33236 25900
rect 33516 26320 33572 26332
rect 33516 26268 33518 26320
rect 33570 26268 33572 26320
rect 33516 25956 33572 26268
rect 33516 25890 33572 25900
rect 33068 25506 33124 25518
rect 33068 25454 33070 25506
rect 33122 25454 33124 25506
rect 33068 25172 33124 25454
rect 33068 25106 33124 25116
rect 32844 24892 33348 24948
rect 32396 24724 32452 24734
rect 32172 23202 32228 23212
rect 32284 23828 32340 23838
rect 31724 23102 31726 23154
rect 31778 23102 31780 23154
rect 31724 23090 31780 23102
rect 32284 23156 32340 23772
rect 32396 23268 32452 24668
rect 33180 24724 33236 24734
rect 33180 24630 33236 24668
rect 33068 24554 33124 24566
rect 33068 24502 33070 24554
rect 33122 24502 33124 24554
rect 33068 24276 33124 24502
rect 33068 24210 33124 24220
rect 33012 23604 33068 23614
rect 32844 23492 32900 23502
rect 32396 23202 32452 23212
rect 32732 23268 32788 23278
rect 32284 23090 32340 23100
rect 32564 23044 32620 23054
rect 32564 22950 32620 22988
rect 32004 22930 32060 22942
rect 32004 22878 32006 22930
rect 32058 22878 32060 22930
rect 31444 22372 31500 22540
rect 31556 22594 31668 22606
rect 31556 22542 31558 22594
rect 31610 22542 31668 22594
rect 31556 22540 31668 22542
rect 31724 22708 31780 22718
rect 31556 22530 31612 22540
rect 31724 22372 31780 22652
rect 32004 22596 32060 22878
rect 32732 22708 32788 23212
rect 32732 22642 32788 22652
rect 32004 22540 32564 22596
rect 31836 22372 31892 22382
rect 31444 22316 31668 22372
rect 31724 22370 31892 22372
rect 31724 22318 31838 22370
rect 31890 22318 31892 22370
rect 31724 22316 31892 22318
rect 30716 21756 30996 21812
rect 30716 21028 30772 21756
rect 30716 20972 31108 21028
rect 30940 20804 30996 20814
rect 30604 20748 30884 20804
rect 30604 20580 30660 20590
rect 30492 20578 30660 20580
rect 30492 20526 30606 20578
rect 30658 20526 30660 20578
rect 30492 20524 30660 20526
rect 30604 20514 30660 20524
rect 30604 20020 30660 20030
rect 30380 19842 30436 19852
rect 30492 20018 30660 20020
rect 30492 19966 30606 20018
rect 30658 19966 30660 20018
rect 30492 19964 30660 19966
rect 30492 19572 30548 19964
rect 30604 19954 30660 19964
rect 30044 19516 30548 19572
rect 30716 19850 30772 19862
rect 30716 19798 30718 19850
rect 30770 19798 30772 19850
rect 30716 19572 30772 19798
rect 30828 19572 30884 20748
rect 30940 20710 30996 20748
rect 31052 19796 31108 20972
rect 31276 20804 31332 20814
rect 31276 20634 31332 20748
rect 31388 20804 31444 20814
rect 31612 20804 31668 22316
rect 31836 22306 31892 22316
rect 32060 22372 32116 22382
rect 32060 22278 32116 22316
rect 32284 22372 32340 22382
rect 32284 22278 32340 22316
rect 32508 22352 32564 22540
rect 32732 22484 32788 22494
rect 32844 22484 32900 23436
rect 33012 23210 33068 23548
rect 33012 23158 33014 23210
rect 33066 23158 33068 23210
rect 33012 23146 33068 23158
rect 33180 23268 33236 23278
rect 33180 23210 33236 23212
rect 33180 23158 33182 23210
rect 33234 23158 33236 23210
rect 33180 23146 33236 23158
rect 32732 22482 32900 22484
rect 32732 22430 32734 22482
rect 32786 22430 32900 22482
rect 32732 22428 32900 22430
rect 32732 22418 32788 22428
rect 32956 22370 33012 22382
rect 33180 22372 33236 22382
rect 33292 22372 33348 24892
rect 33404 24722 33460 24734
rect 33404 24670 33406 24722
rect 33458 24670 33460 24722
rect 33404 23604 33460 24670
rect 33404 23538 33460 23548
rect 33516 23938 33572 23950
rect 33516 23886 33518 23938
rect 33570 23886 33572 23938
rect 33516 23492 33572 23886
rect 33740 23548 33796 26460
rect 33964 26402 34020 26852
rect 33964 26350 33966 26402
rect 34018 26350 34020 26402
rect 33964 26338 34020 26350
rect 34076 26740 34132 26750
rect 34076 25620 34132 26684
rect 34580 26740 34636 26750
rect 35308 26740 35364 27244
rect 35420 27244 36036 27300
rect 35420 27186 35476 27244
rect 35420 27134 35422 27186
rect 35474 27134 35476 27186
rect 35420 27122 35476 27134
rect 35756 27076 35812 27086
rect 35588 27018 35644 27030
rect 35588 26974 35590 27018
rect 34580 26514 34636 26684
rect 34580 26462 34582 26514
rect 34634 26462 34636 26514
rect 34580 26450 34636 26462
rect 35084 26684 35364 26740
rect 35532 26966 35590 26974
rect 35642 26966 35644 27018
rect 35756 26982 35812 27020
rect 35980 27074 36036 27244
rect 35980 27022 35982 27074
rect 36034 27022 36036 27074
rect 35980 27010 36036 27022
rect 35532 26964 35644 26966
rect 35588 26908 35644 26964
rect 35532 26740 35588 26908
rect 35084 26402 35140 26684
rect 35084 26350 35086 26402
rect 35138 26350 35140 26402
rect 35084 26338 35140 26350
rect 34748 25956 34804 25966
rect 34188 25732 34244 25742
rect 34188 25730 34692 25732
rect 34188 25678 34190 25730
rect 34242 25678 34692 25730
rect 34188 25676 34692 25678
rect 34188 25666 34244 25676
rect 34076 25554 34132 25564
rect 33944 25450 34000 25462
rect 33944 25398 33946 25450
rect 33998 25398 34000 25450
rect 33944 25284 34000 25398
rect 33944 25218 34000 25228
rect 34300 24722 34356 25676
rect 34636 25562 34692 25676
rect 34636 25510 34638 25562
rect 34690 25510 34692 25562
rect 34636 25498 34692 25510
rect 34748 25468 34804 25900
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35532 25732 35588 26684
rect 36092 26516 36148 27580
rect 36260 27298 36316 27804
rect 37156 27802 37212 27814
rect 36484 27748 36540 27758
rect 36932 27748 36988 27758
rect 37156 27750 37158 27802
rect 37210 27750 37212 27802
rect 37324 27766 37380 27804
rect 37156 27748 37212 27750
rect 36484 27746 36820 27748
rect 36484 27694 36486 27746
rect 36538 27694 36820 27746
rect 36484 27692 36820 27694
rect 36484 27682 36540 27692
rect 36260 27246 36262 27298
rect 36314 27246 36316 27298
rect 36260 27234 36316 27246
rect 36764 26740 36820 27692
rect 36932 27746 37212 27748
rect 36932 27694 36934 27746
rect 36986 27694 37212 27746
rect 36932 27692 37212 27694
rect 36932 27682 36988 27692
rect 37156 27524 37212 27692
rect 37156 27468 37268 27524
rect 36764 26674 36820 26684
rect 36092 26450 36148 26460
rect 37212 26516 37268 27468
rect 37212 26450 37268 26460
rect 37436 26872 37492 28364
rect 37660 27972 37716 28812
rect 37884 28756 37940 29374
rect 37996 29426 38052 29438
rect 37996 29374 37998 29426
rect 38050 29374 38052 29426
rect 37996 28980 38052 29374
rect 38332 29428 38388 30604
rect 38948 30548 39004 30558
rect 38500 30212 38556 30222
rect 38500 29876 38556 30156
rect 38948 30210 39004 30492
rect 39452 30548 39508 31164
rect 39452 30482 39508 30492
rect 39340 30324 39396 30334
rect 38948 30158 38950 30210
rect 39002 30158 39004 30210
rect 38948 30146 39004 30158
rect 39228 30212 39284 30222
rect 38780 30100 38836 30110
rect 38500 29820 38724 29876
rect 38556 29764 38612 29820
rect 38556 29698 38612 29708
rect 38556 29428 38612 29438
rect 38332 29426 38612 29428
rect 38332 29374 38558 29426
rect 38610 29374 38612 29426
rect 38332 29372 38612 29374
rect 38556 29362 38612 29372
rect 38276 29204 38332 29214
rect 37996 28914 38052 28924
rect 38220 29202 38332 29204
rect 38220 29150 38278 29202
rect 38330 29150 38332 29202
rect 38220 29138 38332 29150
rect 37884 28700 38052 28756
rect 37660 27916 37772 27972
rect 37716 27914 37772 27916
rect 37548 27858 37604 27870
rect 37548 27806 37550 27858
rect 37602 27806 37604 27858
rect 37716 27862 37718 27914
rect 37770 27862 37772 27914
rect 37716 27850 37772 27862
rect 37548 27636 37604 27806
rect 37548 27570 37604 27580
rect 37996 27636 38052 28700
rect 38220 27860 38276 29138
rect 38332 28980 38388 28990
rect 38332 28084 38388 28924
rect 38668 28980 38724 29820
rect 38780 29426 38836 30044
rect 39060 29652 39116 29662
rect 39060 29538 39116 29596
rect 39060 29486 39062 29538
rect 39114 29486 39116 29538
rect 39060 29474 39116 29486
rect 38780 29374 38782 29426
rect 38834 29374 38836 29426
rect 38780 29362 38836 29374
rect 38668 28914 38724 28924
rect 39228 28868 39284 30156
rect 39340 30210 39396 30268
rect 39340 30158 39342 30210
rect 39394 30158 39396 30210
rect 39676 30210 39732 31836
rect 39340 30146 39396 30158
rect 39508 30154 39564 30166
rect 39508 30102 39510 30154
rect 39562 30102 39564 30154
rect 39676 30158 39678 30210
rect 39730 30158 39732 30210
rect 39676 30146 39732 30158
rect 39508 29988 39564 30102
rect 39788 29988 39844 32396
rect 39228 28802 39284 28812
rect 39340 29932 39844 29988
rect 39340 28644 39396 29932
rect 39788 29426 39844 29438
rect 39788 29374 39790 29426
rect 39842 29374 39844 29426
rect 39620 29316 39676 29326
rect 39788 29316 39844 29374
rect 39620 29314 39844 29316
rect 39620 29262 39622 29314
rect 39674 29262 39844 29314
rect 39620 29260 39844 29262
rect 39620 29204 39676 29260
rect 39900 29204 39956 32732
rect 39620 29138 39676 29148
rect 39788 29148 39956 29204
rect 39228 28588 39396 28644
rect 39452 28642 39508 28654
rect 39452 28590 39454 28642
rect 39506 28590 39508 28642
rect 38332 28028 38612 28084
rect 38332 27860 38388 27870
rect 38220 27858 38388 27860
rect 38220 27806 38334 27858
rect 38386 27806 38388 27858
rect 38220 27804 38388 27806
rect 38332 27794 38388 27804
rect 38444 27860 38500 27870
rect 38444 27766 38500 27804
rect 37996 27570 38052 27580
rect 38388 27188 38444 27198
rect 37940 27086 37996 27096
rect 38388 27094 38444 27132
rect 37884 27076 37996 27086
rect 37940 27074 37996 27076
rect 37940 27022 37942 27074
rect 37994 27022 37996 27074
rect 37940 27020 37996 27022
rect 37884 27010 37996 27020
rect 38556 27076 38612 28028
rect 38724 27860 38780 27870
rect 39004 27860 39060 27870
rect 38724 27858 39060 27860
rect 38724 27806 38726 27858
rect 38778 27806 39006 27858
rect 39058 27806 39060 27858
rect 38724 27804 39060 27806
rect 38724 27794 38780 27804
rect 39004 27794 39060 27804
rect 39228 27636 39284 28588
rect 39340 28084 39396 28094
rect 39452 28084 39508 28590
rect 39340 28082 39508 28084
rect 39340 28030 39342 28082
rect 39394 28030 39508 28082
rect 39340 28028 39508 28030
rect 39340 28018 39396 28028
rect 39004 27580 39284 27636
rect 38892 27300 38948 27310
rect 38892 27242 38948 27244
rect 38556 27010 38612 27020
rect 38780 27188 38836 27198
rect 38892 27190 38894 27242
rect 38946 27190 38948 27242
rect 38892 27178 38948 27190
rect 38780 27074 38836 27132
rect 38780 27022 38782 27074
rect 38834 27022 38836 27074
rect 38780 27010 38836 27022
rect 37436 26850 37548 26872
rect 37436 26798 37494 26850
rect 37546 26798 37548 26850
rect 37436 26786 37548 26798
rect 37884 26852 37940 27010
rect 39004 26852 39060 27580
rect 39788 27412 39844 29148
rect 40012 27860 40068 32844
rect 40124 32786 40180 33852
rect 40124 32734 40126 32786
rect 40178 32734 40180 32786
rect 40124 32722 40180 32734
rect 40236 32788 40292 34636
rect 40236 32722 40292 32732
rect 40460 32562 40516 32574
rect 40460 32510 40462 32562
rect 40514 32510 40516 32562
rect 40460 32452 40516 32510
rect 40460 32386 40516 32396
rect 40236 31668 40292 31678
rect 40236 31106 40292 31612
rect 40236 31054 40238 31106
rect 40290 31054 40292 31106
rect 40236 31042 40292 31054
rect 40404 31666 40460 31678
rect 40404 31614 40406 31666
rect 40458 31614 40460 31666
rect 40404 31108 40460 31614
rect 40404 31042 40460 31052
rect 40572 30660 40628 36204
rect 40796 36036 40852 36374
rect 41020 36426 41076 36438
rect 41020 36374 41022 36426
rect 41074 36374 41076 36426
rect 41132 36395 41134 36428
rect 41186 36395 41188 36428
rect 41132 36383 41188 36395
rect 41804 36484 41860 36494
rect 41804 36402 41806 36428
rect 41858 36402 41860 36428
rect 41804 36390 41860 36402
rect 42028 36454 42084 36988
rect 42140 36708 42196 37660
rect 42252 37266 42308 37278
rect 42252 37214 42254 37266
rect 42306 37214 42308 37266
rect 42252 36932 42308 37214
rect 42252 36866 42308 36876
rect 42140 36652 42308 36708
rect 42028 36402 42030 36454
rect 42082 36402 42084 36454
rect 42028 36390 42084 36402
rect 42252 36454 42308 36652
rect 42252 36402 42254 36454
rect 42306 36402 42308 36454
rect 42252 36390 42308 36402
rect 42364 36426 42420 36438
rect 41020 36372 41076 36374
rect 41020 36306 41076 36316
rect 41692 36372 41748 36382
rect 40796 35980 40964 36036
rect 40796 35812 40852 35822
rect 40796 35698 40852 35756
rect 40796 35646 40798 35698
rect 40850 35646 40852 35698
rect 40796 35634 40852 35646
rect 40908 34916 40964 35980
rect 41468 35700 41524 35710
rect 41468 35606 41524 35644
rect 41132 35476 41188 35486
rect 41132 35382 41188 35420
rect 41692 35476 41748 36316
rect 42364 36374 42366 36426
rect 42418 36374 42420 36426
rect 41804 36036 41860 36046
rect 41804 35922 41860 35980
rect 42364 35924 42420 36374
rect 41804 35870 41806 35922
rect 41858 35870 41860 35922
rect 41804 35858 41860 35870
rect 42028 35868 42420 35924
rect 42476 35924 42532 38612
rect 42588 38022 42644 38668
rect 42588 37970 42590 38022
rect 42642 37970 42644 38022
rect 42588 37958 42644 37970
rect 42700 37828 42756 39340
rect 42812 39172 42868 39182
rect 42812 38836 42868 39116
rect 42812 38022 42868 38780
rect 43036 38948 43092 38958
rect 43036 38500 43092 38892
rect 43148 38836 43204 38846
rect 43260 38836 43316 40460
rect 43372 40402 43428 40460
rect 43652 40458 43708 40684
rect 43372 40350 43374 40402
rect 43426 40350 43428 40402
rect 43372 40338 43428 40350
rect 43484 40402 43540 40414
rect 43484 40350 43486 40402
rect 43538 40350 43540 40402
rect 43652 40406 43654 40458
rect 43706 40406 43708 40458
rect 43652 40394 43708 40406
rect 43148 38834 43316 38836
rect 43148 38782 43150 38834
rect 43202 38782 43316 38834
rect 43148 38780 43316 38782
rect 43372 40180 43428 40190
rect 43372 38834 43428 40124
rect 43484 39956 43540 40350
rect 43820 40292 43876 40796
rect 43932 40404 43988 41096
rect 43932 40338 43988 40348
rect 44380 40404 44436 41804
rect 44492 41794 44548 41804
rect 44828 42026 44884 42364
rect 44828 41974 44830 42026
rect 44882 41974 44884 42026
rect 44380 40338 44436 40348
rect 44492 41412 44548 41422
rect 44492 40402 44548 41356
rect 44828 41188 44884 41974
rect 44828 41122 44884 41132
rect 44940 40964 44996 40974
rect 44492 40350 44494 40402
rect 44546 40350 44548 40402
rect 44492 40338 44548 40350
rect 44604 40962 44996 40964
rect 44604 40910 44942 40962
rect 44994 40910 44996 40962
rect 44604 40908 44996 40910
rect 44604 40404 44660 40908
rect 44940 40898 44996 40908
rect 45052 40964 45108 42674
rect 45052 40898 45108 40908
rect 44604 40338 44660 40348
rect 43484 39890 43540 39900
rect 43596 40236 43876 40292
rect 43372 38782 43374 38834
rect 43426 38782 43428 38834
rect 43148 38770 43204 38780
rect 43372 38770 43428 38782
rect 43484 38668 43540 38678
rect 43596 38668 43652 40236
rect 43932 40180 43988 40190
rect 43932 39060 43988 40124
rect 44044 40180 44100 40190
rect 45164 40180 45220 43652
rect 45388 43538 45444 43550
rect 45388 43486 45390 43538
rect 45442 43486 45444 43538
rect 45276 41748 45332 41758
rect 45276 41654 45332 41692
rect 45276 41186 45332 41198
rect 45276 41134 45278 41186
rect 45330 41134 45332 41186
rect 45276 40628 45332 41134
rect 45388 41188 45444 43486
rect 45836 42980 45892 42990
rect 45836 42886 45892 42924
rect 45724 41997 45780 42009
rect 45724 41945 45726 41997
rect 45778 41945 45780 41997
rect 45724 41860 45780 41945
rect 45724 41794 45780 41804
rect 46060 41860 46116 45500
rect 46172 45220 46228 45230
rect 46172 45106 46228 45164
rect 46172 45054 46174 45106
rect 46226 45054 46228 45106
rect 46172 45042 46228 45054
rect 46396 44436 46452 45836
rect 46508 45826 46564 45836
rect 47348 45834 47404 45846
rect 46788 45778 46844 45790
rect 46788 45726 46790 45778
rect 46842 45726 46844 45778
rect 46788 45444 46844 45726
rect 46788 45378 46844 45388
rect 47348 45782 47350 45834
rect 47402 45782 47404 45834
rect 48076 45800 48078 45852
rect 48130 45800 48132 45852
rect 47348 45220 47404 45782
rect 47516 45780 47572 45790
rect 48076 45788 48132 45800
rect 48188 45834 48244 45846
rect 48188 45782 48190 45834
rect 48242 45782 48244 45834
rect 47516 45778 47684 45780
rect 47516 45726 47518 45778
rect 47570 45726 47684 45778
rect 47516 45724 47684 45726
rect 47516 45714 47572 45724
rect 46396 44370 46452 44380
rect 47292 45164 47404 45220
rect 47516 45444 47572 45454
rect 47180 44294 47236 44306
rect 47180 44242 47182 44294
rect 47234 44242 47236 44294
rect 47180 43876 47236 44242
rect 47180 43810 47236 43820
rect 46396 43652 46452 43662
rect 46172 43428 46228 43438
rect 46172 43426 46340 43428
rect 46172 43374 46174 43426
rect 46226 43374 46340 43426
rect 46172 43372 46340 43374
rect 46172 43362 46228 43372
rect 46060 41794 46116 41804
rect 46172 41188 46228 41198
rect 45388 41186 45556 41188
rect 45388 41134 45390 41186
rect 45442 41134 45556 41186
rect 45388 41132 45556 41134
rect 45388 41122 45444 41132
rect 45276 40562 45332 40572
rect 45388 40964 45444 40974
rect 45388 40516 45444 40908
rect 45368 40460 45444 40516
rect 45368 40458 45424 40460
rect 45368 40406 45370 40458
rect 45422 40406 45424 40458
rect 45368 40394 45424 40406
rect 44044 40178 44324 40180
rect 44044 40126 44046 40178
rect 44098 40126 44324 40178
rect 44044 40124 44324 40126
rect 45164 40124 45444 40180
rect 44044 40114 44100 40124
rect 44268 39844 44324 40124
rect 44828 39956 44884 39966
rect 44268 39788 44548 39844
rect 44044 39506 44100 39518
rect 44044 39454 44046 39506
rect 44098 39454 44100 39506
rect 44044 39284 44100 39454
rect 44044 39218 44100 39228
rect 43932 39004 44100 39060
rect 43876 38836 43932 38846
rect 43876 38742 43932 38780
rect 43484 38666 43652 38668
rect 43372 38612 43428 38622
rect 43484 38614 43486 38666
rect 43538 38614 43652 38666
rect 43484 38612 43652 38614
rect 43708 38612 43764 38622
rect 43484 38602 43540 38612
rect 43036 38444 43316 38500
rect 43260 38218 43316 38444
rect 43260 38166 43262 38218
rect 43314 38166 43316 38218
rect 43260 38154 43316 38166
rect 42812 37970 42814 38022
rect 42866 37970 42868 38022
rect 43372 38050 43428 38556
rect 42812 37958 42868 37970
rect 42924 37994 42980 38006
rect 42700 37762 42756 37772
rect 42924 37942 42926 37994
rect 42978 37942 42980 37994
rect 43372 37998 43374 38050
rect 43426 37998 43428 38050
rect 43372 37986 43428 37998
rect 43484 38276 43540 38286
rect 42924 37492 42980 37942
rect 42924 37426 42980 37436
rect 43372 37716 43428 37726
rect 43372 37490 43428 37660
rect 43372 37438 43374 37490
rect 43426 37438 43428 37490
rect 42924 37268 42980 37278
rect 42924 37266 43092 37268
rect 42924 37214 42926 37266
rect 42978 37214 43092 37266
rect 42924 37212 43092 37214
rect 42924 37202 42980 37212
rect 42588 37044 42644 37054
rect 42644 36988 42756 37044
rect 42588 36950 42644 36988
rect 41132 35028 41188 35038
rect 41132 34934 41188 34972
rect 40908 34850 40964 34860
rect 41244 34898 41580 34916
rect 41244 34860 41526 34898
rect 40796 34132 40852 34142
rect 41244 34132 41300 34860
rect 41524 34846 41526 34860
rect 41578 34846 41580 34898
rect 41524 34834 41580 34846
rect 41692 34886 41748 35420
rect 42028 35364 42084 35868
rect 42476 35830 42532 35868
rect 42588 36596 42644 36606
rect 42140 35700 42196 35710
rect 42140 35698 42308 35700
rect 42140 35646 42142 35698
rect 42194 35646 42308 35698
rect 42140 35644 42308 35646
rect 42140 35634 42196 35644
rect 42028 35308 42196 35364
rect 42140 35028 42196 35308
rect 41692 34834 41694 34886
rect 41746 34834 41748 34886
rect 40796 34038 40852 34076
rect 40908 34076 41412 34132
rect 40796 33460 40852 33470
rect 40908 33460 40964 34076
rect 41132 33906 41188 33918
rect 41132 33854 41134 33906
rect 41186 33854 41188 33906
rect 41132 33684 41188 33854
rect 41132 33618 41188 33628
rect 40796 33458 40964 33460
rect 40796 33406 40798 33458
rect 40850 33406 40964 33458
rect 40796 33404 40964 33406
rect 41244 33572 41300 33582
rect 40796 33394 40852 33404
rect 41020 32788 41076 32798
rect 41020 32618 41076 32732
rect 40852 32578 40908 32590
rect 40852 32564 40854 32578
rect 40684 32526 40854 32564
rect 40906 32526 40908 32578
rect 41020 32566 41022 32618
rect 41074 32566 41076 32618
rect 41020 32554 41076 32566
rect 41244 32618 41300 33516
rect 41356 33012 41412 34076
rect 41468 34130 41524 34142
rect 41468 34078 41470 34130
rect 41522 34078 41524 34130
rect 41468 33908 41524 34078
rect 41468 33842 41524 33852
rect 41524 33236 41580 33246
rect 41524 33234 41636 33236
rect 41524 33182 41526 33234
rect 41578 33182 41636 33234
rect 41524 33170 41636 33182
rect 41356 32956 41524 33012
rect 41244 32566 41246 32618
rect 41298 32566 41300 32618
rect 40684 32508 40908 32526
rect 40684 31722 40740 32508
rect 41244 32452 41300 32566
rect 40684 31670 40686 31722
rect 40738 31670 40740 31722
rect 40908 32396 41300 32452
rect 41356 32788 41412 32798
rect 40908 31750 40964 32396
rect 41356 32340 41412 32732
rect 41468 32618 41524 32956
rect 41468 32566 41470 32618
rect 41522 32566 41524 32618
rect 41468 32554 41524 32566
rect 40908 31698 40910 31750
rect 40962 31698 40964 31750
rect 40908 31686 40964 31698
rect 41132 32284 41412 32340
rect 41132 31750 41188 32284
rect 41580 32116 41636 33170
rect 41692 32788 41748 34834
rect 41916 34916 41972 34926
rect 41916 34834 41918 34860
rect 41970 34834 41972 34860
rect 41804 34356 41860 34366
rect 41916 34356 41972 34834
rect 42140 34886 42196 34972
rect 42140 34834 42142 34886
rect 42194 34834 42196 34886
rect 42140 34822 42196 34834
rect 41804 34354 41972 34356
rect 41804 34302 41806 34354
rect 41858 34302 41972 34354
rect 41804 34300 41972 34302
rect 41804 33572 41860 34300
rect 42252 33582 42308 35644
rect 42420 35252 42476 35262
rect 42420 35138 42476 35196
rect 42420 35086 42422 35138
rect 42474 35086 42476 35138
rect 42420 35074 42476 35086
rect 42588 34130 42644 36540
rect 42588 34078 42590 34130
rect 42642 34078 42644 34130
rect 42588 34066 42644 34078
rect 42420 34020 42476 34030
rect 42420 33926 42476 33964
rect 42588 33908 42644 33918
rect 42700 33908 42756 36988
rect 43036 36932 43092 37212
rect 42868 36596 42924 36606
rect 42868 36502 42924 36540
rect 42644 33852 42756 33908
rect 42812 35924 42868 35934
rect 42252 33570 42364 33582
rect 42252 33518 42310 33570
rect 42362 33518 42364 33570
rect 42252 33516 42364 33518
rect 41804 33506 41860 33516
rect 42308 33506 42364 33516
rect 41804 33348 41860 33358
rect 41804 33254 41860 33292
rect 41916 33346 41972 33358
rect 41916 33294 41918 33346
rect 41970 33294 41972 33346
rect 41692 32722 41748 32732
rect 41748 32564 41804 32574
rect 41748 32470 41804 32508
rect 41580 32060 41748 32116
rect 41132 31698 41134 31750
rect 41186 31698 41188 31750
rect 41132 31686 41188 31698
rect 41244 32004 41300 32014
rect 41244 31743 41300 31948
rect 41580 31892 41636 31902
rect 41244 31691 41246 31743
rect 41298 31691 41300 31743
rect 40684 31668 40740 31670
rect 40684 31602 40740 31612
rect 41244 31556 41300 31691
rect 41020 31500 41300 31556
rect 41356 31890 41636 31892
rect 41356 31838 41582 31890
rect 41634 31838 41636 31890
rect 41356 31836 41636 31838
rect 41020 31106 41076 31500
rect 41020 31054 41022 31106
rect 41074 31054 41076 31106
rect 41020 31042 41076 31054
rect 40572 30594 40628 30604
rect 41020 30322 41076 30334
rect 41020 30270 41022 30322
rect 41074 30270 41076 30322
rect 40236 30182 40292 30194
rect 40236 30130 40238 30182
rect 40290 30130 40292 30182
rect 40236 29988 40292 30130
rect 40236 29652 40292 29932
rect 40236 29586 40292 29596
rect 40572 29428 40628 29438
rect 40236 29204 40292 29214
rect 40124 28868 40180 28878
rect 40124 28420 40180 28812
rect 40236 28642 40292 29148
rect 40572 28756 40628 29372
rect 40796 29428 40852 29438
rect 41020 29428 41076 30270
rect 40796 29426 41076 29428
rect 40796 29374 40798 29426
rect 40850 29374 41076 29426
rect 40796 29372 41076 29374
rect 40796 29362 40852 29372
rect 40236 28590 40238 28642
rect 40290 28590 40292 28642
rect 40236 28578 40292 28590
rect 40460 28754 40628 28756
rect 40460 28702 40574 28754
rect 40626 28702 40628 28754
rect 40460 28700 40628 28702
rect 40124 28364 40292 28420
rect 40012 27804 40180 27860
rect 39956 27636 40012 27646
rect 40124 27636 40180 27804
rect 40236 27858 40292 28364
rect 40236 27806 40238 27858
rect 40290 27806 40292 27858
rect 40236 27794 40292 27806
rect 40460 27858 40516 28700
rect 40572 28690 40628 28700
rect 41020 28644 41076 29372
rect 41244 29204 41300 29214
rect 41020 28578 41076 28588
rect 41132 28980 41188 28990
rect 41132 28026 41188 28924
rect 41132 27974 41134 28026
rect 41186 27974 41188 28026
rect 41132 27962 41188 27974
rect 41244 28756 41300 29148
rect 40460 27806 40462 27858
rect 40514 27806 40516 27858
rect 40460 27794 40516 27806
rect 41020 27860 41076 27870
rect 40124 27580 40292 27636
rect 39956 27542 40012 27580
rect 39788 27356 40180 27412
rect 39340 27300 39396 27310
rect 39228 27188 39284 27198
rect 37884 26786 37940 26796
rect 38668 26796 39060 26852
rect 39116 27074 39172 27086
rect 39116 27022 39118 27074
rect 39170 27022 39172 27074
rect 36988 26180 37044 26190
rect 36988 26086 37044 26124
rect 35476 25676 35588 25732
rect 35476 25620 35532 25676
rect 35196 25564 35532 25620
rect 34748 25416 34750 25468
rect 34802 25416 34804 25468
rect 34748 25060 34804 25416
rect 34300 24670 34302 24722
rect 34354 24670 34356 24722
rect 34300 24658 34356 24670
rect 34412 25004 34804 25060
rect 34860 25508 34916 25518
rect 34412 24722 34468 25004
rect 34692 24836 34748 24846
rect 34860 24836 34916 25452
rect 35196 25172 35252 25564
rect 35476 25562 35532 25564
rect 35476 25510 35478 25562
rect 35530 25510 35532 25562
rect 35476 25498 35532 25510
rect 35644 25508 35700 25518
rect 35644 25414 35700 25452
rect 35868 25506 35924 25518
rect 35868 25454 35870 25506
rect 35922 25454 35924 25506
rect 35308 25394 35364 25406
rect 35308 25342 35310 25394
rect 35362 25342 35364 25394
rect 35308 25284 35364 25342
rect 35868 25284 35924 25454
rect 36148 25508 36204 25518
rect 36876 25508 36932 25518
rect 36148 25506 36932 25508
rect 36148 25454 36150 25506
rect 36202 25454 36878 25506
rect 36930 25454 36932 25506
rect 36148 25452 36932 25454
rect 36148 25442 36204 25452
rect 36876 25442 36932 25452
rect 35308 25228 35924 25284
rect 37212 25284 37268 25294
rect 37212 25190 37268 25228
rect 35196 25116 35308 25172
rect 35252 24946 35308 25116
rect 35252 24894 35254 24946
rect 35306 24894 35308 24946
rect 35252 24882 35308 24894
rect 35644 25060 35700 25070
rect 34692 24834 34916 24836
rect 34692 24782 34694 24834
rect 34746 24782 34916 24834
rect 34692 24780 34916 24782
rect 35644 24834 35700 25004
rect 35644 24782 35646 24834
rect 35698 24782 35700 24834
rect 34692 24770 34748 24780
rect 35644 24770 35700 24782
rect 34412 24670 34414 24722
rect 34466 24670 34468 24722
rect 34020 24612 34076 24622
rect 34020 24610 34132 24612
rect 34020 24558 34022 24610
rect 34074 24558 34132 24610
rect 34020 24546 34132 24558
rect 34076 23940 34132 24546
rect 34300 23940 34356 23950
rect 34076 23938 34356 23940
rect 34076 23886 34302 23938
rect 34354 23886 34356 23938
rect 34076 23884 34356 23886
rect 33516 23426 33572 23436
rect 33628 23492 33796 23548
rect 34300 23604 34356 23884
rect 34300 23538 34356 23548
rect 33404 23193 33460 23205
rect 33404 23141 33406 23193
rect 33458 23141 33460 23193
rect 33404 22606 33460 23141
rect 33404 22596 33516 22606
rect 33404 22540 33460 22596
rect 33460 22502 33516 22540
rect 32508 22340 32620 22352
rect 32508 22288 32566 22340
rect 32618 22288 32620 22340
rect 32508 22286 32620 22288
rect 32564 22276 32620 22286
rect 32956 22318 32958 22370
rect 33010 22318 33012 22370
rect 32396 21700 32452 21710
rect 32956 21700 33012 22318
rect 32396 21698 33012 21700
rect 32396 21646 32398 21698
rect 32450 21646 33012 21698
rect 32396 21644 33012 21646
rect 33068 22370 33348 22372
rect 33068 22318 33182 22370
rect 33234 22318 33348 22370
rect 33068 22316 33348 22318
rect 32396 21634 32452 21644
rect 32060 21588 32116 21598
rect 32060 21364 32116 21532
rect 31388 20802 31668 20804
rect 31388 20750 31390 20802
rect 31442 20750 31668 20802
rect 31388 20748 31668 20750
rect 31724 20916 31780 20926
rect 31724 20775 31780 20860
rect 31388 20738 31444 20748
rect 31724 20723 31726 20775
rect 31778 20723 31780 20775
rect 31724 20711 31780 20723
rect 32060 20802 32116 21308
rect 32396 20916 32452 20926
rect 32396 20822 32452 20860
rect 32060 20750 32062 20802
rect 32114 20750 32116 20802
rect 32732 20802 32788 21644
rect 31276 20582 31278 20634
rect 31330 20582 31332 20634
rect 31276 20570 31332 20582
rect 31220 20356 31276 20366
rect 31220 20130 31276 20300
rect 32060 20356 32116 20750
rect 32564 20746 32620 20758
rect 32564 20694 32566 20746
rect 32618 20694 32620 20746
rect 32732 20750 32734 20802
rect 32786 20750 32788 20802
rect 32732 20738 32788 20750
rect 32564 20692 32620 20694
rect 32564 20636 32676 20692
rect 32620 20580 32676 20636
rect 33068 20580 33124 22316
rect 33180 22306 33236 22316
rect 33516 21812 33572 21822
rect 33236 21588 33292 21598
rect 33236 21494 33292 21532
rect 33404 21586 33460 21598
rect 33404 21534 33406 21586
rect 33458 21534 33460 21586
rect 33292 20970 33348 20982
rect 33292 20918 33294 20970
rect 33346 20918 33348 20970
rect 32620 20524 33124 20580
rect 33180 20802 33236 20814
rect 33180 20750 33182 20802
rect 33234 20750 33236 20802
rect 33180 20468 33236 20750
rect 32060 20290 32116 20300
rect 32732 20412 33236 20468
rect 31220 20078 31222 20130
rect 31274 20078 31276 20130
rect 31220 20066 31276 20078
rect 32060 20132 32116 20142
rect 31724 20020 31780 20030
rect 31836 20020 31892 20030
rect 31724 20018 31836 20020
rect 31724 19966 31726 20018
rect 31778 19966 31836 20018
rect 31724 19964 31836 19966
rect 31724 19954 31780 19964
rect 31556 19796 31612 19806
rect 31052 19740 31220 19796
rect 31052 19572 31108 19582
rect 30828 19516 30996 19572
rect 30044 17780 30100 19516
rect 30716 19506 30772 19516
rect 30940 18116 30996 19516
rect 30044 17714 30100 17724
rect 30548 18060 30996 18116
rect 30548 17780 30604 18060
rect 30716 17892 30772 17902
rect 30548 17778 30660 17780
rect 30548 17726 30550 17778
rect 30602 17726 30660 17778
rect 30548 17714 30660 17726
rect 28868 16942 28870 16994
rect 28922 16942 28980 16994
rect 28868 16940 28980 16942
rect 29820 16940 29988 16996
rect 28868 16930 28924 16940
rect 29652 16548 29708 16558
rect 28700 16380 28868 16436
rect 27972 15362 28028 15372
rect 27692 15262 27694 15314
rect 27746 15262 27748 15314
rect 27692 15250 27748 15262
rect 28140 15316 28196 15484
rect 28140 15250 28196 15260
rect 28364 16324 28420 16334
rect 28364 15148 28420 16268
rect 28700 16098 28756 16110
rect 28700 16046 28702 16098
rect 28754 16046 28756 16098
rect 28532 15988 28588 15998
rect 28532 15930 28588 15932
rect 28532 15878 28534 15930
rect 28586 15878 28588 15930
rect 28532 15866 28588 15878
rect 28700 15764 28756 16046
rect 28700 15698 28756 15708
rect 28532 15316 28588 15326
rect 28532 15222 28588 15260
rect 28364 15092 28588 15148
rect 27356 13356 27636 13412
rect 27692 14980 27748 14990
rect 27692 13412 27748 14924
rect 28532 14754 28588 15092
rect 28812 14980 28868 16380
rect 29652 16154 29708 16492
rect 29148 16100 29204 16110
rect 29148 15540 29204 16044
rect 29484 16098 29540 16110
rect 29484 16046 29486 16098
rect 29538 16046 29540 16098
rect 29652 16102 29654 16154
rect 29706 16102 29708 16154
rect 29652 16090 29708 16102
rect 29820 16100 29876 16940
rect 29932 16772 29988 16782
rect 29932 16770 30100 16772
rect 29932 16718 29934 16770
rect 29986 16718 30100 16770
rect 29932 16716 30100 16718
rect 29932 16706 29988 16716
rect 29484 15876 29540 16046
rect 29820 16006 29876 16044
rect 29932 16098 29988 16110
rect 29932 16046 29934 16098
rect 29986 16046 29988 16098
rect 29932 15876 29988 16046
rect 29484 15820 29876 15876
rect 29148 15428 29204 15484
rect 29148 15372 29316 15428
rect 28924 15314 28980 15326
rect 28924 15262 28926 15314
rect 28978 15262 28980 15314
rect 29260 15314 29316 15372
rect 28924 15092 28980 15262
rect 29092 15258 29148 15270
rect 29092 15206 29094 15258
rect 29146 15206 29148 15258
rect 29260 15262 29262 15314
rect 29314 15262 29316 15314
rect 29260 15250 29316 15262
rect 29372 15316 29428 15326
rect 29372 15222 29428 15260
rect 29092 15092 29148 15206
rect 29652 15204 29708 15242
rect 29652 15138 29708 15148
rect 28924 15026 28980 15036
rect 29036 15036 29148 15092
rect 29820 15092 29876 15820
rect 29932 15316 29988 15820
rect 30044 15764 30100 16716
rect 30604 16212 30660 17714
rect 30716 17666 30772 17836
rect 30716 17614 30718 17666
rect 30770 17614 30772 17666
rect 30716 17602 30772 17614
rect 31052 17220 31108 19516
rect 31164 17332 31220 19740
rect 31556 19794 31668 19796
rect 31556 19742 31558 19794
rect 31610 19742 31668 19794
rect 31556 19730 31668 19742
rect 31612 18116 31668 19730
rect 31724 19348 31780 19358
rect 31724 19254 31780 19292
rect 31724 18564 31780 18574
rect 31836 18564 31892 19964
rect 31724 18562 31892 18564
rect 31724 18510 31726 18562
rect 31778 18510 31892 18562
rect 31724 18508 31892 18510
rect 32060 20018 32116 20076
rect 32732 20132 32788 20412
rect 33292 20356 33348 20918
rect 32732 20066 32788 20076
rect 32844 20300 33348 20356
rect 32060 19966 32062 20018
rect 32114 19966 32116 20018
rect 32060 19348 32116 19966
rect 32284 20018 32340 20030
rect 32284 19966 32286 20018
rect 32338 19966 32340 20018
rect 32284 19908 32340 19966
rect 32284 19842 32340 19852
rect 32396 19850 32452 19862
rect 31724 18498 31780 18508
rect 32060 18452 32116 19292
rect 32396 19798 32398 19850
rect 32450 19798 32452 19850
rect 32396 19348 32452 19798
rect 32396 19282 32452 19292
rect 32620 19206 32676 19218
rect 32620 19154 32622 19206
rect 32674 19154 32676 19206
rect 32340 19122 32396 19134
rect 32340 19070 32342 19122
rect 32394 19070 32396 19122
rect 32340 18676 32396 19070
rect 32620 19012 32676 19154
rect 32844 19206 32900 20300
rect 33404 20244 33460 21534
rect 33516 20802 33572 21756
rect 33516 20750 33518 20802
rect 33570 20750 33572 20802
rect 33516 20738 33572 20750
rect 33292 20188 33460 20244
rect 33628 20244 33684 23492
rect 34412 23380 34468 24670
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 36092 24052 36148 24062
rect 35308 23938 35364 23950
rect 35308 23886 35310 23938
rect 35362 23886 35364 23938
rect 35308 23828 35364 23886
rect 35756 23938 35812 23950
rect 35756 23886 35758 23938
rect 35810 23886 35812 23938
rect 35308 23772 35700 23828
rect 35644 23770 35700 23772
rect 34972 23714 35028 23726
rect 34972 23662 34974 23714
rect 35026 23662 35028 23714
rect 35644 23718 35646 23770
rect 35698 23718 35700 23770
rect 35644 23706 35700 23718
rect 33964 23324 34468 23380
rect 34636 23492 34692 23502
rect 34636 23378 34692 23436
rect 34636 23326 34638 23378
rect 34690 23326 34692 23378
rect 33964 23266 34020 23324
rect 34636 23314 34692 23326
rect 34972 23380 35028 23662
rect 34972 23314 35028 23324
rect 35084 23604 35140 23614
rect 35756 23604 35812 23886
rect 36092 23911 36148 23996
rect 36988 24052 37044 24062
rect 36988 23958 37044 23996
rect 36092 23859 36094 23911
rect 36146 23859 36148 23911
rect 36428 23940 36484 23950
rect 37100 23940 37156 23950
rect 36428 23938 36932 23940
rect 36428 23886 36430 23938
rect 36482 23886 36932 23938
rect 36428 23884 36932 23886
rect 36428 23874 36484 23884
rect 36092 23847 36148 23859
rect 36876 23828 36932 23884
rect 35756 23548 36036 23604
rect 33964 23214 33966 23266
rect 34018 23214 34020 23266
rect 33964 23202 34020 23214
rect 34300 23154 34356 23166
rect 34300 23102 34302 23154
rect 34354 23102 34356 23154
rect 34300 23044 34356 23102
rect 34972 23156 35028 23166
rect 35084 23156 35140 23548
rect 34972 23154 35140 23156
rect 34972 23102 34974 23154
rect 35026 23102 35140 23154
rect 34972 23100 35140 23102
rect 35756 23380 35812 23390
rect 35756 23154 35812 23324
rect 35756 23102 35758 23154
rect 35810 23102 35812 23154
rect 34972 23090 35028 23100
rect 35756 23090 35812 23102
rect 34300 22978 34356 22988
rect 33964 22932 34020 22942
rect 33964 22594 34020 22876
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 33964 22542 33966 22594
rect 34018 22542 34020 22594
rect 33964 22530 34020 22542
rect 34300 22372 34356 22382
rect 34076 22370 34356 22372
rect 34076 22318 34302 22370
rect 34354 22318 34356 22370
rect 34076 22316 34356 22318
rect 33012 20020 33068 20030
rect 33012 19926 33068 19964
rect 33180 19906 33236 19918
rect 33180 19854 33182 19906
rect 33234 19854 33236 19906
rect 33180 19572 33236 19854
rect 32844 19154 32846 19206
rect 32898 19154 32900 19206
rect 32844 19142 32900 19154
rect 32956 19516 33236 19572
rect 32956 19012 33012 19516
rect 33180 19348 33236 19358
rect 33180 19199 33236 19292
rect 32620 18956 33012 19012
rect 33068 19178 33124 19190
rect 33068 19126 33070 19178
rect 33122 19126 33124 19178
rect 33180 19147 33182 19199
rect 33234 19147 33236 19199
rect 33180 19135 33236 19147
rect 33068 18788 33124 19126
rect 33068 18732 33236 18788
rect 32340 18610 32396 18620
rect 33180 18562 33236 18732
rect 33012 18506 33068 18518
rect 32396 18452 32452 18462
rect 32060 18450 32452 18452
rect 32060 18398 32398 18450
rect 32450 18398 32452 18450
rect 32060 18396 32452 18398
rect 32396 18386 32452 18396
rect 33012 18454 33014 18506
rect 33066 18454 33068 18506
rect 33180 18510 33182 18562
rect 33234 18510 33236 18562
rect 33180 18498 33236 18510
rect 32228 18228 32284 18238
rect 32228 18134 32284 18172
rect 31612 18050 31668 18060
rect 33012 18116 33068 18454
rect 33012 18050 33068 18060
rect 33292 18004 33348 20188
rect 33628 20178 33684 20188
rect 33740 21700 33796 21710
rect 33740 20074 33796 21644
rect 34076 21476 34132 22316
rect 34300 22306 34356 22316
rect 34412 22370 34468 22382
rect 34412 22318 34414 22370
rect 34466 22318 34468 22370
rect 34412 21812 34468 22318
rect 34636 22370 34692 22382
rect 34636 22318 34638 22370
rect 34690 22318 34692 22370
rect 34636 22148 34692 22318
rect 34916 22372 34972 22382
rect 34916 22278 34972 22316
rect 35644 22372 35700 22382
rect 35644 22278 35700 22316
rect 35868 22372 35924 22382
rect 35868 22278 35924 22316
rect 35364 22260 35420 22270
rect 35364 22258 35588 22260
rect 35364 22206 35366 22258
rect 35418 22206 35588 22258
rect 35364 22204 35588 22206
rect 35364 22194 35420 22204
rect 34636 22082 34692 22092
rect 34412 21746 34468 21756
rect 34076 21410 34132 21420
rect 34188 21476 34244 21486
rect 34188 21474 34468 21476
rect 34188 21422 34190 21474
rect 34242 21422 34468 21474
rect 34188 21420 34468 21422
rect 34188 21410 34244 21420
rect 34412 21028 34468 21420
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 34524 21028 34580 21038
rect 35532 21028 35588 22204
rect 35980 22148 36036 23548
rect 36260 22484 36316 22494
rect 36876 22484 36932 23772
rect 37100 23871 37102 23884
rect 37154 23871 37156 23884
rect 37100 23380 37156 23871
rect 37324 23938 37380 23950
rect 37324 23886 37326 23938
rect 37378 23886 37380 23938
rect 37324 23492 37380 23886
rect 37436 23828 37492 26786
rect 37660 26740 37716 26750
rect 37660 26292 37716 26684
rect 37772 26292 37828 26302
rect 38164 26292 38220 26302
rect 37660 26290 38220 26292
rect 37660 26238 37774 26290
rect 37826 26238 38166 26290
rect 38218 26238 38220 26290
rect 37660 26236 38220 26238
rect 37660 25506 37716 26236
rect 37772 26226 37828 26236
rect 38164 26226 38220 26236
rect 37660 25454 37662 25506
rect 37714 25454 37716 25506
rect 37548 25284 37604 25294
rect 37548 24722 37604 25228
rect 37548 24670 37550 24722
rect 37602 24670 37604 24722
rect 37548 24658 37604 24670
rect 37660 24724 37716 25454
rect 37660 24658 37716 24668
rect 37772 26068 37828 26078
rect 38556 26068 38612 26078
rect 37436 23762 37492 23772
rect 37772 23492 37828 26012
rect 38444 26066 38612 26068
rect 38444 26014 38558 26066
rect 38610 26014 38612 26066
rect 38444 26012 38612 26014
rect 38444 25618 38500 26012
rect 38556 26002 38612 26012
rect 38444 25566 38446 25618
rect 38498 25566 38500 25618
rect 38444 25554 38500 25566
rect 38668 24948 38724 26796
rect 39116 26628 39172 27022
rect 38780 26572 39172 26628
rect 39228 26740 39284 27132
rect 39340 27074 39396 27244
rect 39340 27022 39342 27074
rect 39394 27022 39396 27074
rect 39340 27010 39396 27022
rect 39564 27074 39620 27086
rect 39564 27022 39566 27074
rect 39618 27022 39620 27074
rect 39564 26852 39620 27022
rect 39564 26786 39620 26796
rect 39844 26962 39900 26974
rect 39844 26910 39846 26962
rect 39898 26910 39900 26962
rect 38780 26292 38836 26572
rect 38780 26226 38836 26236
rect 38892 26404 38948 26414
rect 38892 26290 38948 26348
rect 38892 26238 38894 26290
rect 38946 26238 38948 26290
rect 38892 26226 38948 26238
rect 39116 26292 39172 26302
rect 39116 26198 39172 26236
rect 39228 26290 39284 26684
rect 39844 26404 39900 26910
rect 40124 26908 40180 27356
rect 40236 27300 40292 27580
rect 41020 27524 41076 27804
rect 41132 27858 41188 27870
rect 41132 27806 41134 27858
rect 41186 27806 41188 27858
rect 41132 27748 41188 27806
rect 41132 27682 41188 27692
rect 41020 27468 41188 27524
rect 40236 27244 40516 27300
rect 40348 27076 40404 27086
rect 40348 26994 40350 27020
rect 40402 26994 40404 27020
rect 40348 26982 40404 26994
rect 40124 26852 40292 26908
rect 40068 26740 40124 26750
rect 40068 26514 40124 26684
rect 40068 26462 40070 26514
rect 40122 26462 40124 26514
rect 40068 26450 40124 26462
rect 39844 26338 39900 26348
rect 39228 26238 39230 26290
rect 39282 26238 39284 26290
rect 39228 26226 39284 26238
rect 39508 26180 39564 26190
rect 39508 26086 39564 26124
rect 39564 25956 39620 25966
rect 38668 24882 38724 24892
rect 38780 25284 38836 25294
rect 38332 24724 38388 24734
rect 38220 24164 38276 24174
rect 38220 24070 38276 24108
rect 37884 23938 37940 23950
rect 37884 23886 37886 23938
rect 37938 23886 37940 23938
rect 37884 23716 37940 23886
rect 37940 23660 38052 23716
rect 37884 23650 37940 23660
rect 37324 23436 37492 23492
rect 37100 23324 37380 23380
rect 36260 22482 36932 22484
rect 36260 22430 36262 22482
rect 36314 22430 36932 22482
rect 36260 22428 36932 22430
rect 36260 22418 36316 22428
rect 37324 22370 37380 23324
rect 37324 22318 37326 22370
rect 37378 22318 37380 22370
rect 37324 22306 37380 22318
rect 37436 22372 37492 23436
rect 37660 23042 37716 23054
rect 37660 22990 37662 23042
rect 37714 22990 37716 23042
rect 37660 22372 37716 22990
rect 37436 22370 37716 22372
rect 37436 22318 37438 22370
rect 37490 22318 37716 22370
rect 37436 22316 37716 22318
rect 37044 22258 37100 22270
rect 37044 22206 37046 22258
rect 37098 22206 37100 22258
rect 35980 22082 36036 22092
rect 36876 22148 36932 22158
rect 37044 22148 37100 22206
rect 36932 22092 37100 22148
rect 36092 21812 36148 21822
rect 36092 21698 36148 21756
rect 36092 21646 36094 21698
rect 36146 21646 36148 21698
rect 36092 21634 36148 21646
rect 36540 21812 36596 21822
rect 36540 21586 36596 21756
rect 36540 21534 36542 21586
rect 36594 21534 36596 21586
rect 36540 21522 36596 21534
rect 36876 21586 36932 22092
rect 37436 21700 37492 22316
rect 37436 21634 37492 21644
rect 36876 21534 36878 21586
rect 36930 21534 36932 21586
rect 36876 21522 36932 21534
rect 37212 21586 37268 21598
rect 37212 21534 37214 21586
rect 37266 21534 37268 21586
rect 37212 21476 37268 21534
rect 36652 21418 36708 21430
rect 36652 21366 36654 21418
rect 36706 21366 36708 21418
rect 36652 21028 36708 21366
rect 37100 21420 37212 21476
rect 34412 21026 34580 21028
rect 34412 20974 34526 21026
rect 34578 20974 34580 21026
rect 34412 20972 34580 20974
rect 34524 20962 34580 20972
rect 35420 20972 35588 21028
rect 35644 20972 36708 21028
rect 36764 21252 36820 21262
rect 34860 20804 34916 20814
rect 35140 20804 35196 20814
rect 34860 20802 35196 20804
rect 34860 20750 34862 20802
rect 34914 20750 35142 20802
rect 35194 20750 35196 20802
rect 34860 20748 35196 20750
rect 34860 20738 34916 20748
rect 35140 20738 35196 20748
rect 35420 20802 35476 20972
rect 35644 20804 35700 20972
rect 36316 20804 36372 20814
rect 35420 20750 35422 20802
rect 35474 20750 35476 20802
rect 35420 20738 35476 20750
rect 35532 20802 35700 20804
rect 35532 20750 35646 20802
rect 35698 20750 35700 20802
rect 35532 20748 35700 20750
rect 34132 20580 34188 20590
rect 35532 20580 35588 20748
rect 35644 20738 35700 20748
rect 36092 20802 36372 20804
rect 36092 20750 36318 20802
rect 36370 20750 36372 20802
rect 36092 20748 36372 20750
rect 35980 20580 36036 20590
rect 34132 20486 34188 20524
rect 35288 20524 35588 20580
rect 35756 20578 36036 20580
rect 35756 20526 35982 20578
rect 36034 20526 36036 20578
rect 35756 20524 36036 20526
rect 33404 20018 33460 20030
rect 33404 19966 33406 20018
rect 33458 19966 33460 20018
rect 33740 20022 33742 20074
rect 33794 20022 33796 20074
rect 35084 20468 35140 20478
rect 33740 20010 33796 20022
rect 34412 20020 34468 20030
rect 33852 20018 34468 20020
rect 33404 18450 33460 19966
rect 33852 19966 34414 20018
rect 34466 19966 34468 20018
rect 33852 19964 34468 19966
rect 33852 19348 33908 19964
rect 34412 19954 34468 19964
rect 35084 19572 35140 20412
rect 35288 20074 35344 20524
rect 35288 20022 35290 20074
rect 35342 20022 35344 20074
rect 35288 20010 35344 20022
rect 35532 20020 35588 20030
rect 35532 19926 35588 19964
rect 33404 18398 33406 18450
rect 33458 18398 33460 18450
rect 33740 19346 33908 19348
rect 33740 19294 33854 19346
rect 33906 19294 33908 19346
rect 33740 19292 33908 19294
rect 33740 18506 33796 19292
rect 33852 19282 33908 19292
rect 34524 19516 35140 19572
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 33740 18454 33742 18506
rect 33794 18454 33796 18506
rect 34524 18462 34580 19516
rect 35756 19346 35812 20524
rect 35980 20514 36036 20524
rect 36092 20142 36148 20748
rect 36316 20738 36372 20748
rect 36036 20130 36148 20142
rect 36036 20078 36038 20130
rect 36090 20078 36148 20130
rect 36036 20076 36148 20078
rect 36540 20580 36596 20590
rect 36764 20580 36820 21196
rect 37100 20914 37156 21420
rect 37212 21410 37268 21420
rect 37100 20862 37102 20914
rect 37154 20862 37156 20914
rect 37100 20850 37156 20862
rect 37324 21364 37380 21374
rect 36596 20524 36820 20580
rect 36036 20066 36092 20076
rect 36316 20020 36372 20030
rect 36316 19926 36372 19964
rect 36540 20018 36596 20524
rect 36876 20132 36932 20142
rect 36876 20038 36932 20076
rect 36540 19966 36542 20018
rect 36594 19966 36596 20018
rect 36540 19954 36596 19966
rect 37212 20020 37268 20030
rect 37212 19926 37268 19964
rect 35756 19294 35758 19346
rect 35810 19294 35812 19346
rect 35756 19282 35812 19294
rect 36540 19236 36596 19246
rect 36316 19234 36596 19236
rect 36316 19182 36542 19234
rect 36594 19182 36596 19234
rect 36316 19180 36596 19182
rect 33740 18442 33796 18454
rect 34468 18450 34580 18462
rect 35196 18452 35252 18462
rect 33404 18228 33460 18398
rect 34468 18398 34470 18450
rect 34522 18398 34580 18450
rect 34468 18386 34580 18398
rect 33404 18162 33460 18172
rect 33292 17938 33348 17948
rect 32172 17892 32228 17902
rect 32172 17666 32228 17836
rect 32172 17614 32174 17666
rect 32226 17614 32228 17666
rect 32172 17602 32228 17614
rect 32620 17892 32676 17902
rect 31164 17266 31220 17276
rect 31052 17154 31108 17164
rect 32620 16882 32676 17836
rect 32956 17668 33012 17678
rect 32956 17666 33236 17668
rect 32956 17614 32958 17666
rect 33010 17614 33236 17666
rect 32956 17612 33236 17614
rect 32956 17602 33012 17612
rect 33180 16994 33236 17612
rect 34412 17444 34468 17454
rect 33180 16942 33182 16994
rect 33234 16942 33236 16994
rect 33180 16930 33236 16942
rect 33628 17220 33684 17230
rect 33628 16938 33684 17164
rect 34244 17050 34300 17062
rect 34244 16998 34246 17050
rect 34298 16998 34300 17050
rect 34244 16996 34300 16998
rect 32620 16830 32622 16882
rect 32674 16830 32676 16882
rect 31836 16772 31892 16782
rect 31836 16678 31892 16716
rect 32508 16324 32564 16334
rect 32620 16324 32676 16830
rect 33012 16884 33068 16894
rect 33012 16790 33068 16828
rect 33628 16886 33630 16938
rect 33682 16886 33684 16938
rect 33628 16884 33684 16886
rect 33852 16940 34300 16996
rect 33852 16938 33908 16940
rect 33852 16886 33854 16938
rect 33906 16886 33908 16938
rect 33852 16874 33908 16886
rect 34412 16882 34468 17388
rect 33628 16808 33684 16828
rect 34412 16830 34414 16882
rect 34466 16830 34468 16882
rect 34412 16818 34468 16830
rect 33740 16772 33796 16782
rect 32508 16322 33012 16324
rect 32508 16270 32510 16322
rect 32562 16270 33012 16322
rect 32508 16268 33012 16270
rect 32508 16258 32564 16268
rect 30604 16146 30660 16156
rect 30940 16212 30996 16222
rect 30212 16100 30268 16110
rect 30212 16006 30268 16044
rect 30044 15698 30100 15708
rect 29932 15250 29988 15260
rect 30044 15428 30100 15438
rect 28812 14914 28868 14924
rect 28532 14702 28534 14754
rect 28586 14702 28588 14754
rect 28532 14690 28588 14702
rect 28364 14644 28420 14654
rect 27804 14532 27860 14542
rect 28252 14530 28308 14542
rect 27804 14438 27860 14476
rect 27972 14474 28028 14486
rect 27972 14422 27974 14474
rect 28026 14422 28028 14474
rect 28252 14478 28254 14530
rect 28306 14478 28308 14530
rect 27972 13860 28028 14422
rect 28140 14420 28196 14430
rect 28140 14196 28196 14364
rect 28140 14130 28196 14140
rect 27076 13188 27132 13198
rect 27076 13094 27132 13132
rect 27356 13020 27412 13356
rect 27692 13346 27748 13356
rect 27804 13804 28028 13860
rect 28252 14084 28308 14478
rect 27804 13188 27860 13804
rect 28252 13636 28308 14028
rect 28252 13570 28308 13580
rect 27804 13122 27860 13132
rect 28364 13524 28420 14588
rect 28868 14308 28924 14318
rect 28868 13970 28924 14252
rect 28868 13918 28870 13970
rect 28922 13918 28924 13970
rect 28868 13906 28924 13918
rect 27356 12964 27524 13020
rect 26908 12910 26910 12962
rect 26962 12910 26964 12962
rect 26460 12236 26628 12292
rect 26348 12180 26404 12190
rect 26348 12178 26516 12180
rect 26348 12126 26350 12178
rect 26402 12126 26516 12178
rect 26348 12124 26516 12126
rect 26348 12114 26404 12124
rect 26236 10948 26292 11340
rect 26068 10892 26292 10948
rect 26348 11508 26404 11518
rect 26348 10948 26404 11452
rect 26460 11394 26516 12124
rect 26460 11342 26462 11394
rect 26514 11342 26516 11394
rect 26460 11172 26516 11342
rect 26572 11396 26628 12236
rect 26684 11954 26740 11966
rect 26684 11902 26686 11954
rect 26738 11902 26740 11954
rect 26684 11620 26740 11902
rect 26908 11788 26964 12910
rect 27300 12068 27356 12078
rect 27300 12066 27412 12068
rect 27300 12014 27302 12066
rect 27354 12014 27412 12066
rect 27300 12002 27412 12014
rect 26908 11732 27076 11788
rect 27020 11620 27076 11732
rect 26684 11554 26740 11564
rect 26908 11562 26964 11574
rect 26908 11510 26910 11562
rect 26962 11510 26964 11562
rect 27020 11554 27076 11564
rect 26572 11330 26628 11340
rect 26684 11394 26740 11406
rect 26684 11342 26686 11394
rect 26738 11342 26740 11394
rect 26460 11106 26516 11116
rect 26348 10892 26572 10948
rect 26068 10834 26124 10892
rect 26068 10782 26070 10834
rect 26122 10782 26124 10834
rect 26068 10770 26124 10782
rect 26236 10612 26292 10892
rect 26516 10666 26572 10892
rect 26348 10612 26404 10622
rect 26236 10610 26404 10612
rect 26236 10558 26350 10610
rect 26402 10558 26404 10610
rect 26236 10556 26404 10558
rect 26348 10546 26404 10556
rect 26516 10614 26518 10666
rect 26570 10614 26572 10666
rect 26684 10836 26740 11342
rect 26684 10722 26740 10780
rect 26684 10670 26686 10722
rect 26738 10670 26740 10722
rect 26684 10658 26740 10670
rect 26796 11396 26852 11406
rect 26516 10612 26572 10614
rect 26516 10536 26572 10556
rect 26796 10610 26852 11340
rect 26796 10558 26798 10610
rect 26850 10558 26852 10610
rect 26796 10546 26852 10558
rect 26908 9828 26964 11510
rect 27020 11396 27076 11406
rect 27020 11302 27076 11340
rect 27356 11060 27412 12002
rect 27356 10994 27412 11004
rect 27076 10388 27132 10398
rect 27076 10294 27132 10332
rect 27468 10052 27524 12964
rect 27636 12740 27692 12750
rect 27580 12738 27692 12740
rect 27580 12686 27638 12738
rect 27690 12686 27692 12738
rect 27580 12674 27692 12686
rect 27580 11508 27636 12674
rect 28364 12292 28420 13468
rect 28364 12226 28420 12236
rect 28700 13412 28756 13422
rect 27692 12180 27748 12190
rect 28476 12180 28532 12190
rect 27692 12178 27860 12180
rect 27692 12126 27694 12178
rect 27746 12126 27860 12178
rect 27692 12124 27860 12126
rect 27692 12114 27748 12124
rect 27580 11442 27636 11452
rect 27636 11170 27692 11182
rect 27636 11118 27638 11170
rect 27690 11118 27692 11170
rect 27636 11060 27692 11118
rect 27636 10994 27692 11004
rect 27636 10612 27692 10622
rect 27636 10518 27692 10556
rect 27804 10612 27860 12124
rect 28476 12086 28532 12124
rect 28700 11844 28756 13356
rect 29036 12740 29092 15036
rect 29820 15026 29876 15036
rect 29316 14980 29372 14990
rect 29316 14586 29372 14924
rect 29148 14532 29204 14542
rect 29316 14534 29318 14586
rect 29370 14534 29372 14586
rect 29316 14522 29372 14534
rect 29596 14530 29652 14542
rect 29148 14438 29204 14476
rect 29596 14478 29598 14530
rect 29650 14478 29652 14530
rect 29316 14420 29372 14430
rect 29316 13970 29372 14364
rect 29484 14418 29540 14430
rect 29484 14366 29486 14418
rect 29538 14366 29540 14418
rect 29484 14196 29540 14366
rect 29484 14130 29540 14140
rect 29596 14084 29652 14478
rect 29876 14420 29932 14430
rect 29876 14326 29932 14364
rect 29596 14018 29652 14028
rect 29316 13918 29318 13970
rect 29370 13918 29372 13970
rect 29316 13748 29372 13918
rect 29484 13748 29540 13758
rect 29316 13746 29540 13748
rect 29316 13694 29486 13746
rect 29538 13694 29540 13746
rect 29316 13692 29540 13694
rect 29484 13682 29540 13692
rect 29820 13522 29876 13534
rect 29820 13470 29822 13522
rect 29874 13470 29876 13522
rect 29820 13412 29876 13470
rect 29820 13346 29876 13356
rect 30044 13188 30100 15372
rect 30380 15341 30436 15353
rect 30380 15289 30382 15341
rect 30434 15289 30436 15341
rect 30156 14530 30212 14542
rect 30156 14478 30158 14530
rect 30210 14478 30212 14530
rect 30156 13972 30212 14478
rect 30380 14532 30436 15289
rect 30380 14466 30436 14476
rect 30492 15092 30548 15102
rect 30492 14754 30548 15036
rect 30492 14702 30494 14754
rect 30546 14702 30548 14754
rect 30492 14308 30548 14702
rect 30156 13906 30212 13916
rect 30268 14252 30548 14308
rect 30940 14502 30996 16156
rect 31164 16212 31220 16222
rect 31164 16070 31220 16156
rect 31164 16018 31166 16070
rect 31218 16018 31220 16070
rect 31164 16006 31220 16018
rect 30940 14450 30942 14502
rect 30994 14450 30996 14502
rect 30940 14308 30996 14450
rect 30268 13748 30324 14252
rect 30940 14242 30996 14252
rect 31836 15316 31892 15326
rect 30604 14196 30660 14206
rect 30268 13654 30324 13692
rect 30436 13972 30492 13982
rect 30436 13802 30492 13916
rect 30436 13750 30438 13802
rect 30490 13750 30492 13802
rect 30604 13858 30660 14140
rect 30604 13806 30606 13858
rect 30658 13806 30660 13858
rect 30604 13794 30660 13806
rect 30716 14084 30772 14094
rect 30436 13524 30492 13750
rect 30716 13746 30772 14028
rect 30716 13694 30718 13746
rect 30770 13694 30772 13746
rect 30716 13682 30772 13694
rect 31276 13972 31332 13982
rect 31164 13636 31220 13646
rect 30436 13458 30492 13468
rect 30996 13524 31052 13534
rect 30996 13430 31052 13468
rect 29484 13132 30100 13188
rect 30156 13412 30212 13422
rect 29484 12964 29540 13132
rect 29428 12908 29540 12964
rect 29596 12962 29652 12974
rect 29596 12910 29598 12962
rect 29650 12910 29652 12962
rect 29428 12906 29484 12908
rect 29428 12854 29430 12906
rect 29482 12854 29484 12906
rect 29428 12842 29484 12854
rect 29596 12852 29652 12910
rect 29596 12786 29652 12796
rect 29036 12674 29092 12684
rect 28700 11788 28980 11844
rect 28028 11172 28084 11182
rect 28028 10612 28084 11116
rect 28644 11170 28700 11182
rect 28644 11118 28646 11170
rect 28698 11118 28700 11170
rect 27804 10610 28084 10612
rect 27804 10558 28030 10610
rect 28082 10558 28084 10610
rect 27804 10556 28084 10558
rect 26908 9762 26964 9772
rect 27132 9996 27524 10052
rect 27580 10388 27636 10398
rect 26516 9716 26572 9726
rect 25788 9042 25956 9044
rect 25788 8990 25790 9042
rect 25842 8990 25956 9042
rect 25788 8988 25956 8990
rect 26012 9604 26068 9614
rect 26012 9042 26068 9548
rect 26516 9602 26572 9660
rect 26516 9550 26518 9602
rect 26570 9550 26572 9602
rect 26516 9380 26572 9550
rect 26964 9602 27020 9614
rect 26964 9550 26966 9602
rect 27018 9550 27020 9602
rect 26964 9492 27020 9550
rect 26964 9426 27020 9436
rect 26012 8990 26014 9042
rect 26066 8990 26068 9042
rect 25788 8978 25844 8988
rect 25676 8874 25732 8886
rect 25676 8822 25678 8874
rect 25730 8822 25732 8874
rect 25676 8708 25732 8822
rect 26012 8820 26068 8990
rect 25676 8642 25732 8652
rect 25788 8764 26012 8820
rect 25788 8258 25844 8764
rect 26012 8726 26068 8764
rect 26348 9324 26572 9380
rect 25564 8202 25676 8214
rect 25564 8150 25622 8202
rect 25674 8150 25676 8202
rect 25788 8206 25790 8258
rect 25842 8206 25844 8258
rect 25788 8194 25844 8206
rect 25900 8260 25956 8270
rect 25900 8166 25956 8204
rect 25564 8148 25676 8150
rect 26180 8148 26236 8158
rect 25564 8092 25732 8148
rect 25340 7980 25542 8036
rect 25340 7812 25396 7822
rect 25228 7474 25284 7486
rect 25228 7422 25230 7474
rect 25282 7422 25284 7474
rect 25228 7140 25284 7422
rect 25340 7474 25396 7756
rect 25340 7422 25342 7474
rect 25394 7422 25396 7474
rect 25486 7512 25542 7980
rect 25486 7460 25488 7512
rect 25540 7460 25542 7512
rect 25486 7448 25542 7460
rect 25340 7410 25396 7422
rect 23324 6610 23326 6636
rect 23378 6610 23380 6636
rect 23324 6598 23380 6610
rect 23548 6692 23604 6702
rect 23940 6694 23942 6746
rect 23994 6694 23996 6746
rect 23940 6682 23996 6694
rect 24108 6860 24388 6916
rect 24780 7084 25284 7140
rect 25676 7140 25732 8092
rect 26180 8054 26236 8092
rect 26348 7924 26404 9324
rect 26460 9042 26516 9054
rect 26460 8990 26462 9042
rect 26514 8990 26516 9042
rect 26460 8484 26516 8990
rect 26628 9044 26684 9054
rect 26628 8950 26684 8988
rect 26796 9042 26852 9054
rect 26796 8990 26798 9042
rect 26850 8990 26852 9042
rect 26796 8820 26852 8990
rect 26908 9044 26964 9054
rect 27132 9044 27188 9996
rect 27580 9940 27636 10332
rect 27524 9884 27636 9940
rect 27244 9826 27300 9838
rect 27244 9774 27246 9826
rect 27298 9774 27300 9826
rect 27244 9380 27300 9774
rect 27244 9314 27300 9324
rect 27356 9828 27412 9838
rect 27524 9782 27580 9884
rect 26908 9042 27188 9044
rect 26908 8990 26910 9042
rect 26962 8990 27188 9042
rect 26908 8988 27188 8990
rect 26908 8978 26964 8988
rect 26796 8484 26852 8764
rect 26516 8428 26628 8484
rect 26796 8428 26964 8484
rect 26460 8418 26516 8428
rect 26572 8258 26628 8428
rect 26684 8372 26740 8382
rect 26740 8316 26796 8372
rect 26684 8314 26796 8316
rect 26684 8306 26742 8314
rect 26572 8206 26574 8258
rect 26626 8206 26628 8258
rect 26740 8262 26742 8306
rect 26794 8262 26796 8314
rect 26740 8250 26796 8262
rect 26908 8258 26964 8428
rect 26572 8194 26628 8206
rect 26908 8206 26910 8258
rect 26962 8206 26964 8258
rect 26908 8194 26964 8206
rect 27020 8260 27076 8988
rect 27188 8820 27244 8830
rect 27020 8166 27076 8204
rect 27132 8818 27244 8820
rect 27132 8766 27190 8818
rect 27242 8766 27244 8818
rect 27132 8754 27244 8766
rect 26124 7868 26404 7924
rect 26460 8148 26516 8158
rect 25900 7476 25956 7486
rect 25900 7362 25956 7420
rect 25900 7310 25902 7362
rect 25954 7310 25956 7362
rect 25900 7298 25956 7310
rect 23548 6598 23604 6636
rect 23772 6578 23828 6590
rect 23772 6526 23774 6578
rect 23826 6526 23828 6578
rect 22820 6468 22876 6478
rect 22764 6466 22876 6468
rect 22764 6414 22822 6466
rect 22874 6414 22876 6466
rect 22764 6402 22876 6414
rect 22652 5908 22708 5918
rect 22652 5814 22708 5852
rect 22652 4340 22708 4350
rect 22652 4246 22708 4284
rect 22764 4116 22820 6402
rect 23772 5908 23828 6526
rect 23772 5842 23828 5852
rect 22876 5460 22932 5470
rect 22876 5122 22932 5404
rect 23212 5290 23268 5302
rect 23212 5238 23214 5290
rect 23266 5238 23268 5290
rect 22876 5070 22878 5122
rect 22930 5070 22932 5122
rect 22876 5058 22932 5070
rect 23100 5124 23156 5134
rect 23100 5030 23156 5068
rect 23212 5012 23268 5238
rect 23436 5236 23492 5246
rect 23436 5124 23492 5180
rect 23212 4946 23268 4956
rect 23324 5122 23492 5124
rect 23324 5070 23438 5122
rect 23490 5070 23492 5122
rect 23324 5068 23492 5070
rect 23156 4452 23212 4462
rect 23156 4358 23212 4396
rect 22764 4050 22820 4060
rect 22876 4338 22932 4350
rect 22876 4286 22878 4338
rect 22930 4286 22932 4338
rect 22876 4004 22932 4286
rect 22876 3938 22932 3948
rect 23324 3678 23380 5068
rect 23436 5058 23492 5068
rect 23996 4900 24052 4910
rect 23436 4338 23492 4350
rect 23436 4286 23438 4338
rect 23490 4286 23492 4338
rect 23436 3892 23492 4286
rect 23772 4114 23828 4126
rect 23772 4062 23774 4114
rect 23826 4062 23828 4114
rect 23772 4004 23828 4062
rect 23772 3938 23828 3948
rect 23436 3826 23492 3836
rect 23996 3892 24052 4844
rect 22540 3602 22596 3612
rect 22764 3668 22820 3678
rect 21980 3469 21982 3521
rect 22034 3469 22036 3521
rect 22764 3554 22820 3612
rect 23268 3666 23380 3678
rect 23268 3614 23270 3666
rect 23322 3614 23380 3666
rect 23268 3612 23380 3614
rect 23268 3602 23324 3612
rect 22764 3502 22766 3554
rect 22818 3502 22820 3554
rect 22764 3490 22820 3502
rect 21980 3457 22036 3469
rect 23996 3454 24052 3836
rect 24108 3668 24164 6860
rect 24276 6692 24332 6702
rect 24276 6522 24332 6636
rect 24276 6470 24278 6522
rect 24330 6470 24332 6522
rect 24276 6458 24332 6470
rect 24444 6690 24500 6702
rect 24444 6638 24446 6690
rect 24498 6638 24500 6690
rect 24444 6020 24500 6638
rect 24780 6690 24836 7084
rect 25676 7074 25732 7084
rect 25452 6916 25508 6926
rect 24780 6638 24782 6690
rect 24834 6638 24836 6690
rect 24780 6626 24836 6638
rect 24892 6690 24948 6702
rect 24892 6638 24894 6690
rect 24946 6638 24948 6690
rect 24892 6580 24948 6638
rect 24892 6356 24948 6524
rect 25060 6634 25116 6646
rect 25060 6582 25062 6634
rect 25114 6582 25116 6634
rect 25060 6580 25116 6582
rect 25060 6514 25116 6524
rect 24892 6300 25396 6356
rect 25116 6132 25172 6142
rect 24556 6020 24612 6030
rect 24444 6018 24612 6020
rect 24444 5966 24558 6018
rect 24610 5966 24612 6018
rect 24444 5964 24612 5966
rect 24556 5908 24612 5964
rect 24556 5842 24612 5852
rect 24444 5684 24500 5694
rect 24220 5122 24276 5134
rect 24220 5070 24222 5122
rect 24274 5070 24276 5122
rect 24220 4452 24276 5070
rect 24220 4386 24276 4396
rect 24444 5124 24500 5628
rect 25116 5460 25172 6076
rect 25228 5908 25284 5918
rect 25228 5814 25284 5852
rect 25340 5906 25396 6300
rect 25452 6132 25508 6860
rect 25900 6802 25956 6814
rect 25900 6750 25902 6802
rect 25954 6750 25956 6802
rect 25900 6468 25956 6750
rect 26012 6646 26068 6658
rect 26012 6594 26014 6646
rect 26066 6594 26068 6646
rect 26012 6580 26068 6594
rect 26012 6514 26068 6524
rect 25900 6402 25956 6412
rect 26124 6356 26180 7868
rect 25452 6066 25508 6076
rect 26012 6300 26180 6356
rect 26236 6690 26292 6702
rect 26236 6638 26238 6690
rect 26290 6638 26292 6690
rect 25340 5854 25342 5906
rect 25394 5854 25396 5906
rect 25340 5842 25396 5854
rect 25526 5943 25582 5955
rect 25526 5908 25528 5943
rect 25580 5908 25582 5943
rect 25526 5842 25582 5852
rect 25900 5684 25956 5694
rect 25900 5590 25956 5628
rect 25172 5404 25396 5460
rect 25116 5394 25172 5404
rect 24332 4340 24388 4350
rect 24444 4340 24500 5068
rect 25340 4900 25396 5404
rect 26012 5348 26068 6300
rect 26236 6244 26292 6638
rect 24780 4844 25396 4900
rect 25900 5292 26068 5348
rect 26124 6188 26292 6244
rect 26348 6468 26404 6478
rect 26124 5908 26180 6188
rect 25900 4900 25956 5292
rect 24556 4340 24612 4350
rect 24444 4338 24612 4340
rect 24444 4286 24558 4338
rect 24610 4286 24612 4338
rect 24444 4284 24612 4286
rect 24332 4238 24388 4284
rect 24556 4274 24612 4284
rect 24780 4338 24836 4844
rect 25900 4834 25956 4844
rect 26012 5012 26068 5022
rect 25228 4452 25284 4462
rect 25228 4358 25284 4396
rect 26012 4394 26068 4956
rect 25408 4371 25464 4383
rect 24780 4286 24782 4338
rect 24834 4286 24836 4338
rect 24780 4274 24836 4286
rect 25408 4319 25410 4371
rect 25462 4319 25464 4371
rect 24276 4226 24388 4238
rect 24276 4174 24278 4226
rect 24330 4174 24388 4226
rect 24276 4172 24388 4174
rect 24276 4162 24332 4172
rect 25408 4116 25464 4319
rect 25564 4374 25620 4386
rect 25564 4340 25566 4374
rect 25618 4340 25620 4374
rect 26012 4342 26014 4394
rect 26066 4342 26068 4394
rect 26012 4330 26068 4342
rect 26124 5010 26180 5852
rect 26124 4958 26126 5010
rect 26178 4958 26180 5010
rect 25564 4274 25620 4284
rect 25408 4060 25956 4116
rect 25452 3892 25508 3902
rect 24108 3602 24164 3612
rect 24836 3668 24892 3678
rect 24836 3574 24892 3612
rect 25172 3556 25228 3566
rect 25172 3462 25228 3500
rect 25452 3554 25508 3836
rect 25900 3722 25956 4060
rect 25900 3670 25902 3722
rect 25954 3670 25956 3722
rect 25900 3658 25956 3670
rect 25452 3502 25454 3554
rect 25506 3502 25508 3554
rect 25452 3490 25508 3502
rect 25676 3556 25732 3566
rect 26012 3556 26068 3566
rect 25676 3554 25956 3556
rect 25676 3502 25678 3554
rect 25730 3502 25956 3554
rect 25676 3500 25956 3502
rect 25676 3490 25732 3500
rect 21084 3444 21140 3446
rect 23996 3442 24108 3454
rect 23996 3390 24054 3442
rect 24106 3390 24108 3442
rect 23996 3388 24108 3390
rect 21084 3378 21140 3388
rect 24052 3378 24108 3388
rect 19460 3330 19516 3332
rect 19460 3278 19462 3330
rect 19514 3278 19516 3330
rect 19460 3266 19516 3278
rect 25900 3332 25956 3500
rect 26012 3462 26068 3500
rect 26124 3332 26180 4958
rect 26236 4788 26292 4798
rect 26236 3668 26292 4732
rect 26348 4394 26404 6412
rect 26460 6132 26516 8092
rect 26740 8036 26796 8046
rect 26740 7698 26796 7980
rect 26740 7646 26742 7698
rect 26794 7646 26796 7698
rect 26740 7634 26796 7646
rect 26908 7588 26964 7598
rect 26908 7474 26964 7532
rect 26908 7422 26910 7474
rect 26962 7422 26964 7474
rect 26908 7410 26964 7422
rect 27132 7364 27188 8754
rect 27356 8484 27412 9772
rect 27522 9770 27580 9782
rect 27522 9718 27524 9770
rect 27576 9718 27580 9770
rect 27522 9716 27580 9718
rect 27522 9706 27578 9716
rect 27804 9044 27860 10556
rect 28028 10546 28084 10556
rect 28364 11060 28420 11070
rect 27916 9940 27972 9950
rect 27916 9938 28196 9940
rect 27916 9886 27918 9938
rect 27970 9886 28196 9938
rect 27916 9884 28196 9886
rect 27916 9874 27972 9884
rect 27692 9042 27860 9044
rect 27692 8990 27806 9042
rect 27858 8990 27860 9042
rect 27692 8988 27860 8990
rect 27580 8484 27636 8494
rect 27356 8482 27636 8484
rect 27356 8430 27582 8482
rect 27634 8430 27636 8482
rect 27356 8428 27636 8430
rect 27580 8418 27636 8428
rect 27300 8146 27356 8158
rect 27300 8094 27302 8146
rect 27354 8094 27356 8146
rect 27300 7588 27356 8094
rect 27020 7308 27188 7364
rect 27244 7532 27356 7588
rect 27692 7588 27748 8988
rect 27804 8978 27860 8988
rect 26852 6468 26908 6478
rect 26852 6374 26908 6412
rect 26460 6076 26740 6132
rect 26348 4342 26350 4394
rect 26402 4342 26404 4394
rect 26348 4116 26404 4342
rect 26460 5906 26516 5918
rect 26460 5854 26462 5906
rect 26514 5854 26516 5906
rect 26460 5124 26516 5854
rect 26460 4340 26516 5068
rect 26684 5012 26740 6076
rect 27020 5908 27076 7308
rect 27244 7252 27300 7532
rect 27692 7522 27748 7532
rect 27804 8482 27860 8494
rect 27804 8430 27806 8482
rect 27858 8430 27860 8482
rect 27692 7364 27748 7374
rect 27188 7196 27300 7252
rect 27356 7362 27748 7364
rect 27356 7310 27694 7362
rect 27746 7310 27748 7362
rect 27356 7308 27748 7310
rect 27188 6746 27244 7196
rect 27188 6694 27190 6746
rect 27242 6694 27244 6746
rect 27356 6802 27412 7308
rect 27692 7298 27748 7308
rect 27356 6750 27358 6802
rect 27410 6750 27412 6802
rect 27356 6738 27412 6750
rect 27188 6682 27244 6694
rect 27580 6692 27636 6702
rect 27580 6598 27636 6636
rect 27804 6662 27860 8430
rect 28140 8258 28196 9884
rect 28140 8206 28142 8258
rect 28194 8206 28196 8258
rect 28140 8194 28196 8206
rect 28252 9604 28308 9614
rect 27972 8036 28028 8046
rect 27972 7942 28028 7980
rect 28252 7700 28308 9548
rect 28364 8708 28420 11004
rect 28644 9602 28700 11118
rect 28812 10498 28868 10510
rect 28812 10446 28814 10498
rect 28866 10446 28868 10498
rect 28812 9940 28868 10446
rect 28924 9940 28980 11788
rect 29708 11396 29764 13132
rect 29988 12906 30044 12918
rect 29820 12850 29876 12862
rect 29820 12798 29822 12850
rect 29874 12798 29876 12850
rect 29820 12180 29876 12798
rect 29988 12854 29990 12906
rect 30042 12854 30044 12906
rect 29988 12404 30044 12854
rect 29988 12338 30044 12348
rect 29820 12114 29876 12124
rect 30156 12180 30212 13356
rect 30268 13188 30324 13198
rect 30268 12628 30324 13132
rect 30548 13076 30604 13086
rect 30548 13018 30604 13020
rect 30548 12966 30550 13018
rect 30602 12966 30604 13018
rect 30548 12954 30604 12966
rect 30940 12962 30996 12974
rect 30940 12910 30942 12962
rect 30994 12910 30996 12962
rect 30716 12852 30772 12862
rect 30716 12758 30772 12796
rect 30268 12562 30324 12572
rect 30940 12628 30996 12910
rect 31164 12934 31220 13580
rect 31164 12882 31166 12934
rect 31218 12882 31220 12934
rect 31164 12870 31220 12882
rect 30940 12562 30996 12572
rect 30828 12180 30884 12190
rect 30156 12114 30212 12124
rect 30492 12178 30884 12180
rect 30492 12126 30830 12178
rect 30882 12126 30884 12178
rect 30492 12124 30884 12126
rect 30380 12068 30436 12078
rect 30380 11974 30436 12012
rect 30492 11630 30548 12124
rect 30828 12114 30884 12124
rect 30940 12178 30996 12190
rect 30940 12126 30942 12178
rect 30994 12126 30996 12178
rect 30436 11618 30548 11630
rect 30436 11566 30438 11618
rect 30490 11566 30548 11618
rect 30436 11564 30548 11566
rect 30604 11956 30660 11966
rect 30436 11554 30492 11564
rect 29708 11340 29988 11396
rect 29652 11172 29708 11182
rect 29652 11078 29708 11116
rect 29932 10612 29988 11340
rect 30604 11373 30660 11900
rect 30604 11321 30606 11373
rect 30658 11321 30660 11373
rect 30604 11309 30660 11321
rect 30716 11394 30772 11406
rect 30716 11342 30718 11394
rect 30770 11342 30772 11394
rect 30100 11284 30156 11294
rect 30100 11190 30156 11228
rect 30268 11172 30324 11182
rect 29932 10556 30212 10612
rect 29988 10388 30044 10398
rect 29820 9940 29876 9950
rect 28924 9884 29204 9940
rect 28812 9874 28868 9884
rect 29148 9882 29204 9884
rect 29148 9830 29150 9882
rect 29202 9830 29204 9882
rect 29820 9846 29876 9884
rect 29988 9882 30044 10332
rect 29148 9818 29204 9830
rect 29988 9830 29990 9882
rect 30042 9830 30044 9882
rect 29988 9818 30044 9830
rect 29428 9770 29484 9782
rect 29428 9718 29430 9770
rect 29482 9718 29484 9770
rect 29428 9716 29484 9718
rect 29428 9660 29540 9716
rect 28644 9550 28646 9602
rect 28698 9550 28700 9602
rect 28644 9156 28700 9550
rect 29484 9604 29540 9660
rect 30156 9604 30212 10556
rect 29484 9548 30212 9604
rect 28644 9100 28868 9156
rect 28588 8932 28644 8942
rect 28364 8642 28420 8652
rect 28476 8930 28644 8932
rect 28476 8878 28590 8930
rect 28642 8878 28644 8930
rect 28476 8876 28644 8878
rect 28476 8370 28532 8876
rect 28588 8866 28644 8876
rect 28476 8318 28478 8370
rect 28530 8318 28532 8370
rect 28476 8306 28532 8318
rect 27804 6610 27806 6662
rect 27858 6610 27860 6662
rect 27804 6468 27860 6610
rect 26908 5852 27076 5908
rect 27468 6412 27860 6468
rect 27916 7644 28308 7700
rect 28812 8036 28868 9100
rect 26908 5796 26964 5852
rect 27244 5796 27300 5806
rect 26852 5740 26964 5796
rect 27020 5794 27300 5796
rect 27020 5742 27246 5794
rect 27298 5742 27300 5794
rect 27020 5740 27300 5742
rect 26852 5178 26908 5740
rect 26852 5126 26854 5178
rect 26906 5126 26908 5178
rect 27020 5234 27076 5740
rect 27244 5730 27300 5740
rect 27020 5182 27022 5234
rect 27074 5182 27076 5234
rect 27020 5170 27076 5182
rect 26852 5114 26908 5126
rect 27468 5094 27524 6412
rect 27916 6132 27972 7644
rect 28812 7476 28868 7980
rect 28812 7410 28868 7420
rect 28924 8708 28980 8718
rect 29708 8708 29764 9548
rect 28588 6690 28644 6702
rect 28588 6638 28590 6690
rect 28642 6638 28644 6690
rect 28420 6468 28476 6478
rect 27916 6066 27972 6076
rect 28364 6466 28476 6468
rect 28364 6414 28422 6466
rect 28474 6414 28476 6466
rect 28364 6402 28476 6414
rect 28364 5572 28420 6402
rect 28588 6244 28644 6638
rect 28588 6178 28644 6188
rect 27692 5516 28420 5572
rect 27692 5178 27748 5516
rect 27692 5126 27694 5178
rect 27746 5126 27748 5178
rect 27692 5114 27748 5126
rect 27916 5348 27972 5358
rect 27916 5122 27972 5292
rect 28812 5348 28868 5358
rect 27468 5042 27470 5094
rect 27522 5042 27524 5094
rect 27916 5070 27918 5122
rect 27970 5070 27972 5122
rect 27916 5058 27972 5070
rect 28252 5122 28308 5134
rect 28252 5070 28254 5122
rect 28306 5070 28308 5122
rect 27468 5012 27524 5042
rect 26684 4956 26908 5012
rect 27468 4956 27748 5012
rect 26852 4900 26908 4956
rect 26852 4844 26964 4900
rect 26796 4340 26852 4350
rect 26460 4338 26852 4340
rect 26460 4286 26798 4338
rect 26850 4286 26852 4338
rect 26460 4284 26852 4286
rect 26796 4274 26852 4284
rect 26908 4228 26964 4844
rect 27580 4228 27636 4238
rect 26908 4172 27020 4228
rect 26348 3780 26404 4060
rect 26348 3714 26404 3724
rect 26236 3554 26292 3612
rect 26236 3502 26238 3554
rect 26290 3502 26292 3554
rect 26964 3610 27020 4172
rect 26964 3558 26966 3610
rect 27018 3558 27020 3610
rect 27132 4226 27636 4228
rect 27132 4174 27582 4226
rect 27634 4174 27636 4226
rect 27132 4172 27636 4174
rect 27132 3666 27188 4172
rect 27580 4162 27636 4172
rect 27132 3614 27134 3666
rect 27186 3614 27188 3666
rect 27132 3602 27188 3614
rect 26964 3546 27020 3558
rect 26236 3490 26292 3502
rect 27692 3516 27748 4956
rect 28252 4900 28308 5070
rect 28252 4834 28308 4844
rect 28812 5124 28868 5292
rect 28700 4452 28756 4462
rect 27692 3464 27694 3516
rect 27746 3464 27748 3516
rect 28588 3556 28644 3566
rect 28700 3556 28756 4396
rect 28588 3554 28756 3556
rect 27692 3452 27748 3464
rect 27804 3498 27860 3510
rect 27804 3446 27806 3498
rect 27858 3446 27860 3498
rect 28588 3502 28590 3554
rect 28642 3502 28756 3554
rect 28588 3500 28756 3502
rect 28812 3554 28868 5068
rect 28812 3502 28814 3554
rect 28866 3502 28868 3554
rect 28588 3490 28644 3500
rect 28812 3490 28868 3502
rect 27804 3388 27860 3446
rect 28420 3388 28476 3398
rect 27804 3386 28476 3388
rect 27804 3334 28422 3386
rect 28474 3334 28476 3386
rect 27804 3332 28476 3334
rect 25900 3276 26180 3332
rect 28420 3322 28476 3332
rect 19796 3266 19852 3276
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 28924 2772 28980 8652
rect 29148 8652 29764 8708
rect 29932 9044 29988 9054
rect 29148 8258 29204 8652
rect 29148 8206 29150 8258
rect 29202 8206 29204 8258
rect 29148 8194 29204 8206
rect 29484 8036 29540 8046
rect 29484 7942 29540 7980
rect 29596 7362 29652 7374
rect 29596 7310 29598 7362
rect 29650 7310 29652 7362
rect 29596 7252 29652 7310
rect 29372 7196 29596 7252
rect 29204 6692 29260 6702
rect 29204 6522 29260 6636
rect 29372 6690 29428 7196
rect 29596 7186 29652 7196
rect 29372 6638 29374 6690
rect 29426 6638 29428 6690
rect 29372 6626 29428 6638
rect 29764 6692 29820 6702
rect 29764 6598 29820 6636
rect 29204 6470 29206 6522
rect 29258 6470 29260 6522
rect 29204 6458 29260 6470
rect 29148 6244 29204 6254
rect 29148 6018 29204 6188
rect 29148 5966 29150 6018
rect 29202 5966 29204 6018
rect 29148 5954 29204 5966
rect 29932 5962 29988 8988
rect 30100 8372 30156 8382
rect 30268 8372 30324 11116
rect 30716 11172 30772 11342
rect 30716 10724 30772 11116
rect 30716 10658 30772 10668
rect 30940 11284 30996 12126
rect 31106 12180 31162 12190
rect 31106 12086 31162 12124
rect 31276 11956 31332 13916
rect 31388 13748 31444 13758
rect 31724 13746 31780 13758
rect 31388 13654 31444 13692
rect 31556 13690 31612 13702
rect 31556 13638 31558 13690
rect 31610 13638 31612 13690
rect 31556 13076 31612 13638
rect 31724 13694 31726 13746
rect 31778 13694 31780 13746
rect 31724 13188 31780 13694
rect 31836 13746 31892 15260
rect 32956 15314 33012 16268
rect 33740 16210 33796 16716
rect 33740 16158 33742 16210
rect 33794 16158 33796 16210
rect 33740 16146 33796 16158
rect 34188 16772 34244 16782
rect 33572 16100 33628 16110
rect 33572 16006 33628 16044
rect 33964 16098 34020 16110
rect 33964 16046 33966 16098
rect 34018 16046 34020 16098
rect 33964 15988 34020 16046
rect 34188 16070 34244 16716
rect 34524 16548 34580 18386
rect 35084 18450 35252 18452
rect 35084 18398 35198 18450
rect 35250 18398 35252 18450
rect 35084 18396 35252 18398
rect 34860 18340 34916 18350
rect 34860 18246 34916 18284
rect 35084 17892 35140 18396
rect 35196 18386 35252 18396
rect 35308 18452 35364 18462
rect 35308 18358 35364 18396
rect 36316 18452 36372 19180
rect 36540 19170 36596 19180
rect 37100 19012 37156 19022
rect 37100 19010 37268 19012
rect 37100 18958 37102 19010
rect 37154 18958 37268 19010
rect 37100 18956 37268 18958
rect 37100 18946 37156 18956
rect 36316 18386 36372 18396
rect 36092 18340 36148 18350
rect 36092 18246 36148 18284
rect 36092 18116 36148 18126
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35420 17892 35476 17902
rect 35084 17890 35476 17892
rect 35084 17838 35422 17890
rect 35474 17838 35476 17890
rect 35084 17836 35476 17838
rect 35420 17826 35476 17836
rect 35812 17668 35868 17678
rect 35812 17574 35868 17612
rect 35980 17666 36036 17678
rect 35980 17614 35982 17666
rect 36034 17614 36036 17666
rect 34860 17554 34916 17566
rect 34860 17502 34862 17554
rect 34914 17502 34916 17554
rect 34860 17444 34916 17502
rect 34860 17378 34916 17388
rect 35980 17220 36036 17614
rect 36092 17666 36148 18060
rect 37212 17780 37268 18956
rect 37212 17714 37268 17724
rect 36092 17614 36094 17666
rect 36146 17614 36148 17666
rect 36092 17602 36148 17614
rect 37212 17332 37268 17342
rect 35980 17154 36036 17164
rect 36876 17220 36932 17230
rect 34188 16018 34190 16070
rect 34242 16018 34244 16070
rect 34188 16006 34244 16018
rect 34300 16492 34580 16548
rect 34692 17050 34748 17062
rect 34692 16998 34694 17050
rect 34746 16998 34748 17050
rect 33964 15922 34020 15932
rect 32956 15262 32958 15314
rect 33010 15262 33012 15314
rect 32172 15204 32228 15214
rect 32172 13870 32228 15148
rect 32116 13858 32228 13870
rect 32116 13806 32118 13858
rect 32170 13806 32228 13858
rect 32116 13804 32228 13806
rect 32116 13794 32172 13804
rect 31836 13694 31838 13746
rect 31890 13694 31892 13746
rect 31836 13682 31892 13694
rect 32732 13748 32788 13758
rect 31948 13636 32004 13646
rect 31724 13122 31780 13132
rect 31836 13524 32004 13580
rect 31500 13020 31612 13076
rect 31836 13074 31892 13524
rect 31836 13022 31838 13074
rect 31890 13022 31892 13074
rect 30716 10500 30772 10510
rect 30716 10406 30772 10444
rect 30548 10164 30604 10174
rect 30548 9940 30604 10108
rect 30940 10164 30996 11228
rect 30940 9940 30996 10108
rect 30548 9938 30660 9940
rect 30548 9886 30550 9938
rect 30602 9886 30660 9938
rect 30548 9874 30660 9886
rect 30492 9380 30548 9390
rect 30492 8930 30548 9324
rect 30492 8878 30494 8930
rect 30546 8878 30548 8930
rect 30492 8596 30548 8878
rect 30492 8530 30548 8540
rect 30100 8370 30324 8372
rect 30100 8318 30102 8370
rect 30154 8318 30324 8370
rect 30100 8316 30324 8318
rect 30100 8306 30156 8316
rect 29932 5910 29934 5962
rect 29986 5910 29988 5962
rect 29932 5898 29988 5910
rect 30044 8036 30100 8046
rect 30044 5962 30100 7980
rect 30212 7924 30268 8316
rect 30604 8158 30660 9874
rect 30828 9884 30996 9940
rect 31164 11900 31332 11956
rect 31388 12852 31444 12862
rect 30828 9042 30884 9884
rect 31164 9828 31220 11900
rect 31388 11508 31444 12796
rect 31500 12628 31556 13020
rect 31836 13010 31892 13022
rect 31668 12964 31724 12974
rect 31668 12870 31724 12908
rect 32060 12964 32116 12974
rect 32732 12964 32788 13692
rect 32956 13746 33012 15262
rect 33292 15652 33348 15662
rect 34300 15652 34356 16492
rect 34692 16436 34748 16998
rect 34860 16902 34916 16914
rect 34860 16850 34862 16902
rect 34914 16850 34916 16902
rect 34860 16772 34916 16850
rect 34972 16884 35028 16894
rect 34972 16790 35028 16828
rect 34860 16706 34916 16716
rect 35644 16772 35700 16782
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 34692 16380 35028 16436
rect 35196 16426 35460 16436
rect 34524 16324 34580 16334
rect 34580 16268 34748 16324
rect 34524 16258 34580 16268
rect 34692 16154 34748 16268
rect 34692 16102 34694 16154
rect 34746 16102 34748 16154
rect 34692 16090 34748 16102
rect 34972 16100 35028 16380
rect 35084 16100 35140 16110
rect 34972 16098 35140 16100
rect 34972 16046 35086 16098
rect 35138 16046 35140 16098
rect 34972 16044 35140 16046
rect 35084 16034 35140 16044
rect 35420 16042 35476 16054
rect 33180 14532 33236 14542
rect 33180 14438 33236 14476
rect 32956 13694 32958 13746
rect 33010 13694 33012 13746
rect 32956 13682 33012 13694
rect 33068 13748 33124 13758
rect 33068 13186 33124 13692
rect 33068 13134 33070 13186
rect 33122 13134 33124 13186
rect 33068 13122 33124 13134
rect 32060 12870 32116 12908
rect 32396 12962 32788 12964
rect 32396 12924 32734 12962
rect 32396 12872 32398 12924
rect 32450 12910 32734 12924
rect 32786 12910 32788 12962
rect 32450 12908 32788 12910
rect 32450 12872 32452 12908
rect 32732 12898 32788 12908
rect 32396 12860 32452 12872
rect 32340 12628 32396 12638
rect 31500 12572 31668 12628
rect 31612 12516 31668 12572
rect 31612 12450 31668 12460
rect 31500 12404 31556 12414
rect 31500 12066 31556 12348
rect 32340 12402 32396 12572
rect 33292 12628 33348 15596
rect 33852 15596 34356 15652
rect 34860 15986 34916 15998
rect 34860 15934 34862 15986
rect 34914 15934 34916 15986
rect 33740 15316 33796 15326
rect 33740 15222 33796 15260
rect 33628 14532 33684 14542
rect 33628 14438 33684 14476
rect 33740 13636 33796 13646
rect 33740 13542 33796 13580
rect 33572 12964 33628 12974
rect 33572 12794 33628 12908
rect 33572 12742 33574 12794
rect 33626 12742 33628 12794
rect 33572 12730 33628 12742
rect 33740 12962 33796 12974
rect 33740 12910 33742 12962
rect 33794 12910 33796 12962
rect 33740 12740 33796 12910
rect 33740 12674 33796 12684
rect 33292 12562 33348 12572
rect 33460 12404 33516 12414
rect 33852 12404 33908 15596
rect 34860 15316 34916 15934
rect 34860 15250 34916 15260
rect 35420 15990 35422 16042
rect 35474 15990 35476 16042
rect 35420 15148 35476 15990
rect 35644 15876 35700 16716
rect 35756 16772 35812 16782
rect 35756 16770 36036 16772
rect 35756 16718 35758 16770
rect 35810 16718 36036 16770
rect 35756 16716 36036 16718
rect 35756 16706 35812 16716
rect 35980 16100 36036 16716
rect 36876 16548 36932 17164
rect 36764 16492 36932 16548
rect 36484 16212 36540 16222
rect 36484 16118 36540 16156
rect 35980 16044 36260 16100
rect 36036 15876 36092 15886
rect 35644 15426 35700 15820
rect 35644 15374 35646 15426
rect 35698 15374 35700 15426
rect 35644 15362 35700 15374
rect 35868 15874 36092 15876
rect 35868 15822 36038 15874
rect 36090 15822 36092 15874
rect 35868 15820 36092 15822
rect 35420 15092 35588 15148
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 33964 14532 34020 14542
rect 33964 13076 34020 14476
rect 34412 14530 34468 14542
rect 34412 14478 34414 14530
rect 34466 14478 34468 14530
rect 34412 13972 34468 14478
rect 34412 13906 34468 13916
rect 35532 13748 35588 15092
rect 35868 14532 35924 15820
rect 36036 15810 36092 15820
rect 36204 15426 36260 16044
rect 36204 15374 36206 15426
rect 36258 15374 36260 15426
rect 36204 15362 36260 15374
rect 36764 15370 36820 16492
rect 37212 16098 37268 17276
rect 37212 16046 37214 16098
rect 37266 16046 37268 16098
rect 37212 16034 37268 16046
rect 37044 15876 37100 15886
rect 36764 15318 36766 15370
rect 36818 15318 36820 15370
rect 36764 15306 36820 15318
rect 36876 15874 37100 15876
rect 36876 15822 37046 15874
rect 37098 15822 37100 15874
rect 36876 15820 37100 15822
rect 36876 15370 36932 15820
rect 37044 15810 37100 15820
rect 37324 15652 37380 21308
rect 37548 21362 37604 21374
rect 37548 21310 37550 21362
rect 37602 21310 37604 21362
rect 37548 19908 37604 21310
rect 37772 20244 37828 23436
rect 37996 23156 38052 23660
rect 38332 23604 38388 24668
rect 38332 23538 38388 23548
rect 38556 24722 38612 24734
rect 38556 24670 38558 24722
rect 38610 24670 38612 24722
rect 38556 23938 38612 24670
rect 38780 24164 38836 25228
rect 38892 24948 38948 24986
rect 38892 24882 38948 24892
rect 39564 24724 39620 25900
rect 40236 24948 40292 26852
rect 40348 26292 40404 26302
rect 40348 25618 40404 26236
rect 40460 25956 40516 27244
rect 40964 26852 41020 26862
rect 40964 26402 41020 26796
rect 40964 26350 40966 26402
rect 41018 26350 41020 26402
rect 40964 26338 41020 26350
rect 40460 25890 40516 25900
rect 40684 26292 40740 26302
rect 40348 25566 40350 25618
rect 40402 25566 40404 25618
rect 40348 25554 40404 25566
rect 40684 25506 40740 26236
rect 40684 25454 40686 25506
rect 40738 25454 40740 25506
rect 40684 25442 40740 25454
rect 41132 25396 41188 27468
rect 41244 27300 41300 28700
rect 41356 27914 41412 31836
rect 41580 31826 41636 31836
rect 41692 31892 41748 32060
rect 41916 32004 41972 33294
rect 42588 33346 42644 33852
rect 42588 33294 42590 33346
rect 42642 33294 42644 33346
rect 42588 33282 42644 33294
rect 42700 33460 42756 33470
rect 42700 33346 42756 33404
rect 42700 33294 42702 33346
rect 42754 33294 42756 33346
rect 42700 33282 42756 33294
rect 42812 33348 42868 35868
rect 43036 35812 43092 36876
rect 43372 36484 43428 37438
rect 43204 36372 43260 36382
rect 43204 36370 43316 36372
rect 43204 36318 43206 36370
rect 43258 36318 43316 36370
rect 43204 36306 43316 36318
rect 43036 35746 43092 35756
rect 43036 35476 43092 35486
rect 43036 35382 43092 35420
rect 43148 35028 43204 35038
rect 42924 34914 42980 34926
rect 42924 34862 42926 34914
rect 42978 34862 42980 34914
rect 42924 34468 42980 34862
rect 43148 34914 43204 34972
rect 43148 34862 43150 34914
rect 43202 34862 43204 34914
rect 43148 34850 43204 34862
rect 42924 34402 42980 34412
rect 42868 33292 42980 33348
rect 42812 33282 42868 33292
rect 42252 32452 42308 32462
rect 42252 32450 42420 32452
rect 42252 32398 42254 32450
rect 42306 32398 42420 32450
rect 42252 32396 42420 32398
rect 42252 32386 42308 32396
rect 41916 31938 41972 31948
rect 41692 31826 41748 31836
rect 42028 31778 42084 31790
rect 41692 31734 41748 31746
rect 41692 31682 41694 31734
rect 41746 31682 41748 31734
rect 41692 30212 41748 31682
rect 42028 31726 42030 31778
rect 42082 31726 42084 31778
rect 42028 31220 42084 31726
rect 41692 30146 41748 30156
rect 41804 31164 42084 31220
rect 42252 31778 42308 31790
rect 42252 31726 42254 31778
rect 42306 31726 42308 31778
rect 42252 31220 42308 31726
rect 42364 31780 42420 32396
rect 42924 32116 42980 33292
rect 43148 33346 43204 33358
rect 43148 33294 43150 33346
rect 43202 33294 43204 33346
rect 43148 33012 43204 33294
rect 43148 32946 43204 32956
rect 43260 32788 43316 36306
rect 43372 35698 43428 36428
rect 43484 36454 43540 38220
rect 43708 38050 43764 38556
rect 43932 38612 43988 38622
rect 43708 37998 43710 38050
rect 43762 37998 43764 38050
rect 43708 37986 43764 37998
rect 43820 38164 43876 38174
rect 43484 36402 43486 36454
rect 43538 36402 43540 36454
rect 43484 36390 43540 36402
rect 43596 37828 43652 37838
rect 43372 35646 43374 35698
rect 43426 35646 43428 35698
rect 43372 35634 43428 35646
rect 43428 34916 43484 34954
rect 43428 34850 43484 34860
rect 43372 34692 43428 34702
rect 43372 34130 43428 34636
rect 43372 34078 43374 34130
rect 43426 34078 43428 34130
rect 43372 34066 43428 34078
rect 43484 33514 43540 33526
rect 43484 33462 43486 33514
rect 43538 33462 43540 33514
rect 43036 32732 43316 32788
rect 43372 33346 43428 33358
rect 43372 33294 43374 33346
rect 43426 33294 43428 33346
rect 43372 32788 43428 33294
rect 43484 33348 43540 33462
rect 43484 33282 43540 33292
rect 43596 33236 43652 37772
rect 43708 37268 43764 37278
rect 43820 37268 43876 38108
rect 43708 37266 43876 37268
rect 43708 37214 43710 37266
rect 43762 37214 43876 37266
rect 43708 37212 43876 37214
rect 43708 37202 43764 37212
rect 43820 37156 43876 37212
rect 43820 37090 43876 37100
rect 43932 37268 43988 38556
rect 43708 36426 43764 36438
rect 43708 36374 43710 36426
rect 43762 36374 43764 36426
rect 43708 36260 43764 36374
rect 43708 36194 43764 36204
rect 43932 36426 43988 37212
rect 43932 36374 43934 36426
rect 43986 36374 43988 36426
rect 44044 36447 44100 39004
rect 44156 38862 44212 38874
rect 44156 38810 44158 38862
rect 44210 38810 44212 38862
rect 44156 38276 44212 38810
rect 44380 38862 44436 38874
rect 44380 38810 44382 38862
rect 44434 38810 44436 38862
rect 44380 38724 44436 38810
rect 44380 38658 44436 38668
rect 44156 38210 44212 38220
rect 44212 38052 44268 38062
rect 44212 37958 44268 37996
rect 44492 37828 44548 39788
rect 44604 39172 44660 39182
rect 44604 38890 44660 39116
rect 44604 38838 44606 38890
rect 44658 38838 44660 38890
rect 44604 38826 44660 38838
rect 44716 38948 44772 38958
rect 44716 38890 44772 38892
rect 44716 38838 44718 38890
rect 44770 38838 44772 38890
rect 44716 38826 44772 38838
rect 44492 37762 44548 37772
rect 44828 37492 44884 39900
rect 45276 39620 45332 39630
rect 45164 39618 45332 39620
rect 45164 39566 45278 39618
rect 45330 39566 45332 39618
rect 45164 39564 45332 39566
rect 44940 39396 44996 39406
rect 44940 39302 44996 39340
rect 45052 39284 45108 39294
rect 44940 39172 44996 39182
rect 44940 38724 44996 39116
rect 45052 38890 45108 39228
rect 45164 39172 45220 39564
rect 45276 39554 45332 39564
rect 45388 39618 45444 40124
rect 45388 39566 45390 39618
rect 45442 39566 45444 39618
rect 45388 39554 45444 39566
rect 45500 39620 45556 41132
rect 45948 41186 46228 41188
rect 45948 41134 46174 41186
rect 46226 41134 46228 41186
rect 45948 41132 46228 41134
rect 45724 41076 45780 41086
rect 45724 40516 45780 41020
rect 45724 40450 45780 40460
rect 45836 40740 45892 40750
rect 45612 40404 45668 40414
rect 45612 40310 45668 40348
rect 45836 39732 45892 40684
rect 45948 39956 46004 41132
rect 46172 41122 46228 41132
rect 46060 40964 46116 40974
rect 46060 40402 46116 40908
rect 46284 40628 46340 43372
rect 46396 40964 46452 43596
rect 47180 43204 47236 43214
rect 47292 43204 47348 45164
rect 47516 44322 47572 45388
rect 47516 44270 47518 44322
rect 47570 44270 47572 44322
rect 47516 44258 47572 44270
rect 47236 43148 47348 43204
rect 47404 43876 47460 43886
rect 47180 43138 47236 43148
rect 47404 42756 47460 43820
rect 46732 41860 46788 41870
rect 46732 41766 46788 41804
rect 46396 40908 46676 40964
rect 46284 40562 46340 40572
rect 46060 40350 46062 40402
rect 46114 40350 46116 40402
rect 46060 40338 46116 40350
rect 46172 40516 46228 40526
rect 46172 40414 46228 40460
rect 46396 40516 46452 40526
rect 46396 40422 46452 40460
rect 46620 40516 46676 40908
rect 47404 40740 47460 42700
rect 47516 42754 47572 42766
rect 47516 42702 47518 42754
rect 47570 42702 47572 42754
rect 47516 41972 47572 42702
rect 47516 41906 47572 41916
rect 47404 40674 47460 40684
rect 47516 41076 47572 41086
rect 46620 40450 46676 40460
rect 46172 40402 46284 40414
rect 46172 40350 46230 40402
rect 46282 40350 46284 40402
rect 46172 40348 46284 40350
rect 46228 40338 46284 40348
rect 46508 40404 46564 40414
rect 46508 40310 46564 40348
rect 47124 40404 47180 40414
rect 47124 40310 47180 40348
rect 47516 40402 47572 41020
rect 47516 40350 47518 40402
rect 47570 40350 47572 40402
rect 47516 40338 47572 40350
rect 47292 40290 47348 40302
rect 47292 40238 47294 40290
rect 47346 40238 47348 40290
rect 46788 40180 46844 40190
rect 46284 40178 46844 40180
rect 46284 40126 46790 40178
rect 46842 40126 46844 40178
rect 46284 40124 46844 40126
rect 45948 39900 46116 39956
rect 45836 39676 46004 39732
rect 45164 39106 45220 39116
rect 45052 38838 45054 38890
rect 45106 38838 45108 38890
rect 45052 38826 45108 38838
rect 45164 38862 45220 38874
rect 45164 38810 45166 38862
rect 45218 38810 45220 38862
rect 45164 38724 45220 38810
rect 44940 38668 45220 38724
rect 45388 38862 45444 38874
rect 45388 38810 45390 38862
rect 45442 38810 45444 38862
rect 45388 38724 45444 38810
rect 45388 38658 45444 38668
rect 45276 38050 45332 38062
rect 45276 37998 45278 38050
rect 45330 37998 45332 38050
rect 44268 37436 44884 37492
rect 44940 37826 44996 37838
rect 44940 37774 44942 37826
rect 44994 37774 44996 37826
rect 44268 37281 44324 37436
rect 44268 37229 44270 37281
rect 44322 37229 44324 37281
rect 44156 37156 44212 37166
rect 44156 37062 44212 37100
rect 44044 36395 44046 36447
rect 44098 36395 44100 36447
rect 44044 36383 44100 36395
rect 43932 35700 43988 36374
rect 44044 35700 44100 35710
rect 43932 35698 44100 35700
rect 43932 35646 44046 35698
rect 44098 35646 44100 35698
rect 43932 35644 44100 35646
rect 43708 35588 43764 35598
rect 43708 35494 43764 35532
rect 43708 34916 43764 34926
rect 43708 34822 43764 34860
rect 44044 34916 44100 35644
rect 44268 35364 44324 37229
rect 44604 37268 44660 37278
rect 44604 37266 44884 37268
rect 44604 37214 44606 37266
rect 44658 37214 44884 37266
rect 44604 37212 44884 37214
rect 44604 37202 44660 37212
rect 44716 36484 44772 36494
rect 44716 36390 44772 36428
rect 44604 36260 44660 36270
rect 44436 35812 44492 35822
rect 44436 35718 44492 35756
rect 44268 35308 44548 35364
rect 44044 34850 44100 34860
rect 44044 34692 44100 34702
rect 44044 34598 44100 34636
rect 43932 33572 43988 33582
rect 43932 33514 43988 33516
rect 43932 33462 43934 33514
rect 43986 33462 43988 33514
rect 43932 33450 43988 33462
rect 43596 33170 43652 33180
rect 43932 33346 43988 33358
rect 43932 33294 43934 33346
rect 43986 33294 43988 33346
rect 43036 32228 43092 32732
rect 43372 32722 43428 32732
rect 43932 32452 43988 33294
rect 44156 33348 44212 33358
rect 44156 33254 44212 33292
rect 44156 33124 44212 33134
rect 44156 32562 44212 33068
rect 44156 32510 44158 32562
rect 44210 32510 44212 32562
rect 44156 32498 44212 32510
rect 43932 32386 43988 32396
rect 43596 32228 43652 32238
rect 43036 32172 43428 32228
rect 42924 32060 43204 32116
rect 42364 31714 42420 31724
rect 43036 31780 43092 31790
rect 43036 31691 43038 31724
rect 43090 31691 43092 31724
rect 43036 31679 43092 31691
rect 43148 31750 43204 32060
rect 43148 31698 43150 31750
rect 43202 31698 43204 31750
rect 43148 31686 43204 31698
rect 43372 31750 43428 32172
rect 43372 31698 43374 31750
rect 43426 31698 43428 31750
rect 43372 31686 43428 31698
rect 43596 31750 43652 32172
rect 43876 32004 43932 32014
rect 43876 31910 43932 31948
rect 43596 31698 43598 31750
rect 43650 31698 43652 31750
rect 43596 31686 43652 31698
rect 44044 31780 44100 31790
rect 42588 31556 42644 31566
rect 42588 31554 42980 31556
rect 42588 31502 42590 31554
rect 42642 31502 42980 31554
rect 42588 31500 42980 31502
rect 42588 31490 42644 31500
rect 41804 29428 41860 31164
rect 42252 31154 42308 31164
rect 42700 31332 42756 31342
rect 42588 30660 42644 30670
rect 42196 29652 42252 29662
rect 42196 29558 42252 29596
rect 41804 29362 41860 29372
rect 42476 28868 42532 28878
rect 42476 28754 42532 28812
rect 42476 28702 42478 28754
rect 42530 28702 42532 28754
rect 42476 28690 42532 28702
rect 41356 27862 41358 27914
rect 41410 27862 41412 27914
rect 42028 28420 42084 28430
rect 41356 27850 41412 27862
rect 41804 27860 41860 27870
rect 41804 27766 41860 27804
rect 42028 27858 42084 28364
rect 42028 27806 42030 27858
rect 42082 27806 42084 27858
rect 41356 27300 41412 27310
rect 41244 27298 41412 27300
rect 41244 27246 41358 27298
rect 41410 27246 41412 27298
rect 41244 27244 41412 27246
rect 41356 27234 41412 27244
rect 42028 26908 42084 27806
rect 42028 26852 42532 26908
rect 41916 26516 41972 26526
rect 41468 26514 41972 26516
rect 41468 26462 41918 26514
rect 41970 26462 41972 26514
rect 41468 26460 41972 26462
rect 41244 26290 41300 26302
rect 41244 26238 41246 26290
rect 41298 26238 41300 26290
rect 41244 26180 41300 26238
rect 41244 26114 41300 26124
rect 41356 26290 41412 26302
rect 41356 26238 41358 26290
rect 41410 26238 41412 26290
rect 41356 25844 41412 26238
rect 41356 25778 41412 25788
rect 41468 25618 41524 26460
rect 41916 26450 41972 26460
rect 41468 25566 41470 25618
rect 41522 25566 41524 25618
rect 41468 25554 41524 25566
rect 41580 26290 41636 26302
rect 41580 26238 41582 26290
rect 41634 26238 41636 26290
rect 41132 25340 41524 25396
rect 39004 24668 39620 24724
rect 39900 24892 40292 24948
rect 38892 24164 38948 24174
rect 38780 24162 38948 24164
rect 38780 24110 38894 24162
rect 38946 24110 38948 24162
rect 38780 24108 38948 24110
rect 38556 23886 38558 23938
rect 38610 23886 38612 23938
rect 37996 23154 38164 23156
rect 37996 23102 37998 23154
rect 38050 23102 38164 23154
rect 37996 23100 38164 23102
rect 37996 23090 38052 23100
rect 37940 22372 37996 22382
rect 38108 22372 38164 23100
rect 38332 22932 38388 22942
rect 38556 22932 38612 23886
rect 38780 23604 38836 23614
rect 38332 22930 38612 22932
rect 38332 22878 38334 22930
rect 38386 22878 38612 22930
rect 38332 22876 38612 22878
rect 38668 23156 38724 23166
rect 38108 22316 38220 22372
rect 37940 22278 37996 22316
rect 38164 21810 38220 22316
rect 38164 21758 38166 21810
rect 38218 21758 38220 21810
rect 38164 21700 38220 21758
rect 38164 21634 38220 21644
rect 38332 21476 38388 22876
rect 38444 22370 38500 22382
rect 38444 22318 38446 22370
rect 38498 22318 38500 22370
rect 38444 21812 38500 22318
rect 38668 22148 38724 23100
rect 38668 22082 38724 22092
rect 38444 21746 38500 21756
rect 37884 21420 38388 21476
rect 37884 20580 37940 21420
rect 38556 21364 38612 21374
rect 38556 21270 38612 21308
rect 38780 20580 38836 23548
rect 38892 22260 38948 24108
rect 38892 22194 38948 22204
rect 39004 23378 39060 24668
rect 39788 24500 39844 24510
rect 39004 23326 39006 23378
rect 39058 23326 39060 23378
rect 38892 21586 38948 21598
rect 38892 21534 38894 21586
rect 38946 21534 38948 21586
rect 38892 20804 38948 21534
rect 39004 21252 39060 23326
rect 39228 24498 39844 24500
rect 39228 24446 39790 24498
rect 39842 24446 39844 24498
rect 39228 24444 39844 24446
rect 39228 22482 39284 24444
rect 39788 24434 39844 24444
rect 39228 22430 39230 22482
rect 39282 22430 39284 22482
rect 39228 22418 39284 22430
rect 39340 24164 39396 24174
rect 39340 23154 39396 24108
rect 39900 23828 39956 24892
rect 41356 24761 41412 24773
rect 40124 24724 40180 24734
rect 40348 24724 40404 24734
rect 40124 24722 40292 24724
rect 40124 24670 40126 24722
rect 40178 24670 40292 24722
rect 40124 24668 40292 24670
rect 40124 24658 40180 24668
rect 40124 23940 40180 23950
rect 40124 23846 40180 23884
rect 39340 23102 39342 23154
rect 39394 23102 39396 23154
rect 39004 21186 39060 21196
rect 39116 22148 39172 22158
rect 38892 20738 38948 20748
rect 39004 20802 39060 20814
rect 39004 20750 39006 20802
rect 39058 20750 39060 20802
rect 37884 20524 38052 20580
rect 37772 20178 37828 20188
rect 37716 20074 37772 20086
rect 37716 20022 37718 20074
rect 37770 20022 37772 20074
rect 37716 20020 37772 20022
rect 37716 19964 37828 20020
rect 37436 19234 37492 19246
rect 37436 19182 37438 19234
rect 37490 19182 37492 19234
rect 37436 18564 37492 19182
rect 37548 19234 37604 19852
rect 37548 19182 37550 19234
rect 37602 19182 37604 19234
rect 37548 19170 37604 19182
rect 37772 19234 37828 19964
rect 37884 20018 37940 20030
rect 37884 19966 37886 20018
rect 37938 19966 37940 20018
rect 37884 19908 37940 19966
rect 37996 20020 38052 20524
rect 38556 20524 38836 20580
rect 38108 20468 38164 20478
rect 38108 20130 38164 20412
rect 38108 20078 38110 20130
rect 38162 20078 38164 20130
rect 38108 20066 38164 20078
rect 38444 20244 38500 20254
rect 37996 19954 38052 19964
rect 38276 19962 38332 19974
rect 37884 19842 37940 19852
rect 38276 19910 38278 19962
rect 38330 19910 38332 19962
rect 38276 19908 38332 19910
rect 38276 19842 38332 19852
rect 38052 19460 38108 19470
rect 38052 19366 38108 19404
rect 37772 19182 37774 19234
rect 37826 19182 37828 19234
rect 37772 19124 37828 19182
rect 38444 19124 38500 20188
rect 38556 19358 38612 20524
rect 39004 20468 39060 20750
rect 39004 20402 39060 20412
rect 39116 20188 39172 22092
rect 39340 21924 39396 23102
rect 39676 23772 39956 23828
rect 39676 23378 39732 23772
rect 40236 23770 40292 24668
rect 40236 23718 40238 23770
rect 40290 23718 40292 23770
rect 40348 23828 40404 24668
rect 40908 24724 40964 24734
rect 40908 24630 40964 24668
rect 41356 24709 41358 24761
rect 41410 24709 41412 24761
rect 41356 24612 41412 24709
rect 41356 24546 41412 24556
rect 41244 24500 41300 24510
rect 40572 24108 41188 24164
rect 40572 23940 40628 24108
rect 41132 24050 41188 24108
rect 41132 23998 41134 24050
rect 41186 23998 41188 24050
rect 41132 23986 41188 23998
rect 40516 23884 40628 23940
rect 40684 23938 40740 23950
rect 40684 23886 40686 23938
rect 40738 23886 40740 23938
rect 40516 23882 40572 23884
rect 40516 23830 40518 23882
rect 40570 23830 40572 23882
rect 40516 23818 40572 23830
rect 40684 23828 40740 23886
rect 40908 23940 40964 23950
rect 40348 23762 40404 23772
rect 40740 23772 40852 23828
rect 40684 23762 40740 23772
rect 40236 23706 40292 23718
rect 39676 23326 39678 23378
rect 39730 23326 39732 23378
rect 39676 23156 39732 23326
rect 40292 23604 40348 23614
rect 40292 23378 40348 23548
rect 40292 23326 40294 23378
rect 40346 23326 40348 23378
rect 40292 23314 40348 23326
rect 40684 23492 40740 23502
rect 39676 23090 39732 23100
rect 39340 21858 39396 21868
rect 40572 22820 40628 22830
rect 40572 21924 40628 22764
rect 39788 21812 39844 21822
rect 39340 21586 39396 21598
rect 39340 21534 39342 21586
rect 39394 21534 39396 21586
rect 39340 20580 39396 21534
rect 39676 21588 39732 21598
rect 39676 21494 39732 21532
rect 39788 20802 39844 21756
rect 40292 21700 40348 21710
rect 40292 21606 40348 21644
rect 40124 21476 40180 21486
rect 39788 20750 39790 20802
rect 39842 20750 39844 20802
rect 39788 20692 39844 20750
rect 39788 20626 39844 20636
rect 39900 21252 39956 21262
rect 40124 21252 40180 21420
rect 40124 21196 40292 21252
rect 39900 20802 39956 21196
rect 39900 20750 39902 20802
rect 39954 20750 39956 20802
rect 39340 20514 39396 20524
rect 39900 20580 39956 20750
rect 39900 20514 39956 20524
rect 40124 20692 40180 20702
rect 39116 20132 39396 20188
rect 38780 20020 38836 20030
rect 38780 19926 38836 19964
rect 39116 19796 39172 19806
rect 38892 19684 38948 19694
rect 38556 19346 38668 19358
rect 38556 19294 38614 19346
rect 38666 19294 38668 19346
rect 38556 19292 38668 19294
rect 38612 19282 38668 19292
rect 37772 19058 37828 19068
rect 38388 19068 38500 19124
rect 38668 19124 38724 19134
rect 38388 18676 38444 19068
rect 37436 18498 37492 18508
rect 37548 18620 38444 18676
rect 37548 17108 37604 18620
rect 38388 18506 38444 18620
rect 38220 18452 38276 18462
rect 38388 18454 38390 18506
rect 38442 18454 38444 18506
rect 38388 18442 38444 18454
rect 38556 18452 38612 18462
rect 37996 18338 38052 18350
rect 37996 18286 37998 18338
rect 38050 18286 38052 18338
rect 37996 18116 38052 18286
rect 37996 18050 38052 18060
rect 37772 17668 37828 17678
rect 36876 15318 36878 15370
rect 36930 15318 36932 15370
rect 36876 15306 36932 15318
rect 36988 15596 37380 15652
rect 37436 17052 37604 17108
rect 37660 17332 37716 17342
rect 36036 15258 36092 15270
rect 36036 15206 36038 15258
rect 36090 15206 36092 15258
rect 36036 15204 36092 15206
rect 36036 15138 36092 15148
rect 36316 14644 36372 14654
rect 36316 14550 36372 14588
rect 36988 14532 37044 15596
rect 37436 15438 37492 17052
rect 37660 16994 37716 17276
rect 37660 16942 37662 16994
rect 37714 16942 37716 16994
rect 37660 16930 37716 16942
rect 37380 15426 37492 15438
rect 37380 15374 37382 15426
rect 37434 15374 37492 15426
rect 37380 15372 37492 15374
rect 37548 16884 37604 16894
rect 37380 15148 37436 15372
rect 37548 15314 37604 16828
rect 37660 16100 37716 16110
rect 37772 16100 37828 17612
rect 38108 17666 38164 17678
rect 38108 17614 38110 17666
rect 38162 17614 38164 17666
rect 38108 16884 38164 17614
rect 38220 17668 38276 18396
rect 38556 18358 38612 18396
rect 38220 17574 38276 17612
rect 38556 17556 38612 17566
rect 38108 16818 38164 16828
rect 38220 17220 38276 17230
rect 38220 16670 38276 17164
rect 38444 16884 38500 16894
rect 38164 16658 38276 16670
rect 38164 16606 38166 16658
rect 38218 16606 38276 16658
rect 38164 16604 38276 16606
rect 38332 16882 38500 16884
rect 38332 16830 38446 16882
rect 38498 16830 38500 16882
rect 38332 16828 38500 16830
rect 38164 16594 38220 16604
rect 37660 16098 37828 16100
rect 37660 16046 37662 16098
rect 37714 16046 37828 16098
rect 37660 16044 37828 16046
rect 37884 16548 37940 16558
rect 37660 16034 37716 16044
rect 37548 15262 37550 15314
rect 37602 15262 37604 15314
rect 37548 15250 37604 15262
rect 37884 15148 37940 16492
rect 37324 15092 37436 15148
rect 37716 15092 37940 15148
rect 38108 16100 38164 16110
rect 35868 14466 35924 14476
rect 36764 14476 37044 14532
rect 37212 14644 37268 14654
rect 37212 14530 37268 14588
rect 37212 14478 37214 14530
rect 37266 14478 37268 14530
rect 36652 14308 36708 14318
rect 36316 14084 36372 14094
rect 36204 13972 36260 13982
rect 36036 13860 36092 13870
rect 36036 13802 36092 13804
rect 36036 13750 36038 13802
rect 36090 13750 36092 13802
rect 36204 13858 36260 13916
rect 36204 13806 36206 13858
rect 36258 13806 36260 13858
rect 36204 13794 36260 13806
rect 36036 13738 36092 13750
rect 35532 13682 35588 13692
rect 35644 13634 35700 13646
rect 35644 13582 35646 13634
rect 35698 13582 35700 13634
rect 35196 13356 35460 13366
rect 34692 13300 34748 13310
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 34692 13186 34748 13244
rect 34692 13134 34694 13186
rect 34746 13134 34748 13186
rect 34692 13122 34748 13134
rect 34132 13076 34188 13086
rect 33964 13074 34188 13076
rect 33964 13022 34134 13074
rect 34186 13022 34188 13074
rect 33964 13020 34188 13022
rect 32340 12350 32342 12402
rect 32394 12350 32396 12402
rect 32340 12338 32396 12350
rect 33292 12348 33460 12404
rect 31500 12014 31502 12066
rect 31554 12014 31556 12066
rect 31500 12002 31556 12014
rect 31612 12180 31668 12190
rect 31500 11508 31556 11518
rect 31388 11506 31556 11508
rect 31388 11454 31502 11506
rect 31554 11454 31556 11506
rect 31388 11452 31556 11454
rect 31500 11442 31556 11452
rect 31612 10724 31668 12124
rect 32508 12178 32564 12190
rect 32508 12126 32510 12178
rect 32562 12126 32564 12178
rect 32508 11956 32564 12126
rect 32508 11890 32564 11900
rect 33292 11732 33348 12348
rect 33460 12310 33516 12348
rect 33628 12348 33908 12404
rect 34076 13010 34188 13020
rect 33292 11666 33348 11676
rect 33404 11844 33460 11854
rect 33404 11506 33460 11788
rect 33404 11454 33406 11506
rect 33458 11454 33460 11506
rect 33404 11442 33460 11454
rect 32620 11172 32676 11182
rect 32340 10778 32396 10790
rect 32340 10726 32342 10778
rect 32394 10726 32396 10778
rect 31388 10668 31706 10724
rect 31276 10388 31332 10398
rect 31276 10294 31332 10332
rect 31276 9828 31332 9838
rect 31164 9826 31332 9828
rect 30828 8990 30830 9042
rect 30882 8990 30884 9042
rect 30828 8978 30884 8990
rect 30940 9770 30996 9782
rect 31164 9774 31278 9826
rect 31330 9774 31332 9826
rect 31164 9772 31332 9774
rect 30940 9718 30942 9770
rect 30994 9718 30996 9770
rect 31276 9762 31332 9772
rect 30940 8596 30996 9718
rect 31164 8820 31220 8830
rect 31164 8726 31220 8764
rect 30828 8540 30996 8596
rect 30548 8146 30660 8158
rect 30548 8094 30550 8146
rect 30602 8094 30660 8146
rect 30548 8092 30660 8094
rect 30716 8258 30772 8270
rect 30716 8206 30718 8258
rect 30770 8206 30772 8258
rect 30548 8082 30604 8092
rect 30716 7924 30772 8206
rect 30212 7868 30772 7924
rect 30828 8036 30884 8540
rect 30212 7700 30268 7868
rect 30212 7698 30324 7700
rect 30212 7646 30214 7698
rect 30266 7646 30324 7698
rect 30212 7634 30324 7646
rect 30044 5910 30046 5962
rect 30098 5910 30100 5962
rect 30044 5898 30100 5910
rect 30268 6692 30324 7634
rect 30828 7588 30884 7980
rect 30772 7530 30884 7588
rect 30772 7478 30774 7530
rect 30826 7478 30884 7530
rect 30772 7466 30884 7478
rect 29596 5796 29652 5806
rect 29316 5460 29372 5470
rect 29316 5234 29372 5404
rect 29316 5182 29318 5234
rect 29370 5182 29372 5234
rect 29316 5170 29372 5182
rect 29484 5348 29540 5358
rect 29484 5122 29540 5292
rect 29484 5070 29486 5122
rect 29538 5070 29540 5122
rect 29484 5058 29540 5070
rect 29484 4452 29540 4462
rect 29484 4358 29540 4396
rect 29596 3666 29652 5740
rect 30268 5348 30324 6636
rect 30828 6580 30884 7466
rect 30940 8372 30996 8382
rect 30940 7474 30996 8316
rect 31388 7700 31444 10668
rect 31650 10648 31706 10668
rect 31650 10596 31652 10648
rect 31704 10596 31706 10648
rect 31650 10584 31706 10596
rect 31836 10610 31892 10622
rect 31836 10558 31838 10610
rect 31890 10558 31892 10610
rect 31836 10164 31892 10558
rect 31948 10612 32004 10622
rect 32340 10612 32396 10726
rect 31948 10610 32396 10612
rect 31948 10558 31950 10610
rect 32002 10558 32396 10610
rect 31948 10556 32396 10558
rect 32508 10610 32564 10622
rect 32508 10558 32510 10610
rect 32562 10558 32564 10610
rect 31948 10546 32004 10556
rect 32508 10500 32564 10558
rect 32508 10276 32564 10444
rect 32508 10210 32564 10220
rect 31836 10098 31892 10108
rect 31836 9940 31892 9950
rect 31836 9826 31892 9884
rect 31668 9770 31724 9782
rect 31500 9714 31556 9726
rect 31500 9662 31502 9714
rect 31554 9662 31556 9714
rect 31500 8370 31556 9662
rect 31668 9718 31670 9770
rect 31722 9718 31724 9770
rect 31836 9774 31838 9826
rect 31890 9774 31892 9826
rect 31836 9762 31892 9774
rect 31668 9156 31724 9718
rect 32620 9716 32676 11116
rect 32956 10724 33012 10734
rect 32956 10612 33012 10668
rect 32844 10610 33012 10612
rect 32844 10558 32958 10610
rect 33010 10558 33012 10610
rect 32844 10556 33012 10558
rect 32844 9950 32900 10556
rect 32956 10546 33012 10556
rect 32788 9940 32900 9950
rect 33236 9940 33292 9950
rect 32788 9938 33292 9940
rect 32788 9886 32790 9938
rect 32842 9886 33238 9938
rect 33290 9886 33292 9938
rect 32788 9884 33292 9886
rect 32788 9874 32844 9884
rect 33236 9874 33292 9884
rect 33628 9828 33684 12348
rect 33852 12193 33908 12205
rect 33852 12141 33854 12193
rect 33906 12141 33908 12193
rect 33740 12066 33796 12078
rect 33740 12014 33742 12066
rect 33794 12014 33796 12066
rect 33740 10610 33796 12014
rect 33852 11620 33908 12141
rect 33852 11554 33908 11564
rect 34076 11518 34132 13010
rect 34860 12964 34916 12974
rect 34860 12290 34916 12908
rect 34860 12238 34862 12290
rect 34914 12238 34916 12290
rect 34860 12226 34916 12238
rect 34972 12962 35028 12974
rect 34972 12910 34974 12962
rect 35026 12910 35028 12962
rect 34020 11506 34132 11518
rect 34020 11454 34022 11506
rect 34074 11454 34132 11506
rect 34020 11452 34132 11454
rect 34188 12178 34244 12190
rect 34188 12126 34190 12178
rect 34242 12126 34244 12178
rect 34020 10724 34076 11452
rect 34188 11396 34244 12126
rect 34524 12180 34580 12190
rect 34972 12178 35028 12910
rect 35196 12964 35252 12974
rect 35196 12870 35252 12908
rect 35644 12740 35700 13582
rect 36204 13412 36260 13422
rect 36204 13186 36260 13356
rect 36204 13134 36206 13186
rect 36258 13134 36260 13186
rect 35812 13076 35868 13086
rect 35812 12740 35868 13020
rect 36204 12964 36260 13134
rect 36204 12898 36260 12908
rect 35644 12674 35700 12684
rect 35756 12738 35868 12740
rect 35756 12686 35814 12738
rect 35866 12686 35868 12738
rect 35756 12674 35868 12686
rect 35756 12404 35812 12674
rect 35756 12310 35812 12348
rect 36204 12628 36260 12638
rect 34524 12086 34580 12124
rect 34692 12122 34748 12134
rect 34692 12070 34694 12122
rect 34746 12070 34748 12122
rect 34692 12068 34748 12070
rect 34692 12002 34748 12012
rect 34972 12126 34974 12178
rect 35026 12126 35028 12178
rect 34300 11732 34356 11742
rect 34300 11450 34356 11676
rect 34972 11620 35028 12126
rect 35644 12180 35700 12190
rect 36092 12180 36148 12190
rect 35252 11956 35308 11966
rect 34300 11398 34302 11450
rect 34354 11398 34356 11450
rect 34300 11386 34356 11398
rect 34860 11564 35028 11620
rect 35084 11954 35308 11956
rect 35084 11902 35254 11954
rect 35306 11902 35308 11954
rect 35084 11900 35308 11902
rect 35084 11620 35140 11900
rect 35252 11890 35308 11900
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35476 11620 35532 11630
rect 35084 11564 35196 11620
rect 34188 11330 34244 11340
rect 34524 11338 34580 11350
rect 34524 11286 34526 11338
rect 34578 11286 34580 11338
rect 34524 11284 34580 11286
rect 34524 11218 34580 11228
rect 33740 10558 33742 10610
rect 33794 10558 33796 10610
rect 33740 10546 33796 10558
rect 33964 10668 34020 10724
rect 33964 10658 34076 10668
rect 32620 9650 32676 9660
rect 33516 9772 33684 9828
rect 32172 9604 32228 9614
rect 32172 9602 32284 9604
rect 32172 9550 32174 9602
rect 32226 9550 32284 9602
rect 32172 9538 32284 9550
rect 31668 9100 31892 9156
rect 31836 8930 31892 9100
rect 31836 8878 31838 8930
rect 31890 8878 31892 8930
rect 31836 8866 31892 8878
rect 32228 9054 32284 9538
rect 33516 9380 33572 9772
rect 33684 9604 33740 9614
rect 33740 9548 33908 9604
rect 33684 9510 33740 9548
rect 33852 9380 33908 9548
rect 33516 9324 33740 9380
rect 33628 9266 33740 9324
rect 33964 9380 34020 10658
rect 34412 10276 34468 10286
rect 34860 10276 34916 11564
rect 35140 11450 35196 11564
rect 35476 11526 35532 11564
rect 34972 11396 35028 11434
rect 34972 11330 35028 11340
rect 35140 11398 35142 11450
rect 35194 11398 35196 11450
rect 35140 11396 35196 11398
rect 35140 11320 35196 11340
rect 34132 10164 34188 10174
rect 34132 9938 34188 10108
rect 34132 9886 34134 9938
rect 34186 9886 34188 9938
rect 34132 9874 34188 9886
rect 34412 9826 34468 10220
rect 34412 9774 34414 9826
rect 34466 9774 34468 9826
rect 34412 9762 34468 9774
rect 34524 10220 34916 10276
rect 35532 11284 35588 11294
rect 35196 10220 35460 10230
rect 34524 9826 34580 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35084 9940 35140 9950
rect 34972 9938 35140 9940
rect 34972 9886 35086 9938
rect 35138 9886 35140 9938
rect 34972 9884 35140 9886
rect 34524 9774 34526 9826
rect 34578 9774 34580 9826
rect 33964 9324 34188 9380
rect 33852 9314 33908 9324
rect 33628 9214 33686 9266
rect 33738 9214 33740 9266
rect 33628 9202 33740 9214
rect 34132 9266 34188 9324
rect 34132 9214 34134 9266
rect 34186 9214 34188 9266
rect 34132 9202 34188 9214
rect 32228 9042 32286 9054
rect 32228 8990 32232 9042
rect 32284 8990 32286 9042
rect 32228 8978 32286 8990
rect 32396 9042 32452 9054
rect 32396 8990 32398 9042
rect 32450 8990 32452 9042
rect 32228 8932 32284 8978
rect 32228 8866 32284 8876
rect 32396 8820 32452 8990
rect 32508 9044 32564 9054
rect 33292 9044 33348 9054
rect 32508 9042 33180 9044
rect 32508 8990 32510 9042
rect 32562 8990 33180 9042
rect 32508 8988 33180 8990
rect 32508 8978 32564 8988
rect 33124 8874 33180 8988
rect 33292 9042 33460 9044
rect 33292 8990 33294 9042
rect 33346 8990 33460 9042
rect 33292 8988 33460 8990
rect 33292 8978 33348 8988
rect 33124 8822 33126 8874
rect 33178 8822 33180 8874
rect 33124 8810 33180 8822
rect 32396 8596 32452 8764
rect 32396 8540 32676 8596
rect 31500 8318 31502 8370
rect 31554 8318 31556 8370
rect 31500 8306 31556 8318
rect 31388 7634 31444 7644
rect 32138 8036 32194 8046
rect 32620 8036 32676 8540
rect 32138 7512 32194 7980
rect 30940 7422 30942 7474
rect 30994 7422 30996 7474
rect 30940 7410 30996 7422
rect 31332 7474 31388 7486
rect 31332 7422 31334 7474
rect 31386 7422 31388 7474
rect 32138 7460 32140 7512
rect 32192 7460 32194 7512
rect 32138 7448 32194 7460
rect 32284 7980 32676 8036
rect 33404 8146 33460 8988
rect 33404 8094 33406 8146
rect 33458 8094 33460 8146
rect 32284 7474 32340 7980
rect 33404 7812 33460 8094
rect 33628 8932 33684 9202
rect 34524 9044 34580 9774
rect 34692 9828 34748 9838
rect 34692 9734 34748 9772
rect 34972 9086 35028 9884
rect 35084 9874 35140 9884
rect 35532 9716 35588 11228
rect 35644 10722 35700 12124
rect 35868 12178 36148 12180
rect 35868 12126 36094 12178
rect 36146 12126 36148 12178
rect 35868 12124 36148 12126
rect 35868 11620 35924 12124
rect 36092 12114 36148 12124
rect 36204 12068 36260 12572
rect 35868 11554 35924 11564
rect 36036 11732 36092 11742
rect 36036 11450 36092 11676
rect 35756 11396 35812 11406
rect 36036 11398 36038 11450
rect 36090 11398 36092 11450
rect 36036 11386 36092 11398
rect 36204 11394 36260 12012
rect 35756 11302 35812 11340
rect 36204 11342 36206 11394
rect 36258 11342 36260 11394
rect 35868 11284 35924 11294
rect 35868 11190 35924 11228
rect 35644 10670 35646 10722
rect 35698 10670 35700 10722
rect 35644 9826 35700 10670
rect 35980 10612 36036 10622
rect 35644 9774 35646 9826
rect 35698 9774 35700 9826
rect 35644 9762 35700 9774
rect 35868 10556 35980 10612
rect 33628 8036 33684 8876
rect 34076 8988 34580 9044
rect 34636 9042 34692 9054
rect 34636 8990 34638 9042
rect 34690 8990 34692 9042
rect 33628 7970 33684 7980
rect 33740 8260 33796 8270
rect 34076 8260 34132 8988
rect 34636 8932 34692 8990
rect 34972 9044 34974 9086
rect 35026 9044 35028 9086
rect 34972 8956 35028 8988
rect 35084 9660 35588 9716
rect 34636 8484 34692 8876
rect 34300 8428 34692 8484
rect 35084 8930 35140 9660
rect 35868 9156 35924 10556
rect 35980 10518 36036 10556
rect 36204 10052 36260 11342
rect 36316 10388 36372 14028
rect 36652 13774 36708 14252
rect 36652 13748 36654 13774
rect 36706 13748 36708 13774
rect 36652 13682 36708 13692
rect 36764 13076 36820 14476
rect 37212 14466 37268 14478
rect 37044 14308 37100 14318
rect 36876 14306 37100 14308
rect 36876 14254 37046 14306
rect 37098 14254 37100 14306
rect 36876 14252 37100 14254
rect 36876 13802 36932 14252
rect 37044 14242 37100 14252
rect 36876 13750 36878 13802
rect 36930 13750 36932 13802
rect 36876 13738 36932 13750
rect 37212 13690 37268 13702
rect 37212 13638 37214 13690
rect 37266 13638 37268 13690
rect 37212 13636 37268 13638
rect 37100 13580 37268 13636
rect 36540 13020 36820 13076
rect 36540 12962 36596 13020
rect 36540 12910 36542 12962
rect 36594 12910 36596 12962
rect 36540 12898 36596 12910
rect 36484 12628 36540 12638
rect 36484 12402 36540 12572
rect 36484 12350 36486 12402
rect 36538 12350 36540 12402
rect 36484 12338 36540 12350
rect 36764 11844 36820 13020
rect 36876 13412 36932 13422
rect 36876 12180 36932 13356
rect 37100 13076 37156 13580
rect 37324 13412 37380 15092
rect 37716 14306 37772 15092
rect 38108 14642 38164 16044
rect 38332 15428 38388 16828
rect 38444 16818 38500 16828
rect 38556 16882 38612 17500
rect 38556 16830 38558 16882
rect 38610 16830 38612 16882
rect 38556 16818 38612 16830
rect 38444 16100 38500 16110
rect 38444 16006 38500 16044
rect 38668 15540 38724 19068
rect 38780 18452 38836 18462
rect 38892 18452 38948 19628
rect 39116 19124 39172 19740
rect 39116 19058 39172 19068
rect 39228 19206 39284 19218
rect 39228 19154 39230 19206
rect 39282 19154 39284 19206
rect 38780 18450 38948 18452
rect 38780 18398 38782 18450
rect 38834 18398 38948 18450
rect 38780 18396 38948 18398
rect 38780 18386 38836 18396
rect 38780 17668 38836 17678
rect 38780 16882 38836 17612
rect 38780 16830 38782 16882
rect 38834 16830 38836 16882
rect 38780 16818 38836 16830
rect 38892 16548 38948 18396
rect 39116 18488 39172 18500
rect 39116 18436 39118 18488
rect 39170 18436 39172 18488
rect 39116 18340 39172 18436
rect 39116 18274 39172 18284
rect 39004 17780 39060 17790
rect 39004 17686 39060 17724
rect 38892 16482 38948 16492
rect 39228 16884 39284 19154
rect 39340 18004 39396 20132
rect 39452 20132 39508 20142
rect 39452 19684 39508 20076
rect 40012 20018 40068 20030
rect 40012 19966 40014 20018
rect 40066 19966 40068 20018
rect 39900 19908 39956 19918
rect 39900 19850 39956 19852
rect 39900 19798 39902 19850
rect 39954 19798 39956 19850
rect 39900 19786 39956 19798
rect 39452 19618 39508 19628
rect 40012 19460 40068 19966
rect 40012 19394 40068 19404
rect 40124 19460 40180 20636
rect 40236 20580 40292 21196
rect 40236 20486 40292 20524
rect 40572 20802 40628 21868
rect 40684 21588 40740 23436
rect 40796 22260 40852 23772
rect 40908 23278 40964 23884
rect 41244 23923 41300 24444
rect 41468 24388 41524 25340
rect 41580 24890 41636 26238
rect 42476 26292 42532 26852
rect 42588 26740 42644 30604
rect 42700 30100 42756 31276
rect 42924 30994 42980 31500
rect 42924 30942 42926 30994
rect 42978 30942 42980 30994
rect 42924 30930 42980 30942
rect 43596 31220 43652 31230
rect 43484 30548 43540 30558
rect 42700 29538 42756 30044
rect 42700 29486 42702 29538
rect 42754 29486 42756 29538
rect 42700 29474 42756 29486
rect 43036 30210 43092 30222
rect 43036 30158 43038 30210
rect 43090 30158 43092 30210
rect 42812 29092 42868 29102
rect 42812 27858 42868 29036
rect 42812 27806 42814 27858
rect 42866 27806 42868 27858
rect 42812 27794 42868 27806
rect 43036 27860 43092 30158
rect 43484 30171 43540 30492
rect 43484 30119 43486 30171
rect 43538 30119 43540 30171
rect 43484 30107 43540 30119
rect 43596 30042 43652 31164
rect 43708 30996 43764 31006
rect 43708 30994 43876 30996
rect 43708 30942 43710 30994
rect 43762 30942 43876 30994
rect 43708 30940 43876 30942
rect 43708 30930 43764 30940
rect 43596 29990 43598 30042
rect 43650 29990 43652 30042
rect 43596 29978 43652 29990
rect 43708 30210 43764 30222
rect 43708 30158 43710 30210
rect 43762 30158 43764 30210
rect 43708 29988 43764 30158
rect 43820 30212 43876 30940
rect 44044 30994 44100 31724
rect 44044 30942 44046 30994
rect 44098 30942 44100 30994
rect 44044 30930 44100 30942
rect 43932 30826 43988 30838
rect 43932 30774 43934 30826
rect 43986 30774 43988 30826
rect 43932 30548 43988 30774
rect 43932 30482 43988 30492
rect 44492 30436 44548 35308
rect 44604 35028 44660 36204
rect 44604 33908 44660 34972
rect 44604 33842 44660 33852
rect 44716 35698 44772 35710
rect 44716 35646 44718 35698
rect 44770 35646 44772 35698
rect 44716 33572 44772 35646
rect 44828 35700 44884 37212
rect 44940 37044 44996 37774
rect 45164 37266 45220 37278
rect 45164 37214 45166 37266
rect 45218 37214 45220 37266
rect 45164 37156 45220 37214
rect 45164 37090 45220 37100
rect 44940 36978 44996 36988
rect 45276 36932 45332 37998
rect 45388 38052 45444 38090
rect 45500 38052 45556 39564
rect 45724 39620 45780 39630
rect 45612 39508 45668 39518
rect 45612 38948 45668 39452
rect 45612 38890 45668 38892
rect 45612 38838 45614 38890
rect 45666 38838 45668 38890
rect 45612 38826 45668 38838
rect 45724 38668 45780 39564
rect 45948 38958 46004 39676
rect 45892 38946 46004 38958
rect 45892 38894 45894 38946
rect 45946 38894 46004 38946
rect 45892 38892 46004 38894
rect 45892 38882 45948 38892
rect 45724 38612 45892 38668
rect 45444 37996 45556 38052
rect 45388 37986 45444 37996
rect 45388 37828 45444 37838
rect 45388 37266 45444 37772
rect 45388 37214 45390 37266
rect 45442 37214 45444 37266
rect 45388 37202 45444 37214
rect 45276 36866 45332 36876
rect 45276 36596 45332 36606
rect 45052 36260 45108 36270
rect 45052 36166 45108 36204
rect 44828 34244 44884 35644
rect 45164 35698 45220 35710
rect 45164 35646 45166 35698
rect 45218 35646 45220 35698
rect 44940 35028 44996 35038
rect 44940 34934 44996 34972
rect 45164 34468 45220 35646
rect 45276 34914 45332 36540
rect 45388 36484 45444 36494
rect 45500 36484 45556 37996
rect 45388 36482 45556 36484
rect 45388 36430 45390 36482
rect 45442 36430 45556 36482
rect 45388 36428 45556 36430
rect 45388 36418 45444 36428
rect 45388 35812 45444 35822
rect 45388 35754 45444 35756
rect 45388 35702 45390 35754
rect 45442 35702 45444 35754
rect 45388 35690 45444 35702
rect 45276 34862 45278 34914
rect 45330 34862 45332 34914
rect 45276 34850 45332 34862
rect 45388 35588 45444 35598
rect 45388 34914 45444 35532
rect 45388 34862 45390 34914
rect 45442 34862 45444 34914
rect 45388 34850 45444 34862
rect 45164 34402 45220 34412
rect 44828 34178 44884 34188
rect 45276 34244 45332 34254
rect 45276 34150 45332 34188
rect 45276 34020 45332 34030
rect 45500 34020 45556 36428
rect 45668 37042 45724 37054
rect 45668 36990 45670 37042
rect 45722 36990 45724 37042
rect 45668 36484 45724 36990
rect 45668 36418 45724 36428
rect 45668 35476 45724 35486
rect 45668 35474 45780 35476
rect 45668 35422 45670 35474
rect 45722 35422 45780 35474
rect 45668 35410 45780 35422
rect 45724 35308 45780 35410
rect 45612 35252 45780 35308
rect 45612 35140 45668 35252
rect 45612 35074 45668 35084
rect 45724 35140 45780 35150
rect 45836 35140 45892 38612
rect 45724 35138 45892 35140
rect 45724 35086 45726 35138
rect 45778 35086 45892 35138
rect 45724 35084 45892 35086
rect 45948 38388 46004 38398
rect 45724 35074 45780 35084
rect 45948 34692 46004 38332
rect 46060 37154 46116 39900
rect 46172 39620 46228 39630
rect 46172 39526 46228 39564
rect 46284 39396 46340 40124
rect 46788 40114 46844 40124
rect 46172 39340 46340 39396
rect 46396 39844 46452 39854
rect 46172 38276 46228 39340
rect 46396 38948 46452 39788
rect 46284 38834 46340 38846
rect 46284 38782 46286 38834
rect 46338 38782 46340 38834
rect 46284 38724 46340 38782
rect 46396 38834 46452 38892
rect 46732 39172 46788 39182
rect 46396 38782 46398 38834
rect 46450 38782 46452 38834
rect 46396 38770 46452 38782
rect 46562 38836 46618 38846
rect 46562 38742 46618 38780
rect 46284 38658 46340 38668
rect 46396 38612 46452 38622
rect 46172 38220 46340 38276
rect 46172 38050 46228 38062
rect 46172 37998 46174 38050
rect 46226 37998 46228 38050
rect 46172 37604 46228 37998
rect 46172 37538 46228 37548
rect 46284 37380 46340 38220
rect 46396 37492 46452 38556
rect 46732 38388 46788 39116
rect 46956 38836 47012 38846
rect 46956 38722 47012 38780
rect 46956 38670 46958 38722
rect 47010 38670 47012 38722
rect 46956 38658 47012 38670
rect 46732 38322 46788 38332
rect 46732 37828 46788 37838
rect 46396 37436 46564 37492
rect 46228 37324 46340 37380
rect 46228 37322 46284 37324
rect 46228 37270 46230 37322
rect 46282 37270 46284 37322
rect 46228 37258 46284 37270
rect 46396 37268 46452 37278
rect 46396 37174 46452 37212
rect 46060 37102 46062 37154
rect 46114 37102 46116 37154
rect 46060 37090 46116 37102
rect 46172 37044 46228 37054
rect 46172 36594 46228 36988
rect 46172 36542 46174 36594
rect 46226 36542 46228 36594
rect 46172 36530 46228 36542
rect 46284 36932 46340 36942
rect 46284 35866 46340 36876
rect 46508 36820 46564 37436
rect 46732 37266 46788 37772
rect 46732 37214 46734 37266
rect 46786 37214 46788 37266
rect 46732 37202 46788 37214
rect 46956 37716 47012 37726
rect 46956 37266 47012 37660
rect 47292 37492 47348 40238
rect 47460 39060 47516 39070
rect 47460 38946 47516 39004
rect 47460 38894 47462 38946
rect 47514 38894 47516 38946
rect 47460 38882 47516 38894
rect 47628 38668 47684 45724
rect 48076 44996 48132 45006
rect 47852 44994 48132 44996
rect 47852 44942 48078 44994
rect 48130 44942 48132 44994
rect 47852 44940 48132 44942
rect 47740 44322 47796 44334
rect 47740 44270 47742 44322
rect 47794 44270 47796 44322
rect 47740 43092 47796 44270
rect 47852 43988 47908 44940
rect 48076 44930 48132 44940
rect 47852 43922 47908 43932
rect 48020 44210 48076 44222
rect 48020 44158 48022 44210
rect 48074 44158 48076 44210
rect 48020 43764 48076 44158
rect 48020 43698 48076 43708
rect 48188 43652 48244 45782
rect 48188 43586 48244 43596
rect 48300 43540 48356 45948
rect 48300 43474 48356 43484
rect 47740 43026 47796 43036
rect 48076 43426 48132 43438
rect 48076 43374 48078 43426
rect 48130 43374 48132 43426
rect 48076 42868 48132 43374
rect 48076 42802 48132 42812
rect 47740 42756 47796 42766
rect 47740 42662 47796 42700
rect 48020 42644 48076 42654
rect 47852 42642 48076 42644
rect 47852 42590 48022 42642
rect 48074 42590 48076 42642
rect 47852 42588 48076 42590
rect 47852 41636 47908 42588
rect 48020 42578 48076 42588
rect 47852 41570 47908 41580
rect 48076 41524 48132 41534
rect 48076 41298 48132 41468
rect 48076 41246 48078 41298
rect 48130 41246 48132 41298
rect 48076 41234 48132 41246
rect 47740 40852 47796 40862
rect 47740 40458 47796 40796
rect 47740 40406 47742 40458
rect 47794 40406 47796 40458
rect 47740 40394 47796 40406
rect 48076 39508 48132 39518
rect 48076 39414 48132 39452
rect 47740 38836 47796 38846
rect 47740 38742 47796 38780
rect 47852 38834 47908 38846
rect 47852 38782 47854 38834
rect 47906 38782 47908 38834
rect 47628 38612 47796 38668
rect 47292 37426 47348 37436
rect 46956 37214 46958 37266
rect 47010 37214 47012 37266
rect 46956 37202 47012 37214
rect 47236 37268 47292 37278
rect 47516 37268 47572 37278
rect 47236 37266 47572 37268
rect 47236 37214 47238 37266
rect 47290 37214 47518 37266
rect 47570 37214 47572 37266
rect 47236 37212 47572 37214
rect 47236 37202 47292 37212
rect 47516 37202 47572 37212
rect 47740 37266 47796 38612
rect 47740 37214 47742 37266
rect 47794 37214 47796 37266
rect 47740 37202 47796 37214
rect 47852 37156 47908 38782
rect 48076 38276 48132 38286
rect 48076 38162 48132 38220
rect 48076 38110 48078 38162
rect 48130 38110 48132 38162
rect 48076 38098 48132 38110
rect 47852 37090 47908 37100
rect 46284 35814 46286 35866
rect 46338 35814 46340 35866
rect 46284 35802 46340 35814
rect 46396 36764 46564 36820
rect 48020 37042 48076 37054
rect 48020 36990 48022 37042
rect 48074 36990 48076 37042
rect 46284 35698 46340 35710
rect 46284 35646 46286 35698
rect 46338 35646 46340 35698
rect 46284 35140 46340 35646
rect 46284 35074 46340 35084
rect 46396 35138 46452 36764
rect 48020 36596 48076 36990
rect 48020 36530 48076 36540
rect 48076 36372 48132 36382
rect 47740 36370 48132 36372
rect 47740 36318 48078 36370
rect 48130 36318 48132 36370
rect 47740 36316 48132 36318
rect 46620 35737 46676 35749
rect 46620 35685 46622 35737
rect 46674 35685 46676 35737
rect 47740 35742 47796 36316
rect 48076 36306 48132 36316
rect 46620 35588 46676 35685
rect 46844 35700 46900 35710
rect 47404 35700 47460 35710
rect 46844 35698 47348 35700
rect 46844 35646 46846 35698
rect 46898 35646 47348 35698
rect 46844 35644 47348 35646
rect 46844 35634 46900 35644
rect 46620 35522 46676 35532
rect 47292 35364 47348 35644
rect 47460 35644 47684 35700
rect 47404 35606 47460 35644
rect 46396 35086 46398 35138
rect 46450 35086 46452 35138
rect 46396 35074 46452 35086
rect 47180 35140 47236 35150
rect 46060 34916 46116 34926
rect 46060 34822 46116 34860
rect 47012 34804 47068 34814
rect 46508 34802 47068 34804
rect 46508 34750 47014 34802
rect 47066 34750 47068 34802
rect 46508 34748 47068 34750
rect 45948 34636 46452 34692
rect 46396 34298 46452 34636
rect 46396 34246 46398 34298
rect 46450 34246 46452 34298
rect 46396 34234 46452 34246
rect 46508 34132 46564 34748
rect 47012 34738 47068 34748
rect 46396 34130 46564 34132
rect 46396 34078 46510 34130
rect 46562 34078 46564 34130
rect 46396 34076 46564 34078
rect 45332 33964 45556 34020
rect 45892 34020 45948 34030
rect 44716 33506 44772 33516
rect 44828 33908 44884 33918
rect 44716 33346 44772 33358
rect 44716 33294 44718 33346
rect 44770 33294 44772 33346
rect 44716 32004 44772 33294
rect 44716 31938 44772 31948
rect 44716 31778 44772 31790
rect 44716 31726 44718 31778
rect 44770 31726 44772 31778
rect 44716 31220 44772 31726
rect 44716 31154 44772 31164
rect 44716 30994 44772 31006
rect 44716 30942 44718 30994
rect 44770 30942 44772 30994
rect 44716 30884 44772 30942
rect 44828 30884 44884 33852
rect 45276 33348 45332 33964
rect 45892 33926 45948 33964
rect 45388 33348 45444 33358
rect 45276 33346 45444 33348
rect 45276 33294 45390 33346
rect 45442 33294 45444 33346
rect 45276 33292 45444 33294
rect 45052 33124 45108 33134
rect 45052 33030 45108 33068
rect 44940 32562 44996 32574
rect 44940 32510 44942 32562
rect 44994 32510 44996 32562
rect 44940 32452 44996 32510
rect 45388 32462 45444 33292
rect 46172 33346 46228 33358
rect 46172 33294 46174 33346
rect 46226 33294 46228 33346
rect 46172 33236 46228 33294
rect 46172 33170 46228 33180
rect 46396 33124 46452 34076
rect 46508 34066 46564 34076
rect 46844 34157 46900 34169
rect 46844 34105 46846 34157
rect 46898 34105 46900 34157
rect 46844 34020 46900 34105
rect 46844 33954 46900 33964
rect 47180 34130 47236 35084
rect 47292 34916 47348 35308
rect 47292 34914 47460 34916
rect 47292 34862 47294 34914
rect 47346 34862 47460 34914
rect 47292 34860 47460 34862
rect 47292 34850 47348 34860
rect 47404 34244 47460 34860
rect 47516 34914 47572 34926
rect 47516 34862 47518 34914
rect 47570 34862 47572 34914
rect 47516 34356 47572 34862
rect 47628 34914 47684 35644
rect 47628 34862 47630 34914
rect 47682 34862 47684 34914
rect 47628 34850 47684 34862
rect 47740 35690 47742 35742
rect 47794 35690 47796 35742
rect 47740 34916 47796 35690
rect 47852 35588 47908 35598
rect 47852 35494 47908 35532
rect 48132 35364 48188 35374
rect 48132 35138 48188 35308
rect 48132 35086 48134 35138
rect 48186 35086 48188 35138
rect 48132 35074 48188 35086
rect 47852 34916 47908 34926
rect 47740 34914 47908 34916
rect 47740 34862 47854 34914
rect 47906 34862 47908 34914
rect 47740 34860 47908 34862
rect 47852 34850 47908 34860
rect 47516 34300 47908 34356
rect 47404 34188 47684 34244
rect 47180 34078 47182 34130
rect 47234 34078 47236 34130
rect 47628 34174 47684 34188
rect 47628 34122 47630 34174
rect 47682 34122 47684 34174
rect 47628 34110 47684 34122
rect 47852 34132 47908 34300
rect 47852 34130 48132 34132
rect 47180 33684 47236 34078
rect 47852 34078 47854 34130
rect 47906 34078 48132 34130
rect 47852 34076 48132 34078
rect 47852 34066 47908 34076
rect 47516 34020 47572 34030
rect 47516 33926 47572 33964
rect 47236 33628 47460 33684
rect 47180 33618 47236 33628
rect 46396 33068 46544 33124
rect 45612 33012 45668 33022
rect 45612 32564 45668 32956
rect 46488 32676 46544 33068
rect 46488 32618 46544 32620
rect 45612 32498 45668 32508
rect 46284 32564 46340 32574
rect 46488 32566 46490 32618
rect 46542 32566 46544 32618
rect 46488 32554 46544 32566
rect 47292 32676 47348 32686
rect 47292 32618 47348 32620
rect 47292 32566 47294 32618
rect 47346 32566 47348 32618
rect 47292 32554 47348 32566
rect 45332 32452 45444 32462
rect 44940 32450 45444 32452
rect 44940 32398 45334 32450
rect 45386 32398 45444 32450
rect 44940 32396 45444 32398
rect 45332 32386 45444 32396
rect 45388 31778 45444 32386
rect 45388 31726 45390 31778
rect 45442 31726 45444 31778
rect 45052 31554 45108 31566
rect 45052 31502 45054 31554
rect 45106 31502 45108 31554
rect 44716 30828 44996 30884
rect 44492 30370 44548 30380
rect 43820 30146 43876 30156
rect 44828 30322 44884 30334
rect 44828 30270 44830 30322
rect 44882 30270 44884 30322
rect 44828 29988 44884 30270
rect 44940 30195 44996 30828
rect 44940 30143 44942 30195
rect 44994 30143 44996 30195
rect 44940 30131 44996 30143
rect 43708 29932 44884 29988
rect 45052 29876 45108 31502
rect 45220 30996 45276 31006
rect 45388 30996 45444 31726
rect 45220 30994 45444 30996
rect 45220 30942 45222 30994
rect 45274 30942 45390 30994
rect 45442 30942 45444 30994
rect 45220 30940 45444 30942
rect 45220 30930 45276 30940
rect 45164 30210 45220 30222
rect 45164 30158 45166 30210
rect 45218 30158 45220 30210
rect 45164 30100 45220 30158
rect 45164 30034 45220 30044
rect 45388 30212 45444 30940
rect 45836 32116 45892 32126
rect 45668 30436 45724 30446
rect 45668 30342 45724 30380
rect 44604 29820 45108 29876
rect 44604 29426 44660 29820
rect 44604 29374 44606 29426
rect 44658 29374 44660 29426
rect 44604 29362 44660 29374
rect 45052 29428 45108 29438
rect 44492 29316 44548 29326
rect 43372 28980 43428 28990
rect 43260 28644 43316 28654
rect 43260 28550 43316 28588
rect 43372 28642 43428 28924
rect 43708 28868 43764 28878
rect 43708 28774 43764 28812
rect 44324 28756 44380 28766
rect 44324 28662 44380 28700
rect 43372 28590 43374 28642
rect 43426 28590 43428 28642
rect 43372 28578 43428 28590
rect 43036 27794 43092 27804
rect 42588 26674 42644 26684
rect 43036 27636 43092 27646
rect 42532 26236 42644 26292
rect 42476 26198 42532 26236
rect 41580 24838 41582 24890
rect 41634 24838 41636 24890
rect 41580 24826 41636 24838
rect 41692 25844 41748 25854
rect 41580 24722 41636 24734
rect 41580 24670 41582 24722
rect 41634 24670 41636 24722
rect 41580 24500 41636 24670
rect 41580 24434 41636 24444
rect 41244 23871 41246 23923
rect 41298 23871 41300 23923
rect 40908 23266 41020 23278
rect 40908 23214 40966 23266
rect 41018 23214 41020 23266
rect 40908 23212 41020 23214
rect 40964 23202 41020 23212
rect 41244 23154 41300 23871
rect 41356 24332 41524 24388
rect 41356 23492 41412 24332
rect 41692 24276 41748 25788
rect 42252 24948 42308 24958
rect 42252 24766 42308 24892
rect 42252 24714 42254 24766
rect 42306 24714 42308 24766
rect 42140 24612 42196 24622
rect 42140 24518 42196 24556
rect 41580 24220 41748 24276
rect 41356 23426 41412 23436
rect 41468 23938 41524 23950
rect 41468 23886 41470 23938
rect 41522 23886 41524 23938
rect 41468 23156 41524 23886
rect 41244 23102 41246 23154
rect 41298 23102 41300 23154
rect 41244 23090 41300 23102
rect 41356 23154 41524 23156
rect 41356 23102 41470 23154
rect 41522 23102 41524 23154
rect 41356 23100 41524 23102
rect 41356 22596 41412 23100
rect 41468 23090 41524 23100
rect 41132 22540 41412 22596
rect 41132 22482 41188 22540
rect 41132 22430 41134 22482
rect 41186 22430 41188 22482
rect 41132 22418 41188 22430
rect 40796 22204 41076 22260
rect 40908 21812 40964 21822
rect 40684 21522 40740 21532
rect 40796 21586 40852 21598
rect 40796 21534 40798 21586
rect 40850 21534 40852 21586
rect 40572 20750 40574 20802
rect 40626 20750 40628 20802
rect 40348 20020 40404 20030
rect 40348 19926 40404 19964
rect 40236 19460 40292 19470
rect 40124 19458 40292 19460
rect 40124 19406 40238 19458
rect 40290 19406 40292 19458
rect 40124 19404 40292 19406
rect 39564 18450 39620 18462
rect 39564 18398 39566 18450
rect 39618 18398 39620 18450
rect 39564 18116 39620 18398
rect 39676 18450 39732 18462
rect 39676 18398 39678 18450
rect 39730 18398 39732 18450
rect 39676 18228 39732 18398
rect 39676 18162 39732 18172
rect 39844 18450 39900 18462
rect 39844 18398 39846 18450
rect 39898 18398 39900 18450
rect 39564 18050 39620 18060
rect 39844 18116 39900 18398
rect 39844 18050 39900 18060
rect 39340 17938 39396 17948
rect 40124 17668 40180 19404
rect 40236 19394 40292 19404
rect 40236 18340 40292 18350
rect 40236 18246 40292 18284
rect 40124 17602 40180 17612
rect 40236 18004 40292 18014
rect 40236 17118 40292 17948
rect 40180 17106 40292 17118
rect 40180 17054 40182 17106
rect 40234 17054 40292 17106
rect 40180 17052 40292 17054
rect 40180 17042 40236 17052
rect 39228 16436 39284 16828
rect 39228 16370 39284 16380
rect 39564 16996 39620 17006
rect 38556 15484 38724 15540
rect 38332 15372 38500 15428
rect 38332 15202 38388 15214
rect 38332 15150 38334 15202
rect 38386 15150 38388 15202
rect 38332 14868 38388 15150
rect 38332 14802 38388 14812
rect 38108 14590 38110 14642
rect 38162 14590 38164 14642
rect 38108 14578 38164 14590
rect 38332 14530 38388 14542
rect 37940 14474 37996 14486
rect 37940 14422 37942 14474
rect 37994 14422 37996 14474
rect 37940 14420 37996 14422
rect 37940 14354 37996 14364
rect 38332 14478 38334 14530
rect 38386 14478 38388 14530
rect 38332 14420 38388 14478
rect 38332 14354 38388 14364
rect 37716 14254 37718 14306
rect 37770 14254 37772 14306
rect 37716 14084 37772 14254
rect 37716 14018 37772 14028
rect 38444 13972 38500 15372
rect 38556 14980 38612 15484
rect 38556 14924 38724 14980
rect 38556 14474 38612 14486
rect 38556 14422 38558 14474
rect 38610 14422 38612 14474
rect 38556 14308 38612 14422
rect 38556 14242 38612 14252
rect 38332 13916 38500 13972
rect 37100 13010 37156 13020
rect 37212 13356 37380 13412
rect 37436 13774 37492 13786
rect 37436 13722 37438 13774
rect 37490 13722 37492 13774
rect 37212 12964 37268 13356
rect 37212 12898 37268 12908
rect 37324 13188 37380 13198
rect 37324 12962 37380 13132
rect 37324 12910 37326 12962
rect 37378 12910 37380 12962
rect 37324 12898 37380 12910
rect 37156 12740 37212 12750
rect 37436 12740 37492 13722
rect 38220 13746 38276 13758
rect 38052 13690 38108 13702
rect 37884 13636 37940 13646
rect 37772 13634 37940 13636
rect 37772 13582 37886 13634
rect 37938 13582 37940 13634
rect 37772 13580 37940 13582
rect 37772 13188 37828 13580
rect 37884 13570 37940 13580
rect 38052 13638 38054 13690
rect 38106 13638 38108 13690
rect 37772 13122 37828 13132
rect 37884 13300 37940 13310
rect 37660 13076 37716 13086
rect 37660 12982 37716 13020
rect 37884 12962 37940 13244
rect 38052 13076 38108 13638
rect 38220 13694 38222 13746
rect 38274 13694 38276 13746
rect 38220 13412 38276 13694
rect 38220 13346 38276 13356
rect 36876 12114 36932 12124
rect 36988 12628 37044 12638
rect 36988 12178 37044 12572
rect 36988 12126 36990 12178
rect 37042 12126 37044 12178
rect 37156 12234 37212 12684
rect 37324 12684 37492 12740
rect 37548 12918 37604 12930
rect 37548 12866 37550 12918
rect 37602 12866 37604 12918
rect 37884 12910 37886 12962
rect 37938 12910 37940 12962
rect 37884 12898 37940 12910
rect 37996 13020 38108 13076
rect 37324 12404 37380 12684
rect 37324 12338 37380 12348
rect 37436 12516 37492 12526
rect 37156 12182 37158 12234
rect 37210 12182 37212 12234
rect 37156 12170 37212 12182
rect 37324 12180 37380 12190
rect 36988 12114 37044 12126
rect 37324 12086 37380 12124
rect 37436 12178 37492 12460
rect 37436 12126 37438 12178
rect 37490 12126 37492 12178
rect 37436 12114 37492 12126
rect 37548 11956 37604 12866
rect 37996 12740 38052 13020
rect 37996 12516 38052 12684
rect 37772 12460 38052 12516
rect 37772 12190 37828 12460
rect 37716 12178 37828 12190
rect 37716 12126 37718 12178
rect 37770 12126 37828 12178
rect 37716 12124 37828 12126
rect 37716 12114 37772 12124
rect 38164 11956 38220 11966
rect 37548 11954 38220 11956
rect 37548 11902 38166 11954
rect 38218 11902 38220 11954
rect 37548 11900 38220 11902
rect 38164 11890 38220 11900
rect 36764 11778 36820 11788
rect 37436 11844 37492 11854
rect 37100 11620 37156 11630
rect 37100 11170 37156 11564
rect 37100 11118 37102 11170
rect 37154 11118 37156 11170
rect 36988 10836 37044 10846
rect 36652 10610 36708 10622
rect 36652 10558 36654 10610
rect 36706 10558 36708 10610
rect 36652 10388 36708 10558
rect 36988 10500 37044 10780
rect 37100 10612 37156 11118
rect 37100 10546 37156 10556
rect 37212 11396 37268 11406
rect 36988 10434 37044 10444
rect 36316 10386 36484 10388
rect 36316 10334 36318 10386
rect 36370 10334 36484 10386
rect 36316 10332 36484 10334
rect 36316 10322 36372 10332
rect 36204 9996 36372 10052
rect 36092 9940 36148 9950
rect 36316 9940 36372 9996
rect 36092 9938 36260 9940
rect 36092 9886 36094 9938
rect 36146 9886 36260 9938
rect 36092 9884 36260 9886
rect 36092 9874 36148 9884
rect 35980 9828 36036 9838
rect 35980 9759 35982 9772
rect 36034 9759 36036 9772
rect 35980 9734 36036 9759
rect 35868 9090 35924 9100
rect 35084 8878 35086 8930
rect 35138 8878 35140 8930
rect 35084 8484 35140 8878
rect 35308 9042 35364 9054
rect 35308 8990 35310 9042
rect 35362 8990 35364 9042
rect 35308 8932 35364 8990
rect 35532 9044 35588 9054
rect 35532 8950 35588 8988
rect 35308 8866 35364 8876
rect 35812 8820 35868 8830
rect 35644 8818 35868 8820
rect 35644 8766 35814 8818
rect 35866 8766 35868 8818
rect 35644 8764 35868 8766
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35084 8428 35252 8484
rect 33404 7746 33460 7756
rect 33740 7598 33796 8204
rect 33908 8204 34132 8260
rect 34188 8260 34244 8298
rect 33908 8148 33964 8204
rect 34188 8194 34244 8204
rect 33684 7586 33796 7598
rect 33684 7534 33686 7586
rect 33738 7534 33796 7586
rect 33684 7532 33796 7534
rect 33852 8092 33964 8148
rect 33684 7522 33740 7532
rect 31164 7364 31220 7374
rect 31052 7362 31220 7364
rect 31052 7310 31166 7362
rect 31218 7310 31220 7362
rect 31052 7308 31220 7310
rect 31332 7364 31388 7422
rect 32284 7422 32286 7474
rect 32338 7422 32340 7474
rect 31724 7364 31780 7374
rect 31332 7362 31780 7364
rect 31332 7310 31726 7362
rect 31778 7310 31780 7362
rect 31332 7308 31780 7310
rect 31052 6802 31108 7308
rect 31164 7298 31220 7308
rect 31724 7298 31780 7308
rect 31052 6750 31054 6802
rect 31106 6750 31108 6802
rect 31052 6738 31108 6750
rect 31276 7140 31332 7150
rect 30828 6524 31220 6580
rect 31164 5962 31220 6524
rect 30772 5908 30828 5918
rect 31164 5910 31166 5962
rect 31218 5910 31220 5962
rect 31164 5898 31220 5910
rect 31276 5908 31332 7084
rect 31612 6468 31668 6478
rect 32284 6468 32340 7422
rect 31500 5908 31556 5918
rect 31276 5906 31556 5908
rect 31276 5854 31502 5906
rect 31554 5854 31556 5906
rect 31276 5852 31556 5854
rect 30772 5814 30828 5852
rect 31500 5842 31556 5852
rect 30604 5796 30660 5806
rect 30156 5292 30268 5348
rect 30156 4574 30212 5292
rect 30268 5282 30324 5292
rect 30492 5794 30660 5796
rect 30492 5742 30606 5794
rect 30658 5742 30660 5794
rect 30492 5740 30660 5742
rect 30268 5124 30324 5134
rect 30492 5124 30548 5740
rect 30604 5730 30660 5740
rect 30268 5122 30548 5124
rect 30268 5070 30270 5122
rect 30322 5070 30548 5122
rect 30268 5068 30548 5070
rect 31388 5460 31444 5470
rect 30268 5058 30324 5068
rect 31388 4900 31444 5404
rect 31612 4900 31668 6412
rect 32060 6412 32340 6468
rect 32396 7474 32452 7486
rect 32396 7422 32398 7474
rect 32450 7422 32452 7474
rect 31892 5850 31948 5862
rect 31724 5796 31780 5806
rect 31724 5702 31780 5740
rect 31892 5798 31894 5850
rect 31946 5798 31948 5850
rect 31892 5460 31948 5798
rect 31892 5394 31948 5404
rect 32060 5124 32116 6412
rect 32396 6142 32452 7422
rect 33180 7474 33236 7486
rect 33180 7422 33182 7474
rect 33234 7422 33236 7474
rect 32340 6130 32452 6142
rect 32340 6078 32342 6130
rect 32394 6078 32452 6130
rect 32340 6076 32452 6078
rect 32956 6578 33012 6590
rect 32956 6526 32958 6578
rect 33010 6526 33012 6578
rect 32956 6132 33012 6526
rect 33180 6580 33236 7422
rect 33404 7474 33460 7486
rect 33404 7422 33406 7474
rect 33458 7422 33460 7474
rect 33404 7364 33460 7422
rect 33404 7298 33460 7308
rect 33180 6514 33236 6524
rect 33516 6580 33572 6590
rect 33516 6486 33572 6524
rect 32340 6066 32396 6076
rect 32956 6066 33012 6076
rect 33338 6468 33394 6478
rect 32508 6020 32564 6030
rect 32508 5906 32564 5964
rect 33338 5956 33394 6412
rect 33068 5908 33124 5918
rect 32508 5854 32510 5906
rect 32562 5854 32564 5906
rect 32508 5842 32564 5854
rect 32676 5906 33124 5908
rect 32676 5854 33070 5906
rect 33122 5854 33124 5906
rect 32676 5852 33124 5854
rect 32676 5346 32732 5852
rect 33068 5842 33124 5852
rect 33180 5906 33236 5918
rect 33180 5854 33182 5906
rect 33234 5854 33236 5906
rect 33338 5904 33340 5956
rect 33392 5904 33394 5956
rect 33338 5892 33394 5904
rect 33740 5908 33796 5918
rect 32676 5294 32678 5346
rect 32730 5294 32732 5346
rect 32676 5282 32732 5294
rect 32172 5236 32228 5246
rect 32172 5142 32228 5180
rect 32508 5236 32564 5246
rect 32060 5058 32116 5068
rect 32508 5122 32564 5180
rect 32508 5070 32510 5122
rect 32562 5070 32564 5122
rect 32508 5058 32564 5070
rect 33180 5124 33236 5854
rect 33852 5908 33908 8092
rect 34020 8036 34076 8046
rect 34020 7942 34076 7980
rect 34188 7512 34244 7524
rect 34188 7460 34190 7512
rect 34242 7460 34244 7512
rect 34188 6804 34244 7460
rect 34188 6738 34244 6748
rect 34076 6132 34132 6142
rect 33964 5908 34020 5918
rect 33852 5852 33964 5908
rect 33740 5794 33796 5852
rect 33964 5842 34020 5852
rect 33740 5742 33742 5794
rect 33794 5742 33796 5794
rect 33740 5730 33796 5742
rect 33908 5684 33964 5694
rect 33740 5572 33796 5582
rect 33348 5348 33404 5358
rect 33348 5236 33404 5292
rect 33180 5058 33236 5068
rect 33292 5234 33404 5236
rect 33292 5182 33350 5234
rect 33402 5182 33404 5234
rect 33292 5170 33404 5182
rect 30100 4562 30212 4574
rect 30100 4510 30102 4562
rect 30154 4510 30212 4562
rect 30100 4508 30212 4510
rect 31164 4844 31444 4900
rect 31578 4844 31668 4900
rect 31724 5012 31780 5022
rect 30100 4498 30156 4508
rect 30772 4226 30828 4238
rect 30772 4174 30774 4226
rect 30826 4174 30828 4226
rect 30772 3780 30828 4174
rect 31164 4226 31220 4844
rect 31578 4376 31634 4844
rect 31578 4324 31580 4376
rect 31632 4324 31634 4376
rect 31578 4312 31634 4324
rect 31724 4338 31780 4956
rect 32732 4900 32788 4910
rect 32396 4788 32452 4798
rect 31724 4286 31726 4338
rect 31778 4286 31780 4338
rect 31724 4274 31780 4286
rect 31836 4340 31892 4350
rect 31836 4338 32284 4340
rect 31836 4286 31838 4338
rect 31890 4286 32284 4338
rect 31836 4284 32284 4286
rect 31836 4274 31892 4284
rect 31164 4174 31166 4226
rect 31218 4174 31220 4226
rect 31164 4162 31220 4174
rect 32228 4170 32284 4284
rect 32228 4118 32230 4170
rect 32282 4118 32284 4170
rect 32228 4106 32284 4118
rect 32396 4338 32452 4732
rect 32396 4286 32398 4338
rect 32450 4286 32452 4338
rect 30772 3714 30828 3724
rect 31500 3892 31556 3902
rect 29596 3614 29598 3666
rect 29650 3614 29652 3666
rect 29596 3602 29652 3614
rect 31500 3666 31556 3836
rect 32396 3892 32452 4286
rect 32396 3826 32452 3836
rect 32732 3790 32788 4844
rect 33292 4574 33348 5170
rect 33628 5122 33684 5134
rect 33628 5070 33630 5122
rect 33682 5070 33684 5122
rect 33628 4788 33684 5070
rect 33740 5122 33796 5516
rect 33740 5070 33742 5122
rect 33794 5070 33796 5122
rect 33740 5058 33796 5070
rect 33908 5122 33964 5628
rect 33908 5070 33910 5122
rect 33962 5070 33964 5122
rect 33908 5058 33964 5070
rect 33628 4722 33684 4732
rect 33236 4564 33348 4574
rect 33964 4564 34020 4574
rect 33236 4562 33684 4564
rect 33236 4510 33238 4562
rect 33290 4510 33684 4562
rect 33236 4508 33684 4510
rect 32732 3780 32844 3790
rect 32732 3724 32788 3780
rect 31500 3614 31502 3666
rect 31554 3614 31556 3666
rect 31500 3602 31556 3614
rect 32340 3668 32396 3678
rect 32340 3574 32396 3612
rect 32788 3666 32844 3724
rect 32788 3614 32790 3666
rect 32842 3614 32844 3666
rect 32788 3602 32844 3614
rect 33236 3668 33292 4508
rect 33628 4338 33684 4508
rect 33628 4286 33630 4338
rect 33682 4286 33684 4338
rect 33628 4274 33684 4286
rect 33236 3574 33292 3612
rect 33628 3556 33684 3566
rect 33628 3469 33630 3500
rect 33682 3469 33684 3500
rect 33628 3457 33684 3469
rect 33964 3517 34020 4508
rect 34076 4004 34132 6076
rect 34300 5694 34356 8428
rect 34412 8260 34468 8270
rect 34692 8260 34748 8270
rect 34412 8258 34580 8260
rect 34412 8206 34414 8258
rect 34466 8206 34580 8258
rect 34412 8204 34580 8206
rect 34412 8194 34468 8204
rect 34412 8036 34468 8046
rect 34412 7476 34468 7980
rect 34524 7812 34580 8204
rect 34692 8166 34748 8204
rect 35196 8148 35252 8428
rect 35308 8372 35364 8382
rect 35308 8278 35364 8316
rect 35644 8258 35700 8764
rect 35812 8754 35868 8764
rect 35420 8214 35476 8226
rect 35420 8162 35422 8214
rect 35474 8162 35476 8214
rect 35644 8206 35646 8258
rect 35698 8206 35700 8258
rect 35644 8194 35700 8206
rect 35980 8260 36036 8270
rect 35980 8166 36036 8204
rect 36204 8260 36260 9884
rect 36316 9874 36372 9884
rect 36428 9716 36484 10332
rect 36652 10322 36708 10332
rect 37212 9828 37268 11340
rect 37436 11396 37492 11788
rect 38332 11732 38388 13916
rect 38668 13870 38724 14924
rect 39228 14868 39284 14878
rect 39228 14642 39284 14812
rect 39228 14590 39230 14642
rect 39282 14590 39284 14642
rect 39228 14578 39284 14590
rect 39452 14532 39508 14542
rect 39060 14476 39116 14486
rect 38892 14474 39116 14476
rect 38892 14422 39062 14474
rect 39114 14422 39116 14474
rect 39452 14438 39508 14476
rect 38892 14420 39116 14422
rect 38668 13858 38780 13870
rect 38668 13806 38726 13858
rect 38778 13806 38780 13858
rect 38668 13804 38780 13806
rect 38724 13794 38780 13804
rect 38444 13748 38500 13758
rect 38444 13746 38612 13748
rect 38444 13694 38446 13746
rect 38498 13694 38612 13746
rect 38444 13692 38612 13694
rect 38444 13682 38500 13692
rect 38444 12740 38500 12750
rect 38444 12178 38500 12684
rect 38556 12516 38612 13692
rect 38892 13524 38948 14420
rect 39060 14410 39116 14420
rect 38892 13458 38948 13468
rect 39284 13636 39340 13646
rect 39564 13636 39620 16940
rect 40012 16884 40068 16894
rect 40012 16100 40068 16828
rect 40012 16044 40180 16100
rect 39676 14474 39732 14486
rect 39676 14422 39678 14474
rect 39730 14422 39732 14474
rect 39676 14308 39732 14422
rect 39676 14242 39732 14252
rect 39956 13972 40012 13982
rect 39956 13878 40012 13916
rect 39284 13634 39620 13636
rect 39284 13582 39286 13634
rect 39338 13582 39620 13634
rect 39284 13580 39620 13582
rect 39284 13300 39340 13580
rect 39284 13234 39340 13244
rect 38668 13076 38724 13086
rect 38668 12982 38724 13020
rect 38556 12450 38612 12460
rect 39396 12740 39452 12750
rect 38444 12126 38446 12178
rect 38498 12126 38500 12178
rect 38444 12114 38500 12126
rect 38556 12292 38612 12302
rect 38556 12068 38612 12236
rect 38892 12180 38948 12190
rect 38556 12002 38612 12012
rect 38724 12122 38780 12134
rect 38724 12070 38726 12122
rect 38778 12070 38780 12122
rect 38892 12086 38948 12124
rect 38332 11666 38388 11676
rect 38724 11508 38780 12070
rect 39396 12068 39452 12684
rect 39956 12180 40012 12190
rect 39956 12086 40012 12124
rect 39396 12066 39508 12068
rect 39396 12014 39398 12066
rect 39450 12014 39508 12066
rect 39396 12002 39508 12014
rect 39004 11732 39060 11742
rect 38724 11452 38836 11508
rect 37548 11396 37604 11406
rect 37436 11394 37548 11396
rect 37436 11342 37438 11394
rect 37490 11342 37548 11394
rect 37436 11340 37548 11342
rect 37436 11330 37492 11340
rect 37548 11302 37604 11340
rect 38220 11394 38276 11406
rect 38220 11342 38222 11394
rect 38274 11342 38276 11394
rect 37884 11172 37940 11182
rect 38220 11172 38276 11342
rect 37884 11170 38276 11172
rect 37884 11118 37886 11170
rect 37938 11118 38276 11170
rect 37884 11116 38276 11118
rect 38556 11170 38612 11182
rect 38556 11118 38558 11170
rect 38610 11118 38612 11170
rect 37884 11106 37940 11116
rect 37324 10612 37380 10622
rect 37324 10518 37380 10556
rect 37996 10612 38052 11116
rect 38556 10948 38612 11118
rect 38556 10882 38612 10892
rect 37660 10388 37716 10398
rect 36316 9660 36484 9716
rect 36988 9772 37268 9828
rect 37324 10386 37716 10388
rect 37324 10334 37662 10386
rect 37714 10334 37716 10386
rect 37324 10332 37716 10334
rect 36316 8708 36372 9660
rect 36484 9156 36540 9166
rect 36484 9062 36540 9100
rect 36652 9042 36708 9054
rect 36652 8990 36654 9042
rect 36706 8990 36708 9042
rect 36316 8652 36484 8708
rect 36204 8194 36260 8204
rect 35420 8148 35476 8162
rect 35196 8092 35476 8148
rect 36316 8036 36372 8046
rect 35532 8034 36372 8036
rect 35532 7982 36318 8034
rect 36370 7982 36372 8034
rect 35532 7980 36372 7982
rect 34524 7756 34804 7812
rect 34748 7586 34804 7756
rect 34748 7534 34750 7586
rect 34802 7534 34804 7586
rect 34748 7522 34804 7534
rect 34916 7700 34972 7710
rect 34916 7530 34972 7644
rect 34524 7476 34580 7486
rect 34412 7474 34580 7476
rect 34412 7422 34526 7474
rect 34578 7422 34580 7474
rect 34916 7478 34918 7530
rect 34970 7478 34972 7530
rect 34916 7466 34972 7478
rect 35420 7476 35476 7486
rect 34412 7420 34580 7422
rect 34524 7410 34580 7420
rect 35420 7382 35476 7420
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35420 6804 35476 6814
rect 35532 6804 35588 7980
rect 36316 7970 36372 7980
rect 36428 8036 36484 8652
rect 36428 7812 36484 7980
rect 36204 7756 36484 7812
rect 36204 7588 36260 7756
rect 36652 7700 36708 8990
rect 36204 7522 36260 7532
rect 36428 7644 36708 7700
rect 36988 7700 37044 9772
rect 37156 9602 37212 9614
rect 37156 9550 37158 9602
rect 37210 9550 37212 9602
rect 37156 9156 37212 9550
rect 37156 8370 37212 9100
rect 37156 8318 37158 8370
rect 37210 8318 37212 8370
rect 37156 8306 37212 8318
rect 36316 7476 36372 7486
rect 36428 7476 36484 7644
rect 36988 7634 37044 7644
rect 36372 7420 36484 7476
rect 36204 7362 36260 7374
rect 36204 7310 36206 7362
rect 36258 7310 36260 7362
rect 36204 7028 36260 7310
rect 36204 6962 36260 6972
rect 35420 6802 35588 6804
rect 35420 6750 35422 6802
rect 35474 6750 35588 6802
rect 35420 6748 35588 6750
rect 35420 6738 35476 6748
rect 36204 6692 36260 6702
rect 36316 6692 36372 7420
rect 37324 7140 37380 10332
rect 37660 10322 37716 10332
rect 37604 9940 37660 9950
rect 37604 9846 37660 9884
rect 37772 9828 37828 9838
rect 37996 9828 38052 10556
rect 38668 10612 38724 10622
rect 38668 10518 38724 10556
rect 38332 10388 38388 10398
rect 38332 10294 38388 10332
rect 38780 10388 38836 11452
rect 38892 11396 38948 11406
rect 38892 11302 38948 11340
rect 38780 10322 38836 10332
rect 39004 10834 39060 11676
rect 39228 11172 39284 11182
rect 39228 11078 39284 11116
rect 39004 10782 39006 10834
rect 39058 10782 39060 10834
rect 39004 10164 39060 10782
rect 39452 10836 39508 12002
rect 40124 11518 40180 16044
rect 40348 15988 40404 15998
rect 40348 15894 40404 15932
rect 40236 15202 40292 15214
rect 40236 15150 40238 15202
rect 40290 15150 40292 15202
rect 40236 15148 40292 15150
rect 40236 15092 40516 15148
rect 40292 14532 40348 14542
rect 40292 14362 40348 14476
rect 40292 14310 40294 14362
rect 40346 14310 40348 14362
rect 40292 14298 40348 14310
rect 40460 14530 40516 15092
rect 40460 14478 40462 14530
rect 40514 14478 40516 14530
rect 40460 14308 40516 14478
rect 40460 14242 40516 14252
rect 40404 13636 40460 13646
rect 40572 13636 40628 20750
rect 40796 20692 40852 21534
rect 40908 21026 40964 21756
rect 40908 20974 40910 21026
rect 40962 20974 40964 21026
rect 40908 20962 40964 20974
rect 41020 20916 41076 22204
rect 41468 21924 41524 21934
rect 41468 21140 41524 21868
rect 41580 21812 41636 24220
rect 42084 24052 42140 24062
rect 42084 23604 42140 23996
rect 42084 23538 42140 23548
rect 42140 23154 42196 23166
rect 42140 23102 42142 23154
rect 42194 23102 42196 23154
rect 42028 22370 42084 22382
rect 42028 22318 42030 22370
rect 42082 22318 42084 22370
rect 41580 21746 41636 21756
rect 41692 22146 41748 22158
rect 41692 22094 41694 22146
rect 41746 22094 41748 22146
rect 41580 21588 41636 21598
rect 41692 21588 41748 22094
rect 42028 21812 42084 22318
rect 42140 22372 42196 23102
rect 42252 22484 42308 24714
rect 42476 24836 42532 24846
rect 42476 24722 42532 24780
rect 42476 24670 42478 24722
rect 42530 24670 42532 24722
rect 42476 24658 42532 24670
rect 42588 24724 42644 26236
rect 43036 24724 43092 27580
rect 43148 27074 43204 27086
rect 43148 27022 43150 27074
rect 43202 27022 43204 27074
rect 43820 27074 43876 27086
rect 43148 26964 43204 27022
rect 43484 27018 43540 27030
rect 43484 26966 43486 27018
rect 43538 26966 43540 27018
rect 43148 26898 43204 26908
rect 43372 26906 43428 26918
rect 43372 26854 43374 26906
rect 43426 26854 43428 26906
rect 43260 26178 43316 26190
rect 43260 26126 43262 26178
rect 43314 26126 43316 26178
rect 43260 25732 43316 26126
rect 43372 25956 43428 26854
rect 43484 26292 43540 26966
rect 43820 27022 43822 27074
rect 43874 27022 43876 27074
rect 43820 26852 43876 27022
rect 43820 26786 43876 26796
rect 44380 26964 44436 26974
rect 43484 26226 43540 26236
rect 43372 25900 43764 25956
rect 43260 25666 43316 25676
rect 43708 25506 43764 25900
rect 44044 25732 44100 25742
rect 44044 25638 44100 25676
rect 43708 25454 43710 25506
rect 43762 25454 43764 25506
rect 43708 25442 43764 25454
rect 43372 25394 43428 25406
rect 43372 25342 43374 25394
rect 43426 25342 43428 25394
rect 43260 24948 43316 24958
rect 43036 24668 43204 24724
rect 42588 24062 42644 24668
rect 42980 24500 43036 24510
rect 42980 24406 43036 24444
rect 43148 24500 43204 24668
rect 43260 24722 43316 24892
rect 43260 24670 43262 24722
rect 43314 24670 43316 24722
rect 43260 24658 43316 24670
rect 43372 24836 43428 25342
rect 44380 24958 44436 26908
rect 44324 24946 44436 24958
rect 44324 24894 44326 24946
rect 44378 24894 44436 24946
rect 44324 24892 44436 24894
rect 44324 24882 44380 24892
rect 43372 24722 43428 24780
rect 43372 24670 43374 24722
rect 43426 24670 43428 24722
rect 43372 24658 43428 24670
rect 43876 24724 43932 24734
rect 43876 24630 43932 24668
rect 43148 24434 43204 24444
rect 42532 24052 42644 24062
rect 42588 23996 42644 24052
rect 42532 23958 42644 23996
rect 42476 23716 42532 23726
rect 42252 22418 42308 22428
rect 42364 23268 42420 23278
rect 42140 22306 42196 22316
rect 42364 22370 42420 23212
rect 42364 22318 42366 22370
rect 42418 22318 42420 22370
rect 42364 21924 42420 22318
rect 42364 21858 42420 21868
rect 42476 22596 42532 23660
rect 42588 23044 42644 23958
rect 42588 22978 42644 22988
rect 42700 24220 43316 24276
rect 41580 21586 41748 21588
rect 41580 21534 41582 21586
rect 41634 21534 41748 21586
rect 41580 21532 41748 21534
rect 41804 21756 42084 21812
rect 42476 21812 42532 22540
rect 42700 22372 42756 24220
rect 42924 24052 42980 24062
rect 42700 22306 42756 22316
rect 42812 24050 42980 24052
rect 42812 23998 42926 24050
rect 42978 23998 42980 24050
rect 42812 23996 42980 23998
rect 42812 22331 42868 23996
rect 42924 23986 42980 23996
rect 43260 23938 43316 24220
rect 43596 23940 43652 23950
rect 43036 23894 43092 23906
rect 43036 23842 43038 23894
rect 43090 23842 43092 23894
rect 43260 23886 43262 23938
rect 43314 23886 43316 23938
rect 43260 23874 43316 23886
rect 43372 23938 43652 23940
rect 43372 23886 43598 23938
rect 43650 23886 43652 23938
rect 43372 23884 43652 23886
rect 43036 23716 43092 23842
rect 43036 23650 43092 23660
rect 43372 23380 43428 23884
rect 43596 23874 43652 23884
rect 42812 22279 42814 22331
rect 42866 22279 42868 22331
rect 42812 22267 42868 22279
rect 42924 23324 43428 23380
rect 43932 23714 43988 23726
rect 43932 23662 43934 23714
rect 43986 23662 43988 23714
rect 42924 22202 42980 23324
rect 43932 23156 43988 23662
rect 44044 23156 44100 23166
rect 43932 23154 44100 23156
rect 43932 23102 44046 23154
rect 44098 23102 44100 23154
rect 43932 23100 44100 23102
rect 44044 23090 44100 23100
rect 43036 22484 43092 22494
rect 43652 22484 43708 22494
rect 43092 22482 43708 22484
rect 43092 22430 43654 22482
rect 43706 22430 43708 22482
rect 43092 22428 43708 22430
rect 43036 22370 43092 22428
rect 43652 22418 43708 22428
rect 43932 22484 43988 22494
rect 43036 22318 43038 22370
rect 43090 22318 43092 22370
rect 43036 22306 43092 22318
rect 43932 22370 43988 22428
rect 43932 22318 43934 22370
rect 43986 22318 43988 22370
rect 43932 22306 43988 22318
rect 44044 22372 44100 22382
rect 44044 22278 44100 22316
rect 42924 22150 42926 22202
rect 42978 22150 42980 22202
rect 42924 22138 42980 22150
rect 43260 22260 43316 22270
rect 42476 21756 42756 21812
rect 41580 21522 41636 21532
rect 41804 21252 41860 21756
rect 41804 21196 42084 21252
rect 41020 20850 41076 20860
rect 41132 21084 41860 21140
rect 40796 20626 40852 20636
rect 41132 20188 41188 21084
rect 41524 20916 41580 20926
rect 41524 20822 41580 20860
rect 41804 20802 41860 21084
rect 41804 20750 41806 20802
rect 41858 20750 41860 20802
rect 41804 20738 41860 20750
rect 42028 20634 42084 21196
rect 42700 21140 42756 21756
rect 42476 21084 43148 21140
rect 42252 21028 42308 21038
rect 42252 20763 42308 20972
rect 42252 20711 42254 20763
rect 42306 20711 42308 20763
rect 42476 20802 42532 21084
rect 43092 21026 43148 21084
rect 43092 20974 43094 21026
rect 43146 20974 43148 21026
rect 43092 20962 43148 20974
rect 42476 20750 42478 20802
rect 42530 20750 42532 20802
rect 42476 20738 42532 20750
rect 42252 20699 42308 20711
rect 42028 20582 42030 20634
rect 42082 20582 42084 20634
rect 42028 20570 42084 20582
rect 40684 20132 41188 20188
rect 40684 13972 40740 20132
rect 40908 20020 40964 20030
rect 40796 18450 40852 18462
rect 40796 18398 40798 18450
rect 40850 18398 40852 18450
rect 40796 17220 40852 18398
rect 40908 18228 40964 19964
rect 41132 19906 41188 19918
rect 43036 19908 43092 19918
rect 41132 19854 41134 19906
rect 41186 19854 41188 19906
rect 41020 18452 41076 18462
rect 41020 18358 41076 18396
rect 40908 18172 41076 18228
rect 40908 18004 40964 18014
rect 40908 17778 40964 17948
rect 40908 17726 40910 17778
rect 40962 17726 40964 17778
rect 40908 17556 40964 17726
rect 40908 17490 40964 17500
rect 40796 17154 40852 17164
rect 40908 16909 40964 16922
rect 40908 16884 40910 16909
rect 40962 16884 40964 16909
rect 40908 16818 40964 16828
rect 40908 16660 40964 16670
rect 40908 15540 40964 16604
rect 40908 15314 40964 15484
rect 40908 15262 40910 15314
rect 40962 15262 40964 15314
rect 40908 15250 40964 15262
rect 41020 15148 41076 18172
rect 41132 17780 41188 19854
rect 42924 19906 43092 19908
rect 42924 19854 43038 19906
rect 43090 19854 43092 19906
rect 42924 19852 43092 19854
rect 42786 19684 42842 19694
rect 42786 19201 42842 19628
rect 41804 19178 41860 19190
rect 41804 19126 41806 19178
rect 41858 19126 41860 19178
rect 41804 18676 41860 19126
rect 41804 18610 41860 18620
rect 42140 19178 42196 19190
rect 42140 19126 42142 19178
rect 42194 19126 42196 19178
rect 41300 18564 41356 18574
rect 41300 18450 41356 18508
rect 41300 18398 41302 18450
rect 41354 18398 41356 18450
rect 41300 18386 41356 18398
rect 41692 18450 41748 18462
rect 41692 18398 41694 18450
rect 41746 18398 41748 18450
rect 41692 18340 41748 18398
rect 41692 18274 41748 18284
rect 42028 18450 42084 18462
rect 42028 18398 42030 18450
rect 42082 18398 42084 18450
rect 42028 18116 42084 18398
rect 42140 18282 42196 19126
rect 42588 19178 42644 19190
rect 42588 19126 42590 19178
rect 42642 19126 42644 19178
rect 42786 19149 42788 19201
rect 42840 19149 42842 19201
rect 42786 19137 42842 19149
rect 42588 18900 42644 19126
rect 42924 19122 42980 19852
rect 43036 19842 43092 19852
rect 42924 19070 42926 19122
rect 42978 19070 42980 19122
rect 42924 19058 42980 19070
rect 42588 18844 42980 18900
rect 42140 18230 42142 18282
rect 42194 18230 42196 18282
rect 42364 18450 42420 18462
rect 42364 18398 42366 18450
rect 42418 18398 42420 18450
rect 42364 18340 42420 18398
rect 42364 18274 42420 18284
rect 42588 18450 42644 18462
rect 42588 18398 42590 18450
rect 42642 18398 42644 18450
rect 42140 18218 42196 18230
rect 42588 18116 42644 18398
rect 42028 18060 42644 18116
rect 42700 18452 42756 18462
rect 42028 17890 42084 18060
rect 42028 17838 42030 17890
rect 42082 17838 42084 17890
rect 42028 17826 42084 17838
rect 41132 17714 41188 17724
rect 41634 17780 41690 17790
rect 41356 17666 41412 17678
rect 41356 17614 41358 17666
rect 41410 17614 41412 17666
rect 41356 17332 41412 17614
rect 41356 17266 41412 17276
rect 41468 17668 41524 17678
rect 41356 16042 41412 16054
rect 40684 13906 40740 13916
rect 40796 15092 41076 15148
rect 41132 15988 41188 15998
rect 41132 15316 41188 15932
rect 41356 15990 41358 16042
rect 41410 15990 41412 16042
rect 41356 15428 41412 15990
rect 41356 15362 41412 15372
rect 40404 13634 40628 13636
rect 40404 13582 40406 13634
rect 40458 13582 40628 13634
rect 40404 13580 40628 13582
rect 40404 13570 40516 13580
rect 40236 12292 40292 12302
rect 40236 12178 40292 12236
rect 40236 12126 40238 12178
rect 40290 12126 40292 12178
rect 40236 12114 40292 12126
rect 40348 12178 40404 12190
rect 40348 12126 40350 12178
rect 40402 12126 40404 12178
rect 40348 11956 40404 12126
rect 40348 11890 40404 11900
rect 40068 11506 40180 11518
rect 40068 11454 40070 11506
rect 40122 11454 40180 11506
rect 40068 11452 40180 11454
rect 40348 11732 40404 11742
rect 40068 11442 40124 11452
rect 40236 11396 40292 11406
rect 39620 10836 39676 10846
rect 39452 10834 39676 10836
rect 39452 10782 39622 10834
rect 39674 10782 39676 10834
rect 39452 10780 39676 10782
rect 39620 10770 39676 10780
rect 40236 10610 40292 11340
rect 40236 10558 40238 10610
rect 40290 10558 40292 10610
rect 38780 10108 39060 10164
rect 39956 10386 40012 10398
rect 39956 10334 39958 10386
rect 40010 10334 40012 10386
rect 38668 10052 38724 10062
rect 38556 9994 38612 10006
rect 38108 9940 38164 9950
rect 38108 9846 38164 9884
rect 38556 9942 38558 9994
rect 38610 9942 38612 9994
rect 37772 9826 38052 9828
rect 37772 9774 37774 9826
rect 37826 9774 38052 9826
rect 37772 9772 38052 9774
rect 37772 9762 37828 9772
rect 37436 8932 37492 8942
rect 37436 8930 37716 8932
rect 37436 8878 37438 8930
rect 37490 8878 37716 8930
rect 37436 8876 37716 8878
rect 37436 8866 37492 8876
rect 37660 8484 37716 8876
rect 38556 8708 38612 9942
rect 38668 9826 38724 9996
rect 38668 9774 38670 9826
rect 38722 9774 38724 9826
rect 38668 9762 38724 9774
rect 38276 8652 38612 8708
rect 37660 8428 38164 8484
rect 37548 8372 37604 8382
rect 37548 8220 37604 8316
rect 38108 8370 38164 8428
rect 38108 8318 38110 8370
rect 38162 8318 38164 8370
rect 38108 8306 38164 8318
rect 38276 8314 38332 8652
rect 38780 8596 38836 10108
rect 39732 10052 39788 10062
rect 39732 9958 39788 9996
rect 39004 9826 39060 9838
rect 39004 9774 39006 9826
rect 39058 9774 39060 9826
rect 39004 9716 39060 9774
rect 39004 9650 39060 9660
rect 39228 9828 39284 9838
rect 39228 9156 39284 9772
rect 39452 9828 39508 9838
rect 39452 9734 39508 9772
rect 39956 9828 40012 10334
rect 40236 9940 40292 10558
rect 40348 10610 40404 11676
rect 40348 10558 40350 10610
rect 40402 10558 40404 10610
rect 40348 10546 40404 10558
rect 39956 9762 40012 9772
rect 40124 9884 40236 9940
rect 39340 9156 39396 9166
rect 39228 9154 39396 9156
rect 39228 9102 39342 9154
rect 39394 9102 39396 9154
rect 39228 9100 39396 9102
rect 39340 9090 39396 9100
rect 39452 9156 39508 9166
rect 37548 8168 37550 8220
rect 37602 8168 37604 8220
rect 37548 8156 37604 8168
rect 37884 8260 37940 8270
rect 38276 8262 38278 8314
rect 38330 8262 38332 8314
rect 38276 8250 38332 8262
rect 38556 8540 38836 8596
rect 37884 8166 37940 8204
rect 38108 8036 38164 8046
rect 37996 7924 38052 7934
rect 36204 6690 36372 6692
rect 36204 6638 36206 6690
rect 36258 6638 36372 6690
rect 36204 6636 36372 6638
rect 36204 6626 36260 6636
rect 35084 6132 35140 6142
rect 34244 5684 34356 5694
rect 34076 3938 34132 3948
rect 34188 5682 34356 5684
rect 34188 5630 34246 5682
rect 34298 5630 34356 5682
rect 34188 5628 34356 5630
rect 34524 5906 34580 5918
rect 34524 5854 34526 5906
rect 34578 5854 34580 5906
rect 34188 5618 34300 5628
rect 33964 3465 33966 3517
rect 34018 3465 34020 3517
rect 34188 3556 34244 5618
rect 34524 5460 34580 5854
rect 34748 5908 34804 5918
rect 34748 5814 34804 5852
rect 34972 5906 35028 5918
rect 34972 5854 34974 5906
rect 35026 5854 35028 5906
rect 34972 5684 35028 5854
rect 35084 5906 35140 6076
rect 35084 5854 35086 5906
rect 35138 5854 35140 5906
rect 35084 5842 35140 5854
rect 35196 5908 35252 5918
rect 35196 5684 35252 5852
rect 36204 5908 36260 5918
rect 36204 5814 36260 5852
rect 35868 5796 35924 5806
rect 35868 5702 35924 5740
rect 34972 5618 35028 5628
rect 35084 5628 35252 5684
rect 35364 5684 35420 5694
rect 36204 5684 36260 5694
rect 35364 5682 35700 5684
rect 35364 5630 35366 5682
rect 35418 5630 35700 5682
rect 35364 5628 35700 5630
rect 34300 5404 34916 5460
rect 34300 5346 34356 5404
rect 34300 5294 34302 5346
rect 34354 5294 34356 5346
rect 34300 5282 34356 5294
rect 34748 5290 34804 5302
rect 34748 5238 34750 5290
rect 34802 5238 34804 5290
rect 34636 5124 34692 5134
rect 34412 4226 34468 4238
rect 34412 4174 34414 4226
rect 34466 4174 34468 4226
rect 34412 3668 34468 4174
rect 34636 3892 34692 5068
rect 34748 4564 34804 5238
rect 34860 5122 34916 5404
rect 35084 5348 35140 5628
rect 35364 5618 35420 5628
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35196 5348 35252 5358
rect 35084 5292 35196 5348
rect 34860 5070 34862 5122
rect 34914 5070 34916 5122
rect 34860 5058 34916 5070
rect 35196 5122 35252 5292
rect 35196 5070 35198 5122
rect 35250 5070 35252 5122
rect 35196 5058 35252 5070
rect 35532 5290 35588 5302
rect 35532 5238 35534 5290
rect 35586 5238 35588 5290
rect 35532 5124 35588 5238
rect 35532 5058 35588 5068
rect 35644 5122 35700 5628
rect 35644 5070 35646 5122
rect 35698 5070 35700 5122
rect 35644 5058 35700 5070
rect 35756 5124 35812 5134
rect 34748 4498 34804 4508
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 34636 3836 34804 3892
rect 35196 3882 35460 3892
rect 34636 3668 34692 3678
rect 34412 3666 34692 3668
rect 34412 3614 34638 3666
rect 34690 3614 34692 3666
rect 34412 3612 34692 3614
rect 34636 3602 34692 3612
rect 34188 3500 34300 3556
rect 33964 3453 34020 3465
rect 34244 3498 34300 3500
rect 34244 3446 34246 3498
rect 34298 3446 34300 3498
rect 34244 3434 34300 3446
rect 34610 3514 34666 3526
rect 34610 3462 34612 3514
rect 34664 3462 34666 3514
rect 34610 3444 34666 3462
rect 34748 3444 34804 3836
rect 35756 3780 35812 5068
rect 35476 3724 35812 3780
rect 35980 5122 36036 5134
rect 35980 5070 35982 5122
rect 36034 5070 36036 5122
rect 35980 3780 36036 5070
rect 36204 4452 36260 5628
rect 36316 5460 36372 6636
rect 36988 7084 37380 7140
rect 37436 7700 37492 7710
rect 36764 6468 36820 6478
rect 36652 5796 36708 5806
rect 36652 5702 36708 5740
rect 36316 5404 36708 5460
rect 36484 5124 36540 5134
rect 36484 5030 36540 5068
rect 36316 4452 36372 4462
rect 36204 4450 36372 4452
rect 36204 4398 36318 4450
rect 36370 4398 36372 4450
rect 36204 4396 36372 4398
rect 36316 4386 36372 4396
rect 35476 3666 35532 3724
rect 35980 3714 36036 3724
rect 36652 4338 36708 5404
rect 36764 5124 36820 6412
rect 36988 6356 37044 7084
rect 37436 7028 37492 7644
rect 37268 6972 37492 7028
rect 37268 6746 37324 6972
rect 37268 6694 37270 6746
rect 37322 6694 37324 6746
rect 37268 6468 37324 6694
rect 37660 6690 37716 6702
rect 37660 6638 37662 6690
rect 37714 6638 37716 6690
rect 37268 6402 37324 6412
rect 37436 6578 37492 6590
rect 37436 6526 37438 6578
rect 37490 6526 37492 6578
rect 36988 5906 37044 6300
rect 37268 6132 37324 6142
rect 37268 6018 37324 6076
rect 37268 5966 37270 6018
rect 37322 5966 37324 6018
rect 37268 5954 37324 5966
rect 36988 5854 36990 5906
rect 37042 5854 37044 5906
rect 36988 5842 37044 5854
rect 37100 5908 37156 5918
rect 37436 5908 37492 6526
rect 37548 5908 37604 5918
rect 37436 5906 37604 5908
rect 37436 5854 37550 5906
rect 37602 5854 37604 5906
rect 37436 5852 37604 5854
rect 36764 5058 36820 5068
rect 36876 5796 36932 5806
rect 36652 4286 36654 4338
rect 36706 4286 36708 4338
rect 35476 3614 35478 3666
rect 35530 3614 35532 3666
rect 35476 3602 35532 3614
rect 36372 3668 36428 3678
rect 36372 3574 36428 3612
rect 36652 3668 36708 4286
rect 36652 3602 36708 3612
rect 36876 3892 36932 5740
rect 37100 5084 37156 5852
rect 37548 5842 37604 5852
rect 37660 5572 37716 6638
rect 37996 6652 38052 7868
rect 38108 7586 38164 7980
rect 38108 7534 38110 7586
rect 38162 7534 38164 7586
rect 38108 7522 38164 7534
rect 38444 8036 38500 8046
rect 37996 6600 37998 6652
rect 38050 6600 38052 6652
rect 37996 6588 38052 6600
rect 38220 7364 38276 7374
rect 37772 5908 37828 5918
rect 38052 5908 38108 5918
rect 37772 5906 38108 5908
rect 37772 5854 37774 5906
rect 37826 5854 38054 5906
rect 38106 5854 38108 5906
rect 37772 5852 38108 5854
rect 38220 5908 38276 7308
rect 38332 6690 38388 6702
rect 38332 6638 38334 6690
rect 38386 6638 38388 6690
rect 38332 6132 38388 6638
rect 38332 6066 38388 6076
rect 38332 5908 38388 5918
rect 38220 5906 38388 5908
rect 38220 5854 38334 5906
rect 38386 5854 38388 5906
rect 38220 5852 38388 5854
rect 37772 5842 37828 5852
rect 38052 5842 38108 5852
rect 38332 5842 38388 5852
rect 38444 5906 38500 7980
rect 38556 7364 38612 8540
rect 38892 8484 38948 8494
rect 38892 8258 38948 8428
rect 38892 8206 38894 8258
rect 38946 8206 38948 8258
rect 38892 8194 38948 8206
rect 39004 8258 39060 8270
rect 39004 8206 39006 8258
rect 39058 8206 39060 8258
rect 38892 7812 38948 7822
rect 38780 7588 38836 7598
rect 38780 7384 38836 7532
rect 38556 7298 38612 7308
rect 38724 7362 38836 7384
rect 38724 7310 38726 7362
rect 38778 7310 38836 7362
rect 38724 7298 38836 7310
rect 38668 7028 38724 7038
rect 38668 6690 38724 6972
rect 38668 6638 38670 6690
rect 38722 6638 38724 6690
rect 38668 6626 38724 6638
rect 38444 5854 38446 5906
rect 38498 5854 38500 5906
rect 38444 5842 38500 5854
rect 38556 5908 38612 5918
rect 37660 5506 37716 5516
rect 37996 5572 38052 5582
rect 37100 5032 37102 5084
rect 37154 5032 37156 5084
rect 37100 5020 37156 5032
rect 37324 5348 37380 5358
rect 37324 5124 37380 5292
rect 37660 5348 37716 5358
rect 37324 4004 37380 5068
rect 37436 5236 37492 5246
rect 37436 5122 37492 5180
rect 37660 5234 37716 5292
rect 37660 5182 37662 5234
rect 37714 5182 37716 5234
rect 37660 5170 37716 5182
rect 37996 5236 38052 5516
rect 37996 5170 38052 5180
rect 37436 5070 37438 5122
rect 37490 5070 37492 5122
rect 37436 5058 37492 5070
rect 37828 5124 37884 5134
rect 37828 5030 37884 5068
rect 38556 5084 38612 5852
rect 38780 5460 38836 7298
rect 38780 5394 38836 5404
rect 38556 5032 38558 5084
rect 38610 5032 38612 5084
rect 38556 5020 38612 5032
rect 38668 5124 38724 5134
rect 37436 4228 37492 4238
rect 37436 4226 37604 4228
rect 37436 4174 37438 4226
rect 37490 4174 37604 4226
rect 37436 4172 37604 4174
rect 37436 4162 37492 4172
rect 37324 3948 37492 4004
rect 36764 3556 36820 3566
rect 36876 3556 36932 3836
rect 36820 3500 36932 3556
rect 37100 3556 37156 3566
rect 36764 3469 36766 3500
rect 36818 3469 36820 3500
rect 36764 3457 36820 3469
rect 37100 3465 37102 3500
rect 37154 3465 37156 3500
rect 37100 3453 37156 3465
rect 37436 3521 37492 3948
rect 37548 3668 37604 4172
rect 38108 4004 38164 4014
rect 38668 4004 38724 5068
rect 38892 5122 38948 7756
rect 39004 7140 39060 8206
rect 39170 8202 39226 8214
rect 39170 8150 39172 8202
rect 39224 8150 39226 8202
rect 39170 8036 39226 8150
rect 39170 7970 39226 7980
rect 39340 7474 39396 7486
rect 39340 7422 39342 7474
rect 39394 7422 39396 7474
rect 39004 7084 39284 7140
rect 39116 6690 39172 6702
rect 39116 6638 39118 6690
rect 39170 6638 39172 6690
rect 39116 6132 39172 6638
rect 39228 6580 39284 7084
rect 39340 6692 39396 7422
rect 39340 6626 39396 6636
rect 39452 6663 39508 9100
rect 39900 9156 39956 9166
rect 39900 9042 39956 9100
rect 39900 8990 39902 9042
rect 39954 8990 39956 9042
rect 39900 8978 39956 8990
rect 40012 9044 40068 9054
rect 40124 9044 40180 9884
rect 40236 9874 40292 9884
rect 40460 9828 40516 13570
rect 40572 12850 40628 12862
rect 40572 12798 40574 12850
rect 40626 12798 40628 12850
rect 40572 12628 40628 12798
rect 40572 12562 40628 12572
rect 40684 12852 40740 12862
rect 40684 11844 40740 12796
rect 40684 11778 40740 11788
rect 40796 11620 40852 15092
rect 41132 14530 41188 15260
rect 41244 15204 41300 15214
rect 41244 15110 41300 15148
rect 41468 15204 41524 17612
rect 41634 17666 41690 17724
rect 42700 17678 42756 18396
rect 42924 18360 42980 18844
rect 42868 18338 42980 18360
rect 42868 18286 42870 18338
rect 42922 18286 42980 18338
rect 42868 18274 42980 18286
rect 41634 17614 41636 17666
rect 41688 17614 41690 17666
rect 41634 17602 41690 17614
rect 42476 17666 42532 17678
rect 42476 17614 42478 17666
rect 42530 17614 42532 17666
rect 42476 17444 42532 17614
rect 42588 17668 42644 17678
rect 42700 17666 42810 17678
rect 42700 17614 42756 17666
rect 42808 17614 42810 17666
rect 42700 17612 42810 17614
rect 42588 17574 42644 17612
rect 42754 17602 42810 17612
rect 42924 17556 42980 18274
rect 43148 17778 43204 17790
rect 43148 17726 43150 17778
rect 43202 17726 43204 17778
rect 43148 17668 43204 17726
rect 43148 17602 43204 17612
rect 42924 17490 42980 17500
rect 42476 17378 42532 17388
rect 43148 16996 43204 17006
rect 42812 16884 42868 16894
rect 41580 16098 41636 16110
rect 41580 16046 41582 16098
rect 41634 16046 41636 16098
rect 42252 16098 42308 16110
rect 41580 15876 41636 16046
rect 41972 16042 42028 16054
rect 41580 15810 41636 15820
rect 41804 15986 41860 15998
rect 41804 15934 41806 15986
rect 41858 15934 41860 15986
rect 41468 15138 41524 15148
rect 41692 15652 41748 15662
rect 41132 14478 41134 14530
rect 41186 14478 41188 14530
rect 41132 14466 41188 14478
rect 41692 14530 41748 15596
rect 41692 14478 41694 14530
rect 41746 14478 41748 14530
rect 41692 14466 41748 14478
rect 40964 14420 41020 14430
rect 40964 14362 41020 14364
rect 40964 14310 40966 14362
rect 41018 14310 41020 14362
rect 40964 14298 41020 14310
rect 41412 13972 41468 13982
rect 41412 13878 41468 13916
rect 41804 13748 41860 15934
rect 41972 15990 41974 16042
rect 42026 15990 42028 16042
rect 41972 15652 42028 15990
rect 42252 16046 42254 16098
rect 42306 16046 42308 16098
rect 42252 15764 42308 16046
rect 42252 15698 42308 15708
rect 42364 16098 42420 16110
rect 42364 16046 42366 16098
rect 42418 16046 42420 16098
rect 41972 15586 42028 15596
rect 42140 15428 42196 15438
rect 41804 13682 41860 13692
rect 41916 15314 41972 15326
rect 41916 15262 41918 15314
rect 41970 15262 41972 15314
rect 41916 13636 41972 15262
rect 41916 13570 41972 13580
rect 42028 15092 42084 15102
rect 42028 14474 42084 15036
rect 42028 14422 42030 14474
rect 42082 14422 42084 14474
rect 41804 13522 41860 13534
rect 41804 13470 41806 13522
rect 41858 13470 41860 13522
rect 41692 13076 41748 13086
rect 41468 13074 41748 13076
rect 41468 13022 41694 13074
rect 41746 13022 41748 13074
rect 41468 13020 41748 13022
rect 41020 12962 41076 12974
rect 41020 12910 41022 12962
rect 41074 12910 41076 12962
rect 41020 12404 41076 12910
rect 41132 12962 41188 12974
rect 41132 12910 41134 12962
rect 41186 12910 41188 12962
rect 41132 12516 41188 12910
rect 41298 12906 41354 12918
rect 41298 12854 41300 12906
rect 41352 12854 41354 12906
rect 41298 12852 41354 12854
rect 41298 12786 41354 12796
rect 41468 12516 41524 13020
rect 41692 13010 41748 13020
rect 41132 12450 41188 12460
rect 41244 12460 41524 12516
rect 41804 12516 41860 13470
rect 41020 12338 41076 12348
rect 41244 12292 41300 12460
rect 41804 12450 41860 12460
rect 42028 12404 42084 14422
rect 42140 13748 42196 15372
rect 42252 15314 42308 15326
rect 42252 15262 42254 15314
rect 42306 15262 42308 15314
rect 42252 14084 42308 15262
rect 42364 15204 42420 16046
rect 42532 16100 42588 16110
rect 42532 16006 42588 16044
rect 42364 15138 42420 15148
rect 42476 15540 42532 15550
rect 42364 14530 42420 14542
rect 42364 14478 42366 14530
rect 42418 14478 42420 14530
rect 42364 14196 42420 14478
rect 42476 14362 42532 15484
rect 42812 15428 42868 16828
rect 43148 16882 43204 16940
rect 43148 16830 43150 16882
rect 43202 16830 43204 16882
rect 43148 16818 43204 16830
rect 43260 16436 43316 22204
rect 43596 22148 43652 22158
rect 43372 22036 43428 22046
rect 43372 20804 43428 21980
rect 43372 20710 43428 20748
rect 43484 21588 43540 21598
rect 43484 20802 43540 21532
rect 43484 20750 43486 20802
rect 43538 20750 43540 20802
rect 43484 20738 43540 20750
rect 43484 19236 43540 19246
rect 43372 19234 43540 19236
rect 43372 19182 43486 19234
rect 43538 19182 43540 19234
rect 43372 19180 43540 19182
rect 43372 17780 43428 19180
rect 43484 19170 43540 19180
rect 43372 17714 43428 17724
rect 43484 18452 43540 18462
rect 43260 16370 43316 16380
rect 42924 16212 42980 16222
rect 43372 16212 43428 16222
rect 42924 16118 42980 16156
rect 43148 16210 43428 16212
rect 43148 16158 43374 16210
rect 43426 16158 43428 16210
rect 43148 16156 43428 16158
rect 42644 15372 42868 15428
rect 42644 15370 42700 15372
rect 42644 15318 42646 15370
rect 42698 15318 42700 15370
rect 42644 15306 42700 15318
rect 42924 15316 42980 15326
rect 43148 15316 43204 16156
rect 43372 16146 43428 16156
rect 43484 16083 43540 18396
rect 43484 16031 43486 16083
rect 43538 16031 43540 16083
rect 43484 16019 43540 16031
rect 43596 15540 43652 22092
rect 44044 21601 44100 21613
rect 44044 21549 44046 21601
rect 44098 21549 44100 21601
rect 43932 21474 43988 21486
rect 43932 21422 43934 21474
rect 43986 21422 43988 21474
rect 43932 21028 43988 21422
rect 43932 20962 43988 20972
rect 43820 20916 43876 20926
rect 43820 20822 43876 20860
rect 43932 20758 43988 20770
rect 43932 20706 43934 20758
rect 43986 20706 43988 20758
rect 43820 20692 43876 20702
rect 43820 20018 43876 20636
rect 43932 20580 43988 20706
rect 43932 20514 43988 20524
rect 44044 20244 44100 21549
rect 44268 21588 44324 21598
rect 44268 21494 44324 21532
rect 44268 21364 44324 21374
rect 44268 20802 44324 21308
rect 44268 20750 44270 20802
rect 44322 20750 44324 20802
rect 44268 20738 44324 20750
rect 44044 20178 44100 20188
rect 43820 19966 43822 20018
rect 43874 19966 43876 20018
rect 43820 19954 43876 19966
rect 44156 20018 44212 20030
rect 44156 19966 44158 20018
rect 44210 19966 44212 20018
rect 44044 19850 44100 19862
rect 44044 19798 44046 19850
rect 44098 19798 44100 19850
rect 44044 19684 44100 19798
rect 44044 19618 44100 19628
rect 43988 19460 44044 19470
rect 44156 19460 44212 19966
rect 44492 20018 44548 29260
rect 44940 29092 44996 29102
rect 44940 28866 44996 29036
rect 44940 28814 44942 28866
rect 44994 28814 44996 28866
rect 44940 28802 44996 28814
rect 45052 27972 45108 29372
rect 45388 29426 45444 30156
rect 45836 29988 45892 32060
rect 46284 32004 46340 32508
rect 46732 32340 46788 32350
rect 46060 31948 46340 32004
rect 46396 32338 46788 32340
rect 46396 32286 46734 32338
rect 46786 32286 46788 32338
rect 46396 32284 46788 32286
rect 45948 30212 46004 30222
rect 45948 30118 46004 30156
rect 46060 30210 46116 31948
rect 46172 31778 46228 31790
rect 46172 31726 46174 31778
rect 46226 31726 46228 31778
rect 46172 31108 46228 31726
rect 46172 31042 46228 31052
rect 46172 30882 46228 30894
rect 46172 30830 46174 30882
rect 46226 30830 46228 30882
rect 46172 30324 46228 30830
rect 46396 30660 46452 32284
rect 46732 32274 46788 32284
rect 46396 30604 46564 30660
rect 46396 30324 46452 30334
rect 46172 30322 46452 30324
rect 46172 30270 46398 30322
rect 46450 30270 46452 30322
rect 46172 30268 46452 30270
rect 46396 30258 46452 30268
rect 46060 30158 46062 30210
rect 46114 30158 46116 30210
rect 46060 30146 46116 30158
rect 46508 30195 46564 30604
rect 46508 30143 46510 30195
rect 46562 30143 46564 30195
rect 46844 30212 46900 30222
rect 47180 30212 47236 30222
rect 47404 30212 47460 33628
rect 48076 33458 48132 34076
rect 48076 33406 48078 33458
rect 48130 33406 48132 33458
rect 48076 33394 48132 33406
rect 48020 32788 48076 32798
rect 48020 32618 48076 32732
rect 47628 32564 47684 32574
rect 47628 32470 47684 32508
rect 48020 32566 48022 32618
rect 48074 32566 48076 32618
rect 47852 32452 47908 32462
rect 47740 32450 47908 32452
rect 47740 32398 47854 32450
rect 47906 32398 47908 32450
rect 47740 32396 47908 32398
rect 47740 31332 47796 32396
rect 47852 32386 47908 32396
rect 48020 31902 48076 32566
rect 48188 32564 48244 32574
rect 48020 31892 48132 31902
rect 46844 30210 47460 30212
rect 46844 30158 46846 30210
rect 46898 30158 47182 30210
rect 47234 30158 47460 30210
rect 46844 30156 47460 30158
rect 47516 31276 47796 31332
rect 47964 31890 48132 31892
rect 47964 31838 48078 31890
rect 48130 31838 48132 31890
rect 47964 31836 48132 31838
rect 47516 30195 47572 31276
rect 47628 31108 47684 31118
rect 47628 30322 47684 31052
rect 47628 30270 47630 30322
rect 47682 30270 47684 30322
rect 47628 30258 47684 30270
rect 46844 30146 46900 30156
rect 47180 30146 47236 30156
rect 46508 30131 46564 30143
rect 47516 30143 47518 30195
rect 47570 30143 47572 30195
rect 47964 30212 48020 31836
rect 48076 31826 48132 31836
rect 48076 31108 48132 31118
rect 48188 31108 48244 32508
rect 48076 31106 48244 31108
rect 48076 31054 48078 31106
rect 48130 31054 48244 31106
rect 48076 31052 48244 31054
rect 48300 32340 48356 32350
rect 48076 31042 48132 31052
rect 47964 30146 48020 30156
rect 47516 30131 47572 30143
rect 48132 29988 48188 29998
rect 45836 29932 46004 29988
rect 45388 29374 45390 29426
rect 45442 29374 45444 29426
rect 45388 28756 45444 29374
rect 45948 29426 46004 29932
rect 48132 29986 48244 29988
rect 48132 29934 48134 29986
rect 48186 29934 48244 29986
rect 48132 29922 48244 29934
rect 45948 29374 45950 29426
rect 46002 29374 46004 29426
rect 45780 29316 45836 29326
rect 45948 29316 46004 29374
rect 46172 29428 46228 29438
rect 46452 29428 46508 29438
rect 46732 29428 46788 29438
rect 46172 29426 46340 29428
rect 46172 29374 46174 29426
rect 46226 29374 46340 29426
rect 46172 29372 46340 29374
rect 46172 29362 46228 29372
rect 45780 29314 45892 29316
rect 45780 29262 45782 29314
rect 45834 29262 45892 29314
rect 45780 29250 45892 29262
rect 45948 29250 46004 29260
rect 45388 28690 45444 28700
rect 45276 28644 45332 28654
rect 45052 27906 45108 27916
rect 45164 28642 45332 28644
rect 45164 28590 45278 28642
rect 45330 28590 45332 28642
rect 45164 28588 45332 28590
rect 44716 27748 44772 27758
rect 44604 26068 44660 26078
rect 44604 22036 44660 26012
rect 44716 25506 44772 27692
rect 45164 27310 45220 28588
rect 45276 28578 45332 28588
rect 45836 28644 45892 29250
rect 45836 28578 45892 28588
rect 46172 29204 46228 29214
rect 45612 28532 45668 28542
rect 45500 28530 45668 28532
rect 45500 28478 45614 28530
rect 45666 28478 45668 28530
rect 45500 28476 45668 28478
rect 45388 27860 45444 27898
rect 45500 27860 45556 28476
rect 45612 28466 45668 28476
rect 46172 28084 46228 29148
rect 46284 28420 46340 29372
rect 46452 29426 46788 29428
rect 46452 29374 46454 29426
rect 46506 29374 46734 29426
rect 46786 29374 46788 29426
rect 46452 29372 46788 29374
rect 46452 29362 46508 29372
rect 46732 29362 46788 29372
rect 47068 29204 47124 29214
rect 47964 29204 48020 29214
rect 47068 29202 47572 29204
rect 47068 29150 47070 29202
rect 47122 29150 47572 29202
rect 47068 29148 47572 29150
rect 47068 29138 47124 29148
rect 47516 28754 47572 29148
rect 47964 29110 48020 29148
rect 47516 28702 47518 28754
rect 47570 28702 47572 28754
rect 47516 28690 47572 28702
rect 48188 28644 48244 29922
rect 48300 29428 48356 32284
rect 48300 29334 48356 29372
rect 48300 28644 48356 28654
rect 48188 28588 48300 28644
rect 46284 28364 46564 28420
rect 46172 28028 46452 28084
rect 45444 27804 45556 27860
rect 46060 27860 46116 27870
rect 45388 27794 45444 27804
rect 45108 27298 45220 27310
rect 45108 27246 45110 27298
rect 45162 27246 45220 27298
rect 45108 27244 45220 27246
rect 45612 27412 45668 27422
rect 45108 27234 45164 27244
rect 45388 27074 45444 27086
rect 45388 27022 45390 27074
rect 45442 27022 45444 27074
rect 44716 25454 44718 25506
rect 44770 25454 44772 25506
rect 44716 25442 44772 25454
rect 44940 26852 44996 26862
rect 44940 25620 44996 26796
rect 45388 26628 45444 27022
rect 45612 27074 45668 27356
rect 45612 27022 45614 27074
rect 45666 27022 45668 27074
rect 45612 27010 45668 27022
rect 46060 27076 46116 27804
rect 46264 27858 46320 27870
rect 46264 27806 46266 27858
rect 46318 27806 46320 27858
rect 46264 27412 46320 27806
rect 46396 27748 46452 28028
rect 46508 27970 46564 28364
rect 46508 27918 46510 27970
rect 46562 27918 46564 27970
rect 46508 27906 46564 27918
rect 46844 27860 46900 27870
rect 46396 27692 46564 27748
rect 46264 27346 46320 27356
rect 46172 27076 46228 27086
rect 46060 27074 46228 27076
rect 46060 27022 46174 27074
rect 46226 27022 46228 27074
rect 46060 27020 46228 27022
rect 46172 27010 46228 27020
rect 46396 27018 46452 27030
rect 46396 26966 46398 27018
rect 46450 26966 46452 27018
rect 45388 26572 46060 26628
rect 45164 26404 45220 26414
rect 45164 26310 45220 26348
rect 46004 26402 46060 26572
rect 46004 26350 46006 26402
rect 46058 26350 46060 26402
rect 46004 26338 46060 26350
rect 46396 26404 46452 26966
rect 45500 26290 45556 26302
rect 45500 26238 45502 26290
rect 45554 26238 45556 26290
rect 45500 26180 45556 26238
rect 45500 26114 45556 26124
rect 45612 26292 45668 26302
rect 45220 25732 45276 25742
rect 45220 25638 45276 25676
rect 44940 25506 44996 25564
rect 45612 25618 45668 26236
rect 45724 26290 45780 26302
rect 45724 26238 45726 26290
rect 45778 26238 45780 26290
rect 45724 25732 45780 26238
rect 46284 26290 46340 26302
rect 46284 26238 46286 26290
rect 46338 26238 46340 26290
rect 45724 25666 45780 25676
rect 46172 25956 46228 25966
rect 45612 25566 45614 25618
rect 45666 25566 45668 25618
rect 45612 25554 45668 25566
rect 44940 25454 44942 25506
rect 44994 25454 44996 25506
rect 46060 25508 46116 25518
rect 44940 25442 44996 25454
rect 45780 25450 45836 25462
rect 45780 25398 45782 25450
rect 45834 25398 45836 25450
rect 46060 25414 46116 25452
rect 45780 25396 45836 25398
rect 45780 25340 46004 25396
rect 44828 24836 44884 24846
rect 44828 24722 44884 24780
rect 44828 24670 44830 24722
rect 44882 24670 44884 24722
rect 44828 24658 44884 24670
rect 45052 24737 45108 24749
rect 45052 24685 45054 24737
rect 45106 24685 45108 24737
rect 44940 23714 44996 23726
rect 44940 23662 44942 23714
rect 44994 23662 44996 23714
rect 44828 23154 44884 23166
rect 44828 23102 44830 23154
rect 44882 23102 44884 23154
rect 44828 23044 44884 23102
rect 44940 23156 44996 23662
rect 45052 23268 45108 24685
rect 45388 24724 45444 24734
rect 45388 24630 45444 24668
rect 45164 24612 45220 24622
rect 45164 24518 45220 24556
rect 45836 24612 45892 24622
rect 45276 23938 45332 23950
rect 45276 23886 45278 23938
rect 45330 23886 45332 23938
rect 45276 23380 45332 23886
rect 45500 23940 45556 23950
rect 45500 23846 45556 23884
rect 45836 23911 45892 24556
rect 45836 23859 45838 23911
rect 45890 23859 45892 23911
rect 45948 23940 46004 25340
rect 46172 24722 46228 25900
rect 46172 24670 46174 24722
rect 46226 24670 46228 24722
rect 46172 24658 46228 24670
rect 46172 23940 46228 23950
rect 45948 23938 46228 23940
rect 45948 23886 46174 23938
rect 46226 23886 46228 23938
rect 45948 23884 46228 23886
rect 45836 23847 45892 23859
rect 46172 23604 46228 23884
rect 46284 23770 46340 26238
rect 46396 25508 46452 26348
rect 46508 25732 46564 27692
rect 46620 27076 46676 27086
rect 46620 26906 46676 27020
rect 46844 27074 46900 27804
rect 47068 27860 47124 27870
rect 47292 27860 47348 27870
rect 47068 27858 47236 27860
rect 47068 27806 47070 27858
rect 47122 27806 47236 27858
rect 47068 27804 47236 27806
rect 47068 27794 47124 27804
rect 46956 27690 47012 27702
rect 46956 27638 46958 27690
rect 47010 27638 47012 27690
rect 46956 27412 47012 27638
rect 46956 27346 47012 27356
rect 46844 27022 46846 27074
rect 46898 27022 46900 27074
rect 46844 27010 46900 27022
rect 47068 27074 47124 27086
rect 47068 27022 47070 27074
rect 47122 27022 47124 27074
rect 46620 26854 46622 26906
rect 46674 26854 46676 26906
rect 46620 26842 46676 26854
rect 47068 26852 47124 27022
rect 47068 26786 47124 26796
rect 47180 26404 47236 27804
rect 47292 27766 47348 27804
rect 47964 27634 48020 27646
rect 47964 27582 47966 27634
rect 48018 27582 48020 27634
rect 47964 27524 48020 27582
rect 47964 27458 48020 27468
rect 48188 27198 48244 28588
rect 48300 28550 48356 28588
rect 48300 27858 48356 27870
rect 48300 27806 48302 27858
rect 48354 27806 48356 27858
rect 48300 27636 48356 27806
rect 48300 27570 48356 27580
rect 48132 27186 48244 27198
rect 48132 27134 48134 27186
rect 48186 27134 48244 27186
rect 48132 27122 48244 27134
rect 47292 27076 47348 27114
rect 47292 27010 47348 27020
rect 47572 26962 47628 26974
rect 47572 26910 47574 26962
rect 47626 26910 47628 26962
rect 47572 26908 47628 26910
rect 46788 26348 47236 26404
rect 47292 26852 47348 26862
rect 47572 26852 47796 26908
rect 47292 26628 47348 26796
rect 46620 26066 46676 26078
rect 46620 26014 46622 26066
rect 46674 26014 46676 26066
rect 46620 25956 46676 26014
rect 46620 25890 46676 25900
rect 46508 25676 46676 25732
rect 46396 25414 46452 25452
rect 46508 25506 46564 25518
rect 46508 25454 46510 25506
rect 46562 25454 46564 25506
rect 46508 24948 46564 25454
rect 46620 25060 46676 25676
rect 46788 25730 46844 26348
rect 47124 26068 47180 26078
rect 47124 25974 47180 26012
rect 47292 25844 47348 26572
rect 47404 26740 47460 26750
rect 47404 26318 47460 26684
rect 47740 26404 47796 26852
rect 47740 26348 47852 26404
rect 47796 26346 47852 26348
rect 47404 26292 47406 26318
rect 47458 26292 47460 26318
rect 47404 26226 47460 26236
rect 47628 26318 47684 26330
rect 47628 26266 47630 26318
rect 47682 26266 47684 26318
rect 47796 26294 47798 26346
rect 47850 26294 47852 26346
rect 47796 26282 47852 26294
rect 47964 26325 48020 26337
rect 46788 25678 46790 25730
rect 46842 25678 46844 25730
rect 46788 25620 46844 25678
rect 46788 25554 46844 25564
rect 47180 25788 47348 25844
rect 47180 25506 47236 25788
rect 47628 25742 47684 26266
rect 47964 26273 47966 26325
rect 48018 26273 48020 26325
rect 47628 25730 47740 25742
rect 47628 25678 47686 25730
rect 47738 25678 47740 25730
rect 47628 25676 47740 25678
rect 47684 25666 47740 25676
rect 47404 25508 47460 25518
rect 47964 25508 48020 26273
rect 48188 25630 48244 27122
rect 48412 26292 48468 26302
rect 48188 25618 48300 25630
rect 48188 25566 48246 25618
rect 48298 25566 48300 25618
rect 48188 25564 48300 25566
rect 48244 25554 48300 25564
rect 47180 25454 47182 25506
rect 47234 25454 47236 25506
rect 47180 25396 47236 25454
rect 47180 25330 47236 25340
rect 47292 25506 48020 25508
rect 47292 25454 47406 25506
rect 47458 25454 48020 25506
rect 47292 25452 48020 25454
rect 46620 24994 46676 25004
rect 46284 23718 46286 23770
rect 46338 23718 46340 23770
rect 46284 23706 46340 23718
rect 46396 24892 46564 24948
rect 46396 23604 46452 24892
rect 47180 23940 47236 23950
rect 46172 23548 46452 23604
rect 45276 23314 45332 23324
rect 45612 23492 45668 23502
rect 45052 23202 45108 23212
rect 44940 23090 44996 23100
rect 45612 23154 45668 23436
rect 45724 23380 45780 23390
rect 45724 23322 45780 23324
rect 45724 23270 45726 23322
rect 45778 23270 45780 23322
rect 45724 23258 45780 23270
rect 46284 23268 46340 23278
rect 46396 23268 46452 23548
rect 47068 23938 47236 23940
rect 47068 23886 47182 23938
rect 47234 23886 47236 23938
rect 47068 23884 47236 23886
rect 46900 23268 46956 23278
rect 46396 23266 46956 23268
rect 46396 23214 46902 23266
rect 46954 23214 46956 23266
rect 46396 23212 46956 23214
rect 46060 23193 46116 23205
rect 45612 23102 45614 23154
rect 45666 23102 45668 23154
rect 45612 23090 45668 23102
rect 45836 23156 45892 23166
rect 44828 22596 44884 22988
rect 45220 23042 45276 23054
rect 45220 22990 45222 23042
rect 45274 22990 45276 23042
rect 45220 22820 45276 22990
rect 45220 22754 45276 22764
rect 44828 22540 45220 22596
rect 45052 22372 45108 22382
rect 44604 21970 44660 21980
rect 44716 22370 45108 22372
rect 44716 22318 45054 22370
rect 45106 22318 45108 22370
rect 44716 22316 45108 22318
rect 44604 21812 44660 21822
rect 44604 21586 44660 21756
rect 44604 21534 44606 21586
rect 44658 21534 44660 21586
rect 44604 20188 44660 21534
rect 44716 20804 44772 22316
rect 45052 22306 45108 22316
rect 45164 22260 45220 22540
rect 45836 22482 45892 23100
rect 45836 22430 45838 22482
rect 45890 22430 45892 22482
rect 45836 22418 45892 22430
rect 46060 23141 46062 23193
rect 46114 23141 46116 23193
rect 45164 22204 45780 22260
rect 45612 21586 45668 21598
rect 45612 21534 45614 21586
rect 45666 21534 45668 21586
rect 44716 20710 44772 20748
rect 44940 21362 44996 21374
rect 44940 21310 44942 21362
rect 44994 21310 44996 21362
rect 44604 20132 44772 20188
rect 44492 19966 44494 20018
rect 44546 19966 44548 20018
rect 44492 19908 44548 19966
rect 44716 20018 44772 20132
rect 44716 19966 44718 20018
rect 44770 19966 44772 20018
rect 44716 19954 44772 19966
rect 44492 19842 44548 19852
rect 44940 19908 44996 21310
rect 45612 21364 45668 21534
rect 45612 21298 45668 21308
rect 45612 21140 45668 21150
rect 45500 20916 45556 20926
rect 45500 20822 45556 20860
rect 45276 20804 45332 20814
rect 45276 20020 45332 20748
rect 45500 20356 45556 20366
rect 45388 20020 45444 20030
rect 45276 20018 45444 20020
rect 45276 19966 45390 20018
rect 45442 19966 45444 20018
rect 45276 19964 45444 19966
rect 44940 19842 44996 19852
rect 45052 19796 45108 19806
rect 45052 19702 45108 19740
rect 43988 19458 44212 19460
rect 43988 19406 43990 19458
rect 44042 19406 44212 19458
rect 43988 19404 44212 19406
rect 43988 19394 44044 19404
rect 43708 19236 43764 19246
rect 43708 19142 43764 19180
rect 44828 19234 44884 19246
rect 44828 19182 44830 19234
rect 44882 19182 44884 19234
rect 44690 18900 44746 18910
rect 43708 18676 43764 18686
rect 43708 18506 43764 18620
rect 43708 18454 43710 18506
rect 43762 18454 43764 18506
rect 44268 18676 44324 18686
rect 43708 18442 43764 18454
rect 43932 18483 43988 18495
rect 43932 18431 43934 18483
rect 43986 18431 43988 18483
rect 43932 17834 43988 18431
rect 43820 17780 43876 17790
rect 43932 17782 43934 17834
rect 43986 17782 43988 17834
rect 43932 17770 43988 17782
rect 44044 17892 44100 17902
rect 43708 17666 43764 17678
rect 43708 17614 43710 17666
rect 43762 17614 43764 17666
rect 43708 17556 43764 17614
rect 43708 17490 43764 17500
rect 43820 16926 43876 17724
rect 43932 17668 43988 17678
rect 43932 17574 43988 17612
rect 43708 16884 43764 16894
rect 43820 16874 43822 16926
rect 43874 16874 43876 16926
rect 43820 16862 43876 16874
rect 44044 16882 44100 17836
rect 43708 16770 43764 16828
rect 44044 16830 44046 16882
rect 44098 16830 44100 16882
rect 44044 16818 44100 16830
rect 43708 16718 43710 16770
rect 43762 16718 43764 16770
rect 43708 16706 43764 16718
rect 43708 16548 43764 16558
rect 43708 16100 43764 16492
rect 43708 16006 43764 16044
rect 43820 16212 43876 16222
rect 43596 15484 43764 15540
rect 43372 15428 43428 15438
rect 42924 15314 43204 15316
rect 42924 15262 42926 15314
rect 42978 15262 43204 15314
rect 42924 15260 43204 15262
rect 43260 15316 43316 15326
rect 42924 15250 42980 15260
rect 43260 15222 43316 15260
rect 43372 15314 43428 15372
rect 43372 15262 43374 15314
rect 43426 15262 43428 15314
rect 42476 14310 42478 14362
rect 42530 14310 42532 14362
rect 42476 14298 42532 14310
rect 42588 15202 42644 15214
rect 42588 15150 42590 15202
rect 42642 15150 42644 15202
rect 42588 14196 42644 15150
rect 42812 15204 42868 15214
rect 43372 15148 43428 15262
rect 42364 14140 42644 14196
rect 42700 14644 42756 14654
rect 42252 14028 42644 14084
rect 42476 13784 42532 13796
rect 42476 13748 42478 13784
rect 42140 13746 42478 13748
rect 42140 13694 42142 13746
rect 42194 13732 42478 13746
rect 42530 13732 42532 13784
rect 42194 13694 42532 13732
rect 42140 13692 42532 13694
rect 42140 13682 42196 13692
rect 42588 13074 42644 14028
rect 42588 13022 42590 13074
rect 42642 13022 42644 13074
rect 42588 13010 42644 13022
rect 42140 12962 42196 12974
rect 42140 12910 42142 12962
rect 42194 12910 42196 12962
rect 42140 12628 42196 12910
rect 42140 12562 42196 12572
rect 42476 12918 42532 12930
rect 42476 12866 42478 12918
rect 42530 12866 42532 12918
rect 42028 12348 42196 12404
rect 41244 12222 41300 12236
rect 41020 12178 41076 12190
rect 41020 12126 41022 12178
rect 41074 12126 41076 12178
rect 41244 12170 41246 12222
rect 41298 12170 41300 12222
rect 41244 12158 41300 12170
rect 41804 12193 41860 12205
rect 41020 11956 41076 12126
rect 41804 12141 41806 12193
rect 41858 12141 41860 12193
rect 41356 12068 41412 12078
rect 41692 12068 41748 12078
rect 41356 11974 41412 12012
rect 41580 12066 41748 12068
rect 41580 12014 41694 12066
rect 41746 12014 41748 12066
rect 41580 12012 41748 12014
rect 41020 11890 41076 11900
rect 41020 11676 41524 11732
rect 41020 11620 41076 11676
rect 40796 11564 41076 11620
rect 40908 11452 41244 11508
rect 40796 11394 40852 11406
rect 40572 11338 40628 11350
rect 40572 11286 40574 11338
rect 40626 11286 40628 11338
rect 40572 11284 40628 11286
rect 40572 11218 40628 11228
rect 40796 11342 40798 11394
rect 40850 11342 40852 11394
rect 40796 10836 40852 11342
rect 40684 10780 40852 10836
rect 40684 10388 40740 10780
rect 40684 10322 40740 10332
rect 40796 10610 40852 10622
rect 40796 10558 40798 10610
rect 40850 10558 40852 10610
rect 40684 9828 40740 9838
rect 40460 9826 40740 9828
rect 40460 9774 40686 9826
rect 40738 9774 40740 9826
rect 40460 9772 40740 9774
rect 40348 9604 40404 9614
rect 40348 9602 40516 9604
rect 40348 9550 40350 9602
rect 40402 9550 40516 9602
rect 40348 9548 40516 9550
rect 40348 9538 40404 9548
rect 40460 9380 40516 9548
rect 40292 9268 40348 9278
rect 40292 9154 40348 9212
rect 40292 9102 40294 9154
rect 40346 9102 40348 9154
rect 40292 9090 40348 9102
rect 40012 9042 40180 9044
rect 40012 8990 40014 9042
rect 40066 8990 40180 9042
rect 40012 8988 40180 8990
rect 40460 9044 40516 9324
rect 40012 8978 40068 8988
rect 40460 8978 40516 8988
rect 39564 8370 39620 8382
rect 39564 8318 39566 8370
rect 39618 8318 39620 8370
rect 39564 7924 39620 8318
rect 40012 8370 40068 8382
rect 40012 8318 40014 8370
rect 40066 8318 40068 8370
rect 39564 7858 39620 7868
rect 39676 8148 39732 8158
rect 39676 7474 39732 8092
rect 39676 7422 39678 7474
rect 39730 7422 39732 7474
rect 40012 7530 40068 8318
rect 40460 8258 40516 8270
rect 40124 8214 40180 8226
rect 40124 8162 40126 8214
rect 40178 8162 40180 8214
rect 40124 8036 40180 8162
rect 40124 7970 40180 7980
rect 40460 8206 40462 8258
rect 40514 8206 40516 8258
rect 40012 7478 40014 7530
rect 40066 7478 40068 7530
rect 40012 7466 40068 7478
rect 40348 7476 40404 7486
rect 39676 7410 39732 7422
rect 40348 7382 40404 7420
rect 40012 7364 40068 7374
rect 39228 6522 39284 6524
rect 39228 6470 39230 6522
rect 39282 6470 39284 6522
rect 39228 6458 39284 6470
rect 39452 6611 39454 6663
rect 39506 6611 39508 6663
rect 39788 7362 40068 7364
rect 39788 7310 40014 7362
rect 40066 7310 40068 7362
rect 39788 7308 40068 7310
rect 39788 6690 39844 7308
rect 40012 7298 40068 7308
rect 40460 7028 40516 8206
rect 40460 6962 40516 6972
rect 39788 6638 39790 6690
rect 39842 6638 39844 6690
rect 39788 6626 39844 6638
rect 40236 6690 40292 6702
rect 40236 6638 40238 6690
rect 40290 6638 40292 6690
rect 39452 6244 39508 6611
rect 40236 6580 40292 6638
rect 40236 6514 40292 6524
rect 40572 6468 40628 6478
rect 40572 6374 40628 6412
rect 39116 6066 39172 6076
rect 39302 6188 39508 6244
rect 40684 6244 40740 9772
rect 40796 8372 40852 10558
rect 40908 9994 40964 11452
rect 41188 11450 41244 11452
rect 41188 11398 41190 11450
rect 41242 11398 41244 11450
rect 41188 11386 41244 11398
rect 41020 11282 41076 11294
rect 41020 11230 41022 11282
rect 41074 11230 41076 11282
rect 41020 10612 41076 11230
rect 41020 10546 41076 10556
rect 40908 9942 40910 9994
rect 40962 9942 40964 9994
rect 40908 9930 40964 9942
rect 41020 9828 41076 9838
rect 41020 9734 41076 9772
rect 41356 9828 41412 9838
rect 41468 9828 41524 11676
rect 41580 11284 41636 12012
rect 41692 12002 41748 12012
rect 41804 12068 41860 12141
rect 42028 12180 42084 12190
rect 42028 12086 42084 12124
rect 41804 12002 41860 12012
rect 42140 11620 42196 12348
rect 42476 11844 42532 12866
rect 42700 12852 42756 14588
rect 42812 14530 42868 15148
rect 43148 15092 43428 15148
rect 43518 15351 43574 15363
rect 43518 15299 43520 15351
rect 43572 15299 43574 15351
rect 43518 15204 43574 15299
rect 43518 15138 43574 15148
rect 43148 14754 43204 15092
rect 43708 14980 43764 15484
rect 43148 14702 43150 14754
rect 43202 14702 43204 14754
rect 43148 14690 43204 14702
rect 43596 14924 43764 14980
rect 43596 14532 43652 14924
rect 43820 14868 43876 16156
rect 44044 16100 44100 16110
rect 43932 16098 44100 16100
rect 43932 16046 44046 16098
rect 44098 16046 44100 16098
rect 43932 16044 44100 16046
rect 43932 15202 43988 16044
rect 44044 16034 44100 16044
rect 44268 16100 44324 18620
rect 44492 18486 44548 18498
rect 44492 18434 44494 18486
rect 44546 18434 44548 18486
rect 44492 17892 44548 18434
rect 44690 18490 44746 18844
rect 44690 18438 44692 18490
rect 44744 18438 44746 18490
rect 44690 18426 44746 18438
rect 44828 18452 44884 19182
rect 44828 18386 44884 18396
rect 44940 19236 44996 19246
rect 44716 18340 44772 18350
rect 44716 18246 44772 18284
rect 44492 17836 44884 17892
rect 44380 17556 44436 17566
rect 44380 16882 44436 17500
rect 44380 16830 44382 16882
rect 44434 16830 44436 16882
rect 44380 16818 44436 16830
rect 44268 16034 44324 16044
rect 44380 16436 44436 16446
rect 44212 15876 44268 15886
rect 43932 15150 43934 15202
rect 43986 15150 43988 15202
rect 43932 15138 43988 15150
rect 44044 15874 44268 15876
rect 44044 15822 44214 15874
rect 44266 15822 44268 15874
rect 44044 15820 44268 15822
rect 43820 14812 43988 14868
rect 42812 14478 42814 14530
rect 42866 14478 42868 14530
rect 42812 14466 42868 14478
rect 42924 14476 43652 14532
rect 43932 14530 43988 14812
rect 43932 14478 43934 14530
rect 43986 14478 43988 14530
rect 42812 14308 42868 14318
rect 42812 13746 42868 14252
rect 42812 13694 42814 13746
rect 42866 13694 42868 13746
rect 42812 13682 42868 13694
rect 42924 13636 42980 14476
rect 43932 14466 43988 14478
rect 43036 13860 43092 13870
rect 43036 13766 43092 13804
rect 43204 13804 43652 13860
rect 43204 13802 43316 13804
rect 43204 13750 43206 13802
rect 43258 13750 43316 13802
rect 43204 13738 43316 13750
rect 42924 13580 43092 13636
rect 42588 12796 42756 12852
rect 42588 12178 42644 12796
rect 42588 12126 42590 12178
rect 42642 12126 42644 12178
rect 42588 12114 42644 12126
rect 42700 12516 42756 12526
rect 42700 12178 42756 12460
rect 42700 12126 42702 12178
rect 42754 12126 42756 12178
rect 42886 12404 42942 12414
rect 42886 12216 42942 12348
rect 42886 12164 42888 12216
rect 42940 12164 42942 12216
rect 42886 12152 42942 12164
rect 42700 12114 42756 12126
rect 43036 11956 43092 13580
rect 43260 13524 43316 13738
rect 43596 13790 43652 13804
rect 43596 13738 43598 13790
rect 43650 13738 43652 13790
rect 43596 13726 43652 13738
rect 43820 13746 43876 13758
rect 43820 13694 43822 13746
rect 43874 13694 43876 13746
rect 43484 13636 43540 13646
rect 43484 13542 43540 13580
rect 43260 13458 43316 13468
rect 43391 13412 43447 13422
rect 43820 13412 43876 13694
rect 43391 12962 43447 13356
rect 43391 12910 43393 12962
rect 43445 12910 43447 12962
rect 43391 12898 43447 12910
rect 43596 13356 43876 13412
rect 44044 13412 44100 15820
rect 44212 15810 44268 15820
rect 44380 15652 44436 16380
rect 44156 15596 44436 15652
rect 44156 14698 44212 15596
rect 44492 15316 44548 17836
rect 44604 17668 44660 17678
rect 44604 16882 44660 17612
rect 44604 16830 44606 16882
rect 44658 16830 44660 16882
rect 44604 16818 44660 16830
rect 44828 16894 44884 17836
rect 44940 17668 44996 19180
rect 45220 19236 45276 19246
rect 45220 19142 45276 19180
rect 45052 18452 45108 18462
rect 45388 18452 45444 19964
rect 45500 19012 45556 20300
rect 45612 20020 45668 21084
rect 45724 20188 45780 22204
rect 46060 22148 46116 23141
rect 46284 23154 46340 23212
rect 46900 23202 46956 23212
rect 46284 23102 46286 23154
rect 46338 23102 46340 23154
rect 46284 23090 46340 23102
rect 46956 22260 47012 22270
rect 46060 22092 46564 22148
rect 46116 21700 46172 21710
rect 46116 21606 46172 21644
rect 45836 21586 45892 21598
rect 45836 21534 45838 21586
rect 45890 21534 45892 21586
rect 45836 21140 45892 21534
rect 46508 21474 46564 22092
rect 46620 21601 46676 21626
rect 46620 21588 46622 21601
rect 46674 21588 46676 21601
rect 46620 21522 46676 21532
rect 46956 21586 47012 22204
rect 47068 21700 47124 23884
rect 47180 23874 47236 23884
rect 47292 23770 47348 25452
rect 47404 25442 47460 25452
rect 48188 25396 48244 25406
rect 47740 24836 47796 24846
rect 47740 24052 47796 24780
rect 48076 24836 48132 24846
rect 48076 24742 48132 24780
rect 47292 23718 47294 23770
rect 47346 23718 47348 23770
rect 47292 23706 47348 23718
rect 47404 23996 47796 24052
rect 47180 23268 47236 23278
rect 47180 23154 47236 23212
rect 47180 23102 47182 23154
rect 47234 23102 47236 23154
rect 47180 23090 47236 23102
rect 47404 23154 47460 23996
rect 47740 23938 47796 23996
rect 47572 23882 47628 23894
rect 47572 23830 47574 23882
rect 47626 23830 47628 23882
rect 47740 23886 47742 23938
rect 47794 23886 47796 23938
rect 47740 23874 47796 23886
rect 47572 23828 47628 23830
rect 47572 23772 47684 23828
rect 47404 23102 47406 23154
rect 47458 23102 47460 23154
rect 47404 23090 47460 23102
rect 47628 23154 47684 23772
rect 48020 23268 48076 23278
rect 48020 23174 48076 23212
rect 47628 23102 47630 23154
rect 47682 23102 47684 23154
rect 47628 22260 47684 23102
rect 47740 23156 47796 23166
rect 47740 23154 47908 23156
rect 47740 23102 47742 23154
rect 47794 23102 47908 23154
rect 47740 23100 47908 23102
rect 47740 23090 47796 23100
rect 47740 22260 47796 22270
rect 47628 22204 47740 22260
rect 47740 22166 47796 22204
rect 47628 21700 47684 21710
rect 47068 21634 47124 21644
rect 47180 21644 47404 21700
rect 46956 21534 46958 21586
rect 47010 21534 47012 21586
rect 46956 21522 47012 21534
rect 46508 21422 46510 21474
rect 46562 21422 46564 21474
rect 46508 21410 46564 21422
rect 45836 21074 45892 21084
rect 46396 20580 46452 20590
rect 45724 20132 46116 20188
rect 45612 19954 45668 19964
rect 45948 19796 46004 19806
rect 45500 18946 45556 18956
rect 45612 19402 45668 19414
rect 45612 19350 45614 19402
rect 45666 19350 45668 19402
rect 45612 18900 45668 19350
rect 45724 19236 45780 19246
rect 45724 19142 45780 19180
rect 45948 19234 46004 19740
rect 45948 19182 45950 19234
rect 46002 19182 46004 19234
rect 45612 18834 45668 18844
rect 45948 18788 46004 19182
rect 45948 18722 46004 18732
rect 45052 18450 45444 18452
rect 45052 18398 45054 18450
rect 45106 18398 45444 18450
rect 45052 18396 45444 18398
rect 45052 18386 45108 18396
rect 44940 17612 45220 17668
rect 44940 17442 44996 17454
rect 44940 17390 44942 17442
rect 44994 17390 44996 17442
rect 44940 17108 44996 17390
rect 44940 17042 44996 17052
rect 44828 16882 44940 16894
rect 44828 16830 44886 16882
rect 44938 16830 44940 16882
rect 44828 16828 44940 16830
rect 44884 16818 44940 16828
rect 44996 16324 45052 16334
rect 44996 16230 45052 16268
rect 44156 14646 44158 14698
rect 44210 14646 44212 14698
rect 44156 14634 44212 14646
rect 44268 15314 44548 15316
rect 44268 15262 44494 15314
rect 44546 15262 44548 15314
rect 44716 16100 44772 16110
rect 44716 15358 44772 16044
rect 44828 16100 44884 16110
rect 44828 16098 44996 16100
rect 44828 16046 44830 16098
rect 44882 16046 44996 16098
rect 44828 16044 44996 16046
rect 44828 16034 44884 16044
rect 44716 15306 44718 15358
rect 44770 15306 44772 15358
rect 44716 15294 44772 15306
rect 44268 15260 44548 15262
rect 44268 14530 44324 15260
rect 44492 15250 44548 15260
rect 44828 15202 44884 15214
rect 44828 15150 44830 15202
rect 44882 15150 44884 15202
rect 44268 14478 44270 14530
rect 44322 14478 44324 14530
rect 44268 14466 44324 14478
rect 44380 14980 44436 14990
rect 44380 14308 44436 14924
rect 42476 11778 42532 11788
rect 42700 11900 43092 11956
rect 43148 12850 43204 12862
rect 43148 12798 43150 12850
rect 43202 12798 43204 12850
rect 41580 11218 41636 11228
rect 41692 11564 42196 11620
rect 41692 11394 41748 11564
rect 41692 11342 41694 11394
rect 41746 11342 41748 11394
rect 41692 10724 41748 11342
rect 41804 11396 41860 11406
rect 41804 11302 41860 11340
rect 42588 11396 42644 11406
rect 42700 11396 42756 11900
rect 43148 11732 43204 12798
rect 43596 12404 43652 13356
rect 44044 13346 44100 13356
rect 44268 14252 44436 14308
rect 44492 14532 44548 14542
rect 44268 13300 44324 14252
rect 44380 14084 44436 14094
rect 44380 13300 44436 14028
rect 44492 13748 44548 14476
rect 44828 14530 44884 15150
rect 44828 14478 44830 14530
rect 44882 14478 44884 14530
rect 44828 14084 44884 14478
rect 44940 14308 44996 16044
rect 45164 14980 45220 17612
rect 45276 17666 45332 17678
rect 45276 17614 45278 17666
rect 45330 17614 45332 17666
rect 45276 17556 45332 17614
rect 45388 17666 45444 18396
rect 45836 18340 45892 18350
rect 45836 18246 45892 18284
rect 45388 17614 45390 17666
rect 45442 17614 45444 17666
rect 45388 17602 45444 17614
rect 45276 17490 45332 17500
rect 46060 17108 46116 20132
rect 46172 20020 46228 20030
rect 46396 20020 46452 20524
rect 47180 20188 47236 21644
rect 47348 21615 47404 21644
rect 47348 21563 47350 21615
rect 47402 21563 47404 21615
rect 47348 21551 47404 21563
rect 47292 21474 47348 21486
rect 47292 21422 47294 21474
rect 47346 21422 47348 21474
rect 47292 20580 47348 21422
rect 47292 20514 47348 20524
rect 47404 21364 47460 21374
rect 47404 20690 47460 21308
rect 47404 20638 47406 20690
rect 47458 20638 47460 20690
rect 47180 20132 47348 20188
rect 46172 20018 46452 20020
rect 46172 19966 46174 20018
rect 46226 19966 46452 20018
rect 46172 19964 46452 19966
rect 46172 19954 46228 19964
rect 47292 19684 47348 20132
rect 47180 19628 47348 19684
rect 47180 19402 47236 19628
rect 47180 19350 47182 19402
rect 47234 19350 47236 19402
rect 47180 19338 47236 19350
rect 46844 19236 46900 19246
rect 46844 19142 46900 19180
rect 47068 19234 47124 19246
rect 47068 19182 47070 19234
rect 47122 19182 47124 19234
rect 47068 19012 47124 19182
rect 47404 19234 47460 20638
rect 47628 20188 47684 21644
rect 47740 21588 47796 21598
rect 47852 21588 47908 23100
rect 48188 23044 48244 25340
rect 47796 21532 47908 21588
rect 47964 22988 48244 23044
rect 47740 21494 47796 21532
rect 47964 21364 48020 22988
rect 47852 21308 48020 21364
rect 48076 21588 48132 21598
rect 47852 20188 47908 21308
rect 47964 20578 48020 20590
rect 47964 20526 47966 20578
rect 48018 20526 48020 20578
rect 47964 20356 48020 20526
rect 47964 20290 48020 20300
rect 48076 20188 48132 21532
rect 48244 21474 48300 21486
rect 48244 21422 48246 21474
rect 48298 21422 48300 21474
rect 48244 21252 48300 21422
rect 48244 21186 48300 21196
rect 48300 20804 48356 20814
rect 48300 20710 48356 20748
rect 48412 20188 48468 26236
rect 48748 22484 48804 22494
rect 48748 20804 48804 22428
rect 48748 20188 48804 20748
rect 47404 19182 47406 19234
rect 47458 19182 47460 19234
rect 47404 19170 47460 19182
rect 47516 20132 47684 20188
rect 47740 20132 47908 20188
rect 47964 20132 48132 20188
rect 48188 20132 48468 20188
rect 48524 20132 48804 20188
rect 47516 19012 47572 20132
rect 47628 20020 47684 20030
rect 47628 19234 47684 19964
rect 47628 19182 47630 19234
rect 47682 19182 47684 19234
rect 47628 19170 47684 19182
rect 47068 18956 47572 19012
rect 47292 18788 47348 18798
rect 46172 17668 46228 17678
rect 46172 17666 46452 17668
rect 46172 17614 46174 17666
rect 46226 17614 46452 17666
rect 46172 17612 46452 17614
rect 46172 17602 46228 17612
rect 46396 17332 46452 17612
rect 46396 17276 46564 17332
rect 46060 17052 46228 17108
rect 45500 16996 45556 17006
rect 45388 16915 45444 16927
rect 45388 16863 45390 16915
rect 45442 16863 45444 16915
rect 45388 16042 45444 16863
rect 45388 15990 45390 16042
rect 45442 15990 45444 16042
rect 45164 14914 45220 14924
rect 45276 15204 45332 15214
rect 45164 14644 45220 14682
rect 45164 14578 45220 14588
rect 44940 14242 44996 14252
rect 45164 14474 45220 14486
rect 45164 14422 45166 14474
rect 45218 14422 45220 14474
rect 45164 14084 45220 14422
rect 44828 14028 45108 14084
rect 45052 13860 45108 14028
rect 45164 14018 45220 14028
rect 45276 13870 45332 15148
rect 45388 14980 45444 15990
rect 45388 14914 45444 14924
rect 45500 15316 45556 16940
rect 45612 16915 45668 16927
rect 45612 16863 45614 16915
rect 45666 16863 45668 16915
rect 45612 16436 45668 16863
rect 45612 16370 45668 16380
rect 46060 16915 46116 16927
rect 46060 16863 46062 16915
rect 46114 16863 46116 16915
rect 46060 16324 46116 16863
rect 46060 16258 46116 16268
rect 46172 16212 46228 17052
rect 46508 16994 46564 17276
rect 46508 16942 46510 16994
rect 46562 16942 46564 16994
rect 46508 16930 46564 16942
rect 46370 16915 46426 16927
rect 46370 16863 46372 16915
rect 46424 16884 46426 16915
rect 46956 16884 47012 16894
rect 46424 16863 46452 16884
rect 46370 16828 46452 16863
rect 46396 16772 46452 16828
rect 46956 16790 47012 16828
rect 47292 16884 47348 18732
rect 47740 18564 47796 20132
rect 47964 19470 48020 20132
rect 48076 20020 48132 20030
rect 48076 19926 48132 19964
rect 47908 19458 48020 19470
rect 47908 19406 47910 19458
rect 47962 19406 48020 19458
rect 47908 19404 48020 19406
rect 47908 19394 47964 19404
rect 47740 18508 47908 18564
rect 47740 18340 47796 18350
rect 47740 18246 47796 18284
rect 47684 16884 47740 16894
rect 47292 16882 47572 16884
rect 47292 16830 47294 16882
rect 47346 16830 47572 16882
rect 47292 16828 47572 16830
rect 47292 16818 47348 16828
rect 46396 16716 46900 16772
rect 46844 16714 46900 16716
rect 46844 16662 46846 16714
rect 46898 16662 46900 16714
rect 46844 16650 46900 16662
rect 47516 16212 47572 16828
rect 47684 16790 47740 16828
rect 46172 16156 46340 16212
rect 47516 16156 47796 16212
rect 45612 16100 45668 16110
rect 45612 15652 45668 16044
rect 45612 15426 45668 15596
rect 45612 15374 45614 15426
rect 45666 15374 45668 15426
rect 45612 15362 45668 15374
rect 45724 16042 45780 16054
rect 45724 15990 45726 16042
rect 45778 15990 45780 16042
rect 45500 14756 45556 15260
rect 45724 15204 45780 15990
rect 45724 15138 45780 15148
rect 46172 16042 46228 16054
rect 46172 15990 46174 16042
rect 46226 15990 46228 16042
rect 45052 13804 45164 13860
rect 44828 13748 44884 13758
rect 44492 13654 44548 13692
rect 44660 13690 44716 13702
rect 44660 13638 44662 13690
rect 44714 13638 44716 13690
rect 44828 13654 44884 13692
rect 44940 13746 44996 13758
rect 44940 13694 44942 13746
rect 44994 13694 44996 13746
rect 44660 13636 44716 13638
rect 44660 13570 44716 13580
rect 44940 13412 44996 13694
rect 45108 13636 45164 13804
rect 45220 13858 45332 13870
rect 45220 13806 45222 13858
rect 45274 13806 45332 13858
rect 45220 13804 45332 13806
rect 45388 14700 45556 14756
rect 45612 14980 45668 14990
rect 45220 13794 45276 13804
rect 44940 13346 44996 13356
rect 45052 13580 45164 13636
rect 45276 13636 45332 13646
rect 44604 13300 44660 13310
rect 44380 13244 44548 13300
rect 44268 13234 44324 13244
rect 44268 12962 44324 12974
rect 44268 12910 44270 12962
rect 44322 12910 44324 12962
rect 44268 12740 44324 12910
rect 44268 12674 44324 12684
rect 44492 12516 44548 13244
rect 43596 12338 43652 12348
rect 43876 12460 44548 12516
rect 43876 12402 43932 12460
rect 44604 12404 44660 13244
rect 44716 12964 44772 12974
rect 45052 12964 45108 13580
rect 45276 13524 45332 13580
rect 44716 12962 45108 12964
rect 44716 12910 44718 12962
rect 44770 12910 45108 12962
rect 44716 12908 45108 12910
rect 45164 13468 45332 13524
rect 44716 12898 44772 12908
rect 45052 12740 45108 12750
rect 45164 12740 45220 13468
rect 45052 12738 45220 12740
rect 45052 12686 45054 12738
rect 45106 12686 45220 12738
rect 45052 12684 45220 12686
rect 45276 13300 45332 13310
rect 45052 12674 45108 12684
rect 43876 12350 43878 12402
rect 43930 12350 43932 12402
rect 43876 12338 43932 12350
rect 44492 12348 44660 12404
rect 44268 12292 44324 12302
rect 43260 12180 43316 12190
rect 43260 12066 43316 12124
rect 43260 12014 43262 12066
rect 43314 12014 43316 12066
rect 43260 12002 43316 12014
rect 44268 12078 44324 12236
rect 44268 12066 44380 12078
rect 44268 12014 44326 12066
rect 44378 12014 44380 12066
rect 44268 12002 44380 12014
rect 43148 11666 43204 11676
rect 43484 11844 43540 11854
rect 42924 11562 42980 11574
rect 42924 11510 42926 11562
rect 42978 11510 42980 11562
rect 42924 11508 42980 11510
rect 42924 11452 43260 11508
rect 43204 11450 43260 11452
rect 42644 11340 42756 11396
rect 42812 11394 42868 11406
rect 42812 11342 42814 11394
rect 42866 11342 42868 11394
rect 43204 11398 43206 11450
rect 43258 11398 43260 11450
rect 43204 11386 43260 11398
rect 42588 11302 42644 11340
rect 42084 11284 42140 11294
rect 42084 11282 42308 11284
rect 42084 11230 42086 11282
rect 42138 11230 42308 11282
rect 42084 11228 42308 11230
rect 42084 11218 42140 11228
rect 42252 11172 42308 11228
rect 42812 11172 42868 11342
rect 42252 11116 42868 11172
rect 42924 11284 42980 11294
rect 41692 10658 41748 10668
rect 41580 10612 41636 10650
rect 41580 10546 41636 10556
rect 41356 9826 41468 9828
rect 41356 9774 41358 9826
rect 41410 9774 41468 9826
rect 41356 9772 41468 9774
rect 41356 9762 41412 9772
rect 41468 9734 41524 9772
rect 41580 10388 41636 10398
rect 41132 9156 41188 9166
rect 41132 9062 41188 9100
rect 40796 8306 40852 8316
rect 41580 8260 41636 10332
rect 42644 10276 42700 10286
rect 41916 9994 41972 10006
rect 41916 9942 41918 9994
rect 41970 9942 41972 9994
rect 41692 9828 41748 9838
rect 41692 9734 41748 9772
rect 41804 8932 41860 8942
rect 41804 8370 41860 8876
rect 41916 8708 41972 9942
rect 42644 9938 42700 10220
rect 42644 9886 42646 9938
rect 42698 9886 42700 9938
rect 42644 9874 42700 9886
rect 42028 9826 42084 9838
rect 42028 9774 42030 9826
rect 42082 9774 42084 9826
rect 42028 9268 42084 9774
rect 42924 9828 42980 11228
rect 43372 11282 43428 11294
rect 43372 11230 43374 11282
rect 43426 11230 43428 11282
rect 43372 10612 43428 11230
rect 43484 10722 43540 11788
rect 43820 11732 43876 11742
rect 43484 10670 43486 10722
rect 43538 10670 43540 10722
rect 43484 10658 43540 10670
rect 43596 11394 43652 11406
rect 43596 11342 43598 11394
rect 43650 11342 43652 11394
rect 43372 10546 43428 10556
rect 43372 10388 43428 10398
rect 43596 10388 43652 11342
rect 43820 11366 43876 11676
rect 43820 11314 43822 11366
rect 43874 11314 43876 11366
rect 43820 11302 43876 11314
rect 44044 10724 44100 10734
rect 44044 10630 44100 10668
rect 43428 10332 43652 10388
rect 44100 10500 44156 10510
rect 44268 10500 44324 12002
rect 44156 10444 44324 10500
rect 44492 10948 44548 12348
rect 44940 12180 44996 12190
rect 44940 12086 44996 12124
rect 45164 12180 45220 12190
rect 45276 12180 45332 13244
rect 45388 12964 45444 14700
rect 45500 14530 45556 14542
rect 45500 14478 45502 14530
rect 45554 14478 45556 14530
rect 45500 13412 45556 14478
rect 45500 13346 45556 13356
rect 45388 12962 45556 12964
rect 45388 12910 45390 12962
rect 45442 12910 45556 12962
rect 45388 12908 45556 12910
rect 45388 12898 45444 12908
rect 45164 12178 45332 12180
rect 45164 12126 45166 12178
rect 45218 12126 45332 12178
rect 45164 12124 45332 12126
rect 45388 12292 45444 12302
rect 45388 12234 45444 12236
rect 45388 12182 45390 12234
rect 45442 12182 45444 12234
rect 45164 12068 45220 12124
rect 45164 12002 45220 12012
rect 44660 11956 44716 11966
rect 44660 11862 44716 11900
rect 45388 11361 45444 12182
rect 45500 12068 45556 12908
rect 45612 12292 45668 14924
rect 46172 14644 46228 15990
rect 46284 14756 46340 16156
rect 47068 16100 47124 16110
rect 46440 16058 46496 16070
rect 46440 16006 46442 16058
rect 46494 16006 46496 16058
rect 47068 16006 47124 16044
rect 47292 16100 47348 16110
rect 47292 16006 47348 16044
rect 46440 15540 46496 16006
rect 46620 15986 46676 15998
rect 47572 15988 47628 15998
rect 46620 15934 46622 15986
rect 46674 15934 46676 15986
rect 46620 15652 46676 15934
rect 46620 15586 46676 15596
rect 47404 15986 47628 15988
rect 47404 15934 47574 15986
rect 47626 15934 47628 15986
rect 47404 15932 47628 15934
rect 46396 15484 46496 15540
rect 46396 15204 46452 15484
rect 47404 15204 47460 15932
rect 47572 15922 47628 15932
rect 47516 15652 47572 15662
rect 47516 15314 47572 15596
rect 47516 15262 47518 15314
rect 47570 15262 47572 15314
rect 47516 15250 47572 15262
rect 46396 15138 46452 15148
rect 47292 15148 47460 15204
rect 47740 15148 47796 16156
rect 46844 14980 46900 14990
rect 47292 14980 47348 15148
rect 46284 14700 46620 14756
rect 46172 14578 46228 14588
rect 46564 14642 46620 14700
rect 46564 14590 46566 14642
rect 46618 14590 46620 14642
rect 46844 14698 46900 14924
rect 46844 14646 46846 14698
rect 46898 14646 46900 14698
rect 46844 14634 46900 14646
rect 46956 14924 47348 14980
rect 47516 15092 47796 15148
rect 46564 14578 46620 14590
rect 45836 14532 45892 14542
rect 45836 14438 45892 14476
rect 46956 14530 47012 14924
rect 47516 14644 47572 15092
rect 47852 14654 47908 18508
rect 48076 17554 48132 17566
rect 48076 17502 48078 17554
rect 48130 17502 48132 17554
rect 46956 14478 46958 14530
rect 47010 14478 47012 14530
rect 46956 14466 47012 14478
rect 47292 14588 47572 14644
rect 47796 14642 47908 14654
rect 47796 14590 47798 14642
rect 47850 14590 47908 14642
rect 47796 14588 47908 14590
rect 47964 16882 48020 16894
rect 47964 16830 47966 16882
rect 48018 16830 48020 16882
rect 47964 16100 48020 16830
rect 48076 16882 48132 17502
rect 48076 16830 48078 16882
rect 48130 16830 48132 16882
rect 48076 16548 48132 16830
rect 48076 16482 48132 16492
rect 48188 16222 48244 20132
rect 48132 16210 48244 16222
rect 48132 16158 48134 16210
rect 48186 16158 48244 16210
rect 48132 16156 48244 16158
rect 48300 19908 48356 19918
rect 48132 16146 48188 16156
rect 48300 16085 48356 19852
rect 47292 14530 47348 14588
rect 47796 14578 47852 14588
rect 47292 14478 47294 14530
rect 47346 14478 47348 14530
rect 45948 14308 46004 14318
rect 45724 13860 45780 13870
rect 45724 13746 45780 13804
rect 45724 13694 45726 13746
rect 45778 13694 45780 13746
rect 45724 13682 45780 13694
rect 45948 13748 46004 14252
rect 46508 13860 46564 13870
rect 46284 13748 46340 13758
rect 46004 13746 46340 13748
rect 46004 13694 46286 13746
rect 46338 13694 46340 13746
rect 46004 13692 46340 13694
rect 45948 13654 46004 13692
rect 46284 13682 46340 13692
rect 46508 13746 46564 13804
rect 46508 13694 46510 13746
rect 46562 13694 46564 13746
rect 46508 13682 46564 13694
rect 47292 13746 47348 14478
rect 47964 13860 48020 16044
rect 48188 16029 48356 16085
rect 48412 16212 48468 16222
rect 48188 14476 48244 16029
rect 48300 15316 48356 15326
rect 48300 15222 48356 15260
rect 48132 14420 48244 14476
rect 48132 13970 48188 14420
rect 48244 14308 48300 14318
rect 48412 14308 48468 16156
rect 48244 14306 48468 14308
rect 48244 14254 48246 14306
rect 48298 14254 48468 14306
rect 48244 14252 48468 14254
rect 48244 14242 48300 14252
rect 48132 13918 48134 13970
rect 48186 13918 48188 13970
rect 48132 13906 48188 13918
rect 47852 13804 48020 13860
rect 47292 13694 47294 13746
rect 47346 13694 47348 13746
rect 47292 13682 47348 13694
rect 47516 13746 47572 13758
rect 47516 13694 47518 13746
rect 47570 13694 47572 13746
rect 45724 13578 45780 13590
rect 45724 13526 45726 13578
rect 45778 13526 45780 13578
rect 47292 13578 47348 13590
rect 45724 12740 45780 13526
rect 46788 13524 46844 13534
rect 45724 12674 45780 12684
rect 45836 13522 46844 13524
rect 45836 13470 46790 13522
rect 46842 13470 46844 13522
rect 45836 13468 46844 13470
rect 45612 12226 45668 12236
rect 45836 12234 45892 13468
rect 46788 13458 46844 13468
rect 47292 13526 47294 13578
rect 47346 13526 47348 13578
rect 46172 12964 46228 12974
rect 46172 12962 46340 12964
rect 46172 12910 46174 12962
rect 46226 12910 46340 12962
rect 46172 12908 46340 12910
rect 46172 12898 46228 12908
rect 45836 12182 45838 12234
rect 45890 12182 45892 12234
rect 45836 12170 45892 12182
rect 46172 12740 46228 12750
rect 46172 12234 46228 12684
rect 46172 12182 46174 12234
rect 46226 12182 46228 12234
rect 46172 12170 46228 12182
rect 46284 12068 46340 12908
rect 46482 12628 46538 12638
rect 46482 12218 46538 12572
rect 47292 12628 47348 13526
rect 47292 12562 47348 12572
rect 47516 12516 47572 13694
rect 47516 12450 47572 12460
rect 47628 13524 47684 13534
rect 46482 12166 46484 12218
rect 46536 12166 46538 12218
rect 46482 12154 46538 12166
rect 47068 12180 47124 12190
rect 47068 12086 47124 12124
rect 47292 12180 47348 12190
rect 47292 12086 47348 12124
rect 47628 12178 47684 13468
rect 47852 12180 47908 13804
rect 48076 13524 48132 13534
rect 48076 13074 48132 13468
rect 48076 13022 48078 13074
rect 48130 13022 48132 13074
rect 48076 13010 48132 13022
rect 48300 12628 48356 12638
rect 48132 12516 48188 12526
rect 47628 12126 47630 12178
rect 47682 12126 47684 12178
rect 47628 12114 47684 12126
rect 47740 12178 47908 12180
rect 47740 12126 47854 12178
rect 47906 12126 47908 12178
rect 47740 12124 47908 12126
rect 46508 12068 46564 12078
rect 45500 12012 45780 12068
rect 46284 12066 46564 12068
rect 46284 12014 46510 12066
rect 46562 12014 46564 12066
rect 46284 12012 46564 12014
rect 45388 11309 45390 11361
rect 45442 11309 45444 11361
rect 43372 10050 43428 10332
rect 43372 9998 43374 10050
rect 43426 9998 43428 10050
rect 43372 9986 43428 9998
rect 44100 9938 44156 10444
rect 44100 9886 44102 9938
rect 44154 9886 44156 9938
rect 44100 9874 44156 9886
rect 42924 9762 42980 9772
rect 43708 9826 43764 9838
rect 43708 9774 43710 9826
rect 43762 9774 43764 9826
rect 42028 9202 42084 9212
rect 43708 9716 43764 9774
rect 43036 8932 43092 8942
rect 43036 8838 43092 8876
rect 41916 8652 42028 8708
rect 41804 8318 41806 8370
rect 41858 8318 41860 8370
rect 41804 8306 41860 8318
rect 41972 8314 42028 8652
rect 41412 8202 41468 8214
rect 41412 8150 41414 8202
rect 41466 8150 41468 8202
rect 41972 8262 41974 8314
rect 42026 8262 42028 8314
rect 41972 8250 42028 8262
rect 42364 8372 42420 8382
rect 43708 8372 43764 9660
rect 44492 9278 44548 10892
rect 44996 11170 45052 11182
rect 44996 11118 44998 11170
rect 45050 11118 45052 11170
rect 44996 10948 45052 11118
rect 44996 10882 45052 10892
rect 44828 10836 44884 10846
rect 44828 10052 44884 10780
rect 45388 10836 45444 11309
rect 45388 10770 45444 10780
rect 45388 10276 45444 10286
rect 45052 10052 45108 10062
rect 44828 10050 45108 10052
rect 44828 9998 45054 10050
rect 45106 9998 45108 10050
rect 44828 9996 45108 9998
rect 45052 9986 45108 9996
rect 44716 9826 44772 9838
rect 45388 9828 45444 10220
rect 45724 10276 45780 12012
rect 46508 12002 46564 12012
rect 46956 12010 47012 12022
rect 46172 11956 46228 11966
rect 45836 11844 45892 11854
rect 45836 11357 45892 11788
rect 45836 11305 45838 11357
rect 45890 11305 45892 11357
rect 45836 11293 45892 11305
rect 46172 11361 46228 11900
rect 46956 11958 46958 12010
rect 47010 11958 47012 12010
rect 46956 11844 47012 11958
rect 47740 11956 47796 12124
rect 46956 11778 47012 11788
rect 47180 11900 47796 11956
rect 47180 11618 47236 11900
rect 47180 11566 47182 11618
rect 47234 11566 47236 11618
rect 47180 11554 47236 11566
rect 46508 11508 46564 11518
rect 46172 11309 46174 11361
rect 46226 11309 46228 11361
rect 46172 11297 46228 11309
rect 46284 11506 46564 11508
rect 46284 11454 46510 11506
rect 46562 11454 46564 11506
rect 46284 11452 46564 11454
rect 45724 10210 45780 10220
rect 45836 11172 45892 11182
rect 44716 9774 44718 9826
rect 44770 9774 44772 9826
rect 44716 9716 44772 9774
rect 44716 9650 44772 9660
rect 45164 9826 45444 9828
rect 45164 9774 45390 9826
rect 45442 9774 45444 9826
rect 45164 9772 45444 9774
rect 44940 9492 44996 9502
rect 44492 9266 44604 9278
rect 44492 9214 44550 9266
rect 44602 9214 44604 9266
rect 44492 9212 44604 9214
rect 44548 9202 44604 9212
rect 41580 8166 41636 8204
rect 41412 8148 41468 8150
rect 41412 8092 41524 8148
rect 41020 7474 41076 7486
rect 41020 7422 41022 7474
rect 41074 7422 41076 7474
rect 41020 7252 41076 7422
rect 41020 7186 41076 7196
rect 41132 7474 41188 7486
rect 41132 7422 41134 7474
rect 41186 7422 41188 7474
rect 41132 7028 41188 7422
rect 41020 6972 41188 7028
rect 41300 7474 41356 7486
rect 41300 7422 41302 7474
rect 41354 7422 41356 7474
rect 41300 7028 41356 7422
rect 41020 6468 41076 6972
rect 41300 6962 41356 6972
rect 41356 6692 41412 6702
rect 41020 6402 41076 6412
rect 41188 6466 41244 6478
rect 41188 6414 41190 6466
rect 41242 6414 41244 6466
rect 41188 6244 41244 6414
rect 40684 6188 41244 6244
rect 39004 6020 39060 6030
rect 39004 5906 39060 5964
rect 39302 5944 39358 6188
rect 39004 5854 39006 5906
rect 39058 5854 39060 5906
rect 39004 5842 39060 5854
rect 39116 5908 39172 5918
rect 39302 5892 39304 5944
rect 39356 5892 39358 5944
rect 39302 5880 39358 5892
rect 39452 6020 39508 6030
rect 39116 5814 39172 5852
rect 38892 5070 38894 5122
rect 38946 5070 38948 5122
rect 38892 5058 38948 5070
rect 39004 5460 39060 5470
rect 37772 3668 37828 3678
rect 37548 3666 37828 3668
rect 37548 3614 37774 3666
rect 37826 3614 37828 3666
rect 37548 3612 37828 3614
rect 37772 3602 37828 3612
rect 37436 3469 37438 3521
rect 37490 3469 37492 3521
rect 37436 3457 37492 3469
rect 37746 3514 37802 3526
rect 37746 3462 37748 3514
rect 37800 3462 37802 3514
rect 34610 3388 34804 3444
rect 37746 3444 37802 3462
rect 37746 3378 37802 3388
rect 38108 3388 38164 3948
rect 38220 3948 38724 4004
rect 38780 4340 38836 4350
rect 38220 3554 38276 3948
rect 38780 3892 38836 4284
rect 39004 4228 39060 5404
rect 39284 5460 39340 5470
rect 39284 5178 39340 5404
rect 39116 5122 39172 5134
rect 39116 5070 39118 5122
rect 39170 5070 39172 5122
rect 39284 5126 39286 5178
rect 39338 5126 39340 5178
rect 39284 5114 39340 5126
rect 39452 5124 39508 5964
rect 41244 5921 41300 5933
rect 40012 5906 40068 5918
rect 40012 5854 40014 5906
rect 40066 5854 40068 5906
rect 39676 5796 39732 5806
rect 40012 5796 40068 5854
rect 40908 5906 40964 5918
rect 40908 5854 40910 5906
rect 40962 5854 40964 5906
rect 39676 5794 40068 5796
rect 39676 5742 39678 5794
rect 39730 5742 40068 5794
rect 39676 5740 40068 5742
rect 40180 5796 40236 5806
rect 39676 5730 39732 5740
rect 40180 5738 40236 5740
rect 40180 5686 40182 5738
rect 40234 5686 40236 5738
rect 40180 5684 40236 5686
rect 40124 5628 40236 5684
rect 40572 5796 40628 5806
rect 39116 5012 39172 5070
rect 39116 4946 39172 4956
rect 39340 4452 39396 4462
rect 39452 4452 39508 5068
rect 39788 5124 39844 5134
rect 39788 5030 39844 5068
rect 40124 5122 40180 5628
rect 40236 5460 40292 5470
rect 40236 5236 40292 5404
rect 40460 5236 40516 5246
rect 40236 5234 40516 5236
rect 40236 5182 40462 5234
rect 40514 5182 40516 5234
rect 40236 5180 40516 5182
rect 40460 5170 40516 5180
rect 40124 5070 40126 5122
rect 40178 5070 40180 5122
rect 40124 5058 40180 5070
rect 40348 5066 40404 5078
rect 40348 5014 40350 5066
rect 40402 5014 40404 5066
rect 40348 5012 40404 5014
rect 40404 4956 40516 5012
rect 40348 4946 40404 4956
rect 39340 4450 39508 4452
rect 39340 4398 39342 4450
rect 39394 4398 39508 4450
rect 39340 4396 39508 4398
rect 39340 4386 39396 4396
rect 39900 4340 39956 4350
rect 39900 4246 39956 4284
rect 40236 4338 40292 4350
rect 40236 4286 40238 4338
rect 40290 4286 40292 4338
rect 39004 4172 39228 4228
rect 38612 3836 38836 3892
rect 38612 3778 38668 3836
rect 38612 3726 38614 3778
rect 38666 3726 38668 3778
rect 38612 3714 38668 3726
rect 39172 3666 39228 4172
rect 39172 3614 39174 3666
rect 39226 3614 39228 3666
rect 39172 3602 39228 3614
rect 39788 4170 39844 4182
rect 39788 4118 39790 4170
rect 39842 4118 39844 4170
rect 38220 3502 38222 3554
rect 38274 3502 38276 3554
rect 38220 3490 38276 3502
rect 38332 3554 38388 3566
rect 38332 3502 38334 3554
rect 38386 3502 38388 3554
rect 38332 3388 38388 3502
rect 38108 3332 38388 3388
rect 39788 3444 39844 4118
rect 40236 3780 40292 4286
rect 40236 3714 40292 3724
rect 39956 3668 40012 3678
rect 39956 3574 40012 3612
rect 40292 3556 40348 3566
rect 40292 3462 40348 3500
rect 39788 3378 39844 3388
rect 40460 3388 40516 4956
rect 40572 3554 40628 5740
rect 40908 5684 40964 5854
rect 41244 5869 41246 5921
rect 41298 5869 41300 5921
rect 41244 5684 41300 5869
rect 41356 5794 41412 6636
rect 41356 5742 41358 5794
rect 41410 5742 41412 5794
rect 41356 5730 41412 5742
rect 40908 5618 40964 5628
rect 41132 5628 41300 5684
rect 41132 5460 41188 5628
rect 41468 5572 41524 8092
rect 42364 8046 42420 8316
rect 43596 8316 43764 8372
rect 43820 9042 43876 9054
rect 43820 8990 43822 9042
rect 43874 8990 43876 9042
rect 43820 8372 43876 8990
rect 43036 8202 43092 8214
rect 43036 8150 43038 8202
rect 43090 8150 43092 8202
rect 43036 8148 43092 8150
rect 43316 8202 43372 8214
rect 43316 8150 43318 8202
rect 43370 8150 43372 8202
rect 43316 8148 43372 8150
rect 43036 8082 43092 8092
rect 43148 8092 43372 8148
rect 42364 8034 42476 8046
rect 42364 7982 42422 8034
rect 42474 7982 42476 8034
rect 42364 7970 42476 7982
rect 42252 7924 42308 7934
rect 41580 7476 41636 7486
rect 41580 6802 41636 7420
rect 42252 7476 42308 7868
rect 42252 7382 42308 7420
rect 41692 7364 41748 7374
rect 41692 7270 41748 7308
rect 42364 7252 42420 7970
rect 43148 7700 43204 8092
rect 42700 7644 43204 7700
rect 43428 8036 43484 8046
rect 42588 7474 42644 7486
rect 42588 7422 42590 7474
rect 42642 7422 42644 7474
rect 42588 7364 42644 7422
rect 42588 7298 42644 7308
rect 42700 7306 42756 7644
rect 43428 7586 43484 7980
rect 43428 7534 43430 7586
rect 43482 7534 43484 7586
rect 43428 7522 43484 7534
rect 42924 7476 42980 7486
rect 42924 7382 42980 7420
rect 43148 7474 43204 7486
rect 43148 7422 43150 7474
rect 43202 7422 43204 7474
rect 41580 6750 41582 6802
rect 41634 6750 41636 6802
rect 41580 6738 41636 6750
rect 42252 7196 42420 7252
rect 42700 7254 42702 7306
rect 42754 7254 42756 7306
rect 43148 7364 43204 7422
rect 43596 7364 43652 8316
rect 43820 8306 43876 8316
rect 44130 8596 44186 8606
rect 44130 8225 44186 8540
rect 44716 8372 44772 8382
rect 43764 8202 43820 8214
rect 43764 8150 43766 8202
rect 43818 8150 43820 8202
rect 44130 8173 44132 8225
rect 44184 8173 44186 8225
rect 44130 8161 44186 8173
rect 44268 8260 44324 8270
rect 43764 8036 43820 8150
rect 43148 7298 43204 7308
rect 43484 7308 43652 7364
rect 43708 7980 43764 8036
rect 43708 7970 43820 7980
rect 43932 8148 43988 8158
rect 42700 7242 42756 7254
rect 42028 6690 42084 6702
rect 41692 6646 41748 6658
rect 41692 6594 41694 6646
rect 41746 6594 41748 6646
rect 41692 6580 41748 6594
rect 41692 6514 41748 6524
rect 42028 6638 42030 6690
rect 42082 6638 42084 6690
rect 41804 5908 41860 5918
rect 41804 5814 41860 5852
rect 41132 5394 41188 5404
rect 41244 5516 41524 5572
rect 41580 5796 41636 5806
rect 40684 5348 40740 5358
rect 40684 4452 40740 5292
rect 41244 5346 41300 5516
rect 41244 5294 41246 5346
rect 41298 5294 41300 5346
rect 41244 5282 41300 5294
rect 40796 5236 40852 5246
rect 40796 5122 40852 5180
rect 40796 5070 40798 5122
rect 40850 5070 40852 5122
rect 40796 5058 40852 5070
rect 41020 5124 41076 5134
rect 41580 5124 41636 5740
rect 42028 5572 42084 6638
rect 42140 5908 42196 5918
rect 42140 5814 42196 5852
rect 42252 5796 42308 7196
rect 43036 6802 43092 6814
rect 43036 6750 43038 6802
rect 43090 6750 43092 6802
rect 42364 6690 42420 6702
rect 42364 6638 42366 6690
rect 42418 6638 42420 6690
rect 42364 6244 42420 6638
rect 42364 6178 42420 6188
rect 42476 6690 42532 6702
rect 42476 6638 42478 6690
rect 42530 6638 42532 6690
rect 43036 6692 43092 6750
rect 42476 6468 42532 6638
rect 42644 6634 42700 6646
rect 42644 6582 42646 6634
rect 42698 6582 42700 6634
rect 43036 6626 43092 6636
rect 43148 6804 43204 6814
rect 42644 6580 42700 6582
rect 42644 6514 42700 6524
rect 42476 6020 42532 6412
rect 42476 5954 42532 5964
rect 42812 5908 42868 5918
rect 42532 5796 42588 5806
rect 42252 5794 42644 5796
rect 42252 5742 42534 5794
rect 42586 5742 42644 5794
rect 42252 5740 42644 5742
rect 42532 5730 42644 5740
rect 42028 5506 42084 5516
rect 40684 4386 40740 4396
rect 40852 3892 40908 3902
rect 40852 3610 40908 3836
rect 40572 3502 40574 3554
rect 40626 3502 40628 3554
rect 40572 3490 40628 3502
rect 40684 3556 40740 3566
rect 40852 3558 40854 3610
rect 40906 3558 40908 3610
rect 40852 3546 40908 3558
rect 41020 3554 41076 5068
rect 41487 5091 41636 5124
rect 41487 5039 41489 5091
rect 41541 5068 41636 5091
rect 41692 5124 41748 5134
rect 41541 5039 41543 5068
rect 41487 5027 41543 5039
rect 41412 4452 41468 4462
rect 41412 4394 41468 4396
rect 41412 4342 41414 4394
rect 41466 4342 41468 4394
rect 41412 4330 41468 4342
rect 41692 4394 41748 5068
rect 42364 5124 42420 5134
rect 42364 5030 42420 5068
rect 42476 5012 42532 5022
rect 41692 4342 41694 4394
rect 41746 4342 41748 4394
rect 41356 4228 41412 4238
rect 41356 4134 41412 4172
rect 40684 3442 40740 3500
rect 41020 3502 41022 3554
rect 41074 3502 41076 3554
rect 41020 3490 41076 3502
rect 41468 3892 41524 3902
rect 41468 3554 41524 3836
rect 41692 3722 41748 4342
rect 41692 3670 41694 3722
rect 41746 3670 41748 3722
rect 42196 4394 42252 4406
rect 42196 4342 42198 4394
rect 42250 4342 42252 4394
rect 42196 3778 42252 4342
rect 42476 4394 42532 4956
rect 42476 4342 42478 4394
rect 42530 4342 42532 4394
rect 42476 4330 42532 4342
rect 42588 4340 42644 5730
rect 42700 5348 42756 5358
rect 42700 5122 42756 5292
rect 42700 5070 42702 5122
rect 42754 5070 42756 5122
rect 42700 5058 42756 5070
rect 42812 5122 42868 5852
rect 43036 5684 43092 5694
rect 43148 5684 43204 6748
rect 43372 6356 43428 6366
rect 43484 6356 43540 7308
rect 43708 6692 43764 7970
rect 43932 7507 43988 8092
rect 44268 8146 44324 8204
rect 44716 8258 44772 8316
rect 44716 8206 44718 8258
rect 44770 8206 44772 8258
rect 44716 8194 44772 8206
rect 44268 8094 44270 8146
rect 44322 8094 44324 8146
rect 44268 8082 44324 8094
rect 44940 8148 44996 9436
rect 45164 8942 45220 9772
rect 45388 9762 45444 9772
rect 45836 9716 45892 11116
rect 45948 10612 46004 10622
rect 45948 10518 46004 10556
rect 46172 9940 46228 9950
rect 46284 9940 46340 11452
rect 46508 11442 46564 11452
rect 46844 11396 46900 11406
rect 46482 11354 46538 11366
rect 46482 11302 46484 11354
rect 46536 11302 46538 11354
rect 46482 11284 46538 11302
rect 46482 11218 46538 11228
rect 46732 10610 46788 10622
rect 46732 10558 46734 10610
rect 46786 10558 46788 10610
rect 46732 10276 46788 10558
rect 46732 10210 46788 10220
rect 46844 10164 46900 11340
rect 46956 11284 47012 11294
rect 46956 10442 47012 11228
rect 47068 10612 47124 10622
rect 47068 10518 47124 10556
rect 47292 10610 47348 10622
rect 47292 10558 47294 10610
rect 47346 10558 47348 10610
rect 46956 10390 46958 10442
rect 47010 10390 47012 10442
rect 46956 10378 47012 10390
rect 46844 10098 46900 10108
rect 46172 9938 46340 9940
rect 46172 9886 46174 9938
rect 46226 9886 46340 9938
rect 46172 9884 46340 9886
rect 46172 9874 46228 9884
rect 45724 9660 45892 9716
rect 45276 9044 45332 9054
rect 45276 8950 45332 8988
rect 45612 9044 45668 9054
rect 45612 8950 45668 8988
rect 45108 8930 45220 8942
rect 45108 8878 45110 8930
rect 45162 8878 45220 8930
rect 45108 8876 45220 8878
rect 45108 8372 45164 8876
rect 45108 8306 45164 8316
rect 45500 8260 45556 8270
rect 45500 8166 45556 8204
rect 44940 8082 44996 8092
rect 45724 8036 45780 9660
rect 47124 9268 47180 9278
rect 47124 9174 47180 9212
rect 46284 9044 46340 9054
rect 46620 9044 46676 9054
rect 46284 9042 46452 9044
rect 46284 8990 46286 9042
rect 46338 8990 46452 9042
rect 46284 8988 46452 8990
rect 46284 8978 46340 8988
rect 46172 8874 46228 8886
rect 46172 8822 46174 8874
rect 46226 8822 46228 8874
rect 46172 8596 46228 8822
rect 46396 8596 46452 8988
rect 46620 8950 46676 8988
rect 47292 9044 47348 10558
rect 47740 10610 47796 10622
rect 47740 10558 47742 10610
rect 47794 10558 47796 10610
rect 47740 10388 47796 10558
rect 47852 10610 47908 12124
rect 47964 12404 48020 12414
rect 47964 12068 48020 12348
rect 48132 12290 48188 12460
rect 48132 12238 48134 12290
rect 48186 12238 48188 12290
rect 48132 12226 48188 12238
rect 47964 12012 48132 12068
rect 47964 11508 48020 11518
rect 47964 11414 48020 11452
rect 48076 11284 48132 12012
rect 47852 10558 47854 10610
rect 47906 10558 47908 10610
rect 47852 10546 47908 10558
rect 47964 11228 48132 11284
rect 48300 11394 48356 12572
rect 48300 11342 48302 11394
rect 48354 11342 48356 11394
rect 47964 10388 48020 11228
rect 48300 11172 48356 11342
rect 48300 11106 48356 11116
rect 48132 10612 48188 10622
rect 48132 10518 48188 10556
rect 47740 10332 48020 10388
rect 47628 10164 47684 10174
rect 47684 10108 47796 10164
rect 47628 10098 47684 10108
rect 47572 9828 47628 9838
rect 47572 9266 47628 9772
rect 47572 9214 47574 9266
rect 47626 9214 47628 9266
rect 47572 9202 47628 9214
rect 46396 8540 46676 8596
rect 46172 8530 46228 8540
rect 45724 7980 46116 8036
rect 43932 7455 43934 7507
rect 43986 7455 43988 7507
rect 44212 7530 44268 7542
rect 44212 7478 44214 7530
rect 44266 7478 44268 7530
rect 44212 7476 44268 7478
rect 44660 7530 44716 7542
rect 44660 7478 44662 7530
rect 44714 7478 44716 7530
rect 44660 7476 44716 7478
rect 43932 6804 43988 7455
rect 44044 7420 44268 7476
rect 44380 7420 44716 7476
rect 44940 7514 45040 7588
rect 44940 7462 44986 7514
rect 45038 7462 45040 7514
rect 44940 7450 45040 7462
rect 44044 6858 44100 7420
rect 44044 6806 44046 6858
rect 44098 6806 44100 6858
rect 44044 6794 44100 6806
rect 43932 6738 43988 6748
rect 43428 6300 43540 6356
rect 43596 6690 43764 6692
rect 43596 6638 43710 6690
rect 43762 6638 43764 6690
rect 43596 6636 43764 6638
rect 43372 5906 43428 6300
rect 43372 5854 43374 5906
rect 43426 5854 43428 5906
rect 43372 5842 43428 5854
rect 43596 5906 43652 6636
rect 43708 6626 43764 6636
rect 43820 6692 43876 6702
rect 43596 5854 43598 5906
rect 43650 5854 43652 5906
rect 43596 5842 43652 5854
rect 43708 5908 43764 5918
rect 43820 5908 43876 6636
rect 44044 6692 44100 6702
rect 44044 6598 44100 6636
rect 44380 6132 44436 7420
rect 44940 7140 44996 7450
rect 45052 7364 45108 7374
rect 45052 7270 45108 7308
rect 45612 7364 45668 7374
rect 45612 7362 45780 7364
rect 45612 7310 45614 7362
rect 45666 7310 45780 7362
rect 45612 7308 45780 7310
rect 45612 7298 45668 7308
rect 44940 7074 44996 7084
rect 43988 6076 44436 6132
rect 44716 6804 44772 6814
rect 43988 6018 44044 6076
rect 43988 5966 43990 6018
rect 44042 5966 44044 6018
rect 43988 5954 44044 5966
rect 43708 5906 43876 5908
rect 43708 5854 43710 5906
rect 43762 5854 43876 5906
rect 43708 5852 43876 5854
rect 43708 5842 43764 5852
rect 43036 5682 43204 5684
rect 43036 5630 43038 5682
rect 43090 5630 43204 5682
rect 43036 5628 43204 5630
rect 43036 5618 43092 5628
rect 42812 5070 42814 5122
rect 42866 5070 42868 5122
rect 42812 5058 42868 5070
rect 42924 5572 42980 5582
rect 42924 5134 42980 5516
rect 42924 5122 43034 5134
rect 42924 5070 42980 5122
rect 43032 5070 43034 5122
rect 42924 5068 43034 5070
rect 42978 5058 43034 5068
rect 43148 5012 43204 5628
rect 43372 5234 43428 5246
rect 43372 5182 43374 5234
rect 43426 5182 43428 5234
rect 43372 5124 43428 5182
rect 43820 5236 43876 5246
rect 43820 5142 43876 5180
rect 43372 5058 43428 5068
rect 43932 5124 43988 5134
rect 43932 5055 43934 5068
rect 43986 5055 43988 5068
rect 44268 5124 44324 6076
rect 44716 5962 44772 6748
rect 44828 6692 44884 6702
rect 44828 6690 45220 6692
rect 44828 6638 44830 6690
rect 44882 6638 45220 6690
rect 44828 6636 45220 6638
rect 44828 6626 44884 6636
rect 44996 6468 45052 6478
rect 44996 6374 45052 6412
rect 44716 5910 44718 5962
rect 44770 5910 44772 5962
rect 44716 5898 44772 5910
rect 44996 5962 45052 5974
rect 44996 5910 44998 5962
rect 45050 5910 45052 5962
rect 44996 5908 45052 5910
rect 44828 5852 45052 5908
rect 44716 5236 44772 5246
rect 44268 5122 44660 5124
rect 44268 5070 44270 5122
rect 44322 5070 44660 5122
rect 44268 5068 44660 5070
rect 44268 5058 44324 5068
rect 43932 5030 43988 5055
rect 43148 4946 43204 4956
rect 43708 4452 43764 4462
rect 42700 4340 42756 4350
rect 42588 4338 42756 4340
rect 42588 4286 42702 4338
rect 42754 4286 42756 4338
rect 42588 4284 42756 4286
rect 42196 3726 42198 3778
rect 42250 3726 42252 3778
rect 42196 3714 42252 3726
rect 42588 3892 42644 3902
rect 41692 3658 41748 3670
rect 41468 3502 41470 3554
rect 41522 3502 41524 3554
rect 41468 3490 41524 3502
rect 41692 3556 41748 3566
rect 41692 3462 41748 3500
rect 42476 3556 42532 3566
rect 42476 3462 42532 3500
rect 42588 3554 42644 3836
rect 42700 3668 42756 4284
rect 43484 4228 43540 4238
rect 43484 4134 43540 4172
rect 43708 3722 43764 4396
rect 42700 3602 42756 3612
rect 43092 3668 43148 3678
rect 43708 3670 43710 3722
rect 43762 3670 43764 3722
rect 43708 3658 43764 3670
rect 44044 3780 44100 3790
rect 43092 3574 43148 3612
rect 42588 3502 42590 3554
rect 42642 3502 42644 3554
rect 42588 3490 42644 3502
rect 43708 3556 43764 3566
rect 43708 3462 43764 3500
rect 44044 3554 44100 3724
rect 44044 3502 44046 3554
rect 44098 3502 44100 3554
rect 44044 3490 44100 3502
rect 44492 3556 44548 3566
rect 44604 3556 44660 5068
rect 44716 5122 44772 5180
rect 44716 5070 44718 5122
rect 44770 5070 44772 5122
rect 44716 5058 44772 5070
rect 44828 3722 44884 5852
rect 45052 5348 45108 5358
rect 45164 5348 45220 6636
rect 45388 6690 45444 6702
rect 45388 6638 45390 6690
rect 45442 6638 45444 6690
rect 45388 5572 45444 6638
rect 45612 6692 45668 6702
rect 45612 6598 45668 6636
rect 45500 6468 45556 6478
rect 45500 5962 45556 6412
rect 45724 6468 45780 7308
rect 45724 6402 45780 6412
rect 45892 6578 45948 6590
rect 45892 6526 45894 6578
rect 45946 6526 45948 6578
rect 45892 6244 45948 6526
rect 45892 6178 45948 6188
rect 45500 5910 45502 5962
rect 45554 5910 45556 5962
rect 45948 6018 46004 6030
rect 45948 5966 45950 6018
rect 46002 5966 46004 6018
rect 45500 5898 45556 5910
rect 45810 5939 45866 5951
rect 45810 5908 45812 5939
rect 45864 5908 45866 5939
rect 45810 5842 45866 5852
rect 45444 5516 45668 5572
rect 45388 5506 45444 5516
rect 45052 5346 45220 5348
rect 45052 5294 45054 5346
rect 45106 5294 45220 5346
rect 45052 5292 45220 5294
rect 45388 5348 45444 5358
rect 44828 3670 44830 3722
rect 44882 3670 44884 3722
rect 44828 3658 44884 3670
rect 44940 5124 44996 5134
rect 44492 3554 44660 3556
rect 44492 3502 44494 3554
rect 44546 3502 44660 3554
rect 44492 3500 44660 3502
rect 44716 3556 44772 3566
rect 44940 3556 44996 5068
rect 45052 3892 45108 5292
rect 45388 4452 45444 5292
rect 45612 5234 45668 5516
rect 45612 5182 45614 5234
rect 45666 5182 45668 5234
rect 45612 5170 45668 5182
rect 45948 5236 46004 5966
rect 45948 5170 46004 5180
rect 46060 5086 46116 7980
rect 46620 7700 46676 8540
rect 46396 7644 46676 7700
rect 46396 7140 46452 7644
rect 47068 7140 47124 7150
rect 46396 7084 46732 7140
rect 46284 7028 46340 7038
rect 46284 6690 46340 6972
rect 46284 6638 46286 6690
rect 46338 6638 46340 6690
rect 46284 6626 46340 6638
rect 46396 6692 46452 6702
rect 46452 6636 46564 6692
rect 46396 6598 46452 6636
rect 46396 6468 46452 6478
rect 46396 5906 46452 6412
rect 46396 5854 46398 5906
rect 46450 5854 46452 5906
rect 46396 5842 46452 5854
rect 46508 5572 46564 6636
rect 46676 6690 46732 7084
rect 47068 6858 47124 7084
rect 47068 6806 47070 6858
rect 47122 6806 47124 6858
rect 47068 6794 47124 6806
rect 47180 6692 47236 6702
rect 46676 6638 46678 6690
rect 46730 6638 46732 6690
rect 46676 6626 46732 6638
rect 46956 6690 47236 6692
rect 46956 6638 47182 6690
rect 47234 6638 47236 6690
rect 46956 6636 47236 6638
rect 47292 6692 47348 8988
rect 47404 8146 47460 8158
rect 47404 8094 47406 8146
rect 47458 8094 47460 8146
rect 47404 7028 47460 8094
rect 47516 7364 47572 7374
rect 47516 7270 47572 7308
rect 47404 6962 47460 6972
rect 47516 6692 47572 6702
rect 47292 6690 47572 6692
rect 47292 6638 47518 6690
rect 47570 6638 47572 6690
rect 47292 6636 47572 6638
rect 46956 6030 47012 6636
rect 47180 6626 47236 6636
rect 46900 6018 47012 6030
rect 46900 5966 46902 6018
rect 46954 5966 47012 6018
rect 46900 5964 47012 5966
rect 47404 6244 47460 6254
rect 46900 5954 46956 5964
rect 46620 5906 46676 5918
rect 46620 5854 46622 5906
rect 46674 5854 46676 5906
rect 46620 5572 46676 5854
rect 47292 5908 47348 5918
rect 47292 5738 47348 5852
rect 47404 5906 47460 6188
rect 47404 5854 47406 5906
rect 47458 5854 47460 5906
rect 47404 5842 47460 5854
rect 47516 5908 47572 6636
rect 47628 5908 47684 5918
rect 47516 5906 47684 5908
rect 47516 5854 47630 5906
rect 47682 5854 47684 5906
rect 47516 5852 47684 5854
rect 47628 5842 47684 5852
rect 47292 5686 47294 5738
rect 47346 5686 47348 5738
rect 47292 5674 47348 5686
rect 45836 5030 46116 5086
rect 46396 5516 46676 5572
rect 45388 4450 45780 4452
rect 45388 4398 45390 4450
rect 45442 4398 45780 4450
rect 45388 4396 45780 4398
rect 45388 4386 45444 4396
rect 45724 4338 45780 4396
rect 45724 4286 45726 4338
rect 45778 4286 45780 4338
rect 45724 4274 45780 4286
rect 45052 3826 45108 3836
rect 45836 3678 45892 5030
rect 45948 4340 46004 4350
rect 46396 4340 46452 5516
rect 47516 5236 47572 5246
rect 47516 5142 47572 5180
rect 47740 4900 47796 10108
rect 47852 9940 47908 10332
rect 48076 9940 48132 9950
rect 47852 9938 48132 9940
rect 47852 9886 48078 9938
rect 48130 9886 48132 9938
rect 47852 9884 48132 9886
rect 48076 9874 48132 9884
rect 48244 9268 48300 9278
rect 48524 9268 48580 20132
rect 48244 9266 48580 9268
rect 48244 9214 48246 9266
rect 48298 9214 48580 9266
rect 48244 9212 48580 9214
rect 48636 17556 48692 17566
rect 48244 9202 48300 9212
rect 48636 9044 48692 17500
rect 48188 8988 48692 9044
rect 47964 8034 48020 8046
rect 47964 7982 47966 8034
rect 48018 7982 48020 8034
rect 47964 6916 48020 7982
rect 47964 6850 48020 6860
rect 48188 6702 48244 8988
rect 48300 8258 48356 8270
rect 48300 8206 48302 8258
rect 48354 8206 48356 8258
rect 48300 8148 48356 8206
rect 48300 7700 48356 8092
rect 48300 7634 48356 7644
rect 48132 6690 48244 6702
rect 48132 6638 48134 6690
rect 48186 6638 48244 6690
rect 48132 6636 48244 6638
rect 48300 7474 48356 7486
rect 48300 7422 48302 7474
rect 48354 7422 48356 7474
rect 48132 6626 48188 6636
rect 48300 5806 48356 7422
rect 48244 5794 48356 5806
rect 48244 5742 48246 5794
rect 48298 5742 48356 5794
rect 48244 5730 48356 5742
rect 48300 5122 48356 5730
rect 48300 5070 48302 5122
rect 48354 5070 48356 5122
rect 47068 4844 47964 4900
rect 46732 4340 46788 4350
rect 45948 4338 46788 4340
rect 45948 4286 45950 4338
rect 46002 4286 46734 4338
rect 46786 4286 46788 4338
rect 45948 4284 46788 4286
rect 45948 4274 46004 4284
rect 46732 4274 46788 4284
rect 47068 4338 47124 4844
rect 47908 4562 47964 4844
rect 47908 4510 47910 4562
rect 47962 4510 47964 4562
rect 47908 4498 47964 4510
rect 47068 4286 47070 4338
rect 47122 4286 47124 4338
rect 47068 4274 47124 4286
rect 47460 4226 47516 4238
rect 47460 4174 47462 4226
rect 47514 4174 47516 4226
rect 46228 4114 46284 4126
rect 46228 4062 46230 4114
rect 46282 4062 46284 4114
rect 45332 3668 45388 3678
rect 45332 3574 45388 3612
rect 45780 3666 45892 3678
rect 45780 3614 45782 3666
rect 45834 3614 45892 3666
rect 45780 3612 45892 3614
rect 46060 4004 46116 4014
rect 45780 3602 45836 3612
rect 44716 3554 44996 3556
rect 44716 3502 44718 3554
rect 44770 3502 44996 3554
rect 44716 3500 44996 3502
rect 44492 3490 44548 3500
rect 44716 3490 44772 3500
rect 40684 3390 40686 3442
rect 40738 3390 40740 3442
rect 40684 3388 40740 3390
rect 40460 3332 40740 3388
rect 46060 3332 46116 3948
rect 46228 3556 46284 4062
rect 47460 3780 47516 4174
rect 47460 3714 47516 3724
rect 46676 3668 46732 3678
rect 46676 3574 46732 3612
rect 47572 3668 47628 3678
rect 47572 3574 47628 3612
rect 48020 3668 48076 3678
rect 48020 3574 48076 3612
rect 48300 3668 48356 5070
rect 48300 3602 48356 3612
rect 46228 3490 46284 3500
rect 46228 3332 46284 3342
rect 46060 3330 46284 3332
rect 46060 3278 46230 3330
rect 46282 3278 46284 3330
rect 46060 3276 46284 3278
rect 46228 3266 46284 3276
rect 28924 2706 28980 2716
<< via2 >>
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 2380 45612 2436 45668
rect 3108 45666 3164 45668
rect 3108 45614 3110 45666
rect 3110 45614 3162 45666
rect 3162 45614 3164 45666
rect 3108 45612 3164 45614
rect 4564 45666 4620 45668
rect 2660 45218 2716 45220
rect 2660 45166 2662 45218
rect 2662 45166 2714 45218
rect 2714 45166 2716 45218
rect 2660 45164 2716 45166
rect 1876 43426 1932 43428
rect 1876 43374 1878 43426
rect 1878 43374 1930 43426
rect 1930 43374 1932 43426
rect 1876 43372 1932 43374
rect 1484 42476 1540 42532
rect 28 25228 84 25284
rect 1932 42530 1988 42532
rect 1932 42478 1934 42530
rect 1934 42478 1986 42530
rect 1986 42478 1988 42530
rect 1932 42476 1988 42478
rect 1596 42140 1652 42196
rect 4564 45614 4566 45666
rect 4566 45614 4618 45666
rect 4618 45614 4620 45666
rect 4564 45612 4620 45614
rect 4564 45388 4620 45444
rect 6860 45836 6916 45892
rect 4452 45276 4508 45332
rect 3724 44940 3780 44996
rect 6692 45666 6748 45668
rect 6692 45614 6694 45666
rect 6694 45614 6746 45666
rect 6746 45614 6748 45666
rect 6692 45612 6748 45614
rect 6300 45500 6356 45556
rect 5012 45276 5068 45332
rect 6188 45388 6244 45444
rect 4004 44994 4060 44996
rect 4004 44942 4006 44994
rect 4006 44942 4058 44994
rect 4058 44942 4060 44994
rect 4004 44940 4060 44942
rect 3556 44828 3612 44884
rect 4900 44994 4956 44996
rect 4900 44942 4902 44994
rect 4902 44942 4954 44994
rect 4954 44942 4956 44994
rect 4900 44940 4956 44942
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4284 43932 4340 43988
rect 4732 44044 4788 44100
rect 1988 41298 2044 41300
rect 1988 41246 1990 41298
rect 1990 41246 2042 41298
rect 2042 41246 2044 41298
rect 1988 41244 2044 41246
rect 1988 40514 2044 40516
rect 1988 40462 1990 40514
rect 1990 40462 2042 40514
rect 2042 40462 2044 40514
rect 1988 40460 2044 40462
rect 1820 40236 1876 40292
rect 1596 39004 1652 39060
rect 1596 33346 1652 33348
rect 1596 33294 1598 33346
rect 1598 33294 1650 33346
rect 1650 33294 1652 33346
rect 1596 33292 1652 33294
rect 3052 43596 3108 43652
rect 4060 43650 4116 43652
rect 4060 43598 4062 43650
rect 4062 43598 4114 43650
rect 4114 43598 4116 43650
rect 4060 43596 4116 43598
rect 4396 43596 4452 43652
rect 4956 43708 5012 43764
rect 2604 42924 2660 42980
rect 2772 42924 2828 42980
rect 3668 43260 3724 43316
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 5068 43484 5124 43540
rect 7308 45890 7364 45892
rect 7308 45838 7310 45890
rect 7310 45838 7362 45890
rect 7362 45838 7364 45890
rect 7308 45836 7364 45838
rect 8260 45500 8316 45556
rect 9212 45612 9268 45668
rect 9828 45666 9884 45668
rect 9828 45614 9830 45666
rect 9830 45614 9882 45666
rect 9882 45614 9884 45666
rect 9828 45612 9884 45614
rect 9772 45388 9828 45444
rect 9212 45052 9268 45108
rect 5964 44044 6020 44100
rect 5852 43820 5908 43876
rect 5180 43260 5236 43316
rect 4956 43036 5012 43092
rect 9100 44380 9156 44436
rect 8428 44322 8484 44324
rect 7084 44044 7140 44100
rect 7084 43596 7140 43652
rect 7420 43525 7422 43540
rect 7422 43525 7474 43540
rect 7474 43525 7476 43540
rect 7420 43484 7476 43525
rect 7756 43538 7812 43540
rect 7756 43486 7758 43538
rect 7758 43486 7810 43538
rect 7810 43486 7812 43538
rect 7756 43484 7812 43486
rect 5684 43036 5740 43092
rect 6412 43036 6468 43092
rect 3220 42140 3276 42196
rect 2604 41804 2660 41860
rect 2604 41244 2660 41300
rect 2716 41186 2772 41188
rect 2716 41134 2718 41186
rect 2718 41134 2770 41186
rect 2770 41134 2772 41186
rect 2716 41132 2772 41134
rect 2884 40684 2940 40740
rect 3388 41132 3444 41188
rect 2436 40236 2492 40292
rect 2604 40348 2660 40404
rect 3388 40236 3444 40292
rect 3948 42476 4004 42532
rect 5292 42812 5348 42868
rect 4676 42476 4732 42532
rect 4284 41970 4340 41972
rect 4284 41918 4286 41970
rect 4286 41918 4338 41970
rect 4338 41918 4340 41970
rect 4284 41916 4340 41918
rect 5087 41804 5143 41860
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 5964 42476 6020 42532
rect 5964 41970 6020 41972
rect 5964 41918 5966 41970
rect 5966 41918 6018 41970
rect 6018 41918 6020 41970
rect 5964 41916 6020 41918
rect 6524 42812 6580 42868
rect 7084 43148 7140 43204
rect 7980 44044 8036 44100
rect 8428 44270 8430 44322
rect 8430 44270 8482 44322
rect 8482 44270 8484 44322
rect 8428 44268 8484 44270
rect 8540 43708 8596 43764
rect 7868 43148 7924 43204
rect 8764 43148 8820 43204
rect 8876 43484 8932 43540
rect 6300 41970 6356 41972
rect 6300 41918 6302 41970
rect 6302 41918 6354 41970
rect 6354 41918 6356 41970
rect 6300 41916 6356 41918
rect 6188 41804 6244 41860
rect 6860 41692 6916 41748
rect 7084 41804 7140 41860
rect 6188 41580 6244 41636
rect 3836 40572 3892 40628
rect 4396 40460 4452 40516
rect 4004 40236 4060 40292
rect 4172 40236 4228 40292
rect 5180 40460 5236 40516
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 3500 39116 3556 39172
rect 4060 39564 4116 39620
rect 3948 39116 4004 39172
rect 3444 38220 3500 38276
rect 2996 38162 3052 38164
rect 2996 38110 2998 38162
rect 2998 38110 3050 38162
rect 3050 38110 3052 38162
rect 2996 38108 3052 38110
rect 3836 38220 3892 38276
rect 5068 39676 5124 39732
rect 4844 39564 4900 39620
rect 5348 40402 5404 40404
rect 5348 40350 5350 40402
rect 5350 40350 5402 40402
rect 5402 40350 5404 40402
rect 5348 40348 5404 40350
rect 4676 39004 4732 39060
rect 5180 38946 5236 38948
rect 5180 38894 5182 38946
rect 5182 38894 5234 38946
rect 5234 38894 5236 38946
rect 5180 38892 5236 38894
rect 4676 38722 4732 38724
rect 4676 38670 4678 38722
rect 4678 38670 4730 38722
rect 4730 38670 4732 38722
rect 4676 38668 4732 38670
rect 5516 38668 5572 38724
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 3948 38108 4004 38164
rect 2604 38050 2660 38052
rect 2604 37998 2606 38050
rect 2606 37998 2658 38050
rect 2658 37998 2660 38050
rect 2604 37996 2660 37998
rect 3780 38050 3836 38052
rect 3780 37998 3782 38050
rect 3782 37998 3834 38050
rect 3834 37998 3836 38050
rect 3780 37996 3836 37998
rect 2604 36482 2660 36484
rect 2604 36430 2606 36482
rect 2606 36430 2658 36482
rect 2658 36430 2660 36482
rect 2604 36428 2660 36430
rect 2660 35308 2716 35364
rect 3892 36482 3948 36484
rect 3892 36430 3894 36482
rect 3894 36430 3946 36482
rect 3946 36430 3948 36482
rect 3892 36428 3948 36430
rect 3612 35756 3668 35812
rect 3500 35308 3556 35364
rect 2604 34412 2660 34468
rect 2156 33292 2212 33348
rect 1596 32732 1652 32788
rect 3164 34914 3220 34916
rect 3164 34862 3166 34914
rect 3166 34862 3218 34914
rect 3218 34862 3220 34914
rect 3164 34860 3220 34862
rect 4284 37266 4340 37268
rect 4284 37214 4286 37266
rect 4286 37214 4338 37266
rect 4338 37214 4340 37266
rect 4284 37212 4340 37214
rect 4732 37100 4788 37156
rect 6412 40684 6468 40740
rect 6244 40514 6300 40516
rect 6244 40462 6246 40514
rect 6246 40462 6298 40514
rect 6298 40462 6300 40514
rect 6244 40460 6300 40462
rect 5852 40236 5908 40292
rect 5852 39788 5908 39844
rect 6300 39730 6356 39732
rect 6300 39678 6302 39730
rect 6302 39678 6354 39730
rect 6354 39678 6356 39730
rect 6300 39676 6356 39678
rect 6076 39618 6132 39620
rect 6076 39566 6078 39618
rect 6078 39566 6130 39618
rect 6130 39566 6132 39618
rect 6076 39564 6132 39566
rect 7532 41580 7588 41636
rect 7700 41970 7756 41972
rect 7700 41918 7702 41970
rect 7702 41918 7754 41970
rect 7754 41918 7756 41970
rect 7700 41916 7756 41918
rect 6972 40908 7028 40964
rect 7532 40402 7588 40404
rect 7532 40350 7534 40402
rect 7534 40350 7586 40402
rect 7586 40350 7588 40402
rect 7532 40348 7588 40350
rect 8988 43036 9044 43092
rect 9436 44380 9492 44436
rect 9660 44322 9716 44324
rect 9660 44270 9662 44322
rect 9662 44270 9714 44322
rect 9714 44270 9716 44322
rect 9660 44268 9716 44270
rect 11844 45724 11900 45780
rect 10556 45388 10612 45444
rect 10332 45106 10388 45108
rect 10332 45054 10334 45106
rect 10334 45054 10386 45106
rect 10386 45054 10388 45106
rect 10332 45052 10388 45054
rect 12236 45500 12292 45556
rect 9996 44295 10052 44324
rect 9996 44268 9998 44295
rect 9998 44268 10050 44295
rect 10050 44268 10052 44295
rect 9996 43932 10052 43988
rect 9660 43036 9716 43092
rect 9996 43148 10052 43204
rect 8932 42028 8988 42084
rect 7868 41132 7924 41188
rect 8092 41132 8148 41188
rect 8204 41916 8260 41972
rect 7756 41020 7812 41076
rect 8092 40460 8148 40516
rect 8764 41970 8820 41972
rect 8764 41918 8766 41970
rect 8766 41918 8818 41970
rect 8818 41918 8820 41970
rect 8764 41916 8820 41918
rect 8932 41356 8988 41412
rect 8764 41074 8820 41076
rect 8764 41022 8766 41074
rect 8766 41022 8818 41074
rect 8818 41022 8820 41074
rect 8764 41020 8820 41022
rect 8876 40514 8932 40516
rect 8876 40462 8878 40514
rect 8878 40462 8930 40514
rect 8930 40462 8932 40514
rect 8876 40460 8932 40462
rect 8316 40348 8372 40404
rect 8988 40348 9044 40404
rect 6468 39340 6524 39396
rect 5964 38668 6020 38724
rect 6972 38892 7028 38948
rect 7084 38834 7140 38836
rect 7084 38782 7086 38834
rect 7086 38782 7138 38834
rect 7138 38782 7140 38834
rect 7084 38780 7140 38782
rect 6748 38332 6804 38388
rect 6748 38050 6804 38052
rect 6748 37998 6750 38050
rect 6750 37998 6802 38050
rect 6802 37998 6804 38050
rect 6748 37996 6804 37998
rect 6860 37660 6916 37716
rect 5796 37548 5852 37604
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4956 37100 5012 37156
rect 4228 36482 4284 36484
rect 4228 36430 4230 36482
rect 4230 36430 4282 36482
rect 4282 36430 4284 36482
rect 4228 36428 4284 36430
rect 4844 35684 4846 35700
rect 4846 35684 4898 35700
rect 4898 35684 4900 35700
rect 4844 35644 4900 35684
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 2940 34188 2996 34244
rect 3500 34300 3556 34356
rect 3220 32786 3276 32788
rect 3220 32734 3222 32786
rect 3222 32734 3274 32786
rect 3274 32734 3276 32786
rect 3220 32732 3276 32734
rect 4060 34524 4116 34580
rect 4284 34748 4340 34804
rect 4172 34300 4228 34356
rect 4284 34188 4340 34244
rect 4732 35084 4788 35140
rect 4508 34914 4564 34916
rect 4508 34862 4510 34914
rect 4510 34862 4562 34914
rect 4562 34862 4564 34914
rect 4508 34860 4564 34862
rect 5068 36316 5124 36372
rect 6524 37548 6580 37604
rect 5964 37266 6020 37268
rect 5964 37214 5966 37266
rect 5966 37214 6018 37266
rect 6018 37214 6020 37266
rect 5964 37212 6020 37214
rect 6244 37212 6300 37268
rect 6244 36876 6300 36932
rect 5796 36594 5852 36596
rect 5796 36542 5798 36594
rect 5798 36542 5850 36594
rect 5850 36542 5852 36594
rect 5796 36540 5852 36542
rect 5628 36428 5684 36484
rect 5908 36316 5964 36372
rect 5404 35810 5460 35812
rect 5404 35758 5406 35810
rect 5406 35758 5458 35810
rect 5458 35758 5460 35810
rect 5404 35756 5460 35758
rect 5068 34860 5124 34916
rect 5180 34748 5236 34804
rect 5012 34524 5068 34580
rect 5292 34300 5348 34356
rect 4732 33964 4788 34020
rect 3668 33852 3724 33908
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4116 33292 4172 33348
rect 2940 31836 2996 31892
rect 2604 31778 2660 31780
rect 2604 31726 2606 31778
rect 2606 31726 2658 31778
rect 2658 31726 2660 31778
rect 2604 31724 2660 31726
rect 5124 33346 5180 33348
rect 5124 33294 5126 33346
rect 5126 33294 5178 33346
rect 5178 33294 5180 33346
rect 5124 33292 5180 33294
rect 4116 32786 4172 32788
rect 4116 32734 4118 32786
rect 4118 32734 4170 32786
rect 4170 32734 4172 32786
rect 4116 32732 4172 32734
rect 4172 31948 4228 32004
rect 4284 32172 4340 32228
rect 3500 31836 3556 31892
rect 3052 31724 3108 31780
rect 3612 31612 3668 31668
rect 2492 30604 2548 30660
rect 3052 30604 3108 30660
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4844 32002 4900 32004
rect 4844 31950 4846 32002
rect 4846 31950 4898 32002
rect 4898 31950 4900 32002
rect 4844 31948 4900 31950
rect 5292 31724 5348 31780
rect 4452 31612 4508 31668
rect 5124 31612 5180 31668
rect 3500 30210 3556 30212
rect 3500 30158 3502 30210
rect 3502 30158 3554 30210
rect 3554 30158 3556 30210
rect 3500 30156 3556 30158
rect 4844 30716 4900 30772
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4172 30156 4228 30212
rect 4376 30380 4432 30436
rect 2828 30044 2884 30100
rect 4620 30098 4676 30100
rect 4620 30046 4622 30098
rect 4622 30046 4674 30098
rect 4674 30046 4676 30098
rect 4620 30044 4676 30046
rect 6076 35420 6132 35476
rect 6748 37100 6804 37156
rect 6524 36540 6580 36596
rect 6636 36258 6692 36260
rect 6636 36206 6638 36258
rect 6638 36206 6690 36258
rect 6690 36206 6692 36258
rect 6636 36204 6692 36206
rect 11004 44322 11060 44324
rect 11004 44270 11006 44322
rect 11006 44270 11058 44322
rect 11058 44270 11060 44322
rect 11004 44268 11060 44270
rect 12348 45052 12404 45108
rect 12684 45388 12740 45444
rect 12796 44828 12852 44884
rect 13020 44322 13076 44324
rect 13020 44270 13022 44322
rect 13022 44270 13074 44322
rect 13074 44270 13076 44322
rect 13020 44268 13076 44270
rect 10780 43932 10836 43988
rect 10668 43708 10724 43764
rect 10220 43538 10276 43540
rect 10220 43486 10222 43538
rect 10222 43486 10274 43538
rect 10274 43486 10276 43538
rect 10220 43484 10276 43486
rect 11004 43538 11060 43540
rect 11004 43486 11006 43538
rect 11006 43486 11058 43538
rect 11058 43486 11060 43538
rect 11004 43484 11060 43486
rect 10220 43148 10276 43204
rect 10556 43036 10612 43092
rect 10108 42364 10164 42420
rect 11340 42812 11396 42868
rect 10332 41970 10388 41972
rect 10332 41918 10334 41970
rect 10334 41918 10386 41970
rect 10386 41918 10388 41970
rect 10332 41916 10388 41918
rect 10556 41804 10612 41860
rect 9884 41186 9940 41188
rect 9884 41134 9886 41186
rect 9886 41134 9938 41186
rect 9938 41134 9940 41186
rect 9884 41132 9940 41134
rect 9716 40626 9772 40628
rect 9716 40574 9718 40626
rect 9718 40574 9770 40626
rect 9770 40574 9772 40626
rect 9716 40572 9772 40574
rect 14588 45724 14644 45780
rect 17500 45724 17556 45780
rect 17164 45666 17220 45668
rect 17164 45614 17166 45666
rect 17166 45614 17218 45666
rect 17218 45614 17220 45666
rect 17164 45612 17220 45614
rect 13916 45388 13972 45444
rect 15484 45106 15540 45108
rect 15484 45054 15486 45106
rect 15486 45054 15538 45106
rect 15538 45054 15540 45106
rect 15484 45052 15540 45054
rect 16268 45106 16324 45108
rect 16268 45054 16270 45106
rect 16270 45054 16322 45106
rect 16322 45054 16324 45106
rect 16268 45052 16324 45054
rect 13468 44716 13524 44772
rect 13580 44268 13636 44324
rect 13916 44940 13972 44996
rect 16940 44940 16996 44996
rect 17500 45052 17556 45108
rect 15596 44828 15652 44884
rect 15148 44604 15204 44660
rect 11676 42812 11732 42868
rect 11340 41804 11396 41860
rect 10892 41580 10948 41636
rect 11508 41580 11564 41636
rect 13580 43596 13636 43652
rect 13448 43538 13504 43540
rect 13448 43486 13450 43538
rect 13450 43486 13502 43538
rect 13502 43486 13504 43538
rect 13448 43484 13504 43486
rect 12460 42866 12516 42868
rect 12460 42814 12462 42866
rect 12462 42814 12514 42866
rect 12514 42814 12516 42866
rect 12460 42812 12516 42814
rect 13692 43148 13748 43204
rect 13916 43260 13972 43316
rect 13580 42812 13636 42868
rect 12012 42700 12068 42756
rect 12572 42739 12628 42756
rect 12572 42700 12574 42739
rect 12574 42700 12626 42739
rect 12626 42700 12628 42739
rect 12908 42754 12964 42756
rect 12908 42702 12910 42754
rect 12910 42702 12962 42754
rect 12962 42702 12964 42754
rect 12908 42700 12964 42702
rect 13804 42754 13860 42756
rect 13804 42702 13806 42754
rect 13806 42702 13858 42754
rect 13858 42702 13860 42754
rect 13804 42700 13860 42702
rect 13916 42588 13972 42644
rect 14140 43596 14196 43652
rect 14252 43260 14308 43316
rect 14924 43820 14980 43876
rect 14476 43525 14478 43540
rect 14478 43525 14530 43540
rect 14530 43525 14532 43540
rect 14476 43484 14532 43525
rect 11900 41916 11956 41972
rect 11788 41356 11844 41412
rect 11900 41692 11956 41748
rect 10668 41244 10724 41300
rect 10892 41186 10948 41188
rect 10892 41134 10894 41186
rect 10894 41134 10946 41186
rect 10946 41134 10948 41186
rect 10892 41132 10948 41134
rect 11564 41132 11620 41188
rect 11228 40684 11284 40740
rect 10164 40626 10220 40628
rect 10164 40574 10166 40626
rect 10166 40574 10218 40626
rect 10218 40574 10220 40626
rect 10164 40572 10220 40574
rect 10892 40572 10948 40628
rect 7420 37548 7476 37604
rect 7196 37378 7252 37380
rect 7196 37326 7198 37378
rect 7198 37326 7250 37378
rect 7250 37326 7252 37378
rect 7196 37324 7252 37326
rect 7868 38668 7924 38724
rect 8764 38834 8820 38836
rect 8764 38782 8766 38834
rect 8766 38782 8818 38834
rect 8818 38782 8820 38834
rect 8764 38780 8820 38782
rect 7644 37324 7700 37380
rect 8036 37378 8092 37380
rect 8036 37326 8038 37378
rect 8038 37326 8090 37378
rect 8090 37326 8092 37378
rect 8036 37324 8092 37326
rect 8764 37436 8820 37492
rect 9044 37490 9100 37492
rect 9044 37438 9046 37490
rect 9046 37438 9098 37490
rect 9098 37438 9100 37490
rect 9044 37436 9100 37438
rect 9212 39004 9268 39060
rect 8428 37324 8484 37380
rect 8148 36876 8204 36932
rect 6972 36204 7028 36260
rect 8596 36876 8652 36932
rect 11452 40348 11508 40404
rect 11676 41020 11732 41076
rect 12292 41746 12348 41748
rect 12292 41694 12294 41746
rect 12294 41694 12346 41746
rect 12346 41694 12348 41746
rect 12292 41692 12348 41694
rect 12796 41804 12852 41860
rect 12460 41298 12516 41300
rect 12460 41246 12462 41298
rect 12462 41246 12514 41298
rect 12514 41246 12516 41298
rect 12460 41244 12516 41246
rect 12684 41244 12740 41300
rect 12012 41020 12068 41076
rect 11340 40290 11396 40292
rect 11340 40238 11342 40290
rect 11342 40238 11394 40290
rect 11394 40238 11396 40290
rect 11340 40236 11396 40238
rect 12348 40572 12404 40628
rect 12124 40236 12180 40292
rect 10332 39842 10388 39844
rect 10332 39790 10334 39842
rect 10334 39790 10386 39842
rect 10386 39790 10388 39842
rect 10332 39788 10388 39790
rect 9996 39452 10052 39508
rect 9660 39004 9716 39060
rect 9436 38668 9492 38724
rect 9436 37436 9492 37492
rect 9660 37772 9716 37828
rect 10332 39004 10388 39060
rect 11284 39452 11340 39508
rect 12572 40460 12628 40516
rect 12796 40796 12852 40852
rect 12908 40684 12964 40740
rect 13020 41580 13076 41636
rect 12908 40348 12964 40404
rect 12012 39452 12068 39508
rect 11676 39228 11732 39284
rect 10780 39004 10836 39060
rect 10444 38780 10500 38836
rect 10220 38444 10276 38500
rect 10220 37996 10276 38052
rect 10984 37772 11040 37828
rect 9716 36988 9772 37044
rect 11452 37772 11508 37828
rect 11564 38668 11620 38724
rect 9548 36652 9604 36708
rect 10500 36706 10556 36708
rect 10500 36654 10502 36706
rect 10502 36654 10554 36706
rect 10554 36654 10556 36706
rect 10500 36652 10556 36654
rect 7644 36092 7700 36148
rect 8316 36428 8372 36484
rect 8204 36204 8260 36260
rect 6412 35420 6468 35476
rect 7980 35308 8036 35364
rect 5572 34524 5628 34580
rect 5684 34412 5740 34468
rect 6188 34300 6244 34356
rect 6300 34188 6356 34244
rect 7308 34914 7364 34916
rect 7308 34862 7310 34914
rect 7310 34862 7362 34914
rect 7362 34862 7364 34914
rect 7308 34860 7364 34862
rect 6916 34524 6972 34580
rect 7532 34748 7588 34804
rect 7140 34300 7196 34356
rect 6748 34076 6804 34132
rect 6860 34188 6916 34244
rect 5572 33852 5628 33908
rect 6188 33346 6244 33348
rect 6188 33294 6190 33346
rect 6190 33294 6242 33346
rect 6242 33294 6244 33346
rect 6188 33292 6244 33294
rect 6076 33180 6132 33236
rect 5740 32284 5796 32340
rect 6524 33852 6580 33908
rect 6076 32562 6132 32564
rect 6076 32510 6078 32562
rect 6078 32510 6130 32562
rect 6130 32510 6132 32562
rect 6076 32508 6132 32510
rect 8204 35308 8260 35364
rect 8092 34076 8148 34132
rect 7532 33852 7588 33908
rect 7700 33852 7756 33908
rect 6636 32508 6692 32564
rect 6748 33628 6804 33684
rect 6076 31948 6132 32004
rect 5628 31836 5684 31892
rect 6076 31724 6132 31780
rect 4956 30044 5012 30100
rect 5908 30882 5964 30884
rect 5908 30830 5910 30882
rect 5910 30830 5962 30882
rect 5962 30830 5964 30882
rect 5908 30828 5964 30830
rect 3052 29596 3108 29652
rect 4956 29596 5012 29652
rect 1820 29260 1876 29316
rect 2772 29260 2828 29316
rect 3276 29484 3332 29540
rect 3724 29426 3780 29428
rect 3724 29374 3726 29426
rect 3726 29374 3778 29426
rect 3778 29374 3780 29426
rect 3724 29372 3780 29374
rect 4600 29260 4656 29316
rect 4476 29034 4532 29036
rect 4060 28924 4116 28980
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 1708 28588 1764 28644
rect 3724 28754 3780 28756
rect 3724 28702 3726 28754
rect 3726 28702 3778 28754
rect 3778 28702 3780 28754
rect 3724 28700 3780 28702
rect 2828 27244 2884 27300
rect 3052 27074 3108 27076
rect 3052 27022 3054 27074
rect 3054 27022 3106 27074
rect 3106 27022 3108 27074
rect 3052 27020 3108 27022
rect 1708 26124 1764 26180
rect 2548 26178 2604 26180
rect 2548 26126 2550 26178
rect 2550 26126 2602 26178
rect 2602 26126 2604 26178
rect 2548 26124 2604 26126
rect 1932 26066 1988 26068
rect 1932 26014 1934 26066
rect 1934 26014 1986 26066
rect 1986 26014 1988 26066
rect 1932 26012 1988 26014
rect 2660 25730 2716 25732
rect 2660 25678 2662 25730
rect 2662 25678 2714 25730
rect 2714 25678 2716 25730
rect 2660 25676 2716 25678
rect 1708 24892 1764 24948
rect 2156 25340 2212 25396
rect 3836 26908 3892 26964
rect 4172 28812 4228 28868
rect 4844 28812 4900 28868
rect 4508 28642 4564 28644
rect 4508 28590 4510 28642
rect 4510 28590 4562 28642
rect 4562 28590 4564 28642
rect 4508 28588 4564 28590
rect 5068 29372 5124 29428
rect 4900 27916 4956 27972
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 5516 29596 5572 29652
rect 5740 29708 5796 29764
rect 5348 29484 5404 29540
rect 5628 29484 5684 29540
rect 5516 29260 5572 29316
rect 5516 28924 5572 28980
rect 5180 28364 5236 28420
rect 5852 29484 5908 29540
rect 5628 28588 5684 28644
rect 5740 28812 5796 28868
rect 7700 33628 7756 33684
rect 7084 33068 7140 33124
rect 8428 35196 8484 35252
rect 8428 34748 8484 34804
rect 8428 33740 8484 33796
rect 8988 36092 9044 36148
rect 8876 35810 8932 35812
rect 8876 35758 8878 35810
rect 8878 35758 8930 35810
rect 8930 35758 8932 35810
rect 8876 35756 8932 35758
rect 8652 34914 8708 34916
rect 8652 34862 8654 34914
rect 8654 34862 8706 34914
rect 8706 34862 8708 34914
rect 8652 34860 8708 34862
rect 9548 36482 9604 36484
rect 9548 36430 9550 36482
rect 9550 36430 9602 36482
rect 9602 36430 9604 36482
rect 9548 36428 9604 36430
rect 9304 36316 9360 36372
rect 9212 34914 9268 34916
rect 9212 34862 9214 34914
rect 9214 34862 9266 34914
rect 9266 34862 9268 34914
rect 9212 34860 9268 34862
rect 8988 34300 9044 34356
rect 9100 34748 9156 34804
rect 11284 37154 11340 37156
rect 11284 37102 11286 37154
rect 11286 37102 11338 37154
rect 11338 37102 11340 37154
rect 11284 37100 11340 37102
rect 11452 36764 11508 36820
rect 9492 35756 9548 35812
rect 9455 34914 9511 34916
rect 9455 34862 9457 34914
rect 9457 34862 9509 34914
rect 9509 34862 9511 34914
rect 9455 34860 9511 34862
rect 9884 35308 9940 35364
rect 11452 36092 11508 36148
rect 11676 38050 11732 38052
rect 11676 37998 11678 38050
rect 11678 37998 11730 38050
rect 11730 37998 11732 38050
rect 11676 37996 11732 37998
rect 12292 39618 12348 39620
rect 12292 39566 12294 39618
rect 12294 39566 12346 39618
rect 12346 39566 12348 39618
rect 12292 39564 12348 39566
rect 12460 39506 12516 39508
rect 12460 39454 12462 39506
rect 12462 39454 12514 39506
rect 12514 39454 12516 39506
rect 12460 39452 12516 39454
rect 12124 39004 12180 39060
rect 12728 39004 12784 39060
rect 12124 37996 12180 38052
rect 12572 38050 12628 38052
rect 12572 37998 12574 38050
rect 12574 37998 12626 38050
rect 12626 37998 12628 38050
rect 12572 37996 12628 37998
rect 12012 37884 12068 37940
rect 11676 37772 11732 37828
rect 12460 37324 12516 37380
rect 12348 37100 12404 37156
rect 12012 36764 12068 36820
rect 12572 37266 12628 37268
rect 12572 37214 12574 37266
rect 12574 37214 12626 37266
rect 12626 37214 12628 37266
rect 12572 37212 12628 37214
rect 11788 36204 11844 36260
rect 11116 35756 11172 35812
rect 9660 34860 9716 34916
rect 6412 31052 6468 31108
rect 6188 30994 6244 30996
rect 6188 30942 6190 30994
rect 6190 30942 6242 30994
rect 6242 30942 6244 30994
rect 6188 30940 6244 30942
rect 6748 30994 6804 30996
rect 6748 30942 6750 30994
rect 6750 30942 6802 30994
rect 6802 30942 6804 30994
rect 6748 30940 6804 30942
rect 6972 30994 7028 30996
rect 6972 30942 6974 30994
rect 6974 30942 7026 30994
rect 7026 30942 7028 30994
rect 6972 30940 7028 30942
rect 7756 31948 7812 32004
rect 7980 31763 8036 31780
rect 7980 31724 7982 31763
rect 7982 31724 8034 31763
rect 8034 31724 8036 31763
rect 8316 33180 8372 33236
rect 8876 33234 8932 33236
rect 8876 33182 8878 33234
rect 8878 33182 8930 33234
rect 8930 33182 8932 33234
rect 8876 33180 8932 33182
rect 8316 31948 8372 32004
rect 8540 31778 8596 31780
rect 8540 31726 8542 31778
rect 8542 31726 8594 31778
rect 8594 31726 8596 31778
rect 8540 31724 8596 31726
rect 9100 33404 9156 33460
rect 9324 33516 9380 33572
rect 9212 32732 9268 32788
rect 9660 34354 9716 34356
rect 9660 34302 9662 34354
rect 9662 34302 9714 34354
rect 9714 34302 9716 34354
rect 9660 34300 9716 34302
rect 9548 31778 9604 31780
rect 9548 31726 9550 31778
rect 9550 31726 9602 31778
rect 9602 31726 9604 31778
rect 9548 31724 9604 31726
rect 7812 31106 7868 31108
rect 7812 31054 7814 31106
rect 7814 31054 7866 31106
rect 7866 31054 7868 31106
rect 7812 31052 7868 31054
rect 8204 30994 8260 30996
rect 8204 30942 8206 30994
rect 8206 30942 8258 30994
rect 8258 30942 8260 30994
rect 8204 30940 8260 30942
rect 7084 30492 7140 30548
rect 6300 30322 6356 30324
rect 6300 30270 6302 30322
rect 6302 30270 6354 30322
rect 6354 30270 6356 30322
rect 6300 30268 6356 30270
rect 7420 29932 7476 29988
rect 7756 30604 7812 30660
rect 6076 29148 6132 29204
rect 6076 28364 6132 28420
rect 4508 27074 4564 27076
rect 4508 27022 4510 27074
rect 4510 27022 4562 27074
rect 4562 27022 4564 27074
rect 4508 27020 4564 27022
rect 5292 27468 5348 27524
rect 4844 27020 4900 27076
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 5180 26290 5236 26292
rect 5180 26238 5182 26290
rect 5182 26238 5234 26290
rect 5234 26238 5236 26290
rect 5180 26236 5236 26238
rect 3164 25340 3220 25396
rect 2492 24722 2548 24724
rect 2492 24670 2494 24722
rect 2494 24670 2546 24722
rect 2546 24670 2548 24722
rect 2492 24668 2548 24670
rect 2044 23436 2100 23492
rect 1484 21420 1540 21476
rect 2828 24498 2884 24500
rect 2828 24446 2830 24498
rect 2830 24446 2882 24498
rect 2882 24446 2884 24498
rect 2828 24444 2884 24446
rect 3388 25116 3444 25172
rect 2600 23548 2656 23604
rect 3052 23436 3108 23492
rect 3164 24780 3220 24836
rect 3556 24722 3612 24724
rect 3556 24670 3558 24722
rect 3558 24670 3610 24722
rect 3610 24670 3612 24722
rect 3556 24668 3612 24670
rect 3164 23324 3220 23380
rect 4844 25116 4900 25172
rect 3948 24444 4004 24500
rect 4302 24610 4358 24612
rect 4302 24558 4304 24610
rect 4304 24558 4356 24610
rect 4356 24558 4358 24610
rect 4302 24556 4358 24558
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4396 24050 4452 24052
rect 4396 23998 4398 24050
rect 4398 23998 4450 24050
rect 4450 23998 4452 24050
rect 4396 23996 4452 23998
rect 4172 23938 4228 23940
rect 4172 23886 4174 23938
rect 4174 23886 4226 23938
rect 4226 23886 4228 23938
rect 4172 23884 4228 23886
rect 2156 21756 2212 21812
rect 3164 22764 3220 22820
rect 2828 22428 2884 22484
rect 3332 22764 3388 22820
rect 3500 22428 3556 22484
rect 3276 21756 3332 21812
rect 2604 21586 2660 21588
rect 2604 21534 2606 21586
rect 2606 21534 2658 21586
rect 2658 21534 2660 21586
rect 2604 21532 2660 21534
rect 3836 23772 3892 23828
rect 3892 23100 3948 23156
rect 3724 22204 3780 22260
rect 3500 21756 3556 21812
rect 3612 21698 3668 21700
rect 3612 21646 3614 21698
rect 3614 21646 3666 21698
rect 3666 21646 3668 21698
rect 3612 21644 3668 21646
rect 4056 21756 4112 21812
rect 4564 23772 4620 23828
rect 4284 23548 4340 23604
rect 4844 23100 4900 23156
rect 4788 22930 4844 22932
rect 4788 22878 4790 22930
rect 4790 22878 4842 22930
rect 4842 22878 4844 22930
rect 4788 22876 4844 22878
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4620 22428 4676 22484
rect 4508 22204 4564 22260
rect 4172 21644 4228 21700
rect 4508 21980 4564 22036
rect 5964 27858 6020 27860
rect 5964 27806 5966 27858
rect 5966 27806 6018 27858
rect 6018 27806 6020 27858
rect 5964 27804 6020 27806
rect 5740 27468 5796 27524
rect 5628 27074 5684 27076
rect 5628 27022 5630 27074
rect 5630 27022 5682 27074
rect 5682 27022 5684 27074
rect 5628 27020 5684 27022
rect 6636 29426 6692 29428
rect 6636 29374 6638 29426
rect 6638 29374 6690 29426
rect 6690 29374 6692 29426
rect 6636 29372 6692 29374
rect 6300 28754 6356 28756
rect 6300 28702 6302 28754
rect 6302 28702 6354 28754
rect 6354 28702 6356 28754
rect 6300 28700 6356 28702
rect 6188 27916 6244 27972
rect 6412 28364 6468 28420
rect 6244 27244 6300 27300
rect 5852 26796 5908 26852
rect 5516 24780 5572 24836
rect 5516 24332 5572 24388
rect 5628 23996 5684 24052
rect 5292 23772 5348 23828
rect 5180 23324 5236 23380
rect 4732 22370 4788 22372
rect 4732 22318 4734 22370
rect 4734 22318 4786 22370
rect 4786 22318 4788 22370
rect 4732 22316 4788 22318
rect 5964 25676 6020 25732
rect 6076 25452 6132 25508
rect 6300 25340 6356 25396
rect 6188 24668 6244 24724
rect 5740 23436 5796 23492
rect 5628 23212 5684 23268
rect 5404 22316 5460 22372
rect 5516 22876 5572 22932
rect 4732 21980 4788 22036
rect 4620 21868 4676 21924
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 1596 19964 1652 20020
rect 2156 19740 2212 19796
rect 2268 20018 2324 20020
rect 2268 19966 2270 20018
rect 2270 19966 2322 20018
rect 2322 19966 2324 20018
rect 2268 19964 2324 19966
rect 3052 19906 3108 19908
rect 3052 19854 3054 19906
rect 3054 19854 3106 19906
rect 3106 19854 3108 19906
rect 3052 19852 3108 19854
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 5404 21868 5460 21924
rect 5852 23212 5908 23268
rect 5964 23100 6020 23156
rect 6076 23324 6132 23380
rect 7476 29650 7532 29652
rect 7476 29598 7478 29650
rect 7478 29598 7530 29650
rect 7530 29598 7532 29650
rect 7476 29596 7532 29598
rect 8540 30940 8596 30996
rect 8428 30828 8484 30884
rect 8316 30604 8372 30660
rect 9996 34130 10052 34132
rect 9996 34078 9998 34130
rect 9998 34078 10050 34130
rect 10050 34078 10052 34130
rect 9996 34076 10052 34078
rect 9996 33458 10052 33460
rect 9996 33406 9998 33458
rect 9998 33406 10050 33458
rect 10050 33406 10052 33458
rect 9996 33404 10052 33406
rect 11116 35196 11172 35252
rect 10668 33740 10724 33796
rect 11284 34802 11340 34804
rect 11284 34750 11286 34802
rect 11286 34750 11338 34802
rect 11338 34750 11340 34802
rect 11284 34748 11340 34750
rect 11060 34412 11116 34468
rect 11060 33852 11116 33908
rect 11228 34524 11284 34580
rect 12124 35698 12180 35700
rect 12124 35646 12126 35698
rect 12126 35646 12178 35698
rect 12178 35646 12180 35698
rect 12124 35644 12180 35646
rect 13580 41468 13636 41524
rect 13132 40684 13188 40740
rect 13916 41020 13972 41076
rect 14140 40684 14196 40740
rect 13580 40402 13636 40404
rect 13580 40350 13582 40402
rect 13582 40350 13634 40402
rect 13634 40350 13636 40402
rect 13580 40348 13636 40350
rect 14588 43372 14644 43428
rect 14756 43036 14812 43092
rect 15036 43538 15092 43540
rect 15036 43486 15038 43538
rect 15038 43486 15090 43538
rect 15090 43486 15092 43538
rect 15036 43484 15092 43486
rect 14924 42812 14980 42868
rect 15036 43036 15092 43092
rect 15036 42754 15092 42756
rect 15036 42702 15038 42754
rect 15038 42702 15090 42754
rect 15090 42702 15092 42754
rect 15036 42700 15092 42702
rect 14700 42588 14756 42644
rect 16604 44882 16660 44884
rect 16604 44830 16606 44882
rect 16606 44830 16658 44882
rect 16658 44830 16660 44882
rect 16604 44828 16660 44830
rect 17668 44716 17724 44772
rect 15932 43596 15988 43652
rect 16380 43538 16436 43540
rect 16380 43486 16382 43538
rect 16382 43486 16434 43538
rect 16434 43486 16436 43538
rect 16380 43484 16436 43486
rect 16716 43484 16772 43540
rect 16156 42812 16212 42868
rect 15428 42588 15484 42644
rect 16380 42754 16436 42756
rect 16380 42702 16382 42754
rect 16382 42702 16434 42754
rect 16434 42702 16436 42754
rect 16380 42700 16436 42702
rect 15932 42588 15988 42644
rect 16268 42588 16324 42644
rect 14868 41970 14924 41972
rect 14868 41918 14870 41970
rect 14870 41918 14922 41970
rect 14922 41918 14924 41970
rect 14868 41916 14924 41918
rect 15260 41692 15316 41748
rect 15148 41580 15204 41636
rect 15372 41580 15428 41636
rect 15894 41955 15896 41972
rect 15896 41955 15948 41972
rect 15948 41955 15950 41972
rect 15894 41916 15950 41955
rect 16492 41916 16548 41972
rect 14456 40684 14512 40740
rect 14700 40684 14756 40740
rect 14252 39900 14308 39956
rect 13916 39676 13972 39732
rect 13524 39618 13580 39620
rect 13524 39566 13526 39618
rect 13526 39566 13578 39618
rect 13578 39566 13580 39618
rect 13524 39564 13580 39566
rect 13244 39452 13300 39508
rect 13580 38780 13636 38836
rect 13132 37324 13188 37380
rect 13356 38108 13412 38164
rect 13916 39228 13972 39284
rect 14364 39564 14420 39620
rect 15596 41132 15652 41188
rect 16044 41468 16100 41524
rect 15800 41020 15856 41076
rect 14924 39452 14980 39508
rect 15372 39340 15428 39396
rect 15820 40572 15876 40628
rect 16884 43538 16940 43540
rect 16884 43486 16886 43538
rect 16886 43486 16938 43538
rect 16938 43486 16940 43538
rect 16884 43484 16940 43486
rect 16716 42028 16772 42084
rect 16884 42028 16940 42084
rect 20076 45862 20132 45892
rect 20076 45836 20078 45862
rect 20078 45836 20130 45862
rect 20130 45836 20132 45862
rect 18508 45612 18564 45668
rect 18060 44994 18116 44996
rect 18060 44942 18062 44994
rect 18062 44942 18114 44994
rect 18114 44942 18116 44994
rect 18060 44940 18116 44942
rect 17836 43708 17892 43764
rect 17948 44604 18004 44660
rect 17668 43650 17724 43652
rect 17668 43598 17670 43650
rect 17670 43598 17722 43650
rect 17722 43598 17724 43650
rect 17668 43596 17724 43598
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 19964 44994 20020 44996
rect 19964 44942 19966 44994
rect 19966 44942 20018 44994
rect 20018 44942 20020 44994
rect 19964 44940 20020 44942
rect 20748 45106 20804 45108
rect 20748 45054 20750 45106
rect 20750 45054 20802 45106
rect 20802 45054 20804 45106
rect 20748 45052 20804 45054
rect 20860 44492 20916 44548
rect 19404 44044 19460 44100
rect 19292 43762 19348 43764
rect 19292 43710 19294 43762
rect 19294 43710 19346 43762
rect 19346 43710 19348 43762
rect 19292 43708 19348 43710
rect 17500 42812 17556 42868
rect 17164 42754 17220 42756
rect 17164 42702 17166 42754
rect 17166 42702 17218 42754
rect 17218 42702 17220 42754
rect 17164 42700 17220 42702
rect 17388 42754 17444 42756
rect 17388 42702 17390 42754
rect 17390 42702 17442 42754
rect 17442 42702 17444 42754
rect 17388 42700 17444 42702
rect 17164 42028 17220 42084
rect 16716 41186 16772 41188
rect 16716 41134 16718 41186
rect 16718 41134 16770 41186
rect 16770 41134 16772 41186
rect 16716 41132 16772 41134
rect 16492 40348 16548 40404
rect 16604 40460 16660 40516
rect 14252 38780 14308 38836
rect 13804 38668 13860 38724
rect 14364 38556 14420 38612
rect 13692 37884 13748 37940
rect 13188 37100 13244 37156
rect 13804 37242 13806 37268
rect 13806 37242 13858 37268
rect 13858 37242 13860 37268
rect 13804 37212 13860 37242
rect 13692 37100 13748 37156
rect 14364 38108 14420 38164
rect 15596 39116 15652 39172
rect 15932 38834 15988 38836
rect 14252 38050 14308 38052
rect 14252 37998 14254 38050
rect 14254 37998 14306 38050
rect 14306 37998 14308 38050
rect 14252 37996 14308 37998
rect 15932 38782 15934 38834
rect 15934 38782 15986 38834
rect 15986 38782 15988 38834
rect 15932 38780 15988 38782
rect 14588 37996 14644 38052
rect 15800 38556 15856 38612
rect 14924 38050 14980 38052
rect 14924 37998 14926 38050
rect 14926 37998 14978 38050
rect 14978 37998 14980 38050
rect 14924 37996 14980 37998
rect 16044 38050 16100 38052
rect 16044 37998 16046 38050
rect 16046 37998 16098 38050
rect 16098 37998 16100 38050
rect 16044 37996 16100 37998
rect 15204 37154 15260 37156
rect 15204 37102 15206 37154
rect 15206 37102 15258 37154
rect 15258 37102 15260 37154
rect 15204 37100 15260 37102
rect 12236 35420 12292 35476
rect 12572 35698 12628 35700
rect 12572 35646 12574 35698
rect 12574 35646 12626 35698
rect 12626 35646 12628 35698
rect 12572 35644 12628 35646
rect 11788 34972 11844 35028
rect 10780 33628 10836 33684
rect 9772 31612 9828 31668
rect 11228 33180 11284 33236
rect 10220 31724 10276 31780
rect 9996 31612 10052 31668
rect 9212 30380 9268 30436
rect 8764 30268 8820 30324
rect 9324 30268 9380 30324
rect 8204 30210 8260 30212
rect 8204 30158 8206 30210
rect 8206 30158 8258 30210
rect 8258 30158 8260 30210
rect 8204 30156 8260 30158
rect 8092 30044 8148 30100
rect 8820 30044 8876 30100
rect 9156 30044 9212 30100
rect 9324 30044 9380 30100
rect 8316 29372 8372 29428
rect 8988 29426 9044 29428
rect 8988 29374 8990 29426
rect 8990 29374 9042 29426
rect 9042 29374 9044 29426
rect 8988 29372 9044 29374
rect 6860 28364 6916 28420
rect 7140 28418 7196 28420
rect 7140 28366 7142 28418
rect 7142 28366 7194 28418
rect 7194 28366 7196 28418
rect 7140 28364 7196 28366
rect 6972 28028 7028 28084
rect 6804 27916 6860 27972
rect 6524 27468 6580 27524
rect 6636 27858 6692 27860
rect 6636 27806 6638 27858
rect 6638 27806 6690 27858
rect 6690 27806 6692 27858
rect 6636 27804 6692 27806
rect 7080 27036 7136 27076
rect 7080 27020 7082 27036
rect 7082 27020 7134 27036
rect 7134 27020 7136 27036
rect 7420 28642 7476 28644
rect 7420 28590 7422 28642
rect 7422 28590 7474 28642
rect 7474 28590 7476 28642
rect 7420 28588 7476 28590
rect 10108 31388 10164 31444
rect 10556 31500 10612 31556
rect 9884 30981 9886 30996
rect 9886 30981 9938 30996
rect 9938 30981 9940 30996
rect 9884 30940 9940 30981
rect 10108 30940 10164 30996
rect 9660 29372 9716 29428
rect 9324 29036 9380 29092
rect 8428 28924 8484 28980
rect 8296 28642 8352 28644
rect 8296 28590 8298 28642
rect 8298 28590 8350 28642
rect 8350 28590 8352 28642
rect 8296 28588 8352 28590
rect 7476 28082 7532 28084
rect 7476 28030 7478 28082
rect 7478 28030 7530 28082
rect 7530 28030 7532 28082
rect 7476 28028 7532 28030
rect 7756 27858 7812 27860
rect 7756 27806 7758 27858
rect 7758 27806 7810 27858
rect 7810 27806 7812 27858
rect 7756 27804 7812 27806
rect 8036 27858 8092 27860
rect 8036 27806 8038 27858
rect 8038 27806 8090 27858
rect 8090 27806 8092 27858
rect 8036 27804 8092 27806
rect 7868 27468 7924 27524
rect 7644 27132 7700 27188
rect 9660 28924 9716 28980
rect 9864 28812 9920 28868
rect 11004 32732 11060 32788
rect 10892 32562 10948 32564
rect 10892 32510 10894 32562
rect 10894 32510 10946 32562
rect 10946 32510 10948 32562
rect 10892 32508 10948 32510
rect 11340 32844 11396 32900
rect 11900 33516 11956 33572
rect 12012 34076 12068 34132
rect 11900 33234 11956 33236
rect 11900 33182 11902 33234
rect 11902 33182 11954 33234
rect 11954 33182 11956 33234
rect 11900 33180 11956 33182
rect 11676 32732 11732 32788
rect 11676 32172 11732 32228
rect 11452 31724 11508 31780
rect 10780 30492 10836 30548
rect 10668 29538 10724 29540
rect 10668 29486 10670 29538
rect 10670 29486 10722 29538
rect 10722 29486 10724 29538
rect 10668 29484 10724 29486
rect 10612 28642 10668 28644
rect 10612 28590 10614 28642
rect 10614 28590 10666 28642
rect 10666 28590 10668 28642
rect 10612 28588 10668 28590
rect 11004 30380 11060 30436
rect 12348 35084 12404 35140
rect 12796 35196 12852 35252
rect 12516 34860 12572 34916
rect 12684 34636 12740 34692
rect 12460 34300 12516 34356
rect 12684 34300 12740 34356
rect 12964 34242 13020 34244
rect 12964 34190 12966 34242
rect 12966 34190 13018 34242
rect 13018 34190 13020 34242
rect 12964 34188 13020 34190
rect 12460 33852 12516 33908
rect 12348 33740 12404 33796
rect 12348 33516 12404 33572
rect 12124 31836 12180 31892
rect 12236 31948 12292 32004
rect 12852 33570 12908 33572
rect 12852 33518 12854 33570
rect 12854 33518 12906 33570
rect 12906 33518 12908 33570
rect 12852 33516 12908 33518
rect 12572 33346 12628 33348
rect 12572 33294 12574 33346
rect 12574 33294 12626 33346
rect 12626 33294 12628 33346
rect 12572 33292 12628 33294
rect 12796 32786 12852 32788
rect 12796 32734 12798 32786
rect 12798 32734 12850 32786
rect 12850 32734 12852 32786
rect 12796 32732 12852 32734
rect 12572 32620 12628 32676
rect 12460 31948 12516 32004
rect 12460 31666 12516 31668
rect 12460 31614 12462 31666
rect 12462 31614 12514 31666
rect 12514 31614 12516 31666
rect 12460 31612 12516 31614
rect 12124 31500 12180 31556
rect 11004 30210 11060 30212
rect 11004 30158 11006 30210
rect 11006 30158 11058 30210
rect 11058 30158 11060 30210
rect 11004 30156 11060 30158
rect 13448 35308 13504 35364
rect 13804 36482 13860 36484
rect 13804 36430 13806 36482
rect 13806 36430 13858 36482
rect 13858 36430 13860 36482
rect 13804 36428 13860 36430
rect 13692 35586 13748 35588
rect 13692 35534 13694 35586
rect 13694 35534 13746 35586
rect 13746 35534 13748 35586
rect 13692 35532 13748 35534
rect 13580 35084 13636 35140
rect 15596 36876 15652 36932
rect 15484 35868 15540 35924
rect 13916 35196 13972 35252
rect 15596 35308 15652 35364
rect 15148 35138 15204 35140
rect 15148 35086 15150 35138
rect 15150 35086 15202 35138
rect 15202 35086 15204 35138
rect 15148 35084 15204 35086
rect 13244 31164 13300 31220
rect 14364 34188 14420 34244
rect 13916 34130 13972 34132
rect 13916 34078 13918 34130
rect 13918 34078 13970 34130
rect 13970 34078 13972 34130
rect 13916 34076 13972 34078
rect 13580 33740 13636 33796
rect 13692 33628 13748 33684
rect 13804 33309 13860 33348
rect 13804 33292 13806 33309
rect 13806 33292 13858 33309
rect 13858 33292 13860 33309
rect 14084 33516 14140 33572
rect 14812 34076 14868 34132
rect 14364 33292 14420 33348
rect 14588 33516 14644 33572
rect 14364 32620 14420 32676
rect 13916 32172 13972 32228
rect 14028 32508 14084 32564
rect 15148 34130 15204 34132
rect 15148 34078 15150 34130
rect 15150 34078 15202 34130
rect 15202 34078 15204 34130
rect 15148 34076 15204 34078
rect 14924 33852 14980 33908
rect 15036 33964 15092 34020
rect 15708 34690 15764 34692
rect 15708 34638 15710 34690
rect 15710 34638 15762 34690
rect 15762 34638 15764 34690
rect 15708 34636 15764 34638
rect 15032 33628 15088 33684
rect 13580 32002 13636 32004
rect 13580 31950 13582 32002
rect 13582 31950 13634 32002
rect 13634 31950 13636 32002
rect 13580 31948 13636 31950
rect 13468 31724 13524 31780
rect 13974 31500 14030 31556
rect 11452 29036 11508 29092
rect 11340 28812 11396 28868
rect 8932 27916 8988 27972
rect 9100 27692 9156 27748
rect 9324 27804 9380 27860
rect 6524 26124 6580 26180
rect 6636 25676 6692 25732
rect 6972 25564 7028 25620
rect 7084 25506 7140 25508
rect 7084 25454 7086 25506
rect 7086 25454 7138 25506
rect 7138 25454 7140 25506
rect 7084 25452 7140 25454
rect 6972 24668 7028 24724
rect 6636 23884 6692 23940
rect 6524 23212 6580 23268
rect 6860 24332 6916 24388
rect 6972 23884 7028 23940
rect 6860 22988 6916 23044
rect 7532 26460 7588 26516
rect 7532 25676 7588 25732
rect 7868 26796 7924 26852
rect 7644 24556 7700 24612
rect 7756 25340 7812 25396
rect 7756 24668 7812 24724
rect 8540 27074 8596 27076
rect 8540 27022 8542 27074
rect 8542 27022 8594 27074
rect 8594 27022 8596 27074
rect 8540 27020 8596 27022
rect 8092 26460 8148 26516
rect 8764 26908 8820 26964
rect 8092 26290 8148 26292
rect 8092 26238 8094 26290
rect 8094 26238 8146 26290
rect 8146 26238 8148 26290
rect 8092 26236 8148 26238
rect 8652 26460 8708 26516
rect 8540 25676 8596 25732
rect 8428 25564 8484 25620
rect 7980 25116 8036 25172
rect 8428 25394 8484 25396
rect 8428 25342 8430 25394
rect 8430 25342 8482 25394
rect 8482 25342 8484 25394
rect 8428 25340 8484 25342
rect 8540 25116 8596 25172
rect 9772 27356 9828 27412
rect 9548 27074 9604 27076
rect 9548 27022 9550 27074
rect 9550 27022 9602 27074
rect 9602 27022 9604 27074
rect 9548 27020 9604 27022
rect 8876 26460 8932 26516
rect 9436 26290 9492 26292
rect 9436 26238 9438 26290
rect 9438 26238 9490 26290
rect 9490 26238 9492 26290
rect 9436 26236 9492 26238
rect 8092 24780 8148 24836
rect 8316 24722 8372 24724
rect 8316 24670 8318 24722
rect 8318 24670 8370 24722
rect 8370 24670 8372 24722
rect 8316 24668 8372 24670
rect 7756 23938 7812 23940
rect 7196 23324 7252 23380
rect 7756 23886 7758 23938
rect 7758 23886 7810 23938
rect 7810 23886 7812 23938
rect 7756 23884 7812 23886
rect 8540 24834 8596 24836
rect 8540 24782 8542 24834
rect 8542 24782 8594 24834
rect 8594 24782 8596 24834
rect 8540 24780 8596 24782
rect 8708 24722 8764 24724
rect 8708 24670 8710 24722
rect 8710 24670 8762 24722
rect 8762 24670 8764 24722
rect 8708 24668 8764 24670
rect 10220 28028 10276 28084
rect 9996 27132 10052 27188
rect 10444 27834 10446 27860
rect 10446 27834 10498 27860
rect 10498 27834 10500 27860
rect 10444 27804 10500 27834
rect 10556 27580 10612 27636
rect 10220 27356 10276 27412
rect 11004 28364 11060 28420
rect 10780 27804 10836 27860
rect 10892 27916 10948 27972
rect 10332 27132 10388 27188
rect 10220 26908 10276 26964
rect 9884 25564 9940 25620
rect 10108 25564 10164 25620
rect 8988 24668 9044 24724
rect 9100 25452 9156 25508
rect 8034 23938 8090 23940
rect 8034 23886 8036 23938
rect 8036 23886 8088 23938
rect 8088 23886 8090 23938
rect 8034 23884 8090 23886
rect 7308 23212 7364 23268
rect 5740 21868 5796 21924
rect 5852 21532 5908 21588
rect 5180 20802 5236 20804
rect 5180 20750 5182 20802
rect 5182 20750 5234 20802
rect 5234 20750 5236 20802
rect 5180 20748 5236 20750
rect 6300 22370 6356 22372
rect 6300 22318 6302 22370
rect 6302 22318 6354 22370
rect 6354 22318 6356 22370
rect 6300 22316 6356 22318
rect 6580 22370 6636 22372
rect 6580 22318 6582 22370
rect 6582 22318 6634 22370
rect 6634 22318 6636 22370
rect 6580 22316 6636 22318
rect 6412 22204 6468 22260
rect 6524 21868 6580 21924
rect 5516 20748 5572 20804
rect 4956 19234 5012 19236
rect 4956 19182 4958 19234
rect 4958 19182 5010 19234
rect 5010 19182 5012 19234
rect 4956 19180 5012 19182
rect 4284 18956 4340 19012
rect 5404 18956 5460 19012
rect 4004 18732 4060 18788
rect 2268 18396 2324 18452
rect 3052 18450 3108 18452
rect 3052 18398 3054 18450
rect 3054 18398 3106 18450
rect 3106 18398 3108 18450
rect 3052 18396 3108 18398
rect 5292 18396 5348 18452
rect 3836 18338 3892 18340
rect 3836 18286 3838 18338
rect 3838 18286 3890 18338
rect 3890 18286 3892 18338
rect 3836 18284 3892 18286
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 5124 17778 5180 17780
rect 5124 17726 5126 17778
rect 5126 17726 5178 17778
rect 5178 17726 5180 17778
rect 5124 17724 5180 17726
rect 5292 17612 5348 17668
rect 5516 18396 5572 18452
rect 4228 17554 4284 17556
rect 4228 17502 4230 17554
rect 4230 17502 4282 17554
rect 4282 17502 4284 17554
rect 4228 17500 4284 17502
rect 4676 17554 4732 17556
rect 4676 17502 4678 17554
rect 4678 17502 4730 17554
rect 4730 17502 4732 17554
rect 4676 17500 4732 17502
rect 4340 17106 4396 17108
rect 4340 17054 4342 17106
rect 4342 17054 4394 17106
rect 4394 17054 4396 17106
rect 4340 17052 4396 17054
rect 4732 16770 4788 16772
rect 4732 16718 4734 16770
rect 4734 16718 4786 16770
rect 4786 16718 4788 16770
rect 4732 16716 4788 16718
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 5740 18450 5796 18452
rect 5740 18398 5742 18450
rect 5742 18398 5794 18450
rect 5794 18398 5796 18450
rect 5740 18396 5796 18398
rect 5740 17500 5796 17556
rect 5628 17052 5684 17108
rect 6246 20412 6302 20468
rect 7196 22876 7252 22932
rect 6636 20524 6692 20580
rect 6636 20076 6692 20132
rect 6524 20003 6544 20020
rect 6544 20003 6580 20020
rect 6524 19964 6580 20003
rect 7196 22316 7252 22372
rect 7532 23324 7588 23380
rect 8876 23772 8932 23828
rect 7756 23154 7812 23156
rect 7756 23102 7758 23154
rect 7758 23102 7810 23154
rect 7810 23102 7812 23154
rect 8092 23154 8148 23156
rect 7756 23100 7812 23102
rect 8092 23102 8094 23154
rect 8094 23102 8146 23154
rect 8146 23102 8148 23154
rect 8092 23100 8148 23102
rect 8204 22876 8260 22932
rect 7924 22540 7980 22596
rect 9212 25116 9268 25172
rect 9324 25340 9380 25396
rect 9436 24556 9492 24612
rect 11340 28028 11396 28084
rect 11228 27916 11284 27972
rect 11116 27186 11172 27188
rect 11116 27134 11118 27186
rect 11118 27134 11170 27186
rect 11170 27134 11172 27186
rect 11116 27132 11172 27134
rect 11564 27132 11620 27188
rect 11340 26908 11396 26964
rect 11004 26684 11060 26740
rect 11676 26908 11732 26964
rect 10220 25116 10276 25172
rect 10332 25452 10388 25508
rect 9212 23938 9268 23940
rect 9212 23886 9214 23938
rect 9214 23886 9266 23938
rect 9266 23886 9268 23938
rect 9212 23884 9268 23886
rect 9212 22540 9268 22596
rect 9436 22370 9492 22372
rect 9436 22318 9438 22370
rect 9438 22318 9490 22370
rect 9490 22318 9492 22370
rect 9436 22316 9492 22318
rect 8764 21586 8820 21588
rect 8764 21534 8766 21586
rect 8766 21534 8818 21586
rect 8818 21534 8820 21586
rect 8764 21532 8820 21534
rect 9772 23100 9828 23156
rect 9660 22540 9716 22596
rect 10220 23154 10276 23156
rect 10220 23102 10222 23154
rect 10222 23102 10274 23154
rect 10274 23102 10276 23154
rect 10220 23100 10276 23102
rect 10108 22540 10164 22596
rect 9884 22316 9940 22372
rect 7644 20748 7700 20804
rect 6972 20076 7028 20132
rect 6076 19794 6132 19796
rect 6076 19742 6078 19794
rect 6078 19742 6130 19794
rect 6130 19742 6132 19794
rect 6076 19740 6132 19742
rect 6636 19740 6692 19796
rect 7532 20018 7588 20020
rect 7532 19966 7534 20018
rect 7534 19966 7586 20018
rect 7586 19966 7588 20018
rect 7532 19964 7588 19966
rect 7196 19906 7252 19908
rect 7196 19854 7198 19906
rect 7198 19854 7250 19906
rect 7250 19854 7252 19906
rect 7196 19852 7252 19854
rect 6972 19740 7028 19796
rect 6972 19458 7028 19460
rect 6972 19406 6974 19458
rect 6974 19406 7026 19458
rect 7026 19406 7028 19458
rect 6972 19404 7028 19406
rect 6636 19234 6692 19236
rect 6636 19182 6638 19234
rect 6638 19182 6690 19234
rect 6690 19182 6692 19234
rect 6636 19180 6692 19182
rect 9324 20860 9380 20916
rect 7868 19852 7924 19908
rect 8428 19964 8484 20020
rect 9044 19740 9100 19796
rect 9212 19740 9268 19796
rect 8036 19628 8092 19684
rect 7756 19404 7812 19460
rect 8988 19458 9044 19460
rect 8988 19406 8990 19458
rect 8990 19406 9042 19458
rect 9042 19406 9044 19458
rect 8988 19404 9044 19406
rect 6412 18732 6468 18788
rect 6524 18956 6580 19012
rect 7532 19010 7588 19012
rect 7532 18958 7534 19010
rect 7534 18958 7586 19010
rect 7586 18958 7588 19010
rect 7532 18956 7588 18958
rect 6300 18338 6356 18340
rect 6300 18286 6302 18338
rect 6302 18286 6354 18338
rect 6354 18286 6356 18338
rect 6300 18284 6356 18286
rect 6412 17666 6468 17668
rect 6412 17614 6414 17666
rect 6414 17614 6466 17666
rect 6466 17614 6468 17666
rect 6412 17612 6468 17614
rect 7924 18450 7980 18452
rect 7924 18398 7926 18450
rect 7926 18398 7978 18450
rect 7978 18398 7980 18450
rect 7924 18396 7980 18398
rect 7476 18172 7532 18228
rect 8316 17836 8372 17892
rect 6860 17500 6916 17556
rect 5964 16770 6020 16772
rect 5964 16718 5966 16770
rect 5966 16718 6018 16770
rect 6018 16718 6020 16770
rect 5964 16716 6020 16718
rect 8540 18284 8596 18340
rect 8540 17724 8596 17780
rect 8652 17836 8708 17892
rect 8316 17052 8372 17108
rect 4284 15932 4340 15988
rect 3052 15484 3108 15540
rect 3500 15538 3556 15540
rect 3500 15486 3502 15538
rect 3502 15486 3554 15538
rect 3554 15486 3556 15538
rect 3500 15484 3556 15486
rect 3836 15314 3892 15316
rect 3836 15262 3838 15314
rect 3838 15262 3890 15314
rect 3890 15262 3892 15314
rect 3836 15260 3892 15262
rect 4956 15986 5012 15988
rect 4956 15934 4958 15986
rect 4958 15934 5010 15986
rect 5010 15934 5012 15986
rect 4956 15932 5012 15934
rect 4508 15820 4564 15876
rect 4956 15372 5012 15428
rect 5404 15372 5460 15428
rect 5068 15260 5124 15316
rect 4620 15202 4676 15204
rect 4620 15150 4622 15202
rect 4622 15150 4674 15202
rect 4674 15150 4676 15202
rect 4620 15148 4676 15150
rect 5292 15148 5348 15204
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 2044 13916 2100 13972
rect 4732 14530 4788 14532
rect 4732 14478 4734 14530
rect 4734 14478 4786 14530
rect 4786 14478 4788 14530
rect 4732 14476 4788 14478
rect 5068 14252 5124 14308
rect 3388 13916 3444 13972
rect 4900 13970 4956 13972
rect 4900 13918 4902 13970
rect 4902 13918 4954 13970
rect 4954 13918 4956 13970
rect 4900 13916 4956 13918
rect 3500 13746 3556 13748
rect 3500 13694 3502 13746
rect 3502 13694 3554 13746
rect 3554 13694 3556 13746
rect 3500 13692 3556 13694
rect 6188 15932 6244 15988
rect 5964 15372 6020 15428
rect 6412 16156 6468 16212
rect 5852 14924 5908 14980
rect 6076 14530 6132 14532
rect 6076 14478 6078 14530
rect 6078 14478 6130 14530
rect 6130 14478 6132 14530
rect 6076 14476 6132 14478
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 3388 11676 3444 11732
rect 5964 13692 6020 13748
rect 6300 13356 6356 13412
rect 6300 13020 6356 13076
rect 3948 11676 4004 11732
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 1820 11452 1876 11508
rect 3276 10780 3332 10836
rect 2604 9996 2660 10052
rect 1596 8652 1652 8708
rect 3556 8876 3612 8932
rect 3556 8652 3612 8708
rect 3052 8428 3108 8484
rect 28 8092 84 8148
rect 3836 8258 3892 8260
rect 3836 8206 3838 8258
rect 3838 8206 3890 8258
rect 3890 8206 3892 8258
rect 3836 8204 3892 8206
rect 5124 11564 5180 11620
rect 4508 11394 4564 11396
rect 4508 11342 4510 11394
rect 4510 11342 4562 11394
rect 4562 11342 4564 11394
rect 4508 11340 4564 11342
rect 4396 11228 4452 11284
rect 5292 11116 5348 11172
rect 5068 10780 5124 10836
rect 4508 10498 4564 10500
rect 4508 10446 4510 10498
rect 4510 10446 4562 10498
rect 4562 10446 4564 10498
rect 4508 10444 4564 10446
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4284 9826 4340 9828
rect 4284 9774 4286 9826
rect 4286 9774 4338 9826
rect 4338 9774 4340 9826
rect 4284 9772 4340 9774
rect 4396 9660 4452 9716
rect 5180 10444 5236 10500
rect 5516 11452 5572 11508
rect 7196 16210 7252 16212
rect 7196 16158 7198 16210
rect 7198 16158 7250 16210
rect 7250 16158 7252 16210
rect 7196 16156 7252 16158
rect 10108 20076 10164 20132
rect 9996 19852 10052 19908
rect 9996 18956 10052 19012
rect 9212 17836 9268 17892
rect 8764 17052 8820 17108
rect 6972 15820 7028 15876
rect 7308 15820 7364 15876
rect 7140 15596 7196 15652
rect 8204 15596 8260 15652
rect 6524 14924 6580 14980
rect 6524 14530 6580 14532
rect 6524 14478 6526 14530
rect 6526 14478 6578 14530
rect 6578 14478 6580 14530
rect 6524 14476 6580 14478
rect 6412 12460 6468 12516
rect 6972 14140 7028 14196
rect 7420 15314 7476 15316
rect 7420 15262 7422 15314
rect 7422 15262 7474 15314
rect 7474 15262 7476 15314
rect 7420 15260 7476 15262
rect 7756 15314 7812 15316
rect 7756 15262 7758 15314
rect 7758 15262 7810 15314
rect 7810 15262 7812 15314
rect 7756 15260 7812 15262
rect 8316 15484 8372 15540
rect 8316 15314 8372 15316
rect 8316 15262 8318 15314
rect 8318 15262 8370 15314
rect 8370 15262 8372 15314
rect 8316 15260 8372 15262
rect 8092 15148 8148 15204
rect 6748 13468 6804 13524
rect 6636 12290 6692 12292
rect 6636 12238 6638 12290
rect 6638 12238 6690 12290
rect 6690 12238 6692 12290
rect 6636 12236 6692 12238
rect 6188 11564 6244 11620
rect 5628 11394 5684 11396
rect 5628 11342 5630 11394
rect 5630 11342 5682 11394
rect 5682 11342 5684 11394
rect 5628 11340 5684 11342
rect 5964 11228 6020 11284
rect 6412 11394 6468 11396
rect 6412 11342 6414 11394
rect 6414 11342 6466 11394
rect 6466 11342 6468 11394
rect 6412 11340 6468 11342
rect 6860 13356 6916 13412
rect 6972 12796 7028 12852
rect 6860 11506 6916 11508
rect 6860 11454 6862 11506
rect 6862 11454 6914 11506
rect 6914 11454 6916 11506
rect 6860 11452 6916 11454
rect 6860 11228 6916 11284
rect 5740 9996 5796 10052
rect 6972 10498 7028 10500
rect 6972 10446 6974 10498
rect 6974 10446 7026 10498
rect 7026 10446 7028 10498
rect 6972 10444 7028 10446
rect 4844 9602 4900 9604
rect 4844 9550 4846 9602
rect 4846 9550 4898 9602
rect 4898 9550 4900 9602
rect 4844 9548 4900 9550
rect 5628 9548 5684 9604
rect 6300 9884 6356 9940
rect 6860 9826 6916 9828
rect 6860 9774 6862 9826
rect 6862 9774 6914 9826
rect 6914 9774 6916 9826
rect 6860 9772 6916 9774
rect 5964 9660 6020 9716
rect 6748 9660 6804 9716
rect 5292 9042 5348 9044
rect 5292 8990 5294 9042
rect 5294 8990 5346 9042
rect 5346 8990 5348 9042
rect 5292 8988 5348 8990
rect 5628 8988 5684 9044
rect 4900 8930 4956 8932
rect 4900 8878 4902 8930
rect 4902 8878 4954 8930
rect 4954 8878 4956 8930
rect 4900 8876 4956 8878
rect 4172 8316 4228 8372
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4956 8652 5012 8708
rect 4620 8258 4676 8260
rect 4620 8206 4622 8258
rect 4622 8206 4674 8258
rect 4674 8206 4676 8258
rect 4620 8204 4676 8206
rect 5852 8876 5908 8932
rect 5740 8428 5796 8484
rect 5180 7644 5236 7700
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4508 6860 4564 6916
rect 3948 6636 4004 6692
rect 4956 6636 5012 6692
rect 4844 6466 4900 6468
rect 4844 6414 4846 6466
rect 4846 6414 4898 6466
rect 4898 6414 4900 6466
rect 4844 6412 4900 6414
rect 5740 6860 5796 6916
rect 6860 8930 6916 8932
rect 6860 8878 6862 8930
rect 6862 8878 6914 8930
rect 6914 8878 6916 8930
rect 6860 8876 6916 8878
rect 6076 8316 6132 8372
rect 6860 8370 6916 8372
rect 6860 8318 6862 8370
rect 6862 8318 6914 8370
rect 6914 8318 6916 8370
rect 6860 8316 6916 8318
rect 5796 6690 5852 6692
rect 5796 6638 5798 6690
rect 5798 6638 5850 6690
rect 5850 6638 5852 6690
rect 5796 6636 5852 6638
rect 6748 8204 6804 8260
rect 8540 14812 8596 14868
rect 8316 14364 8372 14420
rect 8428 14306 8484 14308
rect 8428 14254 8430 14306
rect 8430 14254 8482 14306
rect 8482 14254 8484 14306
rect 8428 14252 8484 14254
rect 8876 15260 8932 15316
rect 9996 18060 10052 18116
rect 9436 17052 9492 17108
rect 9324 16828 9380 16884
rect 9996 16940 10052 16996
rect 10220 17948 10276 18004
rect 10108 17666 10164 17668
rect 10108 17614 10110 17666
rect 10110 17614 10162 17666
rect 10162 17614 10164 17666
rect 10108 17612 10164 17614
rect 10108 16828 10164 16884
rect 9492 15314 9548 15316
rect 9492 15262 9494 15314
rect 9494 15262 9546 15314
rect 9546 15262 9548 15314
rect 9492 15260 9548 15262
rect 9660 15148 9716 15204
rect 8764 14812 8820 14868
rect 7420 13522 7476 13524
rect 7420 13470 7422 13522
rect 7422 13470 7474 13522
rect 7474 13470 7476 13522
rect 7420 13468 7476 13470
rect 7980 13468 8036 13524
rect 8092 13356 8148 13412
rect 8092 13074 8148 13076
rect 8092 13022 8094 13074
rect 8094 13022 8146 13074
rect 8146 13022 8148 13074
rect 8092 13020 8148 13022
rect 7196 12236 7252 12292
rect 8540 13746 8596 13748
rect 8540 13694 8542 13746
rect 8542 13694 8594 13746
rect 8594 13694 8596 13746
rect 8540 13692 8596 13694
rect 8876 13634 8932 13636
rect 8876 13582 8878 13634
rect 8878 13582 8930 13634
rect 8930 13582 8932 13634
rect 8876 13580 8932 13582
rect 9100 13468 9156 13524
rect 8428 12684 8484 12740
rect 8652 13356 8708 13412
rect 8652 12796 8708 12852
rect 7252 11788 7308 11844
rect 7868 11394 7924 11396
rect 7868 11342 7870 11394
rect 7870 11342 7922 11394
rect 7922 11342 7924 11394
rect 7868 11340 7924 11342
rect 8316 11340 8372 11396
rect 7756 11228 7812 11284
rect 7532 11116 7588 11172
rect 8204 10444 8260 10500
rect 7308 9938 7364 9940
rect 7308 9886 7310 9938
rect 7310 9886 7362 9938
rect 7362 9886 7364 9938
rect 7308 9884 7364 9886
rect 7084 8652 7140 8708
rect 7308 8930 7364 8932
rect 7308 8878 7310 8930
rect 7310 8878 7362 8930
rect 7362 8878 7364 8930
rect 7308 8876 7364 8878
rect 7420 8652 7476 8708
rect 7308 8316 7364 8372
rect 6972 7420 7028 7476
rect 8764 12738 8820 12740
rect 8764 12686 8766 12738
rect 8766 12686 8818 12738
rect 8818 12686 8820 12738
rect 8764 12684 8820 12686
rect 8988 12178 9044 12180
rect 8988 12126 8990 12178
rect 8990 12126 9042 12178
rect 9042 12126 9044 12178
rect 8988 12124 9044 12126
rect 9436 15036 9492 15092
rect 9548 14924 9604 14980
rect 10892 25340 10948 25396
rect 10780 25116 10836 25172
rect 11340 26236 11396 26292
rect 11116 24892 11172 24948
rect 12236 28812 12292 28868
rect 12348 29372 12404 29428
rect 12180 28364 12236 28420
rect 11788 26684 11844 26740
rect 11900 28028 11956 28084
rect 11676 26572 11732 26628
rect 12012 27845 12014 27860
rect 12014 27845 12066 27860
rect 12066 27845 12068 27860
rect 12012 27804 12068 27845
rect 12124 27356 12180 27412
rect 14476 31778 14532 31780
rect 14476 31726 14478 31778
rect 14478 31726 14530 31778
rect 14530 31726 14532 31778
rect 14476 31724 14532 31726
rect 14868 31948 14924 32004
rect 14588 31276 14644 31332
rect 13804 30604 13860 30660
rect 15820 33516 15876 33572
rect 15708 33346 15764 33348
rect 15708 33294 15710 33346
rect 15710 33294 15762 33346
rect 15762 33294 15764 33346
rect 15708 33292 15764 33294
rect 14140 30994 14196 30996
rect 14140 30942 14142 30994
rect 14142 30942 14194 30994
rect 14194 30942 14196 30994
rect 14140 30940 14196 30942
rect 13468 30210 13524 30212
rect 13468 30158 13470 30210
rect 13470 30158 13522 30210
rect 13522 30158 13524 30210
rect 13468 30156 13524 30158
rect 13244 29596 13300 29652
rect 13356 30044 13412 30100
rect 12796 29372 12852 29428
rect 12684 29036 12740 29092
rect 12460 27804 12516 27860
rect 12684 27804 12740 27860
rect 12460 27020 12516 27076
rect 13020 27834 13022 27860
rect 13022 27834 13074 27860
rect 13074 27834 13076 27860
rect 13020 27804 13076 27834
rect 13244 27020 13300 27076
rect 14344 30210 14400 30212
rect 14344 30158 14346 30210
rect 14346 30158 14398 30210
rect 14398 30158 14400 30210
rect 14344 30156 14400 30158
rect 14140 29036 14196 29092
rect 15260 30380 15316 30436
rect 15484 30604 15540 30660
rect 14252 29932 14308 29988
rect 13468 27970 13524 27972
rect 13468 27918 13470 27970
rect 13470 27918 13522 27970
rect 13522 27918 13524 27970
rect 13468 27916 13524 27918
rect 14028 28476 14084 28532
rect 13804 27916 13860 27972
rect 14028 27844 14030 27860
rect 14030 27844 14082 27860
rect 14082 27844 14084 27860
rect 14028 27804 14084 27844
rect 14140 27692 14196 27748
rect 15036 30210 15092 30212
rect 15036 30158 15038 30210
rect 15038 30158 15090 30210
rect 15090 30158 15092 30210
rect 15036 30156 15092 30158
rect 14588 29372 14644 29428
rect 14364 28604 14420 28644
rect 14364 28588 14366 28604
rect 14366 28588 14418 28604
rect 14418 28588 14420 28604
rect 14476 27916 14532 27972
rect 14924 29426 14980 29428
rect 14924 29374 14926 29426
rect 14926 29374 14978 29426
rect 14978 29374 14980 29426
rect 14924 29372 14980 29374
rect 15036 29036 15092 29092
rect 14756 27858 14812 27860
rect 14756 27806 14758 27858
rect 14758 27806 14810 27858
rect 14810 27806 14812 27858
rect 14756 27804 14812 27806
rect 14364 27580 14420 27636
rect 13636 27244 13692 27300
rect 12348 26572 12404 26628
rect 13468 27020 13524 27076
rect 12124 26178 12180 26180
rect 12124 26126 12126 26178
rect 12126 26126 12178 26178
rect 12178 26126 12180 26178
rect 12124 26124 12180 26126
rect 12012 25676 12068 25732
rect 11564 24668 11620 24724
rect 11676 25116 11732 25172
rect 11228 22652 11284 22708
rect 11340 22092 11396 22148
rect 11788 24892 11844 24948
rect 12236 25564 12292 25620
rect 12460 26290 12516 26292
rect 12460 26238 12462 26290
rect 12462 26238 12514 26290
rect 12514 26238 12516 26290
rect 12460 26236 12516 26238
rect 12840 26276 12842 26292
rect 12842 26276 12894 26292
rect 12894 26276 12896 26292
rect 12840 26236 12896 26276
rect 13860 27074 13916 27076
rect 13860 27022 13862 27074
rect 13862 27022 13914 27074
rect 13914 27022 13916 27074
rect 13860 27020 13916 27022
rect 14420 27132 14476 27188
rect 14140 27074 14196 27076
rect 14140 27022 14142 27074
rect 14142 27022 14194 27074
rect 14194 27022 14196 27074
rect 14140 27020 14196 27022
rect 14252 26962 14308 26964
rect 14252 26910 14254 26962
rect 14254 26910 14306 26962
rect 14306 26910 14308 26962
rect 14252 26908 14308 26910
rect 15036 28476 15092 28532
rect 15148 28364 15204 28420
rect 15484 29596 15540 29652
rect 15596 32732 15652 32788
rect 15484 29426 15540 29428
rect 15484 29374 15486 29426
rect 15486 29374 15538 29426
rect 15538 29374 15540 29426
rect 15484 29372 15540 29374
rect 15951 32732 16007 32788
rect 18004 42754 18060 42756
rect 18004 42702 18006 42754
rect 18006 42702 18058 42754
rect 18058 42702 18060 42754
rect 18004 42700 18060 42702
rect 17724 42588 17780 42644
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 20636 44156 20692 44212
rect 20412 43820 20468 43876
rect 19740 42754 19796 42756
rect 19740 42702 19742 42754
rect 19742 42702 19794 42754
rect 19794 42702 19796 42754
rect 19740 42700 19796 42702
rect 20244 43036 20300 43092
rect 19964 42754 20020 42756
rect 19964 42702 19966 42754
rect 19966 42702 20018 42754
rect 20018 42702 20020 42754
rect 19964 42700 20020 42702
rect 20076 42924 20132 42980
rect 19572 42588 19628 42644
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 19516 41468 19572 41524
rect 17500 41132 17556 41188
rect 17836 40908 17892 40964
rect 17612 40626 17668 40628
rect 17612 40574 17614 40626
rect 17614 40574 17666 40626
rect 17666 40574 17668 40626
rect 17612 40572 17668 40574
rect 17276 40402 17332 40404
rect 17276 40350 17278 40402
rect 17278 40350 17330 40402
rect 17330 40350 17332 40402
rect 17276 40348 17332 40350
rect 17556 39730 17612 39732
rect 17556 39678 17558 39730
rect 17558 39678 17610 39730
rect 17610 39678 17612 39730
rect 17556 39676 17612 39678
rect 19404 41186 19460 41188
rect 19404 41134 19406 41186
rect 19406 41134 19458 41186
rect 19458 41134 19460 41186
rect 19404 41132 19460 41134
rect 18620 40572 18676 40628
rect 20524 43708 20580 43764
rect 20524 43484 20580 43540
rect 21756 45106 21812 45108
rect 21756 45054 21758 45106
rect 21758 45054 21810 45106
rect 21810 45054 21812 45106
rect 21756 45052 21812 45054
rect 21308 44828 21364 44884
rect 20860 43538 20916 43540
rect 20860 43486 20862 43538
rect 20862 43486 20914 43538
rect 20914 43486 20916 43538
rect 20860 43484 20916 43486
rect 21420 42924 21476 42980
rect 20524 42588 20580 42644
rect 19740 41410 19796 41412
rect 19740 41358 19742 41410
rect 19742 41358 19794 41410
rect 19794 41358 19796 41410
rect 19740 41356 19796 41358
rect 20412 41356 20468 41412
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 18228 40514 18284 40516
rect 18228 40462 18230 40514
rect 18230 40462 18282 40514
rect 18282 40462 18284 40514
rect 18228 40460 18284 40462
rect 16940 38834 16996 38836
rect 16940 38782 16942 38834
rect 16942 38782 16994 38834
rect 16994 38782 16996 38834
rect 16940 38780 16996 38782
rect 18396 39900 18452 39956
rect 16940 38108 16996 38164
rect 16604 37660 16660 37716
rect 16380 37378 16436 37380
rect 16380 37326 16382 37378
rect 16382 37326 16434 37378
rect 16434 37326 16436 37378
rect 16380 37324 16436 37326
rect 16716 37266 16772 37268
rect 16716 37214 16718 37266
rect 16718 37214 16770 37266
rect 16770 37214 16772 37266
rect 16716 37212 16772 37214
rect 17332 37212 17388 37268
rect 16492 37100 16548 37156
rect 17780 36876 17836 36932
rect 17836 36316 17892 36372
rect 16268 35196 16324 35252
rect 16716 34972 16772 35028
rect 17220 34972 17276 35028
rect 16268 33404 16324 33460
rect 17052 34860 17108 34916
rect 16772 34802 16828 34804
rect 16772 34750 16774 34802
rect 16774 34750 16826 34802
rect 16826 34750 16828 34802
rect 16772 34748 16828 34750
rect 16940 34130 16996 34132
rect 16940 34078 16942 34130
rect 16942 34078 16994 34130
rect 16994 34078 16996 34130
rect 16940 34076 16996 34078
rect 17500 34412 17556 34468
rect 17052 33628 17108 33684
rect 17836 35420 17892 35476
rect 17948 34748 18004 34804
rect 18284 38220 18340 38276
rect 18228 37826 18284 37828
rect 18228 37774 18230 37826
rect 18230 37774 18282 37826
rect 18282 37774 18284 37826
rect 18228 37772 18284 37774
rect 20300 40402 20356 40404
rect 20300 40350 20302 40402
rect 20302 40350 20354 40402
rect 20354 40350 20356 40402
rect 20300 40348 20356 40350
rect 19292 40124 19348 40180
rect 20132 39564 20188 39620
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 20188 38332 20244 38388
rect 18620 38274 18676 38276
rect 18620 38222 18622 38274
rect 18622 38222 18674 38274
rect 18674 38222 18676 38274
rect 18620 38220 18676 38222
rect 20524 40348 20580 40404
rect 21644 43820 21700 43876
rect 22316 44546 22372 44548
rect 22316 44494 22318 44546
rect 22318 44494 22370 44546
rect 22370 44494 22372 44546
rect 22316 44492 22372 44494
rect 22540 44492 22596 44548
rect 24332 45724 24388 45780
rect 23100 44268 23156 44324
rect 21980 43314 22036 43316
rect 21980 43262 21982 43314
rect 21982 43262 22034 43314
rect 22034 43262 22036 43314
rect 21980 43260 22036 43262
rect 21756 42924 21812 42980
rect 21868 43036 21924 43092
rect 21532 42812 21588 42868
rect 21756 42588 21812 42644
rect 21532 42476 21588 42532
rect 22316 42924 22372 42980
rect 21980 42866 22036 42868
rect 21980 42814 21982 42866
rect 21982 42814 22034 42866
rect 22034 42814 22036 42866
rect 21980 42812 22036 42814
rect 22148 42754 22204 42756
rect 22148 42702 22150 42754
rect 22150 42702 22202 42754
rect 22202 42702 22204 42754
rect 22148 42700 22204 42702
rect 22876 43260 22932 43316
rect 22988 43484 23044 43540
rect 22652 43036 22708 43092
rect 20412 38220 20468 38276
rect 21532 41580 21588 41636
rect 21868 41970 21924 41972
rect 21868 41918 21870 41970
rect 21870 41918 21922 41970
rect 21922 41918 21924 41970
rect 21868 41916 21924 41918
rect 21644 41356 21700 41412
rect 22484 42530 22540 42532
rect 22484 42478 22486 42530
rect 22486 42478 22538 42530
rect 22538 42478 22540 42530
rect 22484 42476 22540 42478
rect 18396 37772 18452 37828
rect 18508 37324 18564 37380
rect 18284 37242 18286 37268
rect 18286 37242 18338 37268
rect 18338 37242 18340 37268
rect 18284 37212 18340 37242
rect 19068 37324 19124 37380
rect 18620 37212 18676 37268
rect 18732 37154 18788 37156
rect 18732 37102 18734 37154
rect 18734 37102 18786 37154
rect 18786 37102 18788 37154
rect 18732 37100 18788 37102
rect 18900 37100 18956 37156
rect 19684 37938 19740 37940
rect 19684 37886 19686 37938
rect 19686 37886 19738 37938
rect 19738 37886 19740 37938
rect 19684 37884 19740 37886
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20188 37660 20244 37716
rect 20412 37660 20468 37716
rect 20580 37660 20636 37716
rect 20044 37604 20100 37606
rect 19292 37266 19348 37268
rect 19292 37214 19294 37266
rect 19294 37214 19346 37266
rect 19346 37214 19348 37266
rect 19292 37212 19348 37214
rect 20300 37212 20356 37268
rect 20076 37100 20132 37156
rect 19180 36652 19236 36708
rect 20916 40572 20972 40628
rect 21980 41020 22036 41076
rect 21532 40572 21588 40628
rect 21308 40402 21364 40404
rect 21308 40350 21310 40402
rect 21310 40350 21362 40402
rect 21362 40350 21364 40402
rect 21308 40348 21364 40350
rect 21588 40402 21644 40404
rect 21588 40350 21590 40402
rect 21590 40350 21642 40402
rect 21642 40350 21644 40402
rect 21588 40348 21644 40350
rect 21420 40236 21476 40292
rect 22764 41970 22820 41972
rect 22764 41918 22766 41970
rect 22766 41918 22818 41970
rect 22818 41918 22820 41970
rect 22764 41916 22820 41918
rect 22708 41468 22764 41524
rect 22428 41020 22484 41076
rect 23436 43260 23492 43316
rect 23548 43372 23604 43428
rect 23660 43036 23716 43092
rect 23212 42700 23268 42756
rect 22988 42476 23044 42532
rect 24220 44322 24276 44324
rect 24220 44270 24222 44322
rect 24222 44270 24274 44322
rect 24274 44270 24276 44322
rect 24220 44268 24276 44270
rect 24780 45890 24836 45892
rect 24780 45838 24782 45890
rect 24782 45838 24834 45890
rect 24834 45838 24836 45890
rect 24780 45836 24836 45838
rect 25228 45106 25284 45108
rect 25228 45054 25230 45106
rect 25230 45054 25282 45106
rect 25282 45054 25284 45106
rect 25228 45052 25284 45054
rect 25004 44546 25060 44548
rect 25004 44494 25006 44546
rect 25006 44494 25058 44546
rect 25058 44494 25060 44546
rect 25004 44492 25060 44494
rect 26012 45612 26068 45668
rect 27132 45724 27188 45780
rect 26796 45666 26852 45668
rect 26796 45614 26798 45666
rect 26798 45614 26850 45666
rect 26850 45614 26852 45666
rect 26796 45612 26852 45614
rect 27244 45500 27300 45556
rect 26236 44492 26292 44548
rect 25900 44380 25956 44436
rect 25340 44322 25396 44324
rect 25340 44270 25342 44322
rect 25342 44270 25394 44322
rect 25394 44270 25396 44322
rect 25340 44268 25396 44270
rect 25228 44044 25284 44100
rect 26908 44716 26964 44772
rect 24556 43314 24612 43316
rect 24556 43262 24558 43314
rect 24558 43262 24610 43314
rect 24610 43262 24612 43314
rect 24556 43260 24612 43262
rect 22876 41132 22932 41188
rect 23324 41916 23380 41972
rect 22092 40348 22148 40404
rect 22204 40236 22260 40292
rect 21308 39618 21364 39620
rect 21308 39566 21310 39618
rect 21310 39566 21362 39618
rect 21362 39566 21364 39618
rect 21308 39564 21364 39566
rect 22316 40124 22372 40180
rect 22184 39564 22240 39620
rect 21084 38892 21140 38948
rect 20860 38834 20916 38836
rect 20860 38782 20862 38834
rect 20862 38782 20914 38834
rect 20914 38782 20916 38834
rect 22184 39004 22240 39060
rect 20860 38780 20916 38782
rect 21196 38722 21252 38724
rect 21196 38670 21198 38722
rect 21198 38670 21250 38722
rect 21250 38670 21252 38722
rect 21196 38668 21252 38670
rect 21980 38668 22036 38724
rect 22428 38780 22484 38836
rect 22820 40402 22876 40404
rect 22820 40350 22822 40402
rect 22822 40350 22874 40402
rect 22874 40350 22876 40402
rect 22820 40348 22876 40350
rect 22540 38892 22596 38948
rect 22092 38556 22148 38612
rect 21084 38332 21140 38388
rect 22932 38722 22988 38724
rect 22932 38670 22934 38722
rect 22934 38670 22986 38722
rect 22986 38670 22988 38722
rect 22932 38668 22988 38670
rect 21084 37548 21140 37604
rect 21308 37660 21364 37716
rect 20748 37212 20804 37268
rect 20412 37100 20468 37156
rect 19292 36540 19348 36596
rect 20412 36540 20468 36596
rect 18284 35756 18340 35812
rect 18452 35868 18508 35924
rect 18788 35756 18844 35812
rect 18172 34972 18228 35028
rect 18284 35420 18340 35476
rect 18172 34802 18228 34804
rect 18172 34750 18174 34802
rect 18174 34750 18226 34802
rect 18226 34750 18228 34802
rect 18172 34748 18228 34750
rect 19068 34914 19124 34916
rect 19068 34862 19070 34914
rect 19070 34862 19122 34914
rect 19122 34862 19124 34914
rect 19068 34860 19124 34862
rect 18060 34130 18116 34132
rect 18060 34078 18062 34130
rect 18062 34078 18114 34130
rect 18114 34078 18116 34130
rect 18060 34076 18116 34078
rect 18284 34412 18340 34468
rect 17612 33740 17668 33796
rect 16492 33180 16548 33236
rect 17500 33180 17556 33236
rect 16828 32562 16884 32564
rect 16828 32510 16830 32562
rect 16830 32510 16882 32562
rect 16882 32510 16884 32562
rect 16828 32508 16884 32510
rect 18264 33315 18320 33348
rect 18264 33292 18266 33315
rect 18266 33292 18318 33315
rect 18318 33292 18320 33315
rect 18060 33180 18116 33236
rect 19964 36204 20020 36260
rect 21512 37436 21568 37492
rect 22540 37884 22596 37940
rect 22428 37436 22484 37492
rect 21644 37324 21700 37380
rect 20748 36764 20804 36820
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19740 35868 19796 35924
rect 20188 35698 20244 35700
rect 20188 35646 20190 35698
rect 20190 35646 20242 35698
rect 20242 35646 20244 35698
rect 20188 35644 20244 35646
rect 19292 35420 19348 35476
rect 19628 35420 19684 35476
rect 19516 35196 19572 35252
rect 19180 34748 19236 34804
rect 18788 34188 18844 34244
rect 18620 33740 18676 33796
rect 18508 33458 18564 33460
rect 18508 33406 18510 33458
rect 18510 33406 18562 33458
rect 18562 33406 18564 33458
rect 18508 33404 18564 33406
rect 17780 32396 17836 32452
rect 17164 32172 17220 32228
rect 17612 32172 17668 32228
rect 15708 31836 15764 31892
rect 16268 32060 16324 32116
rect 15876 31778 15932 31780
rect 15876 31726 15878 31778
rect 15878 31726 15930 31778
rect 15930 31726 15932 31778
rect 15876 31724 15932 31726
rect 16828 31836 16884 31892
rect 16492 31164 16548 31220
rect 16604 31052 16660 31108
rect 16716 31500 16772 31556
rect 17388 31836 17444 31892
rect 17164 31500 17220 31556
rect 16492 29932 16548 29988
rect 16380 29596 16436 29652
rect 15596 29036 15652 29092
rect 15260 28252 15316 28308
rect 15372 28588 15428 28644
rect 15484 28476 15540 28532
rect 15484 28252 15540 28308
rect 15036 27692 15092 27748
rect 15372 27858 15428 27860
rect 15372 27806 15374 27858
rect 15374 27806 15426 27858
rect 15426 27806 15428 27858
rect 15372 27804 15428 27806
rect 15372 27580 15428 27636
rect 13132 25676 13188 25732
rect 13562 25788 13618 25844
rect 12684 25452 12740 25508
rect 13580 25452 13636 25508
rect 13132 25004 13188 25060
rect 12124 24834 12180 24836
rect 12124 24782 12126 24834
rect 12126 24782 12178 24834
rect 12178 24782 12180 24834
rect 12124 24780 12180 24782
rect 12236 24722 12292 24724
rect 12236 24670 12238 24722
rect 12238 24670 12290 24722
rect 12290 24670 12292 24722
rect 12236 24668 12292 24670
rect 11676 23548 11732 23604
rect 12572 23324 12628 23380
rect 12684 24892 12740 24948
rect 12908 23938 12964 23940
rect 12908 23886 12910 23938
rect 12910 23886 12962 23938
rect 12962 23886 12964 23938
rect 12908 23884 12964 23886
rect 11676 22652 11732 22708
rect 10892 21756 10948 21812
rect 10556 21308 10612 21364
rect 11228 21026 11284 21028
rect 11228 20974 11230 21026
rect 11230 20974 11282 21026
rect 11282 20974 11284 21026
rect 11228 20972 11284 20974
rect 11564 20972 11620 21028
rect 11788 22092 11844 22148
rect 13020 23324 13076 23380
rect 12460 22370 12516 22372
rect 12460 22318 12462 22370
rect 12462 22318 12514 22370
rect 12514 22318 12516 22370
rect 12460 22316 12516 22318
rect 11676 20412 11732 20468
rect 10444 19404 10500 19460
rect 14140 26684 14196 26740
rect 13916 25788 13972 25844
rect 13804 25564 13860 25620
rect 14980 27356 15036 27412
rect 14812 27074 14868 27076
rect 14812 27022 14814 27074
rect 14814 27022 14866 27074
rect 14866 27022 14868 27074
rect 14812 27020 14868 27022
rect 15372 26908 15428 26964
rect 14812 26796 14868 26852
rect 18060 31500 18116 31556
rect 17668 30994 17724 30996
rect 17668 30942 17670 30994
rect 17670 30942 17722 30994
rect 17722 30942 17724 30994
rect 17668 30940 17724 30942
rect 17948 31052 18004 31108
rect 17948 30268 18004 30324
rect 18284 32732 18340 32788
rect 18620 32396 18676 32452
rect 18788 32508 18844 32564
rect 21532 37100 21588 37156
rect 20748 36092 20804 36148
rect 20860 36316 20916 36372
rect 20860 35980 20916 36036
rect 21028 36204 21084 36260
rect 20860 35756 20916 35812
rect 20076 34748 20132 34804
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 20300 34524 20356 34580
rect 19292 32508 19348 32564
rect 18956 31948 19012 32004
rect 18284 31164 18340 31220
rect 18620 31750 18676 31780
rect 18620 31724 18622 31750
rect 18622 31724 18674 31750
rect 18674 31724 18676 31750
rect 18396 30882 18452 30884
rect 18396 30830 18398 30882
rect 18398 30830 18450 30882
rect 18450 30830 18452 30882
rect 18396 30828 18452 30830
rect 18620 30994 18676 30996
rect 18620 30942 18622 30994
rect 18622 30942 18674 30994
rect 18674 30942 18676 30994
rect 18620 30940 18676 30942
rect 18732 30828 18788 30884
rect 18340 30156 18396 30212
rect 18508 30268 18564 30324
rect 17500 29932 17556 29988
rect 17556 29148 17612 29204
rect 15596 27804 15652 27860
rect 14308 25506 14364 25508
rect 14308 25454 14310 25506
rect 14310 25454 14362 25506
rect 14362 25454 14364 25506
rect 14308 25452 14364 25454
rect 14924 25506 14980 25508
rect 14924 25454 14926 25506
rect 14926 25454 14978 25506
rect 14978 25454 14980 25506
rect 14924 25452 14980 25454
rect 14476 25394 14532 25396
rect 14476 25342 14478 25394
rect 14478 25342 14530 25394
rect 14530 25342 14532 25394
rect 14476 25340 14532 25342
rect 15484 26124 15540 26180
rect 15372 26012 15428 26068
rect 15148 25788 15204 25844
rect 15036 25340 15092 25396
rect 14028 25116 14084 25172
rect 13356 22316 13412 22372
rect 13468 23548 13524 23604
rect 14140 23938 14196 23940
rect 14140 23886 14142 23938
rect 14142 23886 14194 23938
rect 14194 23886 14196 23938
rect 14140 23884 14196 23886
rect 14364 23884 14420 23940
rect 15484 25452 15540 25508
rect 15596 27468 15652 27524
rect 15708 25506 15764 25508
rect 15708 25454 15710 25506
rect 15710 25454 15762 25506
rect 15762 25454 15764 25506
rect 15708 25452 15764 25454
rect 15148 23884 15204 23940
rect 13916 23324 13972 23380
rect 13748 22652 13804 22708
rect 13692 21868 13748 21924
rect 14196 22876 14252 22932
rect 14140 22316 14196 22372
rect 14028 21980 14084 22036
rect 14700 22594 14756 22596
rect 14700 22542 14702 22594
rect 14702 22542 14754 22594
rect 14754 22542 14756 22594
rect 14700 22540 14756 22542
rect 15372 22428 15428 22484
rect 15092 22370 15148 22372
rect 15092 22318 15094 22370
rect 15094 22318 15146 22370
rect 15146 22318 15148 22370
rect 15092 22316 15148 22318
rect 14588 21644 14644 21700
rect 14700 22092 14756 22148
rect 15372 22092 15428 22148
rect 14812 21756 14868 21812
rect 15186 21644 15242 21700
rect 16940 27804 16996 27860
rect 17720 28476 17776 28532
rect 17612 27020 17668 27076
rect 16212 26012 16268 26068
rect 16604 25900 16660 25956
rect 16492 24892 16548 24948
rect 16380 24498 16436 24500
rect 16380 24446 16382 24498
rect 16382 24446 16434 24498
rect 16434 24446 16436 24498
rect 16380 24444 16436 24446
rect 16940 26290 16996 26292
rect 16940 26238 16942 26290
rect 16942 26238 16994 26290
rect 16994 26238 16996 26290
rect 16940 26236 16996 26238
rect 17556 26178 17612 26180
rect 17556 26126 17558 26178
rect 17558 26126 17610 26178
rect 17610 26126 17612 26178
rect 17556 26124 17612 26126
rect 17948 29596 18004 29652
rect 18172 28924 18228 28980
rect 17948 28476 18004 28532
rect 18284 28476 18340 28532
rect 18284 27858 18340 27860
rect 18284 27806 18286 27858
rect 18286 27806 18338 27858
rect 18338 27806 18340 27858
rect 18284 27804 18340 27806
rect 18844 30492 18900 30548
rect 18844 29708 18900 29764
rect 19404 33068 19460 33124
rect 19404 32060 19460 32116
rect 19404 31052 19460 31108
rect 18620 28924 18676 28980
rect 19964 34300 20020 34356
rect 20076 33404 20132 33460
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19628 31724 19684 31780
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 20188 31052 20244 31108
rect 19516 30828 19572 30884
rect 20132 30882 20188 30884
rect 20132 30830 20134 30882
rect 20134 30830 20186 30882
rect 20186 30830 20188 30882
rect 20132 30828 20188 30830
rect 20076 30492 20132 30548
rect 19516 30268 19572 30324
rect 21084 34860 21140 34916
rect 20748 33740 20804 33796
rect 21364 36482 21420 36484
rect 21364 36430 21366 36482
rect 21366 36430 21418 36482
rect 21418 36430 21420 36482
rect 21364 36428 21420 36430
rect 21308 35980 21364 36036
rect 22316 37324 22372 37380
rect 21756 37266 21812 37268
rect 21756 37214 21758 37266
rect 21758 37214 21810 37266
rect 21810 37214 21812 37266
rect 21756 37212 21812 37214
rect 21644 35980 21700 36036
rect 21756 36988 21812 37044
rect 21308 35532 21364 35588
rect 21308 34300 21364 34356
rect 20972 34106 20974 34132
rect 20974 34106 21026 34132
rect 21026 34106 21028 34132
rect 22204 37100 22260 37156
rect 21980 36482 22036 36484
rect 21980 36430 21982 36482
rect 21982 36430 22034 36482
rect 22034 36430 22036 36482
rect 21980 36428 22036 36430
rect 22820 38220 22876 38276
rect 22652 37266 22708 37268
rect 22652 37214 22654 37266
rect 22654 37214 22706 37266
rect 22706 37214 22708 37266
rect 22652 37212 22708 37214
rect 21588 35586 21644 35588
rect 21588 35534 21590 35586
rect 21590 35534 21642 35586
rect 21642 35534 21644 35586
rect 21588 35532 21644 35534
rect 21868 35980 21924 36036
rect 21868 35308 21924 35364
rect 21980 35196 22036 35252
rect 20972 34076 21028 34106
rect 21756 34914 21812 34916
rect 21756 34862 21758 34914
rect 21758 34862 21810 34914
rect 21810 34862 21812 34914
rect 21756 34860 21812 34862
rect 21644 34076 21700 34132
rect 21532 33852 21588 33908
rect 21364 33740 21420 33796
rect 20412 31948 20468 32004
rect 20804 32956 20860 33012
rect 20748 32562 20804 32564
rect 20748 32510 20750 32562
rect 20750 32510 20802 32562
rect 20802 32510 20804 32562
rect 20748 32508 20804 32510
rect 20412 31052 20468 31108
rect 20524 30716 20580 30772
rect 20636 30940 20692 30996
rect 20636 30268 20692 30324
rect 22484 36706 22540 36708
rect 22484 36654 22486 36706
rect 22486 36654 22538 36706
rect 22538 36654 22540 36706
rect 22484 36652 22540 36654
rect 22428 35532 22484 35588
rect 22428 35308 22484 35364
rect 22428 35084 22484 35140
rect 22540 34860 22596 34916
rect 23212 41186 23268 41188
rect 23212 41134 23214 41186
rect 23214 41134 23266 41186
rect 23266 41134 23268 41186
rect 23212 41132 23268 41134
rect 23436 41692 23492 41748
rect 23548 41020 23604 41076
rect 23324 40684 23380 40740
rect 23996 41244 24052 41300
rect 23828 41186 23884 41188
rect 23828 41134 23830 41186
rect 23830 41134 23882 41186
rect 23882 41134 23884 41186
rect 23828 41132 23884 41134
rect 24892 42252 24948 42308
rect 24444 41970 24500 41972
rect 24444 41918 24446 41970
rect 24446 41918 24498 41970
rect 24498 41918 24500 41970
rect 24444 41916 24500 41918
rect 24780 41580 24836 41636
rect 24724 40626 24780 40628
rect 24724 40574 24726 40626
rect 24726 40574 24778 40626
rect 24778 40574 24780 40626
rect 24724 40572 24780 40574
rect 23660 39452 23716 39508
rect 23660 39228 23716 39284
rect 23492 39116 23548 39172
rect 24444 39228 24500 39284
rect 23996 38668 24052 38724
rect 23324 38220 23380 38276
rect 23212 38162 23268 38164
rect 23212 38110 23214 38162
rect 23214 38110 23266 38162
rect 23266 38110 23268 38162
rect 23212 38108 23268 38110
rect 22876 37154 22932 37156
rect 22876 37102 22878 37154
rect 22878 37102 22930 37154
rect 22930 37102 22932 37154
rect 22876 37100 22932 37102
rect 23548 38444 23604 38500
rect 23660 38108 23716 38164
rect 24612 38444 24668 38500
rect 23492 36988 23548 37044
rect 24220 37884 24276 37940
rect 24780 37324 24836 37380
rect 25452 42700 25508 42756
rect 25900 43538 25956 43540
rect 25900 43486 25902 43538
rect 25902 43486 25954 43538
rect 25954 43486 25956 43538
rect 25900 43484 25956 43486
rect 26796 43538 26852 43540
rect 26796 43486 26830 43538
rect 26830 43486 26852 43538
rect 26796 43484 26852 43486
rect 25900 42754 25956 42756
rect 25900 42702 25902 42754
rect 25902 42702 25954 42754
rect 25954 42702 25956 42754
rect 25900 42700 25956 42702
rect 27020 44604 27076 44660
rect 27580 45164 27636 45220
rect 27916 44994 27972 44996
rect 27916 44942 27918 44994
rect 27918 44942 27970 44994
rect 27970 44942 27972 44994
rect 27916 44940 27972 44942
rect 28252 44940 28308 44996
rect 28364 45388 28420 45444
rect 27804 44716 27860 44772
rect 27244 44380 27300 44436
rect 27804 44156 27860 44212
rect 27580 43820 27636 43876
rect 28196 44322 28252 44324
rect 28196 44270 28198 44322
rect 28198 44270 28250 44322
rect 28250 44270 28252 44322
rect 28196 44268 28252 44270
rect 28868 44604 28924 44660
rect 29708 45890 29764 45892
rect 29708 45838 29710 45890
rect 29710 45838 29762 45890
rect 29762 45838 29764 45890
rect 29708 45836 29764 45838
rect 29204 45500 29260 45556
rect 27916 44044 27972 44100
rect 28364 44044 28420 44100
rect 29148 44940 29204 44996
rect 29708 45106 29764 45108
rect 29708 45054 29710 45106
rect 29710 45054 29762 45106
rect 29762 45054 29764 45106
rect 29708 45052 29764 45054
rect 30156 46956 30212 47012
rect 29988 45388 30044 45444
rect 27804 43596 27860 43652
rect 27356 43538 27412 43540
rect 27356 43486 27358 43538
rect 27358 43486 27410 43538
rect 27410 43486 27412 43538
rect 27356 43484 27412 43486
rect 27692 43538 27748 43540
rect 27692 43486 27694 43538
rect 27694 43486 27746 43538
rect 27746 43486 27748 43538
rect 27692 43484 27748 43486
rect 26796 42028 26852 42084
rect 26236 41916 26292 41972
rect 26104 41804 26160 41860
rect 26124 41580 26180 41636
rect 25452 41298 25508 41300
rect 25452 41246 25454 41298
rect 25454 41246 25506 41298
rect 25506 41246 25508 41298
rect 25452 41244 25508 41246
rect 25116 41186 25172 41188
rect 25116 41134 25118 41186
rect 25118 41134 25170 41186
rect 25170 41134 25172 41186
rect 25116 41132 25172 41134
rect 25788 40572 25844 40628
rect 25340 40124 25396 40180
rect 25004 38892 25060 38948
rect 25676 40236 25732 40292
rect 25788 40124 25844 40180
rect 28252 43516 28254 43540
rect 28254 43516 28306 43540
rect 28306 43516 28308 43540
rect 28252 43484 28308 43516
rect 28084 43148 28140 43204
rect 28232 43260 28288 43316
rect 27188 41970 27244 41972
rect 27188 41918 27190 41970
rect 27190 41918 27242 41970
rect 27242 41918 27244 41970
rect 27188 41916 27244 41918
rect 27468 41804 27524 41860
rect 26908 41580 26964 41636
rect 26348 41132 26404 41188
rect 26572 41186 26628 41188
rect 26572 41134 26574 41186
rect 26574 41134 26626 41186
rect 26626 41134 26628 41186
rect 26572 41132 26628 41134
rect 27132 40684 27188 40740
rect 26964 40290 27020 40292
rect 26964 40238 26966 40290
rect 26966 40238 27018 40290
rect 27018 40238 27020 40290
rect 26964 40236 27020 40238
rect 26684 40124 26740 40180
rect 25676 39228 25732 39284
rect 25564 39116 25620 39172
rect 25452 38332 25508 38388
rect 25340 38220 25396 38276
rect 22764 35084 22820 35140
rect 22876 35308 22932 35364
rect 23324 35196 23380 35252
rect 21868 34188 21924 34244
rect 22036 33964 22092 34020
rect 21196 32732 21252 32788
rect 21868 33852 21924 33908
rect 21868 33292 21924 33348
rect 21644 32956 21700 33012
rect 22204 33852 22260 33908
rect 22316 33740 22372 33796
rect 22428 34076 22484 34132
rect 21308 31612 21364 31668
rect 21980 32060 22036 32116
rect 22204 33628 22260 33684
rect 21980 31890 22036 31892
rect 21980 31838 21982 31890
rect 21982 31838 22034 31890
rect 22034 31838 22036 31890
rect 21980 31836 22036 31838
rect 20748 31164 20804 31220
rect 22540 33852 22596 33908
rect 23660 34412 23716 34468
rect 23772 34300 23828 34356
rect 23548 33964 23604 34020
rect 23324 33906 23380 33908
rect 23324 33854 23326 33906
rect 23326 33854 23378 33906
rect 23378 33854 23380 33906
rect 23324 33852 23380 33854
rect 23772 34130 23828 34132
rect 23772 34078 23774 34130
rect 23774 34078 23826 34130
rect 23826 34078 23828 34130
rect 23772 34076 23828 34078
rect 23772 33852 23828 33908
rect 24444 35586 24500 35588
rect 24444 35534 24446 35586
rect 24446 35534 24498 35586
rect 24498 35534 24500 35586
rect 24444 35532 24500 35534
rect 25116 34412 25172 34468
rect 24276 33906 24332 33908
rect 24276 33854 24278 33906
rect 24278 33854 24330 33906
rect 24330 33854 24332 33906
rect 24276 33852 24332 33854
rect 22988 33628 23044 33684
rect 22204 31612 22260 31668
rect 21756 31052 21812 31108
rect 20972 30828 21028 30884
rect 20860 30604 20916 30660
rect 20412 30044 20468 30100
rect 19628 29708 19684 29764
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 18956 29148 19012 29204
rect 19404 29148 19460 29204
rect 19180 28476 19236 28532
rect 18508 27132 18564 27188
rect 18508 26908 18564 26964
rect 18396 26572 18452 26628
rect 17948 26236 18004 26292
rect 16716 25004 16772 25060
rect 16604 24332 16660 24388
rect 17052 24444 17108 24500
rect 15988 22370 16044 22372
rect 15988 22318 15990 22370
rect 15990 22318 16042 22370
rect 16042 22318 16044 22370
rect 15988 22316 16044 22318
rect 15820 22204 15876 22260
rect 15820 21868 15876 21924
rect 16156 21756 16212 21812
rect 13580 20972 13636 21028
rect 11676 19068 11732 19124
rect 12236 18620 12292 18676
rect 11788 16828 11844 16884
rect 11340 15484 11396 15540
rect 11564 16604 11620 16660
rect 10332 15372 10388 15428
rect 10220 15148 10276 15204
rect 10332 15036 10388 15092
rect 10108 14924 10164 14980
rect 10614 14812 10670 14868
rect 10332 14476 10388 14532
rect 10108 14252 10164 14308
rect 9548 13580 9604 13636
rect 9436 12124 9492 12180
rect 10220 13746 10276 13748
rect 10220 13694 10222 13746
rect 10222 13694 10274 13746
rect 10274 13694 10276 13746
rect 10220 13692 10276 13694
rect 13020 19740 13076 19796
rect 14364 20914 14420 20916
rect 14364 20862 14366 20914
rect 14366 20862 14418 20914
rect 14418 20862 14420 20914
rect 14364 20860 14420 20862
rect 14252 20748 14308 20804
rect 13412 20130 13468 20132
rect 13412 20078 13414 20130
rect 13414 20078 13466 20130
rect 13466 20078 13468 20130
rect 13412 20076 13468 20078
rect 12236 17836 12292 17892
rect 13132 18425 13134 18452
rect 13134 18425 13186 18452
rect 13186 18425 13188 18452
rect 13132 18396 13188 18425
rect 12124 16994 12180 16996
rect 12124 16942 12126 16994
rect 12126 16942 12178 16994
rect 12178 16942 12180 16994
rect 12124 16940 12180 16942
rect 12012 15986 12068 15988
rect 12012 15934 12014 15986
rect 12014 15934 12066 15986
rect 12066 15934 12068 15986
rect 12012 15932 12068 15934
rect 10444 14364 10500 14420
rect 10892 14364 10948 14420
rect 12460 17948 12516 18004
rect 12796 17666 12852 17668
rect 12796 17614 12798 17666
rect 12798 17614 12850 17666
rect 12850 17614 12852 17666
rect 12796 17612 12852 17614
rect 13020 17612 13076 17668
rect 12628 16658 12684 16660
rect 12628 16606 12630 16658
rect 12630 16606 12682 16658
rect 12682 16606 12684 16658
rect 12628 16604 12684 16606
rect 12572 15260 12628 15316
rect 12908 16098 12964 16100
rect 12908 16046 12910 16098
rect 12910 16046 12962 16098
rect 12962 16046 12964 16098
rect 12908 16044 12964 16046
rect 12796 15932 12852 15988
rect 13356 17052 13412 17108
rect 13972 20524 14028 20580
rect 14756 20802 14812 20804
rect 14756 20750 14758 20802
rect 14758 20750 14810 20802
rect 14810 20750 14812 20802
rect 14756 20748 14812 20750
rect 15484 21308 15540 21364
rect 15148 20972 15204 21028
rect 14924 20636 14980 20692
rect 13692 20076 13748 20132
rect 13804 20018 13860 20020
rect 13804 19966 13806 20018
rect 13806 19966 13858 20018
rect 13858 19966 13860 20018
rect 14364 20076 14420 20132
rect 13804 19964 13860 19966
rect 14532 19906 14588 19908
rect 14532 19854 14534 19906
rect 14534 19854 14586 19906
rect 14586 19854 14588 19906
rect 14532 19852 14588 19854
rect 15036 20524 15092 20580
rect 15036 20188 15092 20244
rect 14812 20076 14868 20132
rect 15540 20972 15596 21028
rect 15708 20076 15764 20132
rect 14924 20018 14980 20020
rect 14924 19966 14926 20018
rect 14926 19966 14978 20018
rect 14978 19966 14980 20018
rect 14924 19964 14980 19966
rect 14140 19292 14196 19348
rect 14028 19234 14084 19236
rect 14028 19182 14030 19234
rect 14030 19182 14082 19234
rect 14082 19182 14084 19234
rect 14028 19180 14084 19182
rect 14308 19122 14364 19124
rect 14308 19070 14310 19122
rect 14310 19070 14362 19122
rect 14362 19070 14364 19122
rect 14308 19068 14364 19070
rect 14700 19516 14756 19572
rect 15036 19516 15092 19572
rect 15260 19404 15316 19460
rect 15036 19292 15092 19348
rect 15148 19068 15204 19124
rect 13916 18284 13972 18340
rect 13580 16098 13636 16100
rect 13580 16046 13582 16098
rect 13582 16046 13634 16098
rect 13634 16046 13636 16098
rect 13580 16044 13636 16046
rect 13412 15820 13468 15876
rect 13580 15538 13636 15540
rect 13580 15486 13582 15538
rect 13582 15486 13634 15538
rect 13634 15486 13636 15538
rect 13580 15484 13636 15486
rect 12348 14924 12404 14980
rect 13468 15148 13524 15204
rect 15428 19628 15484 19684
rect 15988 21308 16044 21364
rect 16044 20412 16100 20468
rect 15932 20018 15988 20020
rect 15932 19966 15934 20018
rect 15934 19966 15986 20018
rect 15986 19966 15988 20018
rect 15932 19964 15988 19966
rect 15820 19740 15876 19796
rect 16436 21474 16492 21476
rect 16436 21422 16438 21474
rect 16438 21422 16490 21474
rect 16490 21422 16492 21474
rect 16436 21420 16492 21422
rect 16268 20300 16324 20356
rect 16604 20748 16660 20804
rect 17500 24946 17556 24948
rect 17500 24894 17502 24946
rect 17502 24894 17554 24946
rect 17554 24894 17556 24946
rect 17500 24892 17556 24894
rect 17948 23548 18004 23604
rect 17500 22988 17556 23044
rect 16996 22540 17052 22596
rect 16996 22370 17052 22372
rect 16996 22318 16998 22370
rect 16998 22318 17050 22370
rect 17050 22318 17052 22370
rect 16996 22316 17052 22318
rect 17388 22092 17444 22148
rect 17276 21756 17332 21812
rect 16884 21586 16940 21588
rect 16884 21534 16886 21586
rect 16886 21534 16938 21586
rect 16938 21534 16940 21586
rect 16884 21532 16940 21534
rect 16716 21084 16772 21140
rect 16492 20578 16548 20580
rect 16492 20526 16494 20578
rect 16494 20526 16546 20578
rect 16546 20526 16548 20578
rect 16492 20524 16548 20526
rect 16604 20412 16660 20468
rect 16716 20300 16772 20356
rect 16380 20018 16436 20020
rect 16380 19966 16382 20018
rect 16382 19966 16434 20018
rect 16434 19966 16436 20018
rect 16380 19964 16436 19966
rect 16268 19740 16324 19796
rect 15708 19068 15764 19124
rect 15820 19180 15876 19236
rect 16156 19404 16212 19460
rect 15596 18956 15652 19012
rect 15932 18956 15988 19012
rect 15820 18844 15876 18900
rect 15260 18396 15316 18452
rect 14198 17836 14254 17892
rect 15932 18450 15988 18452
rect 15932 18398 15934 18450
rect 15934 18398 15986 18450
rect 15986 18398 15988 18450
rect 15932 18396 15988 18398
rect 14476 17666 14532 17668
rect 14476 17614 14478 17666
rect 14478 17614 14530 17666
rect 14530 17614 14532 17666
rect 14476 17612 14532 17614
rect 16044 18172 16100 18228
rect 15092 17052 15148 17108
rect 16380 18844 16436 18900
rect 16828 19964 16884 20020
rect 17164 21532 17220 21588
rect 17164 20802 17220 20804
rect 17164 20750 17166 20802
rect 17166 20750 17218 20802
rect 17218 20750 17220 20802
rect 17164 20748 17220 20750
rect 16940 19852 16996 19908
rect 16772 19404 16828 19460
rect 16604 18844 16660 18900
rect 17164 19346 17220 19348
rect 17164 19294 17166 19346
rect 17166 19294 17218 19346
rect 17218 19294 17220 19346
rect 17164 19292 17220 19294
rect 16940 18508 16996 18564
rect 17052 19180 17108 19236
rect 16492 18060 16548 18116
rect 17780 22428 17836 22484
rect 18060 22370 18116 22372
rect 18060 22318 18062 22370
rect 18062 22318 18114 22370
rect 18114 22318 18116 22370
rect 18060 22316 18116 22318
rect 17612 21644 17668 21700
rect 17836 21868 17892 21924
rect 18396 25618 18452 25620
rect 18396 25566 18398 25618
rect 18398 25566 18450 25618
rect 18450 25566 18452 25618
rect 18396 25564 18452 25566
rect 18956 27186 19012 27188
rect 18956 27134 18958 27186
rect 18958 27134 19010 27186
rect 19010 27134 19012 27186
rect 18956 27132 19012 27134
rect 18732 26796 18788 26852
rect 18844 26908 18900 26964
rect 18620 25676 18676 25732
rect 18732 25788 18788 25844
rect 18508 25452 18564 25508
rect 18956 26572 19012 26628
rect 19516 28812 19572 28868
rect 19740 29596 19796 29652
rect 20020 29426 20076 29428
rect 20020 29374 20022 29426
rect 20022 29374 20074 29426
rect 20074 29374 20076 29426
rect 20020 29372 20076 29374
rect 20524 29372 20580 29428
rect 20412 29314 20468 29316
rect 20412 29262 20414 29314
rect 20414 29262 20466 29314
rect 20466 29262 20468 29314
rect 20412 29260 20468 29262
rect 19852 28812 19908 28868
rect 19740 28642 19796 28644
rect 19740 28590 19742 28642
rect 19742 28590 19794 28642
rect 19794 28590 19796 28642
rect 19740 28588 19796 28590
rect 19516 28476 19572 28532
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19740 28028 19796 28084
rect 20412 28700 20468 28756
rect 20300 28642 20356 28644
rect 20300 28590 20302 28642
rect 20302 28590 20354 28642
rect 20354 28590 20356 28642
rect 20300 28588 20356 28590
rect 20524 28476 20580 28532
rect 19740 27132 19796 27188
rect 19404 27020 19460 27076
rect 20748 29932 20804 29988
rect 21644 30716 21700 30772
rect 21420 30604 21476 30660
rect 21084 29932 21140 29988
rect 21196 29484 21252 29540
rect 20860 29372 20916 29428
rect 21084 29148 21140 29204
rect 20916 28588 20972 28644
rect 20636 27692 20692 27748
rect 20300 27244 20356 27300
rect 20300 27074 20356 27076
rect 20300 27022 20302 27074
rect 20302 27022 20354 27074
rect 20354 27022 20356 27074
rect 20300 27020 20356 27022
rect 19068 25788 19124 25844
rect 18956 25506 19012 25508
rect 18956 25454 18958 25506
rect 18958 25454 19010 25506
rect 19010 25454 19012 25506
rect 18956 25452 19012 25454
rect 18284 23324 18340 23380
rect 18284 23154 18340 23156
rect 18284 23102 18286 23154
rect 18286 23102 18338 23154
rect 18338 23102 18340 23154
rect 18284 23100 18340 23102
rect 19292 25340 19348 25396
rect 18844 23660 18900 23716
rect 18732 23548 18788 23604
rect 19964 26796 20020 26852
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19740 26348 19796 26404
rect 20412 26348 20468 26404
rect 20524 27468 20580 27524
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20972 27244 21028 27300
rect 21420 28924 21476 28980
rect 21420 28700 21476 28756
rect 22540 32060 22596 32116
rect 22988 31948 23044 32004
rect 22428 31724 22484 31780
rect 21980 30492 22036 30548
rect 21868 30044 21924 30100
rect 21756 29820 21812 29876
rect 23212 32620 23268 32676
rect 23548 32674 23604 32676
rect 23548 32622 23550 32674
rect 23550 32622 23602 32674
rect 23602 32622 23604 32674
rect 23548 32620 23604 32622
rect 23772 33628 23828 33684
rect 23772 33404 23828 33460
rect 23772 32956 23828 33012
rect 23100 31388 23156 31444
rect 23772 31948 23828 32004
rect 23212 30994 23268 30996
rect 23212 30942 23214 30994
rect 23214 30942 23266 30994
rect 23266 30942 23268 30994
rect 23212 30940 23268 30942
rect 23604 31388 23660 31444
rect 23548 31052 23604 31108
rect 22540 30210 22596 30212
rect 22540 30158 22542 30210
rect 22542 30158 22594 30210
rect 22594 30158 22596 30210
rect 22540 30156 22596 30158
rect 22540 29596 22596 29652
rect 22764 29596 22820 29652
rect 22316 29484 22372 29540
rect 21812 29426 21868 29428
rect 21812 29374 21814 29426
rect 21814 29374 21866 29426
rect 21866 29374 21868 29426
rect 21812 29372 21868 29374
rect 22204 29426 22260 29428
rect 22204 29374 22206 29426
rect 22206 29374 22258 29426
rect 22258 29374 22260 29426
rect 22204 29372 22260 29374
rect 21532 29148 21588 29204
rect 21308 26908 21364 26964
rect 21196 26796 21252 26852
rect 21700 28866 21756 28868
rect 21700 28814 21702 28866
rect 21702 28814 21754 28866
rect 21754 28814 21756 28866
rect 21700 28812 21756 28814
rect 22260 28642 22316 28644
rect 22260 28590 22262 28642
rect 22262 28590 22314 28642
rect 22314 28590 22316 28642
rect 22260 28588 22316 28590
rect 22428 28812 22484 28868
rect 22652 29260 22708 29316
rect 21700 27186 21756 27188
rect 21700 27134 21702 27186
rect 21702 27134 21754 27186
rect 21754 27134 21756 27186
rect 21700 27132 21756 27134
rect 22260 27074 22316 27076
rect 22260 27022 22262 27074
rect 22262 27022 22314 27074
rect 22314 27022 22316 27074
rect 22260 27020 22316 27022
rect 21980 26908 22036 26964
rect 21196 25452 21252 25508
rect 20804 25394 20860 25396
rect 20804 25342 20806 25394
rect 20806 25342 20858 25394
rect 20858 25342 20860 25394
rect 20804 25340 20860 25342
rect 19404 24220 19460 24276
rect 20188 24332 20244 24388
rect 20188 23884 20244 23940
rect 19180 23660 19236 23716
rect 18620 23100 18676 23156
rect 18396 22316 18452 22372
rect 18172 21756 18228 21812
rect 18284 21868 18340 21924
rect 17948 21586 18004 21588
rect 17948 21534 17950 21586
rect 17950 21534 18002 21586
rect 18002 21534 18004 21586
rect 18844 22370 18900 22372
rect 18844 22318 18846 22370
rect 18846 22318 18898 22370
rect 18898 22318 18900 22370
rect 18844 22316 18900 22318
rect 17948 21532 18004 21534
rect 17668 20972 17724 21028
rect 17612 20802 17668 20804
rect 17612 20750 17614 20802
rect 17614 20750 17666 20802
rect 17666 20750 17668 20802
rect 18116 20972 18172 21028
rect 18340 21308 18396 21364
rect 17612 20748 17668 20750
rect 17500 20524 17556 20580
rect 17780 20524 17836 20580
rect 17780 20188 17836 20244
rect 19292 23548 19348 23604
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 20076 22930 20132 22932
rect 20076 22878 20078 22930
rect 20078 22878 20130 22930
rect 20130 22878 20132 22930
rect 20076 22876 20132 22878
rect 19068 21868 19124 21924
rect 19628 22204 19684 22260
rect 20076 22092 20132 22148
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 21532 25340 21588 25396
rect 23436 29484 23492 29540
rect 22876 28140 22932 28196
rect 22988 29372 23044 29428
rect 23212 29036 23268 29092
rect 23100 28866 23156 28868
rect 23100 28814 23102 28866
rect 23102 28814 23154 28866
rect 23154 28814 23156 28866
rect 23100 28812 23156 28814
rect 26236 39618 26292 39620
rect 26236 39566 26238 39618
rect 26238 39566 26290 39618
rect 26290 39566 26292 39618
rect 26236 39564 26292 39566
rect 26124 39116 26180 39172
rect 26124 38220 26180 38276
rect 25620 37548 25676 37604
rect 25564 37324 25620 37380
rect 25956 37660 26012 37716
rect 25564 36594 25620 36596
rect 25564 36542 25566 36594
rect 25566 36542 25618 36594
rect 25618 36542 25620 36594
rect 25564 36540 25620 36542
rect 25340 35308 25396 35364
rect 25452 35084 25508 35140
rect 25452 34188 25508 34244
rect 25396 34018 25452 34020
rect 25396 33966 25398 34018
rect 25398 33966 25450 34018
rect 25450 33966 25452 34018
rect 25396 33964 25452 33966
rect 25228 33740 25284 33796
rect 25116 33628 25172 33684
rect 25340 33404 25396 33460
rect 25116 33292 25172 33348
rect 25004 32172 25060 32228
rect 23884 31836 23940 31892
rect 23996 31500 24052 31556
rect 23884 31276 23940 31332
rect 24556 31948 24612 32004
rect 24780 31500 24836 31556
rect 24892 31388 24948 31444
rect 24668 31052 24724 31108
rect 23660 30492 23716 30548
rect 24276 30994 24332 30996
rect 24276 30942 24278 30994
rect 24278 30942 24330 30994
rect 24330 30942 24332 30994
rect 24276 30940 24332 30942
rect 23996 29932 24052 29988
rect 23828 29650 23884 29652
rect 23828 29598 23830 29650
rect 23830 29598 23882 29650
rect 23882 29598 23884 29650
rect 23828 29596 23884 29598
rect 23436 28364 23492 28420
rect 22652 27692 22708 27748
rect 23100 27692 23156 27748
rect 23100 27132 23156 27188
rect 22876 27046 22932 27076
rect 22876 27020 22878 27046
rect 22878 27020 22930 27046
rect 22930 27020 22932 27046
rect 23660 27020 23716 27076
rect 22540 26908 22596 26964
rect 23212 26908 23268 26964
rect 22316 24892 22372 24948
rect 23884 28700 23940 28756
rect 24220 29596 24276 29652
rect 24332 29260 24388 29316
rect 24556 29484 24612 29540
rect 24668 30044 24724 30100
rect 24220 28642 24276 28644
rect 24220 28590 24222 28642
rect 24222 28590 24274 28642
rect 24274 28590 24276 28642
rect 24220 28588 24276 28590
rect 24444 28252 24500 28308
rect 24108 27132 24164 27188
rect 23492 26402 23548 26404
rect 23492 26350 23494 26402
rect 23494 26350 23546 26402
rect 23546 26350 23548 26402
rect 23492 26348 23548 26350
rect 22428 25340 22484 25396
rect 22204 24780 22260 24836
rect 22092 24668 22148 24724
rect 20636 24050 20692 24052
rect 20636 23998 20638 24050
rect 20638 23998 20690 24050
rect 20690 23998 20692 24050
rect 20636 23996 20692 23998
rect 20412 23154 20468 23156
rect 20412 23102 20414 23154
rect 20414 23102 20466 23154
rect 20466 23102 20468 23154
rect 20412 23100 20468 23102
rect 21532 23938 21588 23940
rect 21532 23886 21534 23938
rect 21534 23886 21586 23938
rect 21586 23886 21588 23938
rect 21532 23884 21588 23886
rect 21924 23938 21980 23940
rect 21924 23886 21926 23938
rect 21926 23886 21978 23938
rect 21978 23886 21980 23938
rect 21924 23884 21980 23886
rect 21084 23154 21140 23156
rect 21084 23102 21086 23154
rect 21086 23102 21138 23154
rect 21138 23102 21140 23154
rect 21084 23100 21140 23102
rect 18900 21084 18956 21140
rect 18732 20802 18788 20804
rect 18732 20750 18734 20802
rect 18734 20750 18786 20802
rect 18786 20750 18788 20802
rect 18732 20748 18788 20750
rect 19068 20412 19124 20468
rect 20692 21810 20748 21812
rect 20692 21758 20694 21810
rect 20694 21758 20746 21810
rect 20746 21758 20748 21810
rect 20692 21756 20748 21758
rect 20188 20774 20244 20804
rect 20188 20748 20190 20774
rect 20190 20748 20242 20774
rect 20242 20748 20244 20774
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 17500 20018 17556 20020
rect 17500 19966 17502 20018
rect 17502 19966 17554 20018
rect 17554 19966 17556 20018
rect 17500 19964 17556 19966
rect 19572 20130 19628 20132
rect 19572 20078 19574 20130
rect 19574 20078 19626 20130
rect 19626 20078 19628 20130
rect 19572 20076 19628 20078
rect 18340 19628 18396 19684
rect 18060 19234 18116 19236
rect 18060 19182 18062 19234
rect 18062 19182 18114 19234
rect 18114 19182 18116 19234
rect 18060 19180 18116 19182
rect 17780 19122 17836 19124
rect 17780 19070 17782 19122
rect 17782 19070 17834 19122
rect 17834 19070 17836 19122
rect 17780 19068 17836 19070
rect 17276 18396 17332 18452
rect 17388 18284 17444 18340
rect 16604 17388 16660 17444
rect 16268 16940 16324 16996
rect 16156 16828 16212 16884
rect 14364 16380 14420 16436
rect 14924 15932 14980 15988
rect 14756 15820 14812 15876
rect 14196 15314 14252 15316
rect 14196 15262 14198 15314
rect 14198 15262 14250 15314
rect 14250 15262 14252 15314
rect 14196 15260 14252 15262
rect 12460 14530 12516 14532
rect 12460 14478 12462 14530
rect 12462 14478 12514 14530
rect 12514 14478 12516 14530
rect 12460 14476 12516 14478
rect 12852 14924 12908 14980
rect 12348 14364 12404 14420
rect 11900 14140 11956 14196
rect 9100 11394 9156 11396
rect 9100 11342 9102 11394
rect 9102 11342 9154 11394
rect 9154 11342 9156 11394
rect 9100 11340 9156 11342
rect 10780 12684 10836 12740
rect 11900 13244 11956 13300
rect 11564 12684 11620 12740
rect 12964 13356 13020 13412
rect 12124 12684 12180 12740
rect 12516 12738 12572 12740
rect 12516 12686 12518 12738
rect 12518 12686 12570 12738
rect 12570 12686 12572 12738
rect 12516 12684 12572 12686
rect 10108 11788 10164 11844
rect 11564 12066 11620 12068
rect 11564 12014 11566 12066
rect 11566 12014 11618 12066
rect 11618 12014 11620 12066
rect 11564 12012 11620 12014
rect 10780 11788 10836 11844
rect 10892 11228 10948 11284
rect 13356 12684 13412 12740
rect 14924 15148 14980 15204
rect 16492 16716 16548 16772
rect 16268 16268 16324 16324
rect 15820 16098 15876 16100
rect 15820 16046 15822 16098
rect 15822 16046 15874 16098
rect 15874 16046 15876 16098
rect 15820 16044 15876 16046
rect 17052 16268 17108 16324
rect 16604 16044 16660 16100
rect 14028 14530 14084 14532
rect 14028 14478 14030 14530
rect 14030 14478 14082 14530
rect 14082 14478 14084 14530
rect 14028 14476 14084 14478
rect 13692 12908 13748 12964
rect 13804 14028 13860 14084
rect 14364 14028 14420 14084
rect 14476 14476 14532 14532
rect 14252 13746 14308 13748
rect 14252 13694 14254 13746
rect 14254 13694 14306 13746
rect 14306 13694 14308 13746
rect 14252 13692 14308 13694
rect 14476 13692 14532 13748
rect 17388 16044 17444 16100
rect 17276 15932 17332 15988
rect 17612 18508 17668 18564
rect 17948 17666 18004 17668
rect 17948 17614 17950 17666
rect 17950 17614 18002 17666
rect 18002 17614 18004 17666
rect 17948 17612 18004 17614
rect 19068 19852 19124 19908
rect 19180 19740 19236 19796
rect 19068 19404 19124 19460
rect 18172 17612 18228 17668
rect 19740 19964 19796 20020
rect 20188 20076 20244 20132
rect 19292 19516 19348 19572
rect 19628 19628 19684 19684
rect 19516 19404 19572 19460
rect 19292 19292 19348 19348
rect 19180 18732 19236 18788
rect 18732 18450 18788 18452
rect 18732 18398 18734 18450
rect 18734 18398 18786 18450
rect 18786 18398 18788 18450
rect 18732 18396 18788 18398
rect 17948 17388 18004 17444
rect 18060 16940 18116 16996
rect 17612 16268 17668 16324
rect 15484 15036 15540 15092
rect 16212 15426 16268 15428
rect 16212 15374 16214 15426
rect 16214 15374 16266 15426
rect 16266 15374 16268 15426
rect 16212 15372 16268 15374
rect 16212 15148 16268 15204
rect 17388 15260 17444 15316
rect 16604 15148 16660 15204
rect 14924 14418 14980 14420
rect 14924 14366 14926 14418
rect 14926 14366 14978 14418
rect 14978 14366 14980 14418
rect 14924 14364 14980 14366
rect 15092 14364 15148 14420
rect 14700 13916 14756 13972
rect 16044 14642 16100 14644
rect 16044 14590 16046 14642
rect 16046 14590 16098 14642
rect 16098 14590 16100 14642
rect 16044 14588 16100 14590
rect 15372 13746 15428 13748
rect 15372 13694 15374 13746
rect 15374 13694 15426 13746
rect 15426 13694 15428 13746
rect 15372 13692 15428 13694
rect 14924 13580 14980 13636
rect 14812 13132 14868 13188
rect 13636 12236 13692 12292
rect 13804 12684 13860 12740
rect 8652 9660 8708 9716
rect 7756 8204 7812 8260
rect 8204 8258 8260 8260
rect 8204 8206 8206 8258
rect 8206 8206 8258 8258
rect 8258 8206 8260 8258
rect 8204 8204 8260 8206
rect 7532 7644 7588 7700
rect 8428 8876 8484 8932
rect 12796 10668 12852 10724
rect 13356 10892 13412 10948
rect 12124 9996 12180 10052
rect 8988 9660 9044 9716
rect 9772 8316 9828 8372
rect 9100 8258 9156 8260
rect 9100 8206 9102 8258
rect 9102 8206 9154 8258
rect 9154 8206 9156 8258
rect 9100 8204 9156 8206
rect 11452 9042 11508 9044
rect 11452 8990 11454 9042
rect 11454 8990 11506 9042
rect 11506 8990 11508 9042
rect 11452 8988 11508 8990
rect 13244 10610 13300 10612
rect 13244 10558 13246 10610
rect 13246 10558 13298 10610
rect 13298 10558 13300 10610
rect 13244 10556 13300 10558
rect 13916 12236 13972 12292
rect 14140 11340 14196 11396
rect 14476 12572 14532 12628
rect 14028 11116 14084 11172
rect 14364 10892 14420 10948
rect 13962 10668 14018 10724
rect 14364 10556 14420 10612
rect 13804 10332 13860 10388
rect 14588 12066 14644 12068
rect 14588 12014 14590 12066
rect 14590 12014 14642 12066
rect 14642 12014 14644 12066
rect 14588 12012 14644 12014
rect 15148 13468 15204 13524
rect 15764 13746 15820 13748
rect 15764 13694 15766 13746
rect 15766 13694 15818 13746
rect 15818 13694 15820 13746
rect 15764 13692 15820 13694
rect 15596 13634 15652 13636
rect 15596 13582 15598 13634
rect 15598 13582 15650 13634
rect 15650 13582 15652 13634
rect 15596 13580 15652 13582
rect 16156 13468 16212 13524
rect 14812 11361 14868 11396
rect 14812 11340 14814 11361
rect 14814 11340 14866 11361
rect 14866 11340 14868 11361
rect 15122 11361 15178 11396
rect 15122 11340 15124 11361
rect 15124 11340 15176 11361
rect 15176 11340 15178 11361
rect 15260 11282 15316 11284
rect 15260 11230 15262 11282
rect 15262 11230 15314 11282
rect 15314 11230 15316 11282
rect 15260 11228 15316 11230
rect 15372 10780 15428 10836
rect 15484 13020 15540 13076
rect 16380 13692 16436 13748
rect 14588 10332 14644 10388
rect 13020 9996 13076 10052
rect 13524 10050 13580 10052
rect 13524 9998 13526 10050
rect 13526 9998 13578 10050
rect 13578 9998 13580 10050
rect 13524 9996 13580 9998
rect 11844 9436 11900 9492
rect 11676 8988 11732 9044
rect 13468 9436 13524 9492
rect 12908 9212 12964 9268
rect 13356 9324 13412 9380
rect 12572 8764 12628 8820
rect 11004 8370 11060 8372
rect 11004 8318 11006 8370
rect 11006 8318 11058 8370
rect 11058 8318 11060 8370
rect 11004 8316 11060 8318
rect 9884 8204 9940 8260
rect 10892 8204 10948 8260
rect 8316 7532 8372 7588
rect 7084 6690 7140 6692
rect 7084 6638 7086 6690
rect 7086 6638 7138 6690
rect 7138 6638 7140 6690
rect 7084 6636 7140 6638
rect 5628 6412 5684 6468
rect 7644 7474 7700 7476
rect 7644 7422 7646 7474
rect 7646 7422 7698 7474
rect 7698 7422 7700 7474
rect 7644 7420 7700 7422
rect 7868 6076 7924 6132
rect 8988 6748 9044 6804
rect 8148 6636 8204 6692
rect 7980 5740 8036 5796
rect 8540 5794 8596 5796
rect 8540 5742 8542 5794
rect 8542 5742 8594 5794
rect 8594 5742 8596 5794
rect 8540 5740 8596 5742
rect 9548 7532 9604 7588
rect 9660 7420 9716 7476
rect 9660 6748 9716 6804
rect 12180 8370 12236 8372
rect 12180 8318 12182 8370
rect 12182 8318 12234 8370
rect 12234 8318 12236 8370
rect 12180 8316 12236 8318
rect 12516 8258 12572 8260
rect 12516 8206 12518 8258
rect 12518 8206 12570 8258
rect 12570 8206 12572 8258
rect 12516 8204 12572 8206
rect 12068 8092 12124 8148
rect 14476 9324 14532 9380
rect 13804 8764 13860 8820
rect 13580 8258 13636 8260
rect 13580 8206 13582 8258
rect 13582 8206 13634 8258
rect 13634 8206 13636 8258
rect 13580 8204 13636 8206
rect 13804 8092 13860 8148
rect 14252 8092 14308 8148
rect 12796 7644 12852 7700
rect 13860 7644 13916 7700
rect 13468 7532 13524 7588
rect 11116 7474 11172 7476
rect 11116 7422 11118 7474
rect 11118 7422 11170 7474
rect 11170 7422 11172 7474
rect 11116 7420 11172 7422
rect 12684 7308 12740 7364
rect 12796 7420 12852 7476
rect 9660 6130 9716 6132
rect 9660 6078 9662 6130
rect 9662 6078 9714 6130
rect 9714 6078 9716 6130
rect 9660 6076 9716 6078
rect 10108 6690 10164 6692
rect 10108 6638 10110 6690
rect 10110 6638 10162 6690
rect 10162 6638 10164 6690
rect 10108 6636 10164 6638
rect 10388 6636 10444 6692
rect 10388 6130 10444 6132
rect 10388 6078 10390 6130
rect 10390 6078 10442 6130
rect 10442 6078 10444 6130
rect 10388 6076 10444 6078
rect 12404 6636 12460 6692
rect 10892 5964 10948 6020
rect 11900 6076 11956 6132
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 12068 6130 12124 6132
rect 12068 6078 12070 6130
rect 12070 6078 12122 6130
rect 12122 6078 12124 6130
rect 12068 6076 12124 6078
rect 12348 6018 12404 6020
rect 12348 5966 12350 6018
rect 12350 5966 12402 6018
rect 12402 5966 12404 6018
rect 12348 5964 12404 5966
rect 12796 5964 12852 6020
rect 13132 6636 13188 6692
rect 13580 7532 13636 7588
rect 13692 7474 13748 7476
rect 13692 7422 13694 7474
rect 13694 7422 13746 7474
rect 13746 7422 13748 7474
rect 13692 7420 13748 7422
rect 14140 7420 14196 7476
rect 14028 7362 14084 7364
rect 14028 7310 14030 7362
rect 14030 7310 14082 7362
rect 14082 7310 14084 7362
rect 14028 7308 14084 7310
rect 13356 5852 13412 5908
rect 13468 6524 13524 6580
rect 13580 5852 13636 5908
rect 13804 6690 13860 6692
rect 13804 6638 13806 6690
rect 13806 6638 13858 6690
rect 13858 6638 13860 6690
rect 13804 6636 13860 6638
rect 14924 10610 14980 10612
rect 14924 10558 14926 10610
rect 14926 10558 14978 10610
rect 14978 10558 14980 10610
rect 14924 10556 14980 10558
rect 14700 9996 14756 10052
rect 15036 10444 15092 10500
rect 14756 9324 14812 9380
rect 14588 8428 14644 8484
rect 15372 10332 15428 10388
rect 15260 9548 15316 9604
rect 16156 12460 16212 12516
rect 16380 11676 16436 11732
rect 16884 13580 16940 13636
rect 16492 13356 16548 13412
rect 15596 11340 15652 11396
rect 15596 11116 15652 11172
rect 15764 10834 15820 10836
rect 15764 10782 15766 10834
rect 15766 10782 15818 10834
rect 15818 10782 15820 10834
rect 15764 10780 15820 10782
rect 15036 9266 15092 9268
rect 15036 9214 15038 9266
rect 15038 9214 15090 9266
rect 15090 9214 15092 9266
rect 15036 9212 15092 9214
rect 14924 8540 14980 8596
rect 14700 8316 14756 8372
rect 14812 7644 14868 7700
rect 16044 9548 16100 9604
rect 15932 8428 15988 8484
rect 16380 11394 16436 11396
rect 16380 11342 16382 11394
rect 16382 11342 16434 11394
rect 16434 11342 16436 11394
rect 16380 11340 16436 11342
rect 16380 10668 16436 10724
rect 17948 15932 18004 15988
rect 18396 14642 18452 14644
rect 18396 14590 18398 14642
rect 18398 14590 18450 14642
rect 18450 14590 18452 14642
rect 18396 14588 18452 14590
rect 18844 18284 18900 18340
rect 19292 17724 19348 17780
rect 18844 17666 18900 17668
rect 18844 17614 18846 17666
rect 18846 17614 18898 17666
rect 18898 17614 18900 17666
rect 18844 17612 18900 17614
rect 19012 17666 19068 17668
rect 19012 17614 19014 17666
rect 19014 17614 19066 17666
rect 19066 17614 19068 17666
rect 19012 17612 19068 17614
rect 19180 17500 19236 17556
rect 18732 16828 18788 16884
rect 19068 16882 19124 16884
rect 19068 16830 19070 16882
rect 19070 16830 19122 16882
rect 19122 16830 19124 16882
rect 19068 16828 19124 16830
rect 19180 16716 19236 16772
rect 19068 16604 19124 16660
rect 18956 15372 19012 15428
rect 18620 15260 18676 15316
rect 17612 13746 17668 13748
rect 17612 13694 17614 13746
rect 17614 13694 17666 13746
rect 17666 13694 17668 13746
rect 17612 13692 17668 13694
rect 17500 13020 17556 13076
rect 17500 12178 17556 12180
rect 17500 12126 17502 12178
rect 17502 12126 17554 12178
rect 17554 12126 17556 12178
rect 17500 12124 17556 12126
rect 16716 11676 16772 11732
rect 17164 11506 17220 11508
rect 17164 11454 17166 11506
rect 17166 11454 17218 11506
rect 17218 11454 17220 11506
rect 17164 11452 17220 11454
rect 17052 11379 17108 11396
rect 17052 11340 17054 11379
rect 17054 11340 17106 11379
rect 17106 11340 17108 11379
rect 17948 13692 18004 13748
rect 18116 13746 18172 13748
rect 18116 13694 18118 13746
rect 18118 13694 18170 13746
rect 18170 13694 18172 13746
rect 18116 13692 18172 13694
rect 18620 13746 18676 13748
rect 18620 13694 18622 13746
rect 18622 13694 18674 13746
rect 18674 13694 18676 13746
rect 18620 13692 18676 13694
rect 18508 13580 18564 13636
rect 19180 15820 19236 15876
rect 20524 19628 20580 19684
rect 20188 19404 20244 19460
rect 20412 19516 20468 19572
rect 20188 19234 20244 19236
rect 20188 19182 20190 19234
rect 20190 19182 20242 19234
rect 20242 19182 20244 19234
rect 20188 19180 20244 19182
rect 20300 19292 20356 19348
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19628 17612 19684 17668
rect 20076 18450 20132 18452
rect 20076 18398 20078 18450
rect 20078 18398 20130 18450
rect 20130 18398 20132 18450
rect 20076 18396 20132 18398
rect 20076 17724 20132 17780
rect 20748 19852 20804 19908
rect 20412 18508 20468 18564
rect 21532 23154 21588 23156
rect 21532 23102 21534 23154
rect 21534 23102 21586 23154
rect 21586 23102 21588 23154
rect 21532 23100 21588 23102
rect 21308 22092 21364 22148
rect 21532 22594 21588 22596
rect 21532 22542 21534 22594
rect 21534 22542 21586 22594
rect 21586 22542 21588 22594
rect 21532 22540 21588 22542
rect 21532 21980 21588 22036
rect 21700 22092 21756 22148
rect 22316 24722 22372 24724
rect 22316 24670 22318 24722
rect 22318 24670 22370 24722
rect 22370 24670 22372 24722
rect 22316 24668 22372 24670
rect 22652 24946 22708 24948
rect 22652 24894 22654 24946
rect 22654 24894 22706 24946
rect 22706 24894 22708 24946
rect 22652 24892 22708 24894
rect 23884 25452 23940 25508
rect 24108 26012 24164 26068
rect 23772 24892 23828 24948
rect 22876 23938 22932 23940
rect 22876 23886 22878 23938
rect 22878 23886 22930 23938
rect 22930 23886 22932 23938
rect 22876 23884 22932 23886
rect 22876 23548 22932 23604
rect 22204 22764 22260 22820
rect 22540 22876 22596 22932
rect 22764 22764 22820 22820
rect 22652 22652 22708 22708
rect 22764 22204 22820 22260
rect 22652 22092 22708 22148
rect 21868 21756 21924 21812
rect 21420 21586 21476 21588
rect 21420 21534 21422 21586
rect 21422 21534 21474 21586
rect 21474 21534 21476 21586
rect 21420 21532 21476 21534
rect 21980 21562 21982 21588
rect 21982 21562 22034 21588
rect 22034 21562 22036 21588
rect 21980 21532 22036 21562
rect 21420 20748 21476 20804
rect 22428 20860 22484 20916
rect 21644 19852 21700 19908
rect 21028 19180 21084 19236
rect 20300 17627 20356 17668
rect 20300 17612 20302 17627
rect 20302 17612 20354 17627
rect 20354 17612 20356 17627
rect 19964 17388 20020 17444
rect 20188 17500 20244 17556
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 21532 19234 21588 19236
rect 21532 19182 21534 19234
rect 21534 19182 21586 19234
rect 21586 19182 21588 19234
rect 21532 19180 21588 19182
rect 21196 18396 21252 18452
rect 21420 18396 21476 18452
rect 21868 20636 21924 20692
rect 22540 20188 22596 20244
rect 22092 19628 22148 19684
rect 22540 19628 22596 19684
rect 22260 19516 22316 19572
rect 22708 19346 22764 19348
rect 22708 19294 22710 19346
rect 22710 19294 22762 19346
rect 22762 19294 22764 19346
rect 22708 19292 22764 19294
rect 22764 18956 22820 19012
rect 21868 18396 21924 18452
rect 21980 18284 22036 18340
rect 22092 18396 22148 18452
rect 21868 18060 21924 18116
rect 21196 17666 21252 17668
rect 21196 17614 21198 17666
rect 21198 17614 21250 17666
rect 21250 17614 21252 17666
rect 21196 17612 21252 17614
rect 19628 17052 19684 17108
rect 20188 17164 20244 17220
rect 19404 15484 19460 15540
rect 19516 16492 19572 16548
rect 20300 16268 20356 16324
rect 20636 16492 20692 16548
rect 19740 16070 19796 16100
rect 19740 16044 19742 16070
rect 19742 16044 19794 16070
rect 19794 16044 19796 16070
rect 20300 15932 20356 15988
rect 19348 14476 19404 14532
rect 20468 15874 20524 15876
rect 20468 15822 20470 15874
rect 20470 15822 20522 15874
rect 20522 15822 20524 15874
rect 20468 15820 20524 15822
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19740 15484 19796 15540
rect 21364 17500 21420 17556
rect 21196 17106 21252 17108
rect 21196 17054 21198 17106
rect 21198 17054 21250 17106
rect 21250 17054 21252 17106
rect 21196 17052 21252 17054
rect 21756 17052 21812 17108
rect 20972 16716 21028 16772
rect 20972 15372 21028 15428
rect 21756 16716 21812 16772
rect 21532 15932 21588 15988
rect 21364 15596 21420 15652
rect 19628 14476 19684 14532
rect 20636 14924 20692 14980
rect 21196 14924 21252 14980
rect 19348 14306 19404 14308
rect 19348 14254 19350 14306
rect 19350 14254 19402 14306
rect 19402 14254 19404 14306
rect 19348 14252 19404 14254
rect 19404 14028 19460 14084
rect 18788 13074 18844 13076
rect 18788 13022 18790 13074
rect 18790 13022 18842 13074
rect 18842 13022 18844 13074
rect 18788 13020 18844 13022
rect 18060 12348 18116 12404
rect 17836 12124 17892 12180
rect 17612 11788 17668 11844
rect 16492 10610 16548 10612
rect 16492 10558 16494 10610
rect 16494 10558 16546 10610
rect 16546 10558 16548 10610
rect 17724 11452 17780 11508
rect 17612 11116 17668 11172
rect 16492 10556 16548 10558
rect 17500 10556 17556 10612
rect 16268 9100 16324 9156
rect 16380 9548 16436 9604
rect 16772 9154 16828 9156
rect 16772 9102 16774 9154
rect 16774 9102 16826 9154
rect 16826 9102 16828 9154
rect 16772 9100 16828 9102
rect 17668 9436 17724 9492
rect 18564 12402 18620 12404
rect 18564 12350 18566 12402
rect 18566 12350 18618 12402
rect 18618 12350 18620 12402
rect 18564 12348 18620 12350
rect 18172 12012 18228 12068
rect 19836 14138 19892 14140
rect 19516 13746 19572 13748
rect 19516 13694 19518 13746
rect 19518 13694 19570 13746
rect 19570 13694 19572 13746
rect 19516 13692 19572 13694
rect 19628 14028 19684 14084
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 18956 12348 19012 12404
rect 19852 13804 19908 13860
rect 20412 14364 20468 14420
rect 20300 13692 20356 13748
rect 20972 14140 21028 14196
rect 20860 13746 20916 13748
rect 20860 13694 20862 13746
rect 20862 13694 20914 13746
rect 20914 13694 20916 13746
rect 20860 13692 20916 13694
rect 21420 14140 21476 14196
rect 20972 13356 21028 13412
rect 21868 16828 21924 16884
rect 22092 17500 22148 17556
rect 22428 18508 22484 18564
rect 22316 18284 22372 18340
rect 22652 18060 22708 18116
rect 22764 17948 22820 18004
rect 22764 17724 22820 17780
rect 22316 16828 22372 16884
rect 22428 17276 22484 17332
rect 22540 16716 22596 16772
rect 22036 16210 22092 16212
rect 22036 16158 22038 16210
rect 22038 16158 22090 16210
rect 22090 16158 22092 16210
rect 22036 16156 22092 16158
rect 21868 15596 21924 15652
rect 22428 16098 22484 16100
rect 22428 16046 22430 16098
rect 22430 16046 22482 16098
rect 22482 16046 22484 16098
rect 22428 16044 22484 16046
rect 24108 24444 24164 24500
rect 24892 29932 24948 29988
rect 25228 32620 25284 32676
rect 25452 33318 25508 33348
rect 25452 33292 25454 33318
rect 25454 33292 25506 33318
rect 25506 33292 25508 33318
rect 25116 31948 25172 32004
rect 25284 31554 25340 31556
rect 25284 31502 25286 31554
rect 25286 31502 25338 31554
rect 25338 31502 25340 31554
rect 25284 31500 25340 31502
rect 25116 31276 25172 31332
rect 26124 36876 26180 36932
rect 26572 37660 26628 37716
rect 26460 37100 26516 37156
rect 26348 36876 26404 36932
rect 25788 36540 25844 36596
rect 26124 36428 26180 36484
rect 25844 35532 25900 35588
rect 25676 35196 25732 35252
rect 26124 35698 26180 35700
rect 26124 35646 26126 35698
rect 26126 35646 26178 35698
rect 26178 35646 26180 35698
rect 26124 35644 26180 35646
rect 26236 35868 26292 35924
rect 27112 39116 27168 39172
rect 27804 41804 27860 41860
rect 27636 41468 27692 41524
rect 27448 40684 27504 40740
rect 27524 40402 27580 40404
rect 27524 40350 27526 40402
rect 27526 40350 27578 40402
rect 27578 40350 27580 40402
rect 27524 40348 27580 40350
rect 28140 40908 28196 40964
rect 28140 40684 28196 40740
rect 30268 46060 30324 46116
rect 30268 45890 30324 45892
rect 30268 45838 30270 45890
rect 30270 45838 30322 45890
rect 30322 45838 30324 45890
rect 30268 45836 30324 45838
rect 29260 43484 29316 43540
rect 29652 43426 29708 43428
rect 29652 43374 29654 43426
rect 29654 43374 29706 43426
rect 29706 43374 29708 43426
rect 29652 43372 29708 43374
rect 28476 43260 28532 43316
rect 28476 42978 28532 42980
rect 28476 42926 28478 42978
rect 28478 42926 28530 42978
rect 28530 42926 28532 42978
rect 28476 42924 28532 42926
rect 29932 43596 29988 43652
rect 30156 43538 30212 43540
rect 30156 43486 30158 43538
rect 30158 43486 30210 43538
rect 30210 43486 30212 43538
rect 30156 43484 30212 43486
rect 30940 45890 30996 45892
rect 30940 45838 30942 45890
rect 30942 45838 30994 45890
rect 30994 45838 30996 45890
rect 30940 45836 30996 45838
rect 31444 45724 31500 45780
rect 33180 46114 33236 46116
rect 33180 46062 33182 46114
rect 33182 46062 33234 46114
rect 33234 46062 33236 46114
rect 33180 46060 33236 46062
rect 33404 46060 33460 46116
rect 32172 45862 32228 45892
rect 32172 45836 32174 45862
rect 32174 45836 32226 45862
rect 32226 45836 32228 45862
rect 33628 45724 33684 45780
rect 30492 44492 30548 44548
rect 30492 43708 30548 43764
rect 30380 43260 30436 43316
rect 29036 42588 29092 42644
rect 30492 43148 30548 43204
rect 29372 42530 29428 42532
rect 29372 42478 29374 42530
rect 29374 42478 29426 42530
rect 29426 42478 29428 42530
rect 29372 42476 29428 42478
rect 28588 42252 28644 42308
rect 28700 42140 28756 42196
rect 28812 41916 28868 41972
rect 27468 40012 27524 40068
rect 27356 39618 27412 39620
rect 27356 39566 27358 39618
rect 27358 39566 27410 39618
rect 27410 39566 27412 39618
rect 27356 39564 27412 39566
rect 27244 38780 27300 38836
rect 27132 38668 27188 38724
rect 28680 40684 28736 40740
rect 28812 40572 28868 40628
rect 28924 40514 28980 40516
rect 28924 40462 28926 40514
rect 28926 40462 28978 40514
rect 28978 40462 28980 40514
rect 28924 40460 28980 40462
rect 29036 40348 29092 40404
rect 29484 41970 29540 41972
rect 29484 41918 29486 41970
rect 29486 41918 29538 41970
rect 29538 41918 29540 41970
rect 29484 41916 29540 41918
rect 29484 41692 29540 41748
rect 29372 40962 29428 40964
rect 29372 40910 29374 40962
rect 29374 40910 29426 40962
rect 29426 40910 29428 40962
rect 29372 40908 29428 40910
rect 29148 40012 29204 40068
rect 28140 39452 28196 39508
rect 29036 39618 29092 39620
rect 29036 39566 29038 39618
rect 29038 39566 29090 39618
rect 29090 39566 29092 39618
rect 29036 39564 29092 39566
rect 29204 39452 29260 39508
rect 28252 39340 28308 39396
rect 28904 39340 28960 39396
rect 29372 39340 29428 39396
rect 29148 38834 29204 38836
rect 29148 38782 29150 38834
rect 29150 38782 29202 38834
rect 29202 38782 29204 38834
rect 29148 38780 29204 38782
rect 28700 38668 28756 38724
rect 29932 42754 29988 42756
rect 29932 42702 29934 42754
rect 29934 42702 29986 42754
rect 29986 42702 29988 42754
rect 29932 42700 29988 42702
rect 30156 42140 30212 42196
rect 30492 41746 30548 41748
rect 30492 41694 30494 41746
rect 30494 41694 30546 41746
rect 30546 41694 30548 41746
rect 30492 41692 30548 41694
rect 30735 44156 30791 44212
rect 30716 43596 30772 43652
rect 30716 43036 30772 43092
rect 31276 43538 31332 43540
rect 30828 42924 30884 42980
rect 31276 43486 31278 43538
rect 31278 43486 31330 43538
rect 31330 43486 31332 43538
rect 31276 43484 31332 43486
rect 31612 43484 31668 43540
rect 30808 42252 30864 42308
rect 32732 45052 32788 45108
rect 31836 44156 31892 44212
rect 31982 43523 31984 43540
rect 31984 43523 32036 43540
rect 32036 43523 32038 43540
rect 31982 43484 32038 43523
rect 31948 43036 32004 43092
rect 32396 43314 32452 43316
rect 32396 43262 32398 43314
rect 32398 43262 32450 43314
rect 32450 43262 32452 43314
rect 32396 43260 32452 43262
rect 32452 42978 32508 42980
rect 32452 42926 32454 42978
rect 32454 42926 32506 42978
rect 32506 42926 32508 42978
rect 32452 42924 32508 42926
rect 32172 42700 32228 42756
rect 31724 42588 31780 42644
rect 29708 41468 29764 41524
rect 29596 41132 29652 41188
rect 32284 42252 32340 42308
rect 32620 42700 32676 42756
rect 30696 41186 30752 41188
rect 30696 41134 30698 41186
rect 30698 41134 30750 41186
rect 30750 41134 30752 41186
rect 30696 41132 30752 41134
rect 29932 40460 29988 40516
rect 30156 40460 30212 40516
rect 29764 40402 29820 40404
rect 29764 40350 29766 40402
rect 29766 40350 29818 40402
rect 29818 40350 29820 40402
rect 29764 40348 29820 40350
rect 29708 38780 29764 38836
rect 29932 39228 29988 39284
rect 30660 40460 30716 40516
rect 30940 41186 30996 41188
rect 30940 41134 30942 41186
rect 30942 41134 30994 41186
rect 30994 41134 30996 41186
rect 30940 41132 30996 41134
rect 31052 40908 31108 40964
rect 30492 40380 30494 40404
rect 30494 40380 30546 40404
rect 30546 40380 30548 40404
rect 30492 40348 30548 40380
rect 30828 39618 30884 39620
rect 30828 39566 30830 39618
rect 30830 39566 30882 39618
rect 30882 39566 30884 39618
rect 30828 39564 30884 39566
rect 30584 39228 30640 39284
rect 30380 38892 30436 38948
rect 30716 39004 30772 39060
rect 30492 38834 30548 38836
rect 30492 38782 30494 38834
rect 30494 38782 30546 38834
rect 30546 38782 30548 38834
rect 30492 38780 30548 38782
rect 29932 38668 29988 38724
rect 30380 38668 30436 38724
rect 28812 38556 28868 38612
rect 28028 38020 28084 38052
rect 27076 37938 27132 37940
rect 27076 37886 27078 37938
rect 27078 37886 27130 37938
rect 27130 37886 27132 37938
rect 27076 37884 27132 37886
rect 28028 37996 28030 38020
rect 28030 37996 28082 38020
rect 28082 37996 28084 38020
rect 28476 37884 28532 37940
rect 27244 37436 27300 37492
rect 28364 37378 28420 37380
rect 28364 37326 28366 37378
rect 28366 37326 28418 37378
rect 28418 37326 28420 37378
rect 28364 37324 28420 37326
rect 27916 37100 27972 37156
rect 26888 36764 26944 36820
rect 27020 36652 27076 36708
rect 26236 35308 26292 35364
rect 27132 35674 27134 35700
rect 27134 35674 27186 35700
rect 27186 35674 27188 35700
rect 27132 35644 27188 35674
rect 25676 34636 25732 34692
rect 25676 33964 25732 34020
rect 26236 34802 26292 34804
rect 26236 34750 26238 34802
rect 26238 34750 26290 34802
rect 26290 34750 26292 34802
rect 26236 34748 26292 34750
rect 26012 33740 26068 33796
rect 26908 35196 26964 35252
rect 26796 34636 26852 34692
rect 26908 33852 26964 33908
rect 28120 36764 28176 36820
rect 27916 36540 27972 36596
rect 27804 35756 27860 35812
rect 30380 38444 30436 38500
rect 30024 38050 30080 38052
rect 30024 37998 30026 38050
rect 30026 37998 30078 38050
rect 30078 37998 30080 38050
rect 30024 37996 30080 37998
rect 30268 38050 30324 38052
rect 30268 37998 30270 38050
rect 30270 37998 30322 38050
rect 30322 37998 30324 38050
rect 30268 37996 30324 37998
rect 29148 37324 29204 37380
rect 29764 37660 29820 37716
rect 27916 35868 27972 35924
rect 29764 37154 29820 37156
rect 29764 37102 29766 37154
rect 29766 37102 29818 37154
rect 29818 37102 29820 37154
rect 29764 37100 29820 37102
rect 27692 35420 27748 35476
rect 27580 35308 27636 35364
rect 28792 35420 28848 35476
rect 30380 37436 30436 37492
rect 30212 37266 30268 37268
rect 30212 37214 30214 37266
rect 30214 37214 30266 37266
rect 30266 37214 30268 37266
rect 30212 37212 30268 37214
rect 32264 41186 32320 41188
rect 32264 41134 32266 41186
rect 32266 41134 32318 41186
rect 32318 41134 32320 41186
rect 32264 41132 32320 41134
rect 32284 40908 32340 40964
rect 31388 40460 31444 40516
rect 31276 40012 31332 40068
rect 31500 40572 31556 40628
rect 31780 40402 31836 40404
rect 31780 40350 31782 40402
rect 31782 40350 31834 40402
rect 31834 40350 31836 40402
rect 31780 40348 31836 40350
rect 33068 45106 33124 45108
rect 33068 45054 33070 45106
rect 33070 45054 33122 45106
rect 33122 45054 33124 45106
rect 33068 45052 33124 45054
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 35028 45890 35084 45892
rect 35028 45838 35030 45890
rect 35030 45838 35082 45890
rect 35082 45838 35084 45890
rect 35028 45836 35084 45838
rect 33068 43538 33124 43540
rect 33068 43486 33070 43538
rect 33070 43486 33122 43538
rect 33122 43486 33124 43538
rect 33068 43484 33124 43486
rect 33068 43148 33124 43204
rect 33292 43036 33348 43092
rect 33740 43372 33796 43428
rect 34076 43426 34132 43428
rect 34076 43374 34078 43426
rect 34078 43374 34130 43426
rect 34130 43374 34132 43426
rect 34076 43372 34132 43374
rect 33852 43148 33908 43204
rect 35308 45612 35364 45668
rect 34972 43596 35028 43652
rect 35084 45388 35140 45444
rect 34412 43260 34468 43316
rect 34188 43036 34244 43092
rect 33740 42924 33796 42980
rect 34748 42924 34804 42980
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 35980 45388 36036 45444
rect 36428 45500 36484 45556
rect 36988 46114 37044 46116
rect 36988 46062 36990 46114
rect 36990 46062 37042 46114
rect 37042 46062 37044 46114
rect 36988 46060 37044 46062
rect 38108 46060 38164 46116
rect 38668 45890 38724 45892
rect 38668 45838 38670 45890
rect 38670 45838 38722 45890
rect 38722 45838 38724 45890
rect 38668 45836 38724 45838
rect 36540 45276 36596 45332
rect 36652 45612 36708 45668
rect 37660 45388 37716 45444
rect 36652 44940 36708 44996
rect 37212 44882 37268 44884
rect 37212 44830 37214 44882
rect 37214 44830 37266 44882
rect 37266 44830 37268 44882
rect 37212 44828 37268 44830
rect 35756 44492 35812 44548
rect 35551 44322 35607 44324
rect 35551 44270 35553 44322
rect 35553 44270 35605 44322
rect 35605 44270 35607 44322
rect 35551 44268 35607 44270
rect 35308 44210 35364 44212
rect 35308 44158 35310 44210
rect 35310 44158 35362 44210
rect 35362 44158 35364 44210
rect 35308 44156 35364 44158
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 35420 42866 35476 42868
rect 35420 42814 35422 42866
rect 35422 42814 35474 42866
rect 35474 42814 35476 42866
rect 35420 42812 35476 42814
rect 33740 42364 33796 42420
rect 32508 39788 32564 39844
rect 32620 39676 32676 39732
rect 31612 39618 31668 39620
rect 31612 39566 31614 39618
rect 31614 39566 31666 39618
rect 31666 39566 31668 39618
rect 32396 39618 32452 39620
rect 31612 39564 31668 39566
rect 32396 39566 32398 39618
rect 32398 39566 32450 39618
rect 32450 39566 32452 39618
rect 32396 39564 32452 39566
rect 31724 39452 31780 39508
rect 32732 39452 32788 39508
rect 31220 39004 31276 39060
rect 31052 38444 31108 38500
rect 31948 38668 32004 38724
rect 32060 38556 32116 38612
rect 30716 38050 30772 38052
rect 30716 37998 30718 38050
rect 30718 37998 30770 38050
rect 30770 37998 30772 38050
rect 30716 37996 30772 37998
rect 31592 37884 31648 37940
rect 30660 37490 30716 37492
rect 30660 37438 30662 37490
rect 30662 37438 30714 37490
rect 30714 37438 30716 37490
rect 30660 37436 30716 37438
rect 30604 37212 30660 37268
rect 30136 36540 30192 36596
rect 30380 36706 30436 36708
rect 30380 36654 30382 36706
rect 30382 36654 30434 36706
rect 30434 36654 30436 36706
rect 30380 36652 30436 36654
rect 29148 36092 29204 36148
rect 28924 35532 28980 35588
rect 28364 35196 28420 35252
rect 28028 34884 28084 34916
rect 28028 34860 28030 34884
rect 28030 34860 28082 34884
rect 28082 34860 28084 34884
rect 27244 34412 27300 34468
rect 26852 33628 26908 33684
rect 26292 32508 26348 32564
rect 27916 33740 27972 33796
rect 27356 33628 27412 33684
rect 28140 33740 28196 33796
rect 28476 35138 28532 35140
rect 28476 35086 28478 35138
rect 28478 35086 28530 35138
rect 28530 35086 28532 35138
rect 28476 35084 28532 35086
rect 28364 34242 28420 34244
rect 28364 34190 28366 34242
rect 28366 34190 28418 34242
rect 28418 34190 28420 34242
rect 28364 34188 28420 34190
rect 28476 33628 28532 33684
rect 27916 32620 27972 32676
rect 25844 31724 25900 31780
rect 25844 31388 25900 31444
rect 26572 31948 26628 32004
rect 25228 31052 25284 31108
rect 25676 30994 25732 30996
rect 25676 30942 25678 30994
rect 25678 30942 25730 30994
rect 25730 30942 25732 30994
rect 25676 30940 25732 30942
rect 25788 30604 25844 30660
rect 25452 30156 25508 30212
rect 25228 30098 25284 30100
rect 25228 30046 25230 30098
rect 25230 30046 25282 30098
rect 25282 30046 25284 30098
rect 25228 30044 25284 30046
rect 25340 29538 25396 29540
rect 25340 29486 25342 29538
rect 25342 29486 25394 29538
rect 25394 29486 25396 29538
rect 25340 29484 25396 29486
rect 25228 29148 25284 29204
rect 25676 30044 25732 30100
rect 26124 29820 26180 29876
rect 26012 29596 26068 29652
rect 25564 29426 25620 29428
rect 25564 29374 25566 29426
rect 25566 29374 25618 29426
rect 25618 29374 25620 29426
rect 25564 29372 25620 29374
rect 26012 29372 26068 29428
rect 24892 27132 24948 27188
rect 24892 26908 24948 26964
rect 24668 26572 24724 26628
rect 24556 26124 24612 26180
rect 24220 24220 24276 24276
rect 24836 25282 24892 25284
rect 24836 25230 24838 25282
rect 24838 25230 24890 25282
rect 24890 25230 24892 25282
rect 24836 25228 24892 25230
rect 24724 24722 24780 24724
rect 24724 24670 24726 24722
rect 24726 24670 24778 24722
rect 24778 24670 24780 24722
rect 24724 24668 24780 24670
rect 24444 24556 24500 24612
rect 24892 24444 24948 24500
rect 23660 24108 23716 24164
rect 23548 23548 23604 23604
rect 24780 23436 24836 23492
rect 23884 23212 23940 23268
rect 23626 23139 23628 23156
rect 23628 23139 23680 23156
rect 23680 23139 23682 23156
rect 23626 23100 23682 23139
rect 23772 23154 23828 23156
rect 23772 23102 23774 23154
rect 23774 23102 23826 23154
rect 23826 23102 23828 23154
rect 23772 23100 23828 23102
rect 23212 22652 23268 22708
rect 23100 22370 23156 22372
rect 23100 22318 23102 22370
rect 23102 22318 23154 22370
rect 23154 22318 23156 22370
rect 23100 22316 23156 22318
rect 22988 22204 23044 22260
rect 23044 21868 23100 21924
rect 23100 20860 23156 20916
rect 23548 22764 23604 22820
rect 25116 28140 25172 28196
rect 25452 28252 25508 28308
rect 25564 28588 25620 28644
rect 25676 27132 25732 27188
rect 25788 27074 25844 27076
rect 25788 27022 25790 27074
rect 25790 27022 25842 27074
rect 25842 27022 25844 27074
rect 25788 27020 25844 27022
rect 25340 26572 25396 26628
rect 25228 26273 25230 26292
rect 25230 26273 25282 26292
rect 25282 26273 25284 26292
rect 25564 26348 25620 26404
rect 25228 26236 25284 26273
rect 25116 26012 25172 26068
rect 25116 25228 25172 25284
rect 25788 25116 25844 25172
rect 25676 25004 25732 25060
rect 25284 24556 25340 24612
rect 25788 24892 25844 24948
rect 26012 27821 26014 27860
rect 26014 27821 26066 27860
rect 26066 27821 26068 27860
rect 26012 27804 26068 27821
rect 27020 31836 27076 31892
rect 27244 31778 27300 31780
rect 27244 31726 27246 31778
rect 27246 31726 27298 31778
rect 27298 31726 27300 31778
rect 27244 31724 27300 31726
rect 27916 31724 27972 31780
rect 28120 31778 28176 31780
rect 28120 31726 28122 31778
rect 28122 31726 28174 31778
rect 28174 31726 28176 31778
rect 28120 31724 28176 31726
rect 28364 31948 28420 32004
rect 28532 31836 28588 31892
rect 26740 31218 26796 31220
rect 26740 31166 26742 31218
rect 26742 31166 26794 31218
rect 26794 31166 26796 31218
rect 26740 31164 26796 31166
rect 26348 29820 26404 29876
rect 26796 30210 26852 30212
rect 26796 30158 26798 30210
rect 26798 30158 26850 30210
rect 26850 30158 26852 30210
rect 26796 30156 26852 30158
rect 26460 29260 26516 29316
rect 28364 31778 28420 31780
rect 28364 31726 28366 31778
rect 28366 31726 28418 31778
rect 28418 31726 28420 31778
rect 28364 31724 28420 31726
rect 27804 31388 27860 31444
rect 28476 31612 28532 31668
rect 28812 35196 28868 35252
rect 29148 35196 29204 35252
rect 29820 35980 29876 36036
rect 29988 35980 30044 36036
rect 29988 35586 30044 35588
rect 29988 35534 29990 35586
rect 29990 35534 30042 35586
rect 30042 35534 30044 35586
rect 29988 35532 30044 35534
rect 30024 34914 30080 34916
rect 30024 34862 30026 34914
rect 30026 34862 30078 34914
rect 30078 34862 30080 34914
rect 30024 34860 30080 34862
rect 29148 34188 29204 34244
rect 28980 33404 29036 33460
rect 28812 31388 28868 31444
rect 28700 31164 28756 31220
rect 29764 34130 29820 34132
rect 29764 34078 29766 34130
rect 29766 34078 29818 34130
rect 29818 34078 29820 34130
rect 29764 34076 29820 34078
rect 30268 35756 30324 35812
rect 32732 38780 32788 38836
rect 32172 38050 32228 38052
rect 32172 37998 32174 38050
rect 32174 37998 32226 38050
rect 32226 37998 32228 38050
rect 32172 37996 32228 37998
rect 33852 40684 33908 40740
rect 33068 39618 33124 39620
rect 33068 39566 33070 39618
rect 33070 39566 33122 39618
rect 33122 39566 33124 39618
rect 33068 39564 33124 39566
rect 33572 39618 33628 39620
rect 33572 39566 33574 39618
rect 33574 39566 33626 39618
rect 33626 39566 33628 39618
rect 33572 39564 33628 39566
rect 33292 39452 33348 39508
rect 33068 38834 33124 38836
rect 33068 38782 33070 38834
rect 33070 38782 33122 38834
rect 33122 38782 33124 38834
rect 33068 38780 33124 38782
rect 34412 42252 34468 42308
rect 36204 43596 36260 43652
rect 36428 43596 36484 43652
rect 36652 43484 36708 43540
rect 34300 42140 34356 42196
rect 34748 41692 34804 41748
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35532 41244 35588 41300
rect 35084 40572 35140 40628
rect 34860 40348 34916 40404
rect 35420 40124 35476 40180
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35980 42028 36036 42084
rect 35848 41970 35904 41972
rect 35848 41918 35850 41970
rect 35850 41918 35902 41970
rect 35902 41918 35904 41970
rect 35848 41916 35904 41918
rect 36092 41858 36148 41860
rect 36092 41806 36094 41858
rect 36094 41806 36146 41858
rect 36146 41806 36148 41858
rect 36092 41804 36148 41806
rect 36652 42028 36708 42084
rect 36204 41468 36260 41524
rect 36316 41804 36372 41860
rect 35924 41410 35980 41412
rect 35924 41358 35926 41410
rect 35926 41358 35978 41410
rect 35978 41358 35980 41410
rect 35924 41356 35980 41358
rect 36204 41186 36260 41188
rect 36204 41134 36206 41186
rect 36206 41134 36258 41186
rect 36258 41134 36260 41186
rect 36204 41132 36260 41134
rect 36876 42028 36932 42084
rect 37380 42140 37436 42196
rect 37100 42028 37156 42084
rect 36764 41356 36820 41412
rect 36988 41692 37044 41748
rect 37324 41916 37380 41972
rect 37548 41916 37604 41972
rect 37436 41580 37492 41636
rect 36988 41132 37044 41188
rect 35644 40402 35700 40404
rect 35644 40350 35646 40402
rect 35646 40350 35698 40402
rect 35698 40350 35700 40402
rect 35644 40348 35700 40350
rect 34636 39340 34692 39396
rect 33964 39004 34020 39060
rect 35084 39004 35140 39060
rect 33944 38668 34000 38724
rect 34188 38220 34244 38276
rect 34804 38834 34860 38836
rect 34804 38782 34806 38834
rect 34806 38782 34858 38834
rect 34858 38782 34860 38834
rect 34804 38780 34860 38782
rect 36708 40460 36764 40516
rect 36204 40236 36260 40292
rect 36204 39116 36260 39172
rect 35868 39004 35924 39060
rect 36540 40348 36596 40404
rect 37212 41158 37268 41188
rect 37212 41132 37214 41158
rect 37214 41132 37266 41158
rect 37266 41132 37268 41158
rect 39172 45778 39228 45780
rect 39172 45726 39174 45778
rect 39174 45726 39226 45778
rect 39226 45726 39228 45778
rect 39172 45724 39228 45726
rect 38892 45388 38948 45444
rect 37996 45276 38052 45332
rect 39004 44716 39060 44772
rect 38799 44044 38855 44100
rect 38052 43596 38108 43652
rect 37884 43538 37940 43540
rect 37884 43486 37886 43538
rect 37886 43486 37938 43538
rect 37938 43486 37940 43538
rect 37884 43484 37940 43486
rect 38556 43538 38612 43540
rect 38556 43486 38558 43538
rect 38558 43486 38610 43538
rect 38610 43486 38612 43538
rect 38556 43484 38612 43486
rect 38108 42252 38164 42308
rect 37996 42082 38052 42084
rect 37996 42030 37998 42082
rect 37998 42030 38050 42082
rect 38050 42030 38052 42082
rect 37996 42028 38052 42030
rect 38556 42028 38612 42084
rect 37828 41580 37884 41636
rect 38220 41804 38276 41860
rect 38444 41692 38500 41748
rect 37548 41132 37604 41188
rect 38108 41186 38164 41188
rect 38108 41134 38110 41186
rect 38110 41134 38162 41186
rect 38162 41134 38164 41186
rect 38108 41132 38164 41134
rect 37436 41020 37492 41076
rect 37660 40460 37716 40516
rect 36652 40124 36708 40180
rect 37156 39676 37212 39732
rect 37828 40402 37884 40404
rect 37828 40350 37830 40402
rect 37830 40350 37882 40402
rect 37882 40350 37884 40402
rect 37828 40348 37884 40350
rect 37884 40012 37940 40068
rect 36652 39116 36708 39172
rect 37324 39618 37380 39620
rect 37324 39566 37326 39618
rect 37326 39566 37378 39618
rect 37378 39566 37380 39618
rect 37324 39564 37380 39566
rect 36428 39004 36484 39060
rect 36988 38892 37044 38948
rect 36540 38834 36596 38836
rect 36540 38782 36542 38834
rect 36542 38782 36594 38834
rect 36594 38782 36596 38834
rect 36540 38780 36596 38782
rect 34860 38108 34916 38164
rect 32172 37266 32228 37268
rect 32172 37214 32174 37266
rect 32174 37214 32226 37266
rect 32226 37214 32228 37266
rect 32172 37212 32228 37214
rect 30828 36652 30884 36708
rect 31500 36652 31556 36708
rect 32004 36540 32060 36596
rect 31108 35980 31164 36036
rect 30716 35756 30772 35812
rect 31836 36428 31892 36484
rect 31724 35420 31780 35476
rect 30492 35084 30548 35140
rect 31592 35308 31648 35364
rect 31556 34802 31612 34804
rect 31556 34750 31558 34802
rect 31558 34750 31610 34802
rect 31610 34750 31612 34802
rect 31556 34748 31612 34750
rect 31108 34690 31164 34692
rect 31108 34638 31110 34690
rect 31110 34638 31162 34690
rect 31162 34638 31164 34690
rect 31108 34636 31164 34638
rect 31556 34412 31612 34468
rect 30156 33740 30212 33796
rect 30716 34130 30772 34132
rect 30716 34078 30718 34130
rect 30718 34078 30770 34130
rect 30770 34078 30772 34130
rect 30716 34076 30772 34078
rect 30044 33628 30100 33684
rect 29484 33292 29540 33348
rect 30044 33346 30100 33348
rect 30044 33294 30046 33346
rect 30046 33294 30098 33346
rect 30098 33294 30100 33346
rect 30044 33292 30100 33294
rect 29820 33068 29876 33124
rect 29372 32732 29428 32788
rect 30136 32732 30192 32788
rect 29260 32562 29316 32564
rect 29260 32510 29262 32562
rect 29262 32510 29314 32562
rect 29314 32510 29316 32562
rect 30380 32674 30436 32676
rect 30380 32622 30382 32674
rect 30382 32622 30434 32674
rect 30434 32622 30436 32674
rect 30380 32620 30436 32622
rect 29260 32508 29316 32510
rect 29036 31948 29092 32004
rect 29148 32172 29204 32228
rect 29036 31778 29092 31780
rect 29036 31726 29038 31778
rect 29038 31726 29090 31778
rect 29090 31726 29092 31778
rect 29036 31724 29092 31726
rect 29540 32002 29596 32004
rect 29540 31950 29542 32002
rect 29542 31950 29594 32002
rect 29594 31950 29596 32002
rect 29540 31948 29596 31950
rect 29260 31612 29316 31668
rect 30212 31500 30268 31556
rect 29596 31276 29652 31332
rect 28028 30716 28084 30772
rect 27916 30044 27972 30100
rect 27188 29426 27244 29428
rect 27188 29374 27190 29426
rect 27190 29374 27242 29426
rect 27242 29374 27244 29426
rect 27188 29372 27244 29374
rect 27580 29596 27636 29652
rect 26740 29148 26796 29204
rect 26572 28530 26628 28532
rect 26572 28478 26574 28530
rect 26574 28478 26626 28530
rect 26626 28478 26628 28530
rect 26572 28476 26628 28478
rect 26572 28252 26628 28308
rect 26348 27858 26404 27860
rect 26348 27806 26350 27858
rect 26350 27806 26402 27858
rect 26402 27806 26404 27858
rect 26348 27804 26404 27806
rect 27300 28642 27356 28644
rect 27300 28590 27302 28642
rect 27302 28590 27354 28642
rect 27354 28590 27356 28642
rect 27300 28588 27356 28590
rect 27916 29426 27972 29428
rect 27916 29374 27918 29426
rect 27918 29374 27970 29426
rect 27970 29374 27972 29426
rect 27916 29372 27972 29374
rect 27748 29148 27804 29204
rect 27580 28364 27636 28420
rect 26852 27970 26908 27972
rect 26852 27918 26854 27970
rect 26854 27918 26906 27970
rect 26906 27918 26908 27970
rect 26852 27916 26908 27918
rect 27020 27804 27076 27860
rect 27636 27858 27692 27860
rect 27636 27806 27638 27858
rect 27638 27806 27690 27858
rect 27690 27806 27692 27858
rect 27636 27804 27692 27806
rect 27804 27858 27860 27860
rect 27804 27806 27806 27858
rect 27806 27806 27858 27858
rect 27858 27806 27860 27858
rect 27804 27804 27860 27806
rect 28252 30210 28308 30212
rect 28252 30158 28254 30210
rect 28254 30158 28306 30210
rect 28306 30158 28308 30210
rect 28252 30156 28308 30158
rect 28252 27916 28308 27972
rect 27804 27244 27860 27300
rect 27804 27074 27860 27076
rect 27804 27022 27806 27074
rect 27806 27022 27858 27074
rect 27858 27022 27860 27074
rect 27804 27020 27860 27022
rect 26460 26236 26516 26292
rect 26572 26348 26628 26404
rect 26908 26290 26964 26292
rect 26908 26238 26910 26290
rect 26910 26238 26962 26290
rect 26962 26238 26964 26290
rect 26908 26236 26964 26238
rect 26796 26012 26852 26068
rect 26348 25900 26404 25956
rect 25900 24780 25956 24836
rect 26236 25116 26292 25172
rect 25004 24332 25060 24388
rect 26124 24444 26180 24500
rect 26516 24892 26572 24948
rect 28196 27746 28252 27748
rect 28196 27694 28198 27746
rect 28198 27694 28250 27746
rect 28250 27694 28252 27746
rect 28196 27692 28252 27694
rect 28364 27468 28420 27524
rect 28476 28364 28532 28420
rect 28588 28476 28644 28532
rect 29372 30994 29428 30996
rect 29372 30942 29374 30994
rect 29374 30942 29426 30994
rect 29426 30942 29428 30994
rect 29372 30940 29428 30942
rect 30268 31276 30324 31332
rect 29204 30828 29260 30884
rect 29540 30604 29596 30660
rect 29708 30380 29764 30436
rect 29148 30210 29204 30212
rect 29148 30158 29150 30210
rect 29150 30158 29202 30210
rect 29202 30158 29204 30210
rect 29148 30156 29204 30158
rect 28812 28252 28868 28308
rect 28924 30044 28980 30100
rect 28812 27916 28868 27972
rect 29260 30044 29316 30100
rect 29148 29402 29150 29428
rect 29150 29402 29202 29428
rect 29202 29402 29204 29428
rect 29148 29372 29204 29402
rect 29148 28812 29204 28868
rect 31836 34130 31892 34132
rect 31836 34078 31838 34130
rect 31838 34078 31890 34130
rect 31890 34078 31892 34130
rect 31836 34076 31892 34078
rect 31948 34188 32004 34244
rect 32060 34636 32116 34692
rect 31052 33628 31108 33684
rect 30920 33404 30976 33460
rect 30828 33068 30884 33124
rect 31164 33292 31220 33348
rect 31500 33346 31556 33348
rect 31500 33294 31502 33346
rect 31502 33294 31554 33346
rect 31554 33294 31556 33346
rect 31500 33292 31556 33294
rect 30716 31500 30772 31556
rect 30604 31052 30660 31108
rect 30716 30994 30772 30996
rect 30716 30942 30718 30994
rect 30718 30942 30770 30994
rect 30770 30942 30772 30994
rect 30716 30940 30772 30942
rect 31836 33628 31892 33684
rect 31724 33404 31780 33460
rect 31948 33516 32004 33572
rect 32396 37548 32452 37604
rect 32396 37100 32452 37156
rect 32732 37324 32788 37380
rect 33852 37826 33908 37828
rect 33852 37774 33854 37826
rect 33854 37774 33906 37826
rect 33906 37774 33908 37826
rect 33852 37772 33908 37774
rect 33460 37548 33516 37604
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35644 38220 35700 38276
rect 33068 37324 33124 37380
rect 33944 37266 34000 37268
rect 33944 37214 33946 37266
rect 33946 37214 33998 37266
rect 33998 37214 34000 37266
rect 33944 37212 34000 37214
rect 34188 37266 34244 37268
rect 34188 37214 34190 37266
rect 34190 37214 34242 37266
rect 34242 37214 34244 37266
rect 34188 37212 34244 37214
rect 32844 37100 32900 37156
rect 32844 36594 32900 36596
rect 32844 36542 32846 36594
rect 32846 36542 32898 36594
rect 32898 36542 32900 36594
rect 32844 36540 32900 36542
rect 32396 36316 32452 36372
rect 32284 34748 32340 34804
rect 32284 33964 32340 34020
rect 32564 36092 32620 36148
rect 34300 36540 34356 36596
rect 34636 36540 34692 36596
rect 33404 36482 33460 36484
rect 33404 36430 33406 36482
rect 33406 36430 33458 36482
rect 33458 36430 33460 36482
rect 33404 36428 33460 36430
rect 33068 35868 33124 35924
rect 32732 35644 32788 35700
rect 33180 35756 33236 35812
rect 34188 36482 34244 36484
rect 34188 36430 34190 36482
rect 34190 36430 34242 36482
rect 34242 36430 34244 36482
rect 34188 36428 34244 36430
rect 33516 35644 33572 35700
rect 34076 35698 34132 35700
rect 34076 35646 34078 35698
rect 34078 35646 34130 35698
rect 34130 35646 34132 35698
rect 34076 35644 34132 35646
rect 34580 36204 34636 36260
rect 35644 37490 35700 37492
rect 35644 37438 35646 37490
rect 35646 37438 35698 37490
rect 35698 37438 35700 37490
rect 35644 37436 35700 37438
rect 35308 37266 35364 37268
rect 35308 37214 35310 37266
rect 35310 37214 35362 37266
rect 35362 37214 35364 37266
rect 35308 37212 35364 37214
rect 34916 36370 34972 36372
rect 34916 36318 34918 36370
rect 34918 36318 34970 36370
rect 34970 36318 34972 36370
rect 34916 36316 34972 36318
rect 34748 36204 34804 36260
rect 33852 35308 33908 35364
rect 32732 34748 32788 34804
rect 32172 33740 32228 33796
rect 32564 33628 32620 33684
rect 30492 30716 30548 30772
rect 30940 31724 30996 31780
rect 30492 30268 30548 30324
rect 29036 28364 29092 28420
rect 28028 26290 28084 26292
rect 28028 26238 28030 26290
rect 28030 26238 28082 26290
rect 28082 26238 28084 26290
rect 28028 26236 28084 26238
rect 27132 24892 27188 24948
rect 26908 24780 26964 24836
rect 26516 24722 26572 24724
rect 26516 24670 26518 24722
rect 26518 24670 26570 24722
rect 26570 24670 26572 24722
rect 26516 24668 26572 24670
rect 26120 24108 26176 24164
rect 25452 23212 25508 23268
rect 24892 22764 24948 22820
rect 25004 23100 25060 23156
rect 25788 23266 25844 23268
rect 25788 23214 25790 23266
rect 25790 23214 25842 23266
rect 25842 23214 25844 23266
rect 25788 23212 25844 23214
rect 25564 23100 25620 23156
rect 26124 23154 26180 23156
rect 26124 23102 26126 23154
rect 26126 23102 26178 23154
rect 26178 23102 26180 23154
rect 26124 23100 26180 23102
rect 26684 24108 26740 24164
rect 27020 24722 27076 24724
rect 27020 24670 27022 24722
rect 27022 24670 27074 24722
rect 27074 24670 27076 24722
rect 27020 24668 27076 24670
rect 26796 23938 26852 23940
rect 26796 23886 26798 23938
rect 26798 23886 26850 23938
rect 26850 23886 26852 23938
rect 26796 23884 26852 23886
rect 27468 24722 27524 24724
rect 27468 24670 27470 24722
rect 27470 24670 27522 24722
rect 27522 24670 27524 24722
rect 27468 24668 27524 24670
rect 27580 24556 27636 24612
rect 27804 25116 27860 25172
rect 27916 25004 27972 25060
rect 28700 25900 28756 25956
rect 28924 27580 28980 27636
rect 29036 27845 29038 27860
rect 29038 27845 29090 27860
rect 29090 27845 29092 27860
rect 29036 27804 29092 27845
rect 30604 30156 30660 30212
rect 30548 29708 30604 29764
rect 32732 33292 32788 33348
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35644 36876 35700 36932
rect 35196 36652 35252 36708
rect 35364 36540 35420 36596
rect 35532 36204 35588 36260
rect 35980 38332 36036 38388
rect 36988 38220 37044 38276
rect 38108 40572 38164 40628
rect 37604 39058 37660 39060
rect 37604 39006 37606 39058
rect 37606 39006 37658 39058
rect 37658 39006 37660 39058
rect 37604 39004 37660 39006
rect 38332 41468 38388 41524
rect 40796 46114 40852 46116
rect 40796 46062 40798 46114
rect 40798 46062 40850 46114
rect 40850 46062 40852 46114
rect 40796 46060 40852 46062
rect 41132 45836 41188 45892
rect 39788 45500 39844 45556
rect 40460 45724 40516 45780
rect 40348 44940 40404 44996
rect 39676 44492 39732 44548
rect 39900 44044 39956 44100
rect 39228 42364 39284 42420
rect 39452 42028 39508 42084
rect 39228 41804 39284 41860
rect 39228 41580 39284 41636
rect 40236 43148 40292 43204
rect 40236 42364 40292 42420
rect 40012 42028 40068 42084
rect 39564 41468 39620 41524
rect 39844 41804 39900 41860
rect 38780 41132 38836 41188
rect 38332 40572 38388 40628
rect 38332 40402 38388 40404
rect 38332 40350 38334 40402
rect 38334 40350 38386 40402
rect 38386 40350 38388 40402
rect 38332 40348 38388 40350
rect 38220 40124 38276 40180
rect 38220 39618 38276 39620
rect 38220 39566 38222 39618
rect 38222 39566 38274 39618
rect 38274 39566 38276 39618
rect 38220 39564 38276 39566
rect 38108 39004 38164 39060
rect 38444 39452 38500 39508
rect 37212 37884 37268 37940
rect 37884 38892 37940 38948
rect 38332 38892 38388 38948
rect 36988 37772 37044 37828
rect 37436 38050 37492 38052
rect 37436 37998 37438 38050
rect 37438 37998 37490 38050
rect 37490 37998 37492 38050
rect 37436 37996 37492 37998
rect 37996 38668 38052 38724
rect 38108 38444 38164 38500
rect 37884 38332 37940 38388
rect 39452 40460 39508 40516
rect 39004 39900 39060 39956
rect 38892 39116 38948 39172
rect 39004 39004 39060 39060
rect 38444 38220 38500 38276
rect 37324 37436 37380 37492
rect 36260 37154 36316 37156
rect 36260 37102 36262 37154
rect 36262 37102 36314 37154
rect 36314 37102 36316 37154
rect 36260 37100 36316 37102
rect 36652 37154 36708 37156
rect 36652 37102 36654 37154
rect 36654 37102 36706 37154
rect 36706 37102 36708 37154
rect 36652 37100 36708 37102
rect 37046 37266 37102 37268
rect 37046 37214 37048 37266
rect 37048 37214 37100 37266
rect 37100 37214 37102 37266
rect 37046 37212 37102 37214
rect 36876 36316 36932 36372
rect 35924 35868 35980 35924
rect 35644 35532 35700 35588
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 33852 34300 33908 34356
rect 33964 34188 34020 34244
rect 33068 34130 33124 34132
rect 33068 34078 33070 34130
rect 33070 34078 33122 34130
rect 33122 34078 33124 34130
rect 33068 34076 33124 34078
rect 34300 33964 34356 34020
rect 32844 32732 32900 32788
rect 33068 33346 33124 33348
rect 33068 33294 33070 33346
rect 33070 33294 33122 33346
rect 33122 33294 33124 33346
rect 33068 33292 33124 33294
rect 32284 32620 32340 32676
rect 33740 33180 33796 33236
rect 33404 32956 33460 33012
rect 33180 32844 33236 32900
rect 31836 31778 31892 31780
rect 31836 31726 31838 31778
rect 31838 31726 31890 31778
rect 31890 31726 31892 31778
rect 31836 31724 31892 31726
rect 31612 31276 31668 31332
rect 31164 31052 31220 31108
rect 30940 30268 30996 30324
rect 30044 29036 30100 29092
rect 30828 30044 30884 30100
rect 30828 29708 30884 29764
rect 31276 30044 31332 30100
rect 29708 28700 29764 28756
rect 29484 28476 29540 28532
rect 30604 28588 30660 28644
rect 32116 31164 32172 31220
rect 32040 30828 32096 30884
rect 32284 30994 32340 30996
rect 32284 30942 32286 30994
rect 32286 30942 32338 30994
rect 32338 30942 32340 30994
rect 32284 30940 32340 30942
rect 32508 31612 32564 31668
rect 32172 30180 32228 30212
rect 32172 30156 32174 30180
rect 32174 30156 32226 30180
rect 32226 30156 32228 30180
rect 31948 29426 32004 29428
rect 31948 29374 31950 29426
rect 31950 29374 32002 29426
rect 32002 29374 32004 29426
rect 31948 29372 32004 29374
rect 31612 29260 31668 29316
rect 30044 28252 30100 28308
rect 29372 28028 29428 28084
rect 29260 27046 29316 27076
rect 29260 27020 29262 27046
rect 29262 27020 29314 27046
rect 29314 27020 29316 27046
rect 29036 26796 29092 26852
rect 29148 26572 29204 26628
rect 29596 27580 29652 27636
rect 29484 26572 29540 26628
rect 28812 25676 28868 25732
rect 28364 25452 28420 25508
rect 28252 25116 28308 25172
rect 29036 24780 29092 24836
rect 29260 25506 29316 25508
rect 29260 25454 29262 25506
rect 29262 25454 29314 25506
rect 29314 25454 29316 25506
rect 29260 25452 29316 25454
rect 27692 24220 27748 24276
rect 27692 23772 27748 23828
rect 28476 24668 28532 24724
rect 29148 24556 29204 24612
rect 29484 26290 29540 26292
rect 29484 26238 29486 26290
rect 29486 26238 29538 26290
rect 29538 26238 29540 26290
rect 29484 26236 29540 26238
rect 29820 27468 29876 27524
rect 29708 27132 29764 27188
rect 29708 25452 29764 25508
rect 29932 27244 29988 27300
rect 30940 27692 30996 27748
rect 30492 27468 30548 27524
rect 30380 27020 30436 27076
rect 30156 26796 30212 26852
rect 29820 26236 29876 26292
rect 29988 26402 30044 26404
rect 29988 26350 29990 26402
rect 29990 26350 30042 26402
rect 30042 26350 30044 26402
rect 29988 26348 30044 26350
rect 29988 25452 30044 25508
rect 32900 31724 32956 31780
rect 36092 35532 36148 35588
rect 35868 35196 35924 35252
rect 36540 34972 36596 35028
rect 37212 36988 37268 37044
rect 37436 36876 37492 36932
rect 37716 37772 37772 37828
rect 37548 36540 37604 36596
rect 37212 35644 37268 35700
rect 37884 37548 37940 37604
rect 37324 36316 37380 36372
rect 36876 35084 36932 35140
rect 37100 35196 37156 35252
rect 36764 34972 36820 35028
rect 34692 34076 34748 34132
rect 36652 34076 36708 34132
rect 35663 33964 35719 34020
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 33516 35252 33572
rect 34972 33346 35028 33348
rect 34972 33294 34974 33346
rect 34974 33294 35026 33346
rect 35026 33294 35028 33346
rect 34972 33292 35028 33294
rect 35532 33516 35588 33572
rect 36316 33628 36372 33684
rect 36988 34354 37044 34356
rect 36988 34302 36990 34354
rect 36990 34302 37042 34354
rect 37042 34302 37044 34354
rect 36988 34300 37044 34302
rect 36876 33516 36932 33572
rect 36988 34076 37044 34132
rect 37660 35980 37716 36036
rect 37436 35698 37492 35700
rect 37436 35646 37438 35698
rect 37438 35646 37490 35698
rect 37490 35646 37492 35698
rect 37436 35644 37492 35646
rect 37548 35532 37604 35588
rect 38556 38444 38612 38500
rect 38556 37996 38612 38052
rect 38220 37772 38276 37828
rect 39676 40460 39732 40516
rect 40852 44940 40908 44996
rect 40908 44546 40964 44548
rect 40908 44494 40910 44546
rect 40910 44494 40962 44546
rect 40962 44494 40964 44546
rect 40908 44492 40964 44494
rect 41020 44044 41076 44100
rect 41244 45276 41300 45332
rect 41356 45388 41412 45444
rect 41244 44828 41300 44884
rect 42252 45106 42308 45108
rect 42252 45054 42254 45106
rect 42254 45054 42306 45106
rect 42306 45054 42308 45106
rect 42252 45052 42308 45054
rect 41468 44380 41524 44436
rect 41804 44380 41860 44436
rect 42140 44044 42196 44100
rect 42476 43484 42532 43540
rect 42588 45052 42644 45108
rect 42420 43148 42476 43204
rect 41132 42812 41188 42868
rect 40124 39900 40180 39956
rect 39228 38946 39284 38948
rect 39228 38894 39230 38946
rect 39230 38894 39282 38946
rect 39282 38894 39284 38946
rect 39228 38892 39284 38894
rect 39564 39116 39620 39172
rect 39900 39058 39956 39060
rect 39900 39006 39902 39058
rect 39902 39006 39954 39058
rect 39954 39006 39956 39058
rect 39900 39004 39956 39006
rect 39452 38556 39508 38612
rect 38892 37436 38948 37492
rect 37996 37100 38052 37156
rect 40908 42476 40964 42532
rect 40796 41970 40852 41972
rect 40796 41918 40798 41970
rect 40798 41918 40850 41970
rect 40850 41918 40852 41970
rect 40796 41916 40852 41918
rect 40684 39564 40740 39620
rect 40796 38834 40852 38836
rect 40796 38782 40798 38834
rect 40798 38782 40850 38834
rect 40850 38782 40852 38834
rect 40796 38780 40852 38782
rect 40684 38668 40740 38724
rect 40908 38220 40964 38276
rect 40852 37938 40908 37940
rect 40852 37886 40854 37938
rect 40854 37886 40906 37938
rect 40906 37886 40908 37938
rect 40852 37884 40908 37886
rect 40012 37436 40068 37492
rect 39564 36482 39620 36484
rect 39564 36430 39566 36482
rect 39566 36430 39618 36482
rect 39618 36430 39620 36482
rect 39564 36428 39620 36430
rect 38612 35810 38668 35812
rect 38612 35758 38614 35810
rect 38614 35758 38666 35810
rect 38666 35758 38668 35810
rect 38612 35756 38668 35758
rect 37716 35196 37772 35252
rect 38108 35644 38164 35700
rect 38892 35698 38948 35700
rect 38892 35646 38894 35698
rect 38894 35646 38946 35698
rect 38946 35646 38948 35698
rect 38892 35644 38948 35646
rect 37660 35026 37716 35028
rect 37660 34974 37662 35026
rect 37662 34974 37714 35026
rect 37714 34974 37716 35026
rect 37660 34972 37716 34974
rect 37828 34300 37884 34356
rect 37100 33628 37156 33684
rect 36316 33346 36372 33348
rect 34524 32956 34580 33012
rect 33068 30994 33124 30996
rect 33068 30942 33070 30994
rect 33070 30942 33122 30994
rect 33122 30942 33124 30994
rect 33068 30940 33124 30942
rect 32508 30380 32564 30436
rect 32396 30268 32452 30324
rect 32564 30044 32620 30100
rect 33180 30268 33236 30324
rect 33516 30380 33572 30436
rect 33628 30210 33684 30212
rect 33628 30158 33630 30210
rect 33630 30158 33682 30210
rect 33682 30158 33684 30210
rect 33628 30156 33684 30158
rect 33180 29932 33236 29988
rect 32284 29148 32340 29204
rect 31836 28924 31892 28980
rect 32844 28812 32900 28868
rect 31724 28588 31780 28644
rect 32564 28642 32620 28644
rect 32564 28590 32566 28642
rect 32566 28590 32618 28642
rect 32618 28590 32620 28642
rect 32564 28588 32620 28590
rect 31052 26572 31108 26628
rect 32732 28364 32788 28420
rect 30492 26178 30548 26180
rect 30492 26126 30494 26178
rect 30494 26126 30546 26178
rect 30546 26126 30548 26178
rect 30492 26124 30548 26126
rect 29484 24722 29540 24724
rect 29484 24670 29486 24722
rect 29486 24670 29538 24722
rect 29538 24670 29540 24722
rect 29484 24668 29540 24670
rect 28868 24332 28924 24388
rect 28252 23436 28308 23492
rect 27020 23212 27076 23268
rect 27692 23212 27748 23268
rect 26572 22876 26628 22932
rect 23660 21868 23716 21924
rect 24892 22092 24948 22148
rect 24500 21868 24556 21924
rect 25060 21868 25116 21924
rect 23436 21084 23492 21140
rect 23324 20802 23380 20804
rect 23324 20750 23326 20802
rect 23326 20750 23378 20802
rect 23378 20750 23380 20802
rect 23324 20748 23380 20750
rect 24276 21698 24332 21700
rect 24276 21646 24278 21698
rect 24278 21646 24330 21698
rect 24330 21646 24332 21698
rect 24276 21644 24332 21646
rect 25116 21644 25172 21700
rect 23436 20300 23492 20356
rect 23548 20188 23604 20244
rect 24108 20076 24164 20132
rect 23492 19964 23548 20020
rect 23100 19794 23156 19796
rect 23100 19742 23102 19794
rect 23102 19742 23154 19794
rect 23154 19742 23156 19794
rect 23100 19740 23156 19742
rect 23156 19516 23212 19572
rect 24108 19906 24164 19908
rect 24108 19854 24110 19906
rect 24110 19854 24162 19906
rect 24162 19854 24164 19906
rect 24108 19852 24164 19854
rect 23772 19740 23828 19796
rect 23660 19516 23716 19572
rect 22988 18450 23044 18452
rect 22988 18398 22990 18450
rect 22990 18398 23042 18450
rect 23042 18398 23044 18450
rect 24724 21586 24780 21588
rect 24724 21534 24726 21586
rect 24726 21534 24778 21586
rect 24778 21534 24780 21586
rect 24724 21532 24780 21534
rect 24892 20914 24948 20916
rect 24892 20862 24894 20914
rect 24894 20862 24946 20914
rect 24946 20862 24948 20914
rect 24892 20860 24948 20862
rect 25452 21532 25508 21588
rect 26124 21644 26180 21700
rect 26236 22652 26292 22708
rect 26012 21532 26068 21588
rect 25676 20748 25732 20804
rect 25452 20300 25508 20356
rect 25564 20524 25620 20580
rect 26796 22764 26852 22820
rect 27244 22930 27300 22932
rect 27244 22878 27246 22930
rect 27246 22878 27298 22930
rect 27298 22878 27300 22930
rect 27244 22876 27300 22878
rect 26908 22652 26964 22708
rect 27960 23140 27962 23156
rect 27962 23140 28014 23156
rect 28014 23140 28016 23156
rect 27960 23100 28016 23140
rect 28252 23100 28308 23156
rect 28364 23660 28420 23716
rect 28700 23772 28756 23828
rect 29260 23772 29316 23828
rect 29372 23884 29428 23940
rect 28700 22876 28756 22932
rect 30156 25116 30212 25172
rect 30268 24780 30324 24836
rect 30716 26012 30772 26068
rect 30492 25340 30548 25396
rect 30604 25452 30660 25508
rect 28588 22764 28644 22820
rect 27692 22316 27748 22372
rect 27356 22092 27412 22148
rect 26460 21980 26516 22036
rect 26124 21196 26180 21252
rect 25116 20076 25172 20132
rect 24332 19740 24388 19796
rect 24052 19516 24108 19572
rect 25564 20188 25620 20244
rect 25452 20018 25508 20020
rect 25452 19966 25454 20018
rect 25454 19966 25506 20018
rect 25506 19966 25508 20018
rect 25452 19964 25508 19966
rect 27198 21756 27254 21812
rect 27972 21810 28028 21812
rect 27972 21758 27974 21810
rect 27974 21758 28026 21810
rect 28026 21758 28028 21810
rect 27972 21756 28028 21758
rect 29640 22332 29696 22372
rect 29640 22316 29642 22332
rect 29642 22316 29694 22332
rect 29694 22316 29696 22332
rect 30492 24556 30548 24612
rect 30156 24220 30212 24276
rect 30000 23660 30056 23716
rect 29932 23154 29988 23156
rect 29932 23102 29934 23154
rect 29934 23102 29986 23154
rect 29986 23102 29988 23154
rect 29932 23100 29988 23102
rect 30380 24108 30436 24164
rect 29932 22764 29988 22820
rect 30604 24220 30660 24276
rect 30940 25900 30996 25956
rect 30828 25788 30884 25844
rect 31052 25506 31108 25508
rect 31052 25454 31054 25506
rect 31054 25454 31106 25506
rect 31106 25454 31108 25506
rect 31052 25452 31108 25454
rect 32564 28082 32620 28084
rect 32564 28030 32566 28082
rect 32566 28030 32618 28082
rect 32618 28030 32620 28082
rect 32564 28028 32620 28030
rect 32116 27970 32172 27972
rect 32116 27918 32118 27970
rect 32118 27918 32170 27970
rect 32170 27918 32172 27970
rect 32116 27916 32172 27918
rect 32732 27132 32788 27188
rect 31612 27074 31668 27076
rect 31612 27022 31614 27074
rect 31614 27022 31666 27074
rect 31666 27022 31668 27074
rect 31612 27020 31668 27022
rect 31836 26796 31892 26852
rect 31668 26572 31724 26628
rect 32116 26572 32172 26628
rect 32732 26572 32788 26628
rect 31836 26012 31892 26068
rect 31164 25340 31220 25396
rect 31332 25228 31388 25284
rect 32172 25340 32228 25396
rect 32060 24892 32116 24948
rect 31948 24780 32004 24836
rect 31724 24668 31780 24724
rect 30940 24108 30996 24164
rect 31724 24220 31780 24276
rect 30828 23660 30884 23716
rect 29820 21756 29876 21812
rect 26796 21196 26852 21252
rect 26796 20972 26852 21028
rect 29148 21532 29204 21588
rect 26572 20076 26628 20132
rect 23884 19234 23940 19236
rect 23884 19182 23886 19234
rect 23886 19182 23938 19234
rect 23938 19182 23940 19234
rect 23884 19180 23940 19182
rect 24220 18956 24276 19012
rect 23772 18844 23828 18900
rect 25004 19292 25060 19348
rect 24836 19180 24892 19236
rect 24556 18956 24612 19012
rect 22988 18396 23044 18398
rect 23212 18172 23268 18228
rect 22876 16268 22932 16324
rect 23436 17724 23492 17780
rect 23548 17612 23604 17668
rect 23660 18396 23716 18452
rect 24556 18508 24612 18564
rect 25676 19292 25732 19348
rect 25564 19180 25620 19236
rect 25284 19122 25340 19124
rect 25284 19070 25286 19122
rect 25286 19070 25338 19122
rect 25338 19070 25340 19122
rect 25284 19068 25340 19070
rect 24780 18956 24836 19012
rect 23324 17276 23380 17332
rect 23716 17276 23772 17332
rect 23212 17164 23268 17220
rect 23380 17106 23436 17108
rect 23380 17054 23382 17106
rect 23382 17054 23434 17106
rect 23434 17054 23436 17106
rect 23380 17052 23436 17054
rect 23436 16716 23492 16772
rect 21756 15148 21812 15204
rect 22316 15148 22372 15204
rect 22148 15036 22204 15092
rect 22540 15372 22596 15428
rect 22428 14700 22484 14756
rect 21756 13804 21812 13860
rect 21980 13746 22036 13748
rect 21980 13694 21982 13746
rect 21982 13694 22034 13746
rect 22034 13694 22036 13746
rect 21980 13692 22036 13694
rect 21308 13580 21364 13636
rect 20748 13020 20804 13076
rect 20636 12962 20692 12964
rect 20636 12910 20638 12962
rect 20638 12910 20690 12962
rect 20690 12910 20692 12962
rect 20636 12908 20692 12910
rect 22428 13580 22484 13636
rect 22316 13468 22372 13524
rect 22652 14140 22708 14196
rect 22540 13468 22596 13524
rect 22092 13356 22148 13412
rect 21700 13132 21756 13188
rect 21756 12962 21812 12964
rect 21756 12910 21758 12962
rect 21758 12910 21810 12962
rect 21810 12910 21812 12962
rect 21756 12908 21812 12910
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19068 11900 19124 11956
rect 18732 11676 18788 11732
rect 18844 11116 18900 11172
rect 18172 9436 18228 9492
rect 19404 12124 19460 12180
rect 19684 12348 19740 12404
rect 21644 12236 21700 12292
rect 19852 12178 19908 12180
rect 19852 12126 19854 12178
rect 19854 12126 19906 12178
rect 19906 12126 19908 12178
rect 19852 12124 19908 12126
rect 21756 12124 21812 12180
rect 19404 11676 19460 11732
rect 18844 9788 18900 9828
rect 16380 8428 16436 8484
rect 15260 8204 15316 8260
rect 16156 7980 16212 8036
rect 15036 7474 15092 7476
rect 15036 7422 15038 7474
rect 15038 7422 15090 7474
rect 15090 7422 15092 7474
rect 15036 7420 15092 7422
rect 14252 6860 14308 6916
rect 14700 6972 14756 7028
rect 13916 5964 13972 6020
rect 13468 5180 13524 5236
rect 12684 4956 12740 5012
rect 13468 5010 13524 5012
rect 13468 4958 13470 5010
rect 13470 4958 13522 5010
rect 13522 4958 13524 5010
rect 13468 4956 13524 4958
rect 15912 6972 15968 7028
rect 14476 6524 14532 6580
rect 14700 6300 14756 6356
rect 14196 5292 14252 5348
rect 14588 4956 14644 5012
rect 13804 4732 13860 4788
rect 14476 4732 14532 4788
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 12572 3948 12628 4004
rect 13356 3948 13412 4004
rect 4684 3892 4740 3894
rect 13356 3724 13412 3780
rect 15148 6860 15204 6916
rect 14924 6412 14980 6468
rect 15036 6651 15092 6692
rect 15036 6636 15038 6651
rect 15038 6636 15090 6651
rect 15090 6636 15092 6651
rect 15260 6524 15316 6580
rect 15148 5852 15204 5908
rect 18060 8428 18116 8484
rect 16940 7474 16996 7476
rect 16940 7422 16942 7474
rect 16942 7422 16994 7474
rect 16994 7422 16996 7474
rect 16940 7420 16996 7422
rect 17948 7420 18004 7476
rect 18060 7308 18116 7364
rect 16772 6972 16828 7028
rect 16380 6662 16436 6692
rect 16380 6636 16382 6662
rect 16382 6636 16434 6662
rect 16434 6636 16436 6662
rect 17052 6690 17108 6692
rect 17052 6638 17054 6690
rect 17054 6638 17106 6690
rect 17106 6638 17108 6690
rect 17052 6636 17108 6638
rect 17388 6690 17444 6692
rect 17388 6638 17390 6690
rect 17390 6638 17442 6690
rect 17442 6638 17444 6690
rect 17388 6636 17444 6638
rect 15932 6578 15988 6580
rect 15932 6526 15934 6578
rect 15934 6526 15986 6578
rect 15986 6526 15988 6578
rect 15932 6524 15988 6526
rect 17836 6412 17892 6468
rect 15764 6300 15820 6356
rect 17612 6300 17668 6356
rect 14476 3612 14532 3668
rect 15260 5180 15316 5236
rect 15036 4284 15092 4340
rect 15372 4956 15428 5012
rect 15708 5906 15764 5908
rect 15708 5854 15710 5906
rect 15710 5854 15762 5906
rect 15762 5854 15764 5906
rect 15708 5852 15764 5854
rect 16044 5740 16100 5796
rect 16492 5869 16494 5908
rect 16494 5869 16546 5908
rect 16546 5869 16548 5908
rect 16492 5852 16548 5869
rect 18844 9772 18846 9788
rect 18846 9772 18898 9788
rect 18898 9772 18900 9788
rect 20804 12066 20860 12068
rect 20804 12014 20806 12066
rect 20806 12014 20858 12066
rect 20858 12014 20860 12066
rect 20804 12012 20860 12014
rect 20188 11954 20244 11956
rect 20188 11902 20190 11954
rect 20190 11902 20242 11954
rect 20242 11902 20244 11954
rect 20188 11900 20244 11902
rect 19628 11340 19684 11396
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19404 9884 19460 9940
rect 19852 10498 19908 10500
rect 19852 10446 19854 10498
rect 19854 10446 19906 10498
rect 19906 10446 19908 10498
rect 19852 10444 19908 10446
rect 20300 11788 20356 11844
rect 21252 11788 21308 11844
rect 21420 11900 21476 11956
rect 22988 15148 23044 15204
rect 22932 13970 22988 13972
rect 22932 13918 22934 13970
rect 22934 13918 22986 13970
rect 22986 13918 22988 13970
rect 22932 13916 22988 13918
rect 23212 16044 23268 16100
rect 23212 15148 23268 15204
rect 23324 15484 23380 15540
rect 23436 15372 23492 15428
rect 23324 14812 23380 14868
rect 24444 18396 24500 18452
rect 24388 17948 24444 18004
rect 24332 17164 24388 17220
rect 23996 16940 24052 16996
rect 23660 16828 23716 16884
rect 23884 16882 23940 16884
rect 23884 16830 23886 16882
rect 23886 16830 23938 16882
rect 23938 16830 23940 16882
rect 23884 16828 23940 16830
rect 23884 16156 23940 16212
rect 24220 15090 24276 15092
rect 24220 15038 24222 15090
rect 24222 15038 24274 15090
rect 24274 15038 24276 15090
rect 24220 15036 24276 15038
rect 25340 18844 25396 18900
rect 26124 19234 26180 19236
rect 26124 19182 26126 19234
rect 26126 19182 26178 19234
rect 26178 19182 26180 19234
rect 26124 19180 26180 19182
rect 26460 18732 26516 18788
rect 26796 18508 26852 18564
rect 26236 18396 26292 18452
rect 25228 18060 25284 18116
rect 26068 17836 26124 17892
rect 26236 18172 26292 18228
rect 25116 17052 25172 17108
rect 25228 17666 25284 17668
rect 25228 17614 25230 17666
rect 25230 17614 25282 17666
rect 25282 17614 25284 17666
rect 25228 17612 25284 17614
rect 25004 16268 25060 16324
rect 25004 15932 25060 15988
rect 25340 17388 25396 17444
rect 25452 17164 25508 17220
rect 25732 17164 25788 17220
rect 25900 17500 25956 17556
rect 26124 17052 26180 17108
rect 25676 16882 25732 16884
rect 25676 16830 25678 16882
rect 25678 16830 25730 16882
rect 25730 16830 25732 16882
rect 25676 16828 25732 16830
rect 25452 16492 25508 16548
rect 25228 15260 25284 15316
rect 24556 14924 24612 14980
rect 23996 14754 24052 14756
rect 23996 14702 23998 14754
rect 23998 14702 24050 14754
rect 24050 14702 24052 14754
rect 23996 14700 24052 14702
rect 24108 13916 24164 13972
rect 23100 13356 23156 13412
rect 22316 13132 22372 13188
rect 22092 12290 22148 12292
rect 22092 12238 22094 12290
rect 22094 12238 22146 12290
rect 22146 12238 22148 12290
rect 22092 12236 22148 12238
rect 22484 12348 22540 12404
rect 21980 12178 22036 12180
rect 21980 12126 21982 12178
rect 21982 12126 22034 12178
rect 22034 12126 22036 12178
rect 21980 12124 22036 12126
rect 22876 13020 22932 13076
rect 22764 12962 22820 12964
rect 22764 12910 22766 12962
rect 22766 12910 22818 12962
rect 22818 12910 22820 12962
rect 22764 12908 22820 12910
rect 23044 12796 23100 12852
rect 23324 12908 23380 12964
rect 23436 13132 23492 13188
rect 23548 12908 23604 12964
rect 23380 12236 23436 12292
rect 22428 12012 22484 12068
rect 21700 11340 21756 11396
rect 21868 11676 21924 11732
rect 21756 10780 21812 10836
rect 22596 11788 22652 11844
rect 22428 11676 22484 11732
rect 21980 10780 22036 10836
rect 20524 10444 20580 10500
rect 20804 10108 20860 10164
rect 20076 9788 20132 9828
rect 20076 9772 20078 9788
rect 20078 9772 20130 9788
rect 20130 9772 20132 9788
rect 18508 7980 18564 8036
rect 18322 7308 18378 7364
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 22652 10108 22708 10164
rect 23100 12178 23156 12180
rect 23100 12126 23102 12178
rect 23102 12126 23154 12178
rect 23154 12126 23156 12178
rect 23100 12124 23156 12126
rect 23548 12012 23604 12068
rect 23772 12738 23828 12740
rect 23772 12686 23774 12738
rect 23774 12686 23826 12738
rect 23826 12686 23828 12738
rect 23772 12684 23828 12686
rect 23380 11788 23436 11844
rect 23156 11676 23212 11732
rect 22540 9884 22596 9940
rect 22428 9826 22484 9828
rect 22428 9774 22430 9826
rect 22430 9774 22482 9826
rect 22482 9774 22484 9826
rect 22428 9772 22484 9774
rect 22708 9884 22764 9940
rect 23436 10108 23492 10164
rect 23996 12460 24052 12516
rect 23772 11900 23828 11956
rect 23772 10892 23828 10948
rect 23660 9996 23716 10052
rect 24668 14530 24724 14532
rect 24668 14478 24670 14530
rect 24670 14478 24722 14530
rect 24722 14478 24724 14530
rect 24668 14476 24724 14478
rect 24780 13916 24836 13972
rect 24444 12962 24500 12964
rect 24444 12910 24446 12962
rect 24446 12910 24498 12962
rect 24498 12910 24500 12962
rect 24444 12908 24500 12910
rect 24332 12796 24388 12852
rect 24892 13020 24948 13076
rect 24612 12796 24668 12852
rect 24780 12124 24836 12180
rect 24052 11394 24108 11396
rect 24052 11342 24054 11394
rect 24054 11342 24106 11394
rect 24106 11342 24108 11394
rect 24052 11340 24108 11342
rect 24500 11452 24556 11508
rect 24332 11394 24388 11396
rect 24332 11342 24334 11394
rect 24334 11342 24386 11394
rect 24386 11342 24388 11394
rect 25452 16044 25508 16100
rect 25228 14476 25284 14532
rect 26628 18284 26684 18340
rect 26460 18172 26516 18228
rect 26796 18060 26852 18116
rect 26460 17948 26516 18004
rect 26628 17948 26684 18004
rect 26628 17500 26684 17556
rect 27020 20188 27076 20244
rect 28028 20188 28084 20244
rect 27132 20130 27188 20132
rect 27132 20078 27134 20130
rect 27134 20078 27186 20130
rect 27186 20078 27188 20130
rect 27132 20076 27188 20078
rect 28420 20242 28476 20244
rect 28420 20190 28422 20242
rect 28422 20190 28474 20242
rect 28474 20190 28476 20242
rect 28420 20188 28476 20190
rect 28868 20242 28924 20244
rect 28868 20190 28870 20242
rect 28870 20190 28922 20242
rect 28922 20190 28924 20242
rect 28868 20188 28924 20190
rect 28028 20018 28084 20020
rect 28028 19966 28030 20018
rect 28030 19966 28082 20018
rect 28082 19966 28084 20018
rect 28028 19964 28084 19966
rect 27020 18450 27076 18452
rect 27020 18398 27022 18450
rect 27022 18398 27074 18450
rect 27074 18398 27076 18450
rect 27020 18396 27076 18398
rect 27692 19180 27748 19236
rect 27860 19292 27916 19348
rect 27860 19010 27916 19012
rect 27860 18958 27862 19010
rect 27862 18958 27914 19010
rect 27914 18958 27916 19010
rect 27860 18956 27916 18958
rect 28140 19180 28196 19236
rect 29372 21420 29428 21476
rect 29708 21586 29764 21588
rect 29708 21534 29710 21586
rect 29710 21534 29762 21586
rect 29762 21534 29764 21586
rect 29708 21532 29764 21534
rect 29820 19234 29876 19236
rect 29820 19182 29822 19234
rect 29822 19182 29874 19234
rect 29874 19182 29876 19234
rect 29820 19180 29876 19182
rect 28308 19010 28364 19012
rect 28308 18958 28310 19010
rect 28310 18958 28362 19010
rect 28362 18958 28364 19010
rect 28308 18956 28364 18958
rect 27468 18284 27524 18340
rect 26908 17948 26964 18004
rect 26348 17164 26404 17220
rect 26684 17106 26740 17108
rect 26684 17054 26686 17106
rect 26686 17054 26738 17106
rect 26738 17054 26740 17106
rect 26684 17052 26740 17054
rect 26348 16882 26404 16884
rect 26348 16830 26350 16882
rect 26350 16830 26402 16882
rect 26402 16830 26404 16882
rect 26348 16828 26404 16830
rect 25956 16268 26012 16324
rect 26348 16604 26404 16660
rect 26236 16098 26292 16100
rect 26236 16046 26238 16098
rect 26238 16046 26290 16098
rect 26290 16046 26292 16098
rect 26236 16044 26292 16046
rect 26068 15874 26124 15876
rect 26068 15822 26070 15874
rect 26070 15822 26122 15874
rect 26122 15822 26124 15874
rect 26068 15820 26124 15822
rect 25732 15202 25788 15204
rect 25732 15150 25734 15202
rect 25734 15150 25786 15202
rect 25786 15150 25788 15202
rect 25732 15148 25788 15150
rect 25564 14924 25620 14980
rect 25900 15036 25956 15092
rect 25452 14028 25508 14084
rect 25732 14028 25788 14084
rect 25340 13916 25396 13972
rect 25900 13916 25956 13972
rect 25396 13468 25452 13524
rect 25564 13356 25620 13412
rect 25172 12962 25228 12964
rect 25172 12910 25174 12962
rect 25174 12910 25226 12962
rect 25226 12910 25228 12962
rect 25172 12908 25228 12910
rect 24332 11340 24388 11342
rect 24780 10780 24836 10836
rect 24220 10332 24276 10388
rect 23380 9884 23436 9940
rect 23884 9884 23940 9940
rect 23660 9826 23716 9828
rect 23660 9774 23662 9826
rect 23662 9774 23714 9826
rect 23714 9774 23716 9826
rect 23660 9772 23716 9774
rect 22540 9660 22596 9716
rect 23548 9714 23604 9716
rect 23548 9662 23550 9714
rect 23550 9662 23602 9714
rect 23602 9662 23604 9714
rect 23548 9660 23604 9662
rect 22988 9548 23044 9604
rect 21252 8764 21308 8820
rect 19404 8428 19460 8484
rect 20132 8428 20188 8484
rect 18732 8092 18788 8148
rect 19180 7474 19236 7476
rect 19180 7422 19182 7474
rect 19182 7422 19234 7474
rect 19234 7422 19236 7474
rect 19180 7420 19236 7422
rect 18396 6524 18452 6580
rect 18508 6412 18564 6468
rect 16828 5740 16884 5796
rect 18172 5740 18228 5796
rect 17164 5180 17220 5236
rect 16044 4396 16100 4452
rect 16044 3724 16100 3780
rect 17948 5122 18004 5124
rect 17948 5070 17950 5122
rect 17950 5070 18002 5122
rect 18002 5070 18004 5122
rect 17948 5068 18004 5070
rect 17444 4396 17500 4452
rect 17276 4338 17332 4340
rect 17276 4286 17278 4338
rect 17278 4286 17330 4338
rect 17330 4286 17332 4338
rect 17276 4284 17332 4286
rect 17836 3612 17892 3668
rect 16268 3554 16324 3556
rect 16268 3502 16270 3554
rect 16270 3502 16322 3554
rect 16322 3502 16324 3554
rect 16268 3500 16324 3502
rect 17556 3554 17612 3556
rect 17556 3502 17558 3554
rect 17558 3502 17610 3554
rect 17610 3502 17612 3554
rect 17556 3500 17612 3502
rect 12628 3442 12684 3444
rect 12628 3390 12630 3442
rect 12630 3390 12682 3442
rect 12682 3390 12684 3442
rect 12628 3388 12684 3390
rect 18844 6636 18900 6692
rect 18732 5852 18788 5908
rect 18284 4956 18340 5012
rect 18956 5292 19012 5348
rect 18900 5122 18956 5124
rect 18900 5070 18902 5122
rect 18902 5070 18954 5122
rect 18954 5070 18956 5122
rect 18900 5068 18956 5070
rect 19068 5122 19124 5124
rect 19068 5070 19070 5122
rect 19070 5070 19122 5122
rect 19122 5070 19124 5122
rect 19068 5068 19124 5070
rect 21980 8428 22036 8484
rect 21868 8230 21924 8260
rect 21868 8204 21870 8230
rect 21870 8204 21922 8230
rect 21922 8204 21924 8230
rect 20300 8092 20356 8148
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 22316 8428 22372 8484
rect 19292 6636 19348 6692
rect 20020 6636 20076 6692
rect 20468 6690 20524 6692
rect 20468 6638 20470 6690
rect 20470 6638 20522 6690
rect 20522 6638 20524 6690
rect 21756 6662 21812 6692
rect 20468 6636 20524 6638
rect 19628 6524 19684 6580
rect 21756 6636 21758 6662
rect 21758 6636 21810 6662
rect 21810 6636 21812 6662
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 20860 5906 20916 5908
rect 20860 5854 20862 5906
rect 20862 5854 20914 5906
rect 20914 5854 20916 5906
rect 20860 5852 20916 5854
rect 20300 5292 20356 5348
rect 19292 5068 19348 5124
rect 19516 5180 19572 5236
rect 19068 4172 19124 4228
rect 18732 3836 18788 3892
rect 18396 3666 18452 3668
rect 18396 3614 18398 3666
rect 18398 3614 18450 3666
rect 18450 3614 18452 3666
rect 18396 3612 18452 3614
rect 18732 3554 18788 3556
rect 18732 3502 18734 3554
rect 18734 3502 18786 3554
rect 18786 3502 18788 3554
rect 18732 3500 18788 3502
rect 20188 5122 20244 5124
rect 20188 5070 20190 5122
rect 20190 5070 20242 5122
rect 20242 5070 20244 5122
rect 20188 5068 20244 5070
rect 21196 5292 21252 5348
rect 20804 5234 20860 5236
rect 20804 5182 20806 5234
rect 20806 5182 20858 5234
rect 20858 5182 20860 5234
rect 20804 5180 20860 5182
rect 21980 7442 21982 7476
rect 21982 7442 22034 7476
rect 22034 7442 22036 7476
rect 21980 7420 22036 7442
rect 22652 8876 22708 8932
rect 24220 10108 24276 10164
rect 23940 8818 23996 8820
rect 23940 8766 23942 8818
rect 23942 8766 23994 8818
rect 23994 8766 23996 8818
rect 23940 8764 23996 8766
rect 23772 8540 23828 8596
rect 24444 9660 24500 9716
rect 24220 9548 24276 9604
rect 24500 9212 24556 9268
rect 23100 7644 23156 7700
rect 23324 8204 23380 8260
rect 23324 7756 23380 7812
rect 22204 5852 22260 5908
rect 21644 5180 21700 5236
rect 20020 4956 20076 5012
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 20300 4172 20356 4228
rect 19180 3500 19236 3556
rect 19516 3612 19572 3668
rect 18172 3388 18228 3444
rect 21868 4844 21924 4900
rect 21980 4396 22036 4452
rect 21868 4284 21924 4340
rect 21980 4060 22036 4116
rect 21532 3517 21588 3556
rect 21532 3500 21534 3517
rect 21534 3500 21586 3517
rect 21586 3500 21588 3517
rect 22316 4338 22372 4340
rect 22316 4286 22318 4338
rect 22318 4286 22370 4338
rect 22370 4286 22372 4338
rect 22316 4284 22372 4286
rect 22428 3778 22484 3780
rect 22428 3726 22430 3778
rect 22430 3726 22482 3778
rect 22482 3726 22484 3778
rect 22428 3724 22484 3726
rect 23772 7698 23828 7700
rect 23772 7646 23774 7698
rect 23774 7646 23826 7698
rect 23826 7646 23828 7698
rect 23772 7644 23828 7646
rect 24108 7474 24164 7476
rect 24108 7422 24110 7474
rect 24110 7422 24162 7474
rect 24162 7422 24164 7474
rect 24108 7420 24164 7422
rect 24668 8428 24724 8484
rect 25116 9884 25172 9940
rect 25228 9436 25284 9492
rect 25452 12572 25508 12628
rect 25676 13020 25732 13076
rect 26124 14924 26180 14980
rect 25956 13020 26012 13076
rect 26012 12572 26068 12628
rect 26236 14418 26292 14420
rect 26236 14366 26238 14418
rect 26238 14366 26290 14418
rect 26290 14366 26292 14418
rect 26236 14364 26292 14366
rect 25676 12178 25732 12180
rect 25676 12126 25678 12178
rect 25678 12126 25730 12178
rect 25730 12126 25732 12178
rect 25676 12124 25732 12126
rect 25564 11452 25620 11508
rect 25452 10834 25508 10836
rect 25452 10782 25454 10834
rect 25454 10782 25506 10834
rect 25506 10782 25508 10834
rect 25452 10780 25508 10782
rect 25452 9884 25508 9940
rect 25564 9772 25620 9828
rect 25676 9996 25732 10052
rect 25340 9212 25396 9268
rect 25228 8876 25284 8932
rect 25396 8930 25452 8932
rect 25396 8878 25398 8930
rect 25398 8878 25450 8930
rect 25450 8878 25452 8930
rect 25396 8876 25452 8878
rect 25452 8428 25508 8484
rect 25788 9602 25844 9604
rect 25788 9550 25790 9602
rect 25790 9550 25842 9602
rect 25842 9550 25844 9602
rect 25788 9548 25844 9550
rect 25676 8988 25732 9044
rect 26124 11676 26180 11732
rect 26348 13746 26404 13748
rect 26348 13694 26350 13746
rect 26350 13694 26402 13746
rect 26402 13694 26404 13746
rect 26348 13692 26404 13694
rect 26684 16268 26740 16324
rect 27188 17666 27244 17668
rect 27188 17614 27190 17666
rect 27190 17614 27242 17666
rect 27242 17614 27244 17666
rect 27188 17612 27244 17614
rect 26908 17388 26964 17444
rect 27244 17388 27300 17444
rect 26796 16044 26852 16100
rect 26908 16828 26964 16884
rect 26572 15596 26628 15652
rect 26572 15260 26628 15316
rect 27580 17164 27636 17220
rect 28028 18172 28084 18228
rect 28588 18172 28644 18228
rect 28812 18172 28868 18228
rect 29036 17836 29092 17892
rect 29260 18284 29316 18340
rect 28140 17724 28196 17780
rect 28588 17724 28644 17780
rect 28140 17388 28196 17444
rect 28308 17276 28364 17332
rect 28028 16380 28084 16436
rect 28140 17164 28196 17220
rect 28476 17052 28532 17108
rect 29820 18338 29876 18340
rect 29820 18286 29822 18338
rect 29822 18286 29874 18338
rect 29874 18286 29876 18338
rect 29820 18284 29876 18286
rect 29484 18060 29540 18116
rect 29708 17948 29764 18004
rect 27468 15820 27524 15876
rect 27916 15874 27972 15876
rect 27916 15822 27918 15874
rect 27918 15822 27970 15874
rect 27970 15822 27972 15874
rect 27916 15820 27972 15822
rect 27132 14924 27188 14980
rect 27244 14700 27300 14756
rect 27468 14588 27524 14644
rect 26684 14530 26740 14532
rect 26684 14478 26686 14530
rect 26686 14478 26738 14530
rect 26738 14478 26740 14530
rect 26684 14476 26740 14478
rect 27020 14140 27076 14196
rect 26684 14028 26740 14084
rect 26572 13916 26628 13972
rect 26572 13692 26628 13748
rect 26684 13804 26740 13860
rect 26796 13580 26852 13636
rect 27020 13804 27076 13860
rect 27412 13804 27468 13860
rect 27356 13634 27412 13636
rect 27356 13582 27358 13634
rect 27358 13582 27410 13634
rect 27410 13582 27412 13634
rect 27356 13580 27412 13582
rect 28700 17276 28756 17332
rect 29428 17106 29484 17108
rect 29428 17054 29430 17106
rect 29430 17054 29482 17106
rect 29482 17054 29484 17106
rect 29428 17052 29484 17054
rect 31052 23826 31108 23828
rect 31052 23774 31054 23826
rect 31054 23774 31106 23826
rect 31106 23774 31108 23826
rect 31052 23772 31108 23774
rect 31612 23548 31668 23604
rect 30940 23324 30996 23380
rect 31052 22764 31108 22820
rect 31612 23324 31668 23380
rect 31836 23884 31892 23940
rect 31948 23548 32004 23604
rect 32060 23324 32116 23380
rect 33012 28642 33068 28644
rect 33012 28590 33014 28642
rect 33014 28590 33066 28642
rect 33066 28590 33068 28642
rect 33012 28588 33068 28590
rect 32956 26962 33012 26964
rect 32956 26910 32958 26962
rect 32958 26910 33010 26962
rect 33010 26910 33012 26962
rect 32956 26908 33012 26910
rect 33964 32732 34020 32788
rect 35364 32844 35420 32900
rect 36316 33294 36318 33346
rect 36318 33294 36370 33346
rect 36370 33294 36372 33346
rect 36316 33292 36372 33294
rect 37100 33234 37156 33236
rect 37100 33182 37102 33234
rect 37102 33182 37154 33234
rect 37154 33182 37156 33234
rect 37100 33180 37156 33182
rect 35868 33068 35924 33124
rect 35868 32732 35924 32788
rect 37100 32732 37156 32788
rect 36204 32620 36260 32676
rect 35532 32396 35588 32452
rect 36092 32396 36148 32452
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 31778 35252 31780
rect 35196 31726 35198 31778
rect 35198 31726 35250 31778
rect 35250 31726 35252 31778
rect 35196 31724 35252 31726
rect 33944 31164 34000 31220
rect 33740 29820 33796 29876
rect 36316 31836 36372 31892
rect 34188 30994 34244 30996
rect 34188 30942 34190 30994
rect 34190 30942 34242 30994
rect 34242 30942 34244 30994
rect 34188 30940 34244 30942
rect 35512 30994 35568 30996
rect 35512 30942 35514 30994
rect 35514 30942 35566 30994
rect 35566 30942 35568 30994
rect 35512 30940 35568 30942
rect 35196 30602 35252 30604
rect 34748 30492 34804 30548
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 34076 29708 34132 29764
rect 33740 29426 33796 29428
rect 33740 29374 33742 29426
rect 33742 29374 33794 29426
rect 33794 29374 33796 29426
rect 33740 29372 33796 29374
rect 33460 29148 33516 29204
rect 33404 28812 33460 28868
rect 33404 28588 33460 28644
rect 33628 28476 33684 28532
rect 33740 28028 33796 28084
rect 35312 30172 35368 30212
rect 35312 30156 35314 30172
rect 35314 30156 35366 30172
rect 35366 30156 35368 30172
rect 35812 30210 35868 30212
rect 35812 30158 35814 30210
rect 35814 30158 35866 30210
rect 35866 30158 35868 30210
rect 35812 30156 35868 30158
rect 36204 30828 36260 30884
rect 36316 30604 36372 30660
rect 37772 33068 37828 33124
rect 37660 32956 37716 33012
rect 37436 32786 37492 32788
rect 37436 32734 37438 32786
rect 37438 32734 37490 32786
rect 37490 32734 37492 32786
rect 37436 32732 37492 32734
rect 37324 31948 37380 32004
rect 36838 31052 36894 31108
rect 36540 30994 36596 30996
rect 36540 30942 36542 30994
rect 36542 30942 36594 30994
rect 36594 30942 36596 30994
rect 36540 30940 36596 30942
rect 36428 30156 36484 30212
rect 36540 30044 36596 30100
rect 34860 29538 34916 29540
rect 34860 29486 34862 29538
rect 34862 29486 34914 29538
rect 34914 29486 34916 29538
rect 34860 29484 34916 29486
rect 37100 29932 37156 29988
rect 36652 29708 36708 29764
rect 34748 28812 34804 28868
rect 34972 29260 35028 29316
rect 34504 28642 34560 28644
rect 34504 28590 34506 28642
rect 34506 28590 34558 28642
rect 34558 28590 34560 28642
rect 34504 28588 34560 28590
rect 34748 28642 34804 28644
rect 34748 28590 34750 28642
rect 34750 28590 34802 28642
rect 34802 28590 34804 28642
rect 34748 28588 34804 28590
rect 35476 29314 35532 29316
rect 35476 29262 35478 29314
rect 35478 29262 35530 29314
rect 35530 29262 35532 29314
rect 35476 29260 35532 29262
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 36092 29426 36148 29428
rect 36092 29374 36094 29426
rect 36094 29374 36146 29426
rect 36146 29374 36148 29426
rect 36092 29372 36148 29374
rect 37192 29484 37248 29540
rect 37548 29484 37604 29540
rect 37324 29372 37380 29428
rect 37156 29036 37212 29092
rect 36316 28866 36372 28868
rect 36316 28814 36318 28866
rect 36318 28814 36370 28866
rect 36370 28814 36372 28866
rect 36316 28812 36372 28814
rect 37156 28754 37212 28756
rect 37156 28702 37158 28754
rect 37158 28702 37210 28754
rect 37210 28702 37212 28754
rect 37156 28700 37212 28702
rect 36072 28642 36128 28644
rect 36072 28590 36074 28642
rect 36074 28590 36126 28642
rect 36126 28590 36128 28642
rect 36072 28588 36128 28590
rect 38668 34412 38724 34468
rect 39452 35868 39508 35924
rect 39228 35420 39284 35476
rect 39004 34300 39060 34356
rect 38668 32844 38724 32900
rect 38556 32732 38612 32788
rect 39732 35698 39788 35700
rect 39732 35646 39734 35698
rect 39734 35646 39786 35698
rect 39786 35646 39788 35698
rect 39732 35644 39788 35646
rect 40236 37436 40292 37492
rect 40572 37436 40628 37492
rect 40348 37212 40404 37268
rect 40124 36540 40180 36596
rect 41580 42812 41636 42868
rect 42252 43036 42308 43092
rect 42700 44828 42756 44884
rect 42980 45778 43036 45780
rect 42980 45726 42982 45778
rect 42982 45726 43034 45778
rect 43034 45726 43036 45778
rect 42980 45724 43036 45726
rect 43260 45388 43316 45444
rect 42812 44492 42868 44548
rect 42700 43372 42756 43428
rect 46284 45890 46340 45892
rect 46284 45838 46286 45890
rect 46286 45838 46338 45890
rect 46338 45838 46340 45890
rect 46284 45836 46340 45838
rect 44604 45276 44660 45332
rect 43260 44380 43316 44436
rect 43764 44268 43820 44324
rect 44268 44322 44324 44324
rect 44268 44270 44270 44322
rect 44270 44270 44322 44322
rect 44322 44270 44324 44322
rect 44268 44268 44324 44270
rect 44100 44098 44156 44100
rect 44100 44046 44102 44098
rect 44102 44046 44154 44098
rect 44154 44046 44156 44098
rect 44100 44044 44156 44046
rect 43036 43820 43092 43876
rect 43484 43538 43540 43540
rect 43484 43486 43486 43538
rect 43486 43486 43538 43538
rect 43538 43486 43540 43538
rect 43484 43484 43540 43486
rect 45388 45106 45444 45108
rect 45388 45054 45390 45106
rect 45390 45054 45442 45106
rect 45442 45054 45444 45106
rect 45388 45052 45444 45054
rect 44940 44268 44996 44324
rect 45612 44546 45668 44548
rect 45612 44494 45614 44546
rect 45614 44494 45666 44546
rect 45666 44494 45668 44546
rect 45612 44492 45668 44494
rect 45052 43650 45108 43652
rect 45052 43598 45054 43650
rect 45054 43598 45106 43650
rect 45106 43598 45108 43650
rect 45052 43596 45108 43598
rect 44604 42924 44660 42980
rect 44940 43484 44996 43540
rect 41804 42028 41860 42084
rect 42700 41916 42756 41972
rect 41468 41171 41524 41188
rect 41468 41132 41470 41171
rect 41470 41132 41522 41171
rect 41522 41132 41524 41171
rect 41804 41020 41860 41076
rect 41916 40348 41972 40404
rect 41524 40012 41580 40068
rect 41356 39788 41412 39844
rect 41356 39618 41412 39620
rect 41356 39566 41358 39618
rect 41358 39566 41410 39618
rect 41410 39566 41412 39618
rect 41356 39564 41412 39566
rect 41692 39340 41748 39396
rect 41692 38780 41748 38836
rect 41132 38668 41188 38724
rect 41916 38668 41972 38724
rect 41244 38556 41300 38612
rect 41692 38220 41748 38276
rect 41580 37660 41636 37716
rect 43484 42476 43540 42532
rect 43484 41916 43540 41972
rect 42196 41186 42252 41188
rect 42196 41134 42198 41186
rect 42198 41134 42250 41186
rect 42250 41134 42252 41186
rect 42196 41132 42252 41134
rect 42476 41186 42532 41188
rect 42476 41134 42478 41186
rect 42478 41134 42530 41186
rect 42530 41134 42532 41186
rect 42476 41132 42532 41134
rect 42588 40908 42644 40964
rect 42924 40796 42980 40852
rect 42756 40684 42812 40740
rect 42252 40460 42308 40516
rect 43372 41074 43428 41076
rect 43372 41022 43374 41074
rect 43374 41022 43426 41074
rect 43426 41022 43428 41074
rect 43372 41020 43428 41022
rect 43708 42588 43764 42644
rect 44156 42812 44212 42868
rect 43988 42700 44044 42756
rect 44492 42252 44548 42308
rect 45052 43372 45108 43428
rect 44492 41804 44548 41860
rect 43596 41356 43652 41412
rect 43932 41580 43988 41636
rect 43596 40908 43652 40964
rect 43932 41148 43988 41188
rect 43932 41132 43934 41148
rect 43934 41132 43986 41148
rect 43986 41132 43988 41148
rect 43820 40796 43876 40852
rect 43484 40572 43540 40628
rect 43652 40684 43708 40740
rect 42476 40402 42532 40404
rect 42476 40350 42478 40402
rect 42478 40350 42530 40402
rect 42530 40350 42532 40402
rect 42476 40348 42532 40350
rect 42140 39452 42196 39508
rect 42140 39228 42196 39284
rect 42252 38892 42308 38948
rect 42364 40012 42420 40068
rect 42700 39340 42756 39396
rect 42588 38668 42644 38724
rect 42084 38332 42140 38388
rect 42364 38220 42420 38276
rect 42140 37660 42196 37716
rect 41580 37266 41636 37268
rect 41580 37214 41582 37266
rect 41582 37214 41634 37266
rect 41634 37214 41636 37266
rect 41580 37212 41636 37214
rect 41356 36988 41412 37044
rect 42028 36988 42084 37044
rect 41524 36706 41580 36708
rect 41524 36654 41526 36706
rect 41526 36654 41578 36706
rect 41578 36654 41580 36706
rect 41524 36652 41580 36654
rect 41132 36447 41188 36484
rect 38892 33628 38948 33684
rect 40068 34130 40124 34132
rect 40068 34078 40070 34130
rect 40070 34078 40122 34130
rect 40122 34078 40124 34130
rect 40068 34076 40124 34078
rect 39116 32956 39172 33012
rect 38892 32562 38948 32564
rect 38892 32510 38894 32562
rect 38894 32510 38946 32562
rect 38946 32510 38948 32562
rect 38892 32508 38948 32510
rect 39172 32562 39228 32564
rect 39172 32510 39174 32562
rect 39174 32510 39226 32562
rect 39226 32510 39228 32562
rect 39172 32508 39228 32510
rect 39004 32396 39060 32452
rect 40012 32844 40068 32900
rect 39900 32732 39956 32788
rect 39788 32396 39844 32452
rect 38556 32172 38612 32228
rect 39676 31836 39732 31892
rect 39452 31164 39508 31220
rect 38332 30882 38388 30884
rect 38332 30830 38334 30882
rect 38334 30830 38386 30882
rect 38386 30830 38388 30882
rect 38332 30828 38388 30830
rect 38332 30604 38388 30660
rect 37772 29932 37828 29988
rect 37660 29148 37716 29204
rect 37660 28924 37716 28980
rect 35868 28364 35924 28420
rect 37436 28364 37492 28420
rect 34972 28028 35028 28084
rect 33908 27692 33964 27748
rect 33796 27468 33852 27524
rect 34524 27356 34580 27412
rect 33796 27020 33852 27076
rect 34188 27132 34244 27188
rect 33180 26572 33236 26628
rect 37324 27858 37380 27860
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35196 27244 35252 27300
rect 35028 27020 35084 27076
rect 35196 26908 35252 26964
rect 33516 26460 33572 26516
rect 33740 26460 33796 26516
rect 33012 26236 33068 26292
rect 33180 25900 33236 25956
rect 33516 25900 33572 25956
rect 33068 25116 33124 25172
rect 32396 24668 32452 24724
rect 32172 23212 32228 23268
rect 32284 23772 32340 23828
rect 33180 24722 33236 24724
rect 33180 24670 33182 24722
rect 33182 24670 33234 24722
rect 33234 24670 33236 24722
rect 33180 24668 33236 24670
rect 33068 24220 33124 24276
rect 33012 23548 33068 23604
rect 32844 23436 32900 23492
rect 32396 23212 32452 23268
rect 32732 23212 32788 23268
rect 32284 23100 32340 23156
rect 32564 23042 32620 23044
rect 32564 22990 32566 23042
rect 32566 22990 32618 23042
rect 32618 22990 32620 23042
rect 32564 22988 32620 22990
rect 31444 22540 31500 22596
rect 31724 22652 31780 22708
rect 32732 22652 32788 22708
rect 30380 19852 30436 19908
rect 30716 19516 30772 19572
rect 30940 20802 30996 20804
rect 30940 20750 30942 20802
rect 30942 20750 30994 20802
rect 30994 20750 30996 20802
rect 30940 20748 30996 20750
rect 31276 20748 31332 20804
rect 32060 22370 32116 22372
rect 32060 22318 32062 22370
rect 32062 22318 32114 22370
rect 32114 22318 32116 22370
rect 32060 22316 32116 22318
rect 32284 22370 32340 22372
rect 32284 22318 32286 22370
rect 32286 22318 32338 22370
rect 32338 22318 32340 22370
rect 32284 22316 32340 22318
rect 33180 23212 33236 23268
rect 33404 23548 33460 23604
rect 34076 26684 34132 26740
rect 35756 27074 35812 27076
rect 34580 26684 34636 26740
rect 35756 27022 35758 27074
rect 35758 27022 35810 27074
rect 35810 27022 35812 27074
rect 35756 27020 35812 27022
rect 35532 26908 35588 26964
rect 35532 26684 35588 26740
rect 34748 25900 34804 25956
rect 34076 25564 34132 25620
rect 33944 25228 34000 25284
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 37324 27806 37326 27858
rect 37326 27806 37378 27858
rect 37378 27806 37380 27858
rect 37324 27804 37380 27806
rect 36764 26684 36820 26740
rect 36092 26460 36148 26516
rect 37212 26460 37268 26516
rect 38948 30492 39004 30548
rect 38500 30210 38556 30212
rect 38500 30158 38502 30210
rect 38502 30158 38554 30210
rect 38554 30158 38556 30210
rect 38500 30156 38556 30158
rect 39452 30492 39508 30548
rect 39340 30268 39396 30324
rect 39228 30210 39284 30212
rect 39228 30158 39230 30210
rect 39230 30158 39282 30210
rect 39282 30158 39284 30210
rect 39228 30156 39284 30158
rect 38780 30044 38836 30100
rect 38556 29708 38612 29764
rect 37996 28924 38052 28980
rect 37548 27580 37604 27636
rect 38332 28924 38388 28980
rect 39060 29596 39116 29652
rect 38668 28924 38724 28980
rect 39228 28812 39284 28868
rect 39620 29148 39676 29204
rect 38444 27858 38500 27860
rect 38444 27806 38446 27858
rect 38446 27806 38498 27858
rect 38498 27806 38500 27858
rect 38444 27804 38500 27806
rect 37996 27580 38052 27636
rect 38388 27186 38444 27188
rect 38388 27134 38390 27186
rect 38390 27134 38442 27186
rect 38442 27134 38444 27186
rect 38388 27132 38444 27134
rect 37884 27020 37940 27076
rect 38892 27244 38948 27300
rect 38556 27020 38612 27076
rect 38780 27132 38836 27188
rect 40236 32732 40292 32788
rect 40460 32396 40516 32452
rect 40236 31612 40292 31668
rect 40404 31052 40460 31108
rect 41132 36428 41134 36447
rect 41134 36428 41186 36447
rect 41186 36428 41188 36447
rect 41804 36454 41860 36484
rect 41804 36428 41806 36454
rect 41806 36428 41858 36454
rect 41858 36428 41860 36454
rect 42252 36876 42308 36932
rect 41020 36316 41076 36372
rect 41692 36316 41748 36372
rect 40796 35756 40852 35812
rect 41468 35698 41524 35700
rect 41468 35646 41470 35698
rect 41470 35646 41522 35698
rect 41522 35646 41524 35698
rect 41468 35644 41524 35646
rect 41132 35474 41188 35476
rect 41132 35422 41134 35474
rect 41134 35422 41186 35474
rect 41186 35422 41188 35474
rect 41132 35420 41188 35422
rect 41804 35980 41860 36036
rect 42812 39116 42868 39172
rect 42812 38780 42868 38836
rect 43036 38892 43092 38948
rect 43372 40460 43428 40516
rect 43372 40124 43428 40180
rect 43932 40348 43988 40404
rect 44380 40348 44436 40404
rect 44492 41356 44548 41412
rect 44828 41132 44884 41188
rect 45052 40908 45108 40964
rect 44604 40348 44660 40404
rect 43484 39900 43540 39956
rect 43932 40124 43988 40180
rect 45276 41746 45332 41748
rect 45276 41694 45278 41746
rect 45278 41694 45330 41746
rect 45330 41694 45332 41746
rect 45276 41692 45332 41694
rect 45836 42978 45892 42980
rect 45836 42926 45838 42978
rect 45838 42926 45890 42978
rect 45890 42926 45892 42978
rect 45836 42924 45892 42926
rect 45724 41804 45780 41860
rect 46172 45164 46228 45220
rect 46788 45388 46844 45444
rect 46396 44380 46452 44436
rect 47516 45388 47572 45444
rect 47180 43820 47236 43876
rect 46396 43596 46452 43652
rect 46060 41804 46116 41860
rect 45276 40572 45332 40628
rect 45388 40908 45444 40964
rect 44828 39900 44884 39956
rect 44044 39228 44100 39284
rect 43876 38834 43932 38836
rect 43876 38782 43878 38834
rect 43878 38782 43930 38834
rect 43930 38782 43932 38834
rect 43876 38780 43932 38782
rect 43372 38556 43428 38612
rect 43708 38556 43764 38612
rect 42700 37772 42756 37828
rect 43484 38220 43540 38276
rect 42924 37436 42980 37492
rect 43372 37660 43428 37716
rect 42588 37042 42644 37044
rect 42588 36990 42590 37042
rect 42590 36990 42642 37042
rect 42642 36990 42644 37042
rect 42588 36988 42644 36990
rect 42476 35922 42532 35924
rect 42476 35870 42478 35922
rect 42478 35870 42530 35922
rect 42530 35870 42532 35922
rect 42476 35868 42532 35870
rect 41692 35420 41748 35476
rect 41132 35026 41188 35028
rect 41132 34974 41134 35026
rect 41134 34974 41186 35026
rect 41186 34974 41188 35026
rect 41132 34972 41188 34974
rect 40908 34860 40964 34916
rect 42588 36540 42644 36596
rect 42140 34972 42196 35028
rect 40796 34130 40852 34132
rect 40796 34078 40798 34130
rect 40798 34078 40850 34130
rect 40850 34078 40852 34130
rect 40796 34076 40852 34078
rect 41132 33628 41188 33684
rect 41244 33516 41300 33572
rect 41020 32732 41076 32788
rect 41468 33852 41524 33908
rect 41356 32732 41412 32788
rect 41916 34886 41972 34916
rect 41916 34860 41918 34886
rect 41918 34860 41970 34886
rect 41970 34860 41972 34886
rect 41804 33516 41860 33572
rect 42420 35196 42476 35252
rect 42420 34018 42476 34020
rect 42420 33966 42422 34018
rect 42422 33966 42474 34018
rect 42474 33966 42476 34018
rect 42420 33964 42476 33966
rect 43036 36876 43092 36932
rect 42868 36594 42924 36596
rect 42868 36542 42870 36594
rect 42870 36542 42922 36594
rect 42922 36542 42924 36594
rect 42868 36540 42924 36542
rect 42588 33852 42644 33908
rect 42812 35868 42868 35924
rect 41804 33346 41860 33348
rect 41804 33294 41806 33346
rect 41806 33294 41858 33346
rect 41858 33294 41860 33346
rect 41804 33292 41860 33294
rect 41692 32732 41748 32788
rect 41748 32562 41804 32564
rect 41748 32510 41750 32562
rect 41750 32510 41802 32562
rect 41802 32510 41804 32562
rect 41748 32508 41804 32510
rect 41244 31948 41300 32004
rect 40684 31612 40740 31668
rect 40572 30604 40628 30660
rect 40236 29932 40292 29988
rect 40236 29596 40292 29652
rect 40572 29372 40628 29428
rect 40236 29148 40292 29204
rect 40124 28812 40180 28868
rect 39956 27634 40012 27636
rect 39956 27582 39958 27634
rect 39958 27582 40010 27634
rect 40010 27582 40012 27634
rect 39956 27580 40012 27582
rect 41244 29148 41300 29204
rect 41020 28588 41076 28644
rect 41132 28924 41188 28980
rect 41244 28700 41300 28756
rect 41020 27804 41076 27860
rect 39340 27244 39396 27300
rect 39228 27132 39284 27188
rect 37884 26796 37940 26852
rect 36988 26178 37044 26180
rect 36988 26126 36990 26178
rect 36990 26126 37042 26178
rect 37042 26126 37044 26178
rect 36988 26124 37044 26126
rect 34860 25452 34916 25508
rect 35644 25506 35700 25508
rect 35644 25454 35646 25506
rect 35646 25454 35698 25506
rect 35698 25454 35700 25506
rect 35644 25452 35700 25454
rect 37212 25282 37268 25284
rect 37212 25230 37214 25282
rect 37214 25230 37266 25282
rect 37266 25230 37268 25282
rect 37212 25228 37268 25230
rect 35644 25004 35700 25060
rect 33516 23436 33572 23492
rect 34300 23548 34356 23604
rect 33460 22594 33516 22596
rect 33460 22542 33462 22594
rect 33462 22542 33514 22594
rect 33514 22542 33516 22594
rect 33460 22540 33516 22542
rect 32060 21532 32116 21588
rect 32060 21308 32116 21364
rect 31724 20860 31780 20916
rect 32396 20914 32452 20916
rect 32396 20862 32398 20914
rect 32398 20862 32450 20914
rect 32450 20862 32452 20914
rect 32396 20860 32452 20862
rect 31220 20300 31276 20356
rect 33516 21756 33572 21812
rect 33236 21586 33292 21588
rect 33236 21534 33238 21586
rect 33238 21534 33290 21586
rect 33290 21534 33292 21586
rect 33236 21532 33292 21534
rect 32060 20300 32116 20356
rect 32060 20076 32116 20132
rect 31836 19964 31892 20020
rect 30044 17724 30100 17780
rect 31052 19516 31108 19572
rect 30716 17836 30772 17892
rect 29652 16492 29708 16548
rect 28140 15484 28196 15540
rect 28140 15260 28196 15316
rect 28364 16268 28420 16324
rect 28532 15932 28588 15988
rect 28700 15708 28756 15764
rect 28532 15314 28588 15316
rect 28532 15262 28534 15314
rect 28534 15262 28586 15314
rect 28586 15262 28588 15314
rect 28532 15260 28588 15262
rect 27692 14924 27748 14980
rect 29148 16044 29204 16100
rect 29820 16098 29876 16100
rect 29820 16046 29822 16098
rect 29822 16046 29874 16098
rect 29874 16046 29876 16098
rect 29820 16044 29876 16046
rect 29148 15484 29204 15540
rect 29372 15314 29428 15316
rect 29372 15262 29374 15314
rect 29374 15262 29426 15314
rect 29426 15262 29428 15314
rect 29372 15260 29428 15262
rect 29652 15202 29708 15204
rect 29652 15150 29654 15202
rect 29654 15150 29706 15202
rect 29706 15150 29708 15202
rect 29652 15148 29708 15150
rect 28924 15036 28980 15092
rect 29932 15820 29988 15876
rect 31724 19346 31780 19348
rect 31724 19294 31726 19346
rect 31726 19294 31778 19346
rect 31778 19294 31780 19346
rect 31724 19292 31780 19294
rect 32732 20076 32788 20132
rect 32284 19852 32340 19908
rect 32060 19292 32116 19348
rect 32396 19292 32452 19348
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 36092 23996 36148 24052
rect 34636 23436 34692 23492
rect 34972 23324 35028 23380
rect 35084 23548 35140 23604
rect 36988 24050 37044 24052
rect 36988 23998 36990 24050
rect 36990 23998 37042 24050
rect 37042 23998 37044 24050
rect 36988 23996 37044 23998
rect 36876 23772 36932 23828
rect 35756 23324 35812 23380
rect 34300 22988 34356 23044
rect 33964 22876 34020 22932
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 33628 20188 33684 20244
rect 33012 20018 33068 20020
rect 33012 19966 33014 20018
rect 33014 19966 33066 20018
rect 33066 19966 33068 20018
rect 33012 19964 33068 19966
rect 33180 19292 33236 19348
rect 32340 18620 32396 18676
rect 32228 18226 32284 18228
rect 32228 18174 32230 18226
rect 32230 18174 32282 18226
rect 32282 18174 32284 18226
rect 32228 18172 32284 18174
rect 31612 18060 31668 18116
rect 33012 18060 33068 18116
rect 33740 21644 33796 21700
rect 34916 22370 34972 22372
rect 34916 22318 34918 22370
rect 34918 22318 34970 22370
rect 34970 22318 34972 22370
rect 34916 22316 34972 22318
rect 35644 22370 35700 22372
rect 35644 22318 35646 22370
rect 35646 22318 35698 22370
rect 35698 22318 35700 22370
rect 35644 22316 35700 22318
rect 35868 22370 35924 22372
rect 35868 22318 35870 22370
rect 35870 22318 35922 22370
rect 35922 22318 35924 22370
rect 35868 22316 35924 22318
rect 34636 22092 34692 22148
rect 34412 21756 34468 21812
rect 34076 21420 34132 21476
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 37100 23923 37156 23940
rect 37100 23884 37102 23923
rect 37102 23884 37154 23923
rect 37154 23884 37156 23923
rect 37660 26684 37716 26740
rect 37548 25228 37604 25284
rect 37660 24668 37716 24724
rect 37772 26012 37828 26068
rect 37436 23772 37492 23828
rect 39564 26796 39620 26852
rect 39228 26684 39284 26740
rect 38780 26236 38836 26292
rect 38892 26348 38948 26404
rect 39116 26290 39172 26292
rect 39116 26238 39118 26290
rect 39118 26238 39170 26290
rect 39170 26238 39172 26290
rect 39116 26236 39172 26238
rect 41132 27692 41188 27748
rect 40348 27046 40404 27076
rect 40348 27020 40350 27046
rect 40350 27020 40402 27046
rect 40402 27020 40404 27046
rect 40068 26684 40124 26740
rect 39844 26348 39900 26404
rect 39508 26178 39564 26180
rect 39508 26126 39510 26178
rect 39510 26126 39562 26178
rect 39562 26126 39564 26178
rect 39508 26124 39564 26126
rect 39564 25900 39620 25956
rect 38668 24892 38724 24948
rect 38780 25228 38836 25284
rect 38332 24722 38388 24724
rect 38332 24670 38334 24722
rect 38334 24670 38386 24722
rect 38386 24670 38388 24722
rect 38332 24668 38388 24670
rect 38220 24162 38276 24164
rect 38220 24110 38222 24162
rect 38222 24110 38274 24162
rect 38274 24110 38276 24162
rect 38220 24108 38276 24110
rect 37884 23660 37940 23716
rect 37772 23436 37828 23492
rect 35980 22092 36036 22148
rect 36876 22092 36932 22148
rect 36092 21756 36148 21812
rect 36540 21756 36596 21812
rect 37436 21644 37492 21700
rect 37212 21420 37268 21476
rect 36764 21196 36820 21252
rect 34132 20578 34188 20580
rect 34132 20526 34134 20578
rect 34134 20526 34186 20578
rect 34186 20526 34188 20578
rect 34132 20524 34188 20526
rect 35084 20412 35140 20468
rect 35532 20018 35588 20020
rect 35532 19966 35534 20018
rect 35534 19966 35586 20018
rect 35586 19966 35588 20018
rect 35532 19964 35588 19966
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 37324 21308 37380 21364
rect 36540 20524 36596 20580
rect 36316 20018 36372 20020
rect 36316 19966 36318 20018
rect 36318 19966 36370 20018
rect 36370 19966 36372 20018
rect 36316 19964 36372 19966
rect 36876 20130 36932 20132
rect 36876 20078 36878 20130
rect 36878 20078 36930 20130
rect 36930 20078 36932 20130
rect 36876 20076 36932 20078
rect 37212 20018 37268 20020
rect 37212 19966 37214 20018
rect 37214 19966 37266 20018
rect 37266 19966 37268 20018
rect 37212 19964 37268 19966
rect 33404 18172 33460 18228
rect 33292 17948 33348 18004
rect 32172 17836 32228 17892
rect 32620 17836 32676 17892
rect 31164 17276 31220 17332
rect 31052 17164 31108 17220
rect 34412 17388 34468 17444
rect 33628 17164 33684 17220
rect 31836 16770 31892 16772
rect 31836 16718 31838 16770
rect 31838 16718 31890 16770
rect 31890 16718 31892 16770
rect 31836 16716 31892 16718
rect 33012 16882 33068 16884
rect 33012 16830 33014 16882
rect 33014 16830 33066 16882
rect 33066 16830 33068 16882
rect 33012 16828 33068 16830
rect 33628 16828 33684 16884
rect 33740 16716 33796 16772
rect 30604 16156 30660 16212
rect 30940 16156 30996 16212
rect 30212 16098 30268 16100
rect 30212 16046 30214 16098
rect 30214 16046 30266 16098
rect 30266 16046 30268 16098
rect 30212 16044 30268 16046
rect 30044 15708 30100 15764
rect 29932 15260 29988 15316
rect 30044 15372 30100 15428
rect 29820 15036 29876 15092
rect 28812 14924 28868 14980
rect 28364 14588 28420 14644
rect 27804 14530 27860 14532
rect 27804 14478 27806 14530
rect 27806 14478 27858 14530
rect 27858 14478 27860 14530
rect 27804 14476 27860 14478
rect 28140 14418 28196 14420
rect 28140 14366 28142 14418
rect 28142 14366 28194 14418
rect 28194 14366 28196 14418
rect 28140 14364 28196 14366
rect 28140 14140 28196 14196
rect 27692 13356 27748 13412
rect 27076 13186 27132 13188
rect 27076 13134 27078 13186
rect 27078 13134 27130 13186
rect 27130 13134 27132 13186
rect 27076 13132 27132 13134
rect 28252 14028 28308 14084
rect 28252 13580 28308 13636
rect 27804 13132 27860 13188
rect 28868 14252 28924 14308
rect 28364 13468 28420 13524
rect 26236 11340 26292 11396
rect 26348 11452 26404 11508
rect 26684 11564 26740 11620
rect 27020 11564 27076 11620
rect 26572 11340 26628 11396
rect 26460 11116 26516 11172
rect 26684 10780 26740 10836
rect 26796 11340 26852 11396
rect 26516 10556 26572 10612
rect 27020 11394 27076 11396
rect 27020 11342 27022 11394
rect 27022 11342 27074 11394
rect 27074 11342 27076 11394
rect 27020 11340 27076 11342
rect 27356 11004 27412 11060
rect 27076 10386 27132 10388
rect 27076 10334 27078 10386
rect 27078 10334 27130 10386
rect 27130 10334 27132 10386
rect 27076 10332 27132 10334
rect 28364 12236 28420 12292
rect 28700 13356 28756 13412
rect 27580 11452 27636 11508
rect 27636 11004 27692 11060
rect 27636 10610 27692 10612
rect 27636 10558 27638 10610
rect 27638 10558 27690 10610
rect 27690 10558 27692 10610
rect 27636 10556 27692 10558
rect 28476 12178 28532 12180
rect 28476 12126 28478 12178
rect 28478 12126 28530 12178
rect 28530 12126 28532 12178
rect 28476 12124 28532 12126
rect 29316 14924 29372 14980
rect 29148 14530 29204 14532
rect 29148 14478 29150 14530
rect 29150 14478 29202 14530
rect 29202 14478 29204 14530
rect 29148 14476 29204 14478
rect 29316 14364 29372 14420
rect 29484 14140 29540 14196
rect 29876 14418 29932 14420
rect 29876 14366 29878 14418
rect 29878 14366 29930 14418
rect 29930 14366 29932 14418
rect 29876 14364 29932 14366
rect 29596 14028 29652 14084
rect 29820 13356 29876 13412
rect 30380 14476 30436 14532
rect 30492 15036 30548 15092
rect 30156 13916 30212 13972
rect 31164 16156 31220 16212
rect 30940 14252 30996 14308
rect 31836 15260 31892 15316
rect 30604 14140 30660 14196
rect 30268 13746 30324 13748
rect 30268 13694 30270 13746
rect 30270 13694 30322 13746
rect 30322 13694 30324 13746
rect 30268 13692 30324 13694
rect 30436 13916 30492 13972
rect 30716 14028 30772 14084
rect 31276 13916 31332 13972
rect 31164 13580 31220 13636
rect 30436 13468 30492 13524
rect 30996 13522 31052 13524
rect 30996 13470 30998 13522
rect 30998 13470 31050 13522
rect 31050 13470 31052 13522
rect 30996 13468 31052 13470
rect 30156 13356 30212 13412
rect 29596 12796 29652 12852
rect 29036 12684 29092 12740
rect 28028 11116 28084 11172
rect 26908 9772 26964 9828
rect 27580 10332 27636 10388
rect 26516 9660 26572 9716
rect 26012 9548 26068 9604
rect 26964 9436 27020 9492
rect 25676 8652 25732 8708
rect 26012 8764 26068 8820
rect 25900 8258 25956 8260
rect 25900 8206 25902 8258
rect 25902 8206 25954 8258
rect 25954 8206 25956 8258
rect 25900 8204 25956 8206
rect 25340 7756 25396 7812
rect 23324 6662 23380 6692
rect 23324 6636 23326 6662
rect 23326 6636 23378 6662
rect 23378 6636 23380 6662
rect 23548 6690 23604 6692
rect 23548 6638 23550 6690
rect 23550 6638 23602 6690
rect 23602 6638 23604 6690
rect 26180 8146 26236 8148
rect 26180 8094 26182 8146
rect 26182 8094 26234 8146
rect 26234 8094 26236 8146
rect 26180 8092 26236 8094
rect 26628 9042 26684 9044
rect 26628 8990 26630 9042
rect 26630 8990 26682 9042
rect 26682 8990 26684 9042
rect 26628 8988 26684 8990
rect 27244 9324 27300 9380
rect 27356 9826 27412 9828
rect 27356 9774 27358 9826
rect 27358 9774 27410 9826
rect 27410 9774 27412 9826
rect 27356 9772 27412 9774
rect 26796 8764 26852 8820
rect 26460 8428 26516 8484
rect 26684 8316 26740 8372
rect 27020 8258 27076 8260
rect 27020 8206 27022 8258
rect 27022 8206 27074 8258
rect 27074 8206 27076 8258
rect 27020 8204 27076 8206
rect 26460 8092 26516 8148
rect 25900 7420 25956 7476
rect 25676 7084 25732 7140
rect 23548 6636 23604 6638
rect 22652 5906 22708 5908
rect 22652 5854 22654 5906
rect 22654 5854 22706 5906
rect 22706 5854 22708 5906
rect 22652 5852 22708 5854
rect 22652 4338 22708 4340
rect 22652 4286 22654 4338
rect 22654 4286 22706 4338
rect 22706 4286 22708 4338
rect 22652 4284 22708 4286
rect 23772 5852 23828 5908
rect 22876 5404 22932 5460
rect 23100 5122 23156 5124
rect 23100 5070 23102 5122
rect 23102 5070 23154 5122
rect 23154 5070 23156 5122
rect 23100 5068 23156 5070
rect 23436 5180 23492 5236
rect 23212 4956 23268 5012
rect 23156 4450 23212 4452
rect 23156 4398 23158 4450
rect 23158 4398 23210 4450
rect 23210 4398 23212 4450
rect 23156 4396 23212 4398
rect 22764 4060 22820 4116
rect 22876 3948 22932 4004
rect 23996 4844 24052 4900
rect 23772 3948 23828 4004
rect 23436 3836 23492 3892
rect 23996 3836 24052 3892
rect 22540 3612 22596 3668
rect 22764 3612 22820 3668
rect 24276 6636 24332 6692
rect 25452 6914 25508 6916
rect 25452 6862 25454 6914
rect 25454 6862 25506 6914
rect 25506 6862 25508 6914
rect 25452 6860 25508 6862
rect 24892 6524 24948 6580
rect 25060 6524 25116 6580
rect 25116 6076 25172 6132
rect 24556 5852 24612 5908
rect 24444 5628 24500 5684
rect 24220 4396 24276 4452
rect 25228 5906 25284 5908
rect 25228 5854 25230 5906
rect 25230 5854 25282 5906
rect 25282 5854 25284 5906
rect 25228 5852 25284 5854
rect 26012 6524 26068 6580
rect 25900 6412 25956 6468
rect 25452 6076 25508 6132
rect 25526 5891 25528 5908
rect 25528 5891 25580 5908
rect 25580 5891 25582 5908
rect 25526 5852 25582 5891
rect 25900 5682 25956 5684
rect 25900 5630 25902 5682
rect 25902 5630 25954 5682
rect 25954 5630 25956 5682
rect 25900 5628 25956 5630
rect 25116 5404 25172 5460
rect 24444 5068 24500 5124
rect 24332 4284 24388 4340
rect 26348 6412 26404 6468
rect 26124 5852 26180 5908
rect 25900 4844 25956 4900
rect 26012 4956 26068 5012
rect 25228 4450 25284 4452
rect 25228 4398 25230 4450
rect 25230 4398 25282 4450
rect 25282 4398 25284 4450
rect 25228 4396 25284 4398
rect 25564 4322 25566 4340
rect 25566 4322 25618 4340
rect 25618 4322 25620 4340
rect 25564 4284 25620 4322
rect 25452 3836 25508 3892
rect 24108 3612 24164 3668
rect 24836 3666 24892 3668
rect 24836 3614 24838 3666
rect 24838 3614 24890 3666
rect 24890 3614 24892 3666
rect 24836 3612 24892 3614
rect 25172 3554 25228 3556
rect 25172 3502 25174 3554
rect 25174 3502 25226 3554
rect 25226 3502 25228 3554
rect 25172 3500 25228 3502
rect 21084 3388 21140 3444
rect 19796 3276 19852 3332
rect 26012 3554 26068 3556
rect 26012 3502 26014 3554
rect 26014 3502 26066 3554
rect 26066 3502 26068 3554
rect 26012 3500 26068 3502
rect 26236 4732 26292 4788
rect 26740 7980 26796 8036
rect 26908 7532 26964 7588
rect 28364 11004 28420 11060
rect 27692 7532 27748 7588
rect 26852 6466 26908 6468
rect 26852 6414 26854 6466
rect 26854 6414 26906 6466
rect 26906 6414 26908 6466
rect 26852 6412 26908 6414
rect 26460 5068 26516 5124
rect 27580 6690 27636 6692
rect 27580 6638 27582 6690
rect 27582 6638 27634 6690
rect 27634 6638 27636 6690
rect 27580 6636 27636 6638
rect 28252 9548 28308 9604
rect 27972 8034 28028 8036
rect 27972 7982 27974 8034
rect 27974 7982 28026 8034
rect 28026 7982 28028 8034
rect 27972 7980 28028 7982
rect 28812 9884 28868 9940
rect 29988 12348 30044 12404
rect 29820 12124 29876 12180
rect 30268 13132 30324 13188
rect 30548 13020 30604 13076
rect 30716 12850 30772 12852
rect 30716 12798 30718 12850
rect 30718 12798 30770 12850
rect 30770 12798 30772 12850
rect 30716 12796 30772 12798
rect 30268 12572 30324 12628
rect 30940 12572 30996 12628
rect 30156 12124 30212 12180
rect 30380 12066 30436 12068
rect 30380 12014 30382 12066
rect 30382 12014 30434 12066
rect 30434 12014 30436 12066
rect 30380 12012 30436 12014
rect 30604 11900 30660 11956
rect 29652 11170 29708 11172
rect 29652 11118 29654 11170
rect 29654 11118 29706 11170
rect 29706 11118 29708 11170
rect 29652 11116 29708 11118
rect 30100 11282 30156 11284
rect 30100 11230 30102 11282
rect 30102 11230 30154 11282
rect 30154 11230 30156 11282
rect 30100 11228 30156 11230
rect 30268 11116 30324 11172
rect 29988 10332 30044 10388
rect 29820 9938 29876 9940
rect 29820 9886 29822 9938
rect 29822 9886 29874 9938
rect 29874 9886 29876 9938
rect 29820 9884 29876 9886
rect 28364 8652 28420 8708
rect 28812 7980 28868 8036
rect 28812 7420 28868 7476
rect 28924 8652 28980 8708
rect 27916 6076 27972 6132
rect 28588 6188 28644 6244
rect 27916 5292 27972 5348
rect 28812 5292 28868 5348
rect 26348 4060 26404 4116
rect 26348 3724 26404 3780
rect 26236 3612 26292 3668
rect 28252 4844 28308 4900
rect 28812 5068 28868 5124
rect 28700 4396 28756 4452
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 29932 8988 29988 9044
rect 29484 8034 29540 8036
rect 29484 7982 29486 8034
rect 29486 7982 29538 8034
rect 29538 7982 29540 8034
rect 29484 7980 29540 7982
rect 29596 7196 29652 7252
rect 29204 6636 29260 6692
rect 29764 6690 29820 6692
rect 29764 6638 29766 6690
rect 29766 6638 29818 6690
rect 29818 6638 29820 6690
rect 29764 6636 29820 6638
rect 29148 6188 29204 6244
rect 30716 11116 30772 11172
rect 30716 10668 30772 10724
rect 31106 12178 31162 12180
rect 31106 12126 31108 12178
rect 31108 12126 31160 12178
rect 31160 12126 31162 12178
rect 31106 12124 31162 12126
rect 31388 13746 31444 13748
rect 31388 13694 31390 13746
rect 31390 13694 31442 13746
rect 31442 13694 31444 13746
rect 31388 13692 31444 13694
rect 34188 16716 34244 16772
rect 33572 16098 33628 16100
rect 33572 16046 33574 16098
rect 33574 16046 33626 16098
rect 33626 16046 33628 16098
rect 33572 16044 33628 16046
rect 34860 18338 34916 18340
rect 34860 18286 34862 18338
rect 34862 18286 34914 18338
rect 34914 18286 34916 18338
rect 34860 18284 34916 18286
rect 35308 18450 35364 18452
rect 35308 18398 35310 18450
rect 35310 18398 35362 18450
rect 35362 18398 35364 18450
rect 35308 18396 35364 18398
rect 36316 18396 36372 18452
rect 36092 18338 36148 18340
rect 36092 18286 36094 18338
rect 36094 18286 36146 18338
rect 36146 18286 36148 18338
rect 36092 18284 36148 18286
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 36092 18060 36148 18116
rect 35812 17666 35868 17668
rect 35812 17614 35814 17666
rect 35814 17614 35866 17666
rect 35866 17614 35868 17666
rect 35812 17612 35868 17614
rect 34860 17388 34916 17444
rect 37212 17724 37268 17780
rect 37212 17276 37268 17332
rect 35980 17164 36036 17220
rect 36876 17164 36932 17220
rect 33964 15932 34020 15988
rect 32172 15148 32228 15204
rect 32732 13692 32788 13748
rect 31948 13580 32004 13636
rect 31724 13132 31780 13188
rect 30940 11228 30996 11284
rect 30716 10498 30772 10500
rect 30716 10446 30718 10498
rect 30718 10446 30770 10498
rect 30770 10446 30772 10498
rect 30716 10444 30772 10446
rect 30548 10108 30604 10164
rect 30940 10108 30996 10164
rect 30492 9324 30548 9380
rect 30492 8540 30548 8596
rect 30044 7980 30100 8036
rect 31388 12796 31444 12852
rect 31668 12962 31724 12964
rect 31668 12910 31670 12962
rect 31670 12910 31722 12962
rect 31722 12910 31724 12962
rect 31668 12908 31724 12910
rect 34972 16882 35028 16884
rect 34972 16830 34974 16882
rect 34974 16830 35026 16882
rect 35026 16830 35028 16882
rect 34972 16828 35028 16830
rect 34860 16716 34916 16772
rect 35644 16716 35700 16772
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 34524 16268 34580 16324
rect 33292 15596 33348 15652
rect 33180 14530 33236 14532
rect 33180 14478 33182 14530
rect 33182 14478 33234 14530
rect 33234 14478 33236 14530
rect 33180 14476 33236 14478
rect 33068 13692 33124 13748
rect 32060 12962 32116 12964
rect 32060 12910 32062 12962
rect 32062 12910 32114 12962
rect 32114 12910 32116 12962
rect 32060 12908 32116 12910
rect 31612 12460 31668 12516
rect 32340 12572 32396 12628
rect 31500 12348 31556 12404
rect 33740 15314 33796 15316
rect 33740 15262 33742 15314
rect 33742 15262 33794 15314
rect 33794 15262 33796 15314
rect 33740 15260 33796 15262
rect 33628 14530 33684 14532
rect 33628 14478 33630 14530
rect 33630 14478 33682 14530
rect 33682 14478 33684 14530
rect 33628 14476 33684 14478
rect 33740 13634 33796 13636
rect 33740 13582 33742 13634
rect 33742 13582 33794 13634
rect 33794 13582 33796 13634
rect 33740 13580 33796 13582
rect 33572 12908 33628 12964
rect 33740 12684 33796 12740
rect 33292 12572 33348 12628
rect 34860 15260 34916 15316
rect 36484 16210 36540 16212
rect 36484 16158 36486 16210
rect 36486 16158 36538 16210
rect 36538 16158 36540 16210
rect 36484 16156 36540 16158
rect 35644 15820 35700 15876
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 33964 14476 34020 14532
rect 34412 13916 34468 13972
rect 38332 23548 38388 23604
rect 38892 24946 38948 24948
rect 38892 24894 38894 24946
rect 38894 24894 38946 24946
rect 38946 24894 38948 24946
rect 38892 24892 38948 24894
rect 40348 26236 40404 26292
rect 40964 26796 41020 26852
rect 40460 25900 40516 25956
rect 40684 26236 40740 26292
rect 42700 33404 42756 33460
rect 43372 36428 43428 36484
rect 43036 35756 43092 35812
rect 43036 35474 43092 35476
rect 43036 35422 43038 35474
rect 43038 35422 43090 35474
rect 43090 35422 43092 35474
rect 43036 35420 43092 35422
rect 43148 34972 43204 35028
rect 42924 34412 42980 34468
rect 42812 33292 42868 33348
rect 41916 31948 41972 32004
rect 41692 31836 41748 31892
rect 41692 30156 41748 30212
rect 43148 32956 43204 33012
rect 43932 38556 43988 38612
rect 43820 38108 43876 38164
rect 43596 37772 43652 37828
rect 43428 34914 43484 34916
rect 43428 34862 43430 34914
rect 43430 34862 43482 34914
rect 43482 34862 43484 34914
rect 43428 34860 43484 34862
rect 43372 34636 43428 34692
rect 43484 33292 43540 33348
rect 43820 37100 43876 37156
rect 43932 37212 43988 37268
rect 43708 36204 43764 36260
rect 44380 38668 44436 38724
rect 44156 38220 44212 38276
rect 44212 38050 44268 38052
rect 44212 37998 44214 38050
rect 44214 37998 44266 38050
rect 44266 37998 44268 38050
rect 44212 37996 44268 37998
rect 44604 39116 44660 39172
rect 44716 38892 44772 38948
rect 44492 37772 44548 37828
rect 44940 39394 44996 39396
rect 44940 39342 44942 39394
rect 44942 39342 44994 39394
rect 44994 39342 44996 39394
rect 44940 39340 44996 39342
rect 45052 39228 45108 39284
rect 44940 39116 44996 39172
rect 45724 41020 45780 41076
rect 45724 40460 45780 40516
rect 45836 40684 45892 40740
rect 45612 40402 45668 40404
rect 45612 40350 45614 40402
rect 45614 40350 45666 40402
rect 45666 40350 45668 40402
rect 45612 40348 45668 40350
rect 46060 40908 46116 40964
rect 47180 43148 47236 43204
rect 47404 43820 47460 43876
rect 47404 42700 47460 42756
rect 46732 41858 46788 41860
rect 46732 41806 46734 41858
rect 46734 41806 46786 41858
rect 46786 41806 46788 41858
rect 46732 41804 46788 41806
rect 46284 40572 46340 40628
rect 46172 40460 46228 40516
rect 46396 40514 46452 40516
rect 46396 40462 46398 40514
rect 46398 40462 46450 40514
rect 46450 40462 46452 40514
rect 46396 40460 46452 40462
rect 47516 41916 47572 41972
rect 47404 40684 47460 40740
rect 47516 41020 47572 41076
rect 46620 40460 46676 40516
rect 46508 40402 46564 40404
rect 46508 40350 46510 40402
rect 46510 40350 46562 40402
rect 46562 40350 46564 40402
rect 46508 40348 46564 40350
rect 47124 40402 47180 40404
rect 47124 40350 47126 40402
rect 47126 40350 47178 40402
rect 47178 40350 47180 40402
rect 47124 40348 47180 40350
rect 45500 39564 45556 39620
rect 45164 39116 45220 39172
rect 45388 38668 45444 38724
rect 44156 37154 44212 37156
rect 44156 37102 44158 37154
rect 44158 37102 44210 37154
rect 44210 37102 44212 37154
rect 44156 37100 44212 37102
rect 43708 35586 43764 35588
rect 43708 35534 43710 35586
rect 43710 35534 43762 35586
rect 43762 35534 43764 35586
rect 43708 35532 43764 35534
rect 43708 34914 43764 34916
rect 43708 34862 43710 34914
rect 43710 34862 43762 34914
rect 43762 34862 43764 34914
rect 43708 34860 43764 34862
rect 44716 36482 44772 36484
rect 44716 36430 44718 36482
rect 44718 36430 44770 36482
rect 44770 36430 44772 36482
rect 44716 36428 44772 36430
rect 44604 36204 44660 36260
rect 44436 35810 44492 35812
rect 44436 35758 44438 35810
rect 44438 35758 44490 35810
rect 44490 35758 44492 35810
rect 44436 35756 44492 35758
rect 44044 34860 44100 34916
rect 44044 34690 44100 34692
rect 44044 34638 44046 34690
rect 44046 34638 44098 34690
rect 44098 34638 44100 34690
rect 44044 34636 44100 34638
rect 43932 33516 43988 33572
rect 43596 33180 43652 33236
rect 43372 32732 43428 32788
rect 44156 33346 44212 33348
rect 44156 33294 44158 33346
rect 44158 33294 44210 33346
rect 44210 33294 44212 33346
rect 44156 33292 44212 33294
rect 44156 33068 44212 33124
rect 43932 32396 43988 32452
rect 42364 31724 42420 31780
rect 43036 31743 43092 31780
rect 43036 31724 43038 31743
rect 43038 31724 43090 31743
rect 43090 31724 43092 31743
rect 43596 32172 43652 32228
rect 43876 32002 43932 32004
rect 43876 31950 43878 32002
rect 43878 31950 43930 32002
rect 43930 31950 43932 32002
rect 43876 31948 43932 31950
rect 44044 31724 44100 31780
rect 42252 31164 42308 31220
rect 42700 31276 42756 31332
rect 42588 30604 42644 30660
rect 42196 29650 42252 29652
rect 42196 29598 42198 29650
rect 42198 29598 42250 29650
rect 42250 29598 42252 29650
rect 42196 29596 42252 29598
rect 41804 29372 41860 29428
rect 42476 28812 42532 28868
rect 42028 28364 42084 28420
rect 41804 27858 41860 27860
rect 41804 27806 41806 27858
rect 41806 27806 41858 27858
rect 41858 27806 41860 27858
rect 41804 27804 41860 27806
rect 41244 26124 41300 26180
rect 41356 25788 41412 25844
rect 37940 22370 37996 22372
rect 37940 22318 37942 22370
rect 37942 22318 37994 22370
rect 37994 22318 37996 22370
rect 37940 22316 37996 22318
rect 38780 23548 38836 23604
rect 38668 23154 38724 23156
rect 38668 23102 38670 23154
rect 38670 23102 38722 23154
rect 38722 23102 38724 23154
rect 38668 23100 38724 23102
rect 38164 21644 38220 21700
rect 38668 22092 38724 22148
rect 38444 21756 38500 21812
rect 38556 21362 38612 21364
rect 38556 21310 38558 21362
rect 38558 21310 38610 21362
rect 38610 21310 38612 21362
rect 38556 21308 38612 21310
rect 38892 22204 38948 22260
rect 39340 24108 39396 24164
rect 40124 23938 40180 23940
rect 40124 23886 40126 23938
rect 40126 23886 40178 23938
rect 40178 23886 40180 23938
rect 40124 23884 40180 23886
rect 39004 21196 39060 21252
rect 39116 22092 39172 22148
rect 38892 20748 38948 20804
rect 37772 20188 37828 20244
rect 37548 19852 37604 19908
rect 38108 20412 38164 20468
rect 38444 20188 38500 20244
rect 37996 19964 38052 20020
rect 37884 19852 37940 19908
rect 38276 19852 38332 19908
rect 38052 19458 38108 19460
rect 38052 19406 38054 19458
rect 38054 19406 38106 19458
rect 38106 19406 38108 19458
rect 38052 19404 38108 19406
rect 39004 20412 39060 20468
rect 40348 24668 40404 24724
rect 40908 24722 40964 24724
rect 40908 24670 40910 24722
rect 40910 24670 40962 24722
rect 40962 24670 40964 24722
rect 40908 24668 40964 24670
rect 41356 24556 41412 24612
rect 41244 24444 41300 24500
rect 40348 23772 40404 23828
rect 40908 23884 40964 23940
rect 40684 23772 40740 23828
rect 40292 23548 40348 23604
rect 40684 23436 40740 23492
rect 39676 23100 39732 23156
rect 39340 21868 39396 21924
rect 40572 22764 40628 22820
rect 40572 21868 40628 21924
rect 39788 21756 39844 21812
rect 39676 21586 39732 21588
rect 39676 21534 39678 21586
rect 39678 21534 39730 21586
rect 39730 21534 39732 21586
rect 39676 21532 39732 21534
rect 40292 21698 40348 21700
rect 40292 21646 40294 21698
rect 40294 21646 40346 21698
rect 40346 21646 40348 21698
rect 40292 21644 40348 21646
rect 40124 21420 40180 21476
rect 39788 20636 39844 20692
rect 39900 21196 39956 21252
rect 39340 20524 39396 20580
rect 39900 20524 39956 20580
rect 40124 20636 40180 20692
rect 38780 20018 38836 20020
rect 38780 19966 38782 20018
rect 38782 19966 38834 20018
rect 38834 19966 38836 20018
rect 38780 19964 38836 19966
rect 39116 19794 39172 19796
rect 39116 19742 39118 19794
rect 39118 19742 39170 19794
rect 39170 19742 39172 19794
rect 39116 19740 39172 19742
rect 38892 19628 38948 19684
rect 37772 19068 37828 19124
rect 38668 19068 38724 19124
rect 37436 18508 37492 18564
rect 38220 18396 38276 18452
rect 38556 18450 38612 18452
rect 37996 18060 38052 18116
rect 37772 17612 37828 17668
rect 37660 17276 37716 17332
rect 36036 15148 36092 15204
rect 36316 14642 36372 14644
rect 36316 14590 36318 14642
rect 36318 14590 36370 14642
rect 36370 14590 36372 14642
rect 36316 14588 36372 14590
rect 37548 16828 37604 16884
rect 38556 18398 38558 18450
rect 38558 18398 38610 18450
rect 38610 18398 38612 18450
rect 38556 18396 38612 18398
rect 38220 17666 38276 17668
rect 38220 17614 38222 17666
rect 38222 17614 38274 17666
rect 38274 17614 38276 17666
rect 38220 17612 38276 17614
rect 38556 17500 38612 17556
rect 38108 16828 38164 16884
rect 38220 17164 38276 17220
rect 37884 16492 37940 16548
rect 38108 16044 38164 16100
rect 35868 14476 35924 14532
rect 37212 14588 37268 14644
rect 36652 14252 36708 14308
rect 36316 14028 36372 14084
rect 36204 13916 36260 13972
rect 35532 13692 35588 13748
rect 36036 13804 36092 13860
rect 35196 13354 35252 13356
rect 34692 13244 34748 13300
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 33460 12402 33516 12404
rect 33460 12350 33462 12402
rect 33462 12350 33514 12402
rect 33514 12350 33516 12402
rect 33460 12348 33516 12350
rect 31612 12124 31668 12180
rect 32508 11900 32564 11956
rect 33292 11676 33348 11732
rect 33404 11788 33460 11844
rect 32620 11116 32676 11172
rect 31276 10386 31332 10388
rect 31276 10334 31278 10386
rect 31278 10334 31330 10386
rect 31330 10334 31332 10386
rect 31276 10332 31332 10334
rect 31164 8818 31220 8820
rect 31164 8766 31166 8818
rect 31166 8766 31218 8818
rect 31218 8766 31220 8818
rect 31164 8764 31220 8766
rect 30828 7980 30884 8036
rect 30268 6690 30324 6692
rect 30268 6638 30270 6690
rect 30270 6638 30322 6690
rect 30322 6638 30324 6690
rect 30268 6636 30324 6638
rect 29596 5740 29652 5796
rect 29316 5404 29372 5460
rect 29484 5292 29540 5348
rect 29484 4450 29540 4452
rect 29484 4398 29486 4450
rect 29486 4398 29538 4450
rect 29538 4398 29540 4450
rect 29484 4396 29540 4398
rect 30940 8316 30996 8372
rect 32508 10444 32564 10500
rect 32508 10220 32564 10276
rect 31836 10108 31892 10164
rect 31836 9884 31892 9940
rect 32956 10668 33012 10724
rect 33852 11564 33908 11620
rect 34860 12908 34916 12964
rect 34524 12178 34580 12180
rect 34524 12126 34526 12178
rect 34526 12126 34578 12178
rect 34578 12126 34580 12178
rect 35196 12962 35252 12964
rect 35196 12910 35198 12962
rect 35198 12910 35250 12962
rect 35250 12910 35252 12962
rect 35196 12908 35252 12910
rect 36204 13356 36260 13412
rect 35812 13020 35868 13076
rect 36204 12908 36260 12964
rect 35644 12684 35700 12740
rect 35756 12402 35812 12404
rect 35756 12350 35758 12402
rect 35758 12350 35810 12402
rect 35810 12350 35812 12402
rect 35756 12348 35812 12350
rect 36204 12572 36260 12628
rect 34524 12124 34580 12126
rect 34692 12012 34748 12068
rect 34188 11340 34244 11396
rect 34300 11676 34356 11732
rect 35644 12124 35700 12180
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 34524 11228 34580 11284
rect 34020 10668 34076 10724
rect 32620 9660 32676 9716
rect 33684 9602 33740 9604
rect 33684 9550 33686 9602
rect 33686 9550 33738 9602
rect 33738 9550 33740 9602
rect 33684 9548 33740 9550
rect 33852 9324 33908 9380
rect 35476 11618 35532 11620
rect 35476 11566 35478 11618
rect 35478 11566 35530 11618
rect 35530 11566 35532 11618
rect 35476 11564 35532 11566
rect 34972 11394 35028 11396
rect 34972 11342 34974 11394
rect 34974 11342 35026 11394
rect 35026 11342 35028 11394
rect 34972 11340 35028 11342
rect 35140 11340 35196 11396
rect 34412 10220 34468 10276
rect 34132 10108 34188 10164
rect 35532 11228 35588 11284
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 32228 8876 32284 8932
rect 32396 8764 32452 8820
rect 31388 7644 31444 7700
rect 32138 7980 32194 8036
rect 34692 9826 34748 9828
rect 34692 9774 34694 9826
rect 34694 9774 34746 9826
rect 34746 9774 34748 9826
rect 34692 9772 34748 9774
rect 36204 12012 36260 12068
rect 35868 11564 35924 11620
rect 36036 11676 36092 11732
rect 35756 11394 35812 11396
rect 35756 11342 35758 11394
rect 35758 11342 35810 11394
rect 35810 11342 35812 11394
rect 35756 11340 35812 11342
rect 35868 11282 35924 11284
rect 35868 11230 35870 11282
rect 35870 11230 35922 11282
rect 35922 11230 35924 11282
rect 35868 11228 35924 11230
rect 35980 10610 36036 10612
rect 35980 10558 35982 10610
rect 35982 10558 36034 10610
rect 36034 10558 36036 10610
rect 35980 10556 36036 10558
rect 33628 8876 33684 8932
rect 33628 7980 33684 8036
rect 34972 9034 34974 9044
rect 34974 9034 35026 9044
rect 35026 9034 35028 9044
rect 34972 8988 35028 9034
rect 34636 8876 34692 8932
rect 36652 13722 36654 13748
rect 36654 13722 36706 13748
rect 36706 13722 36708 13748
rect 36652 13692 36708 13722
rect 36484 12572 36540 12628
rect 36876 13356 36932 13412
rect 38444 16098 38500 16100
rect 38444 16046 38446 16098
rect 38446 16046 38498 16098
rect 38498 16046 38500 16098
rect 38444 16044 38500 16046
rect 39116 19068 39172 19124
rect 38780 17612 38836 17668
rect 39116 18284 39172 18340
rect 39004 17778 39060 17780
rect 39004 17726 39006 17778
rect 39006 17726 39058 17778
rect 39058 17726 39060 17778
rect 39004 17724 39060 17726
rect 38892 16492 38948 16548
rect 39452 20076 39508 20132
rect 39900 19852 39956 19908
rect 39452 19628 39508 19684
rect 40012 19404 40068 19460
rect 40236 20578 40292 20580
rect 40236 20526 40238 20578
rect 40238 20526 40290 20578
rect 40290 20526 40292 20578
rect 40236 20524 40292 20526
rect 43596 31164 43652 31220
rect 43484 30492 43540 30548
rect 42700 30044 42756 30100
rect 42812 29036 42868 29092
rect 43932 30492 43988 30548
rect 44604 34972 44660 35028
rect 44604 33852 44660 33908
rect 45164 37100 45220 37156
rect 44940 36988 44996 37044
rect 45724 39564 45780 39620
rect 45612 39452 45668 39508
rect 45612 38892 45668 38948
rect 45388 38050 45444 38052
rect 45388 37998 45390 38050
rect 45390 37998 45442 38050
rect 45442 37998 45444 38050
rect 45388 37996 45444 37998
rect 45388 37772 45444 37828
rect 45276 36876 45332 36932
rect 45276 36540 45332 36596
rect 45052 36258 45108 36260
rect 45052 36206 45054 36258
rect 45054 36206 45106 36258
rect 45106 36206 45108 36258
rect 45052 36204 45108 36206
rect 44828 35698 44884 35700
rect 44828 35646 44830 35698
rect 44830 35646 44882 35698
rect 44882 35646 44884 35698
rect 44828 35644 44884 35646
rect 44940 35026 44996 35028
rect 44940 34974 44942 35026
rect 44942 34974 44994 35026
rect 44994 34974 44996 35026
rect 44940 34972 44996 34974
rect 45388 35756 45444 35812
rect 45388 35532 45444 35588
rect 45164 34412 45220 34468
rect 44828 34188 44884 34244
rect 45276 34242 45332 34244
rect 45276 34190 45278 34242
rect 45278 34190 45330 34242
rect 45330 34190 45332 34242
rect 45276 34188 45332 34190
rect 45668 36428 45724 36484
rect 45612 35084 45668 35140
rect 45948 38332 46004 38388
rect 46172 39618 46228 39620
rect 46172 39566 46174 39618
rect 46174 39566 46226 39618
rect 46226 39566 46228 39618
rect 46172 39564 46228 39566
rect 46396 39788 46452 39844
rect 46396 38892 46452 38948
rect 46732 39116 46788 39172
rect 46562 38834 46618 38836
rect 46562 38782 46564 38834
rect 46564 38782 46616 38834
rect 46616 38782 46618 38834
rect 46562 38780 46618 38782
rect 46284 38668 46340 38724
rect 46396 38556 46452 38612
rect 46172 37548 46228 37604
rect 46956 38780 47012 38836
rect 46732 38332 46788 38388
rect 46732 37772 46788 37828
rect 46396 37266 46452 37268
rect 46396 37214 46398 37266
rect 46398 37214 46450 37266
rect 46450 37214 46452 37266
rect 46396 37212 46452 37214
rect 46172 36988 46228 37044
rect 46284 36876 46340 36932
rect 46956 37660 47012 37716
rect 47460 39004 47516 39060
rect 47852 43932 47908 43988
rect 48020 43708 48076 43764
rect 48188 43596 48244 43652
rect 48300 43484 48356 43540
rect 47740 43036 47796 43092
rect 48076 42812 48132 42868
rect 47740 42754 47796 42756
rect 47740 42702 47742 42754
rect 47742 42702 47794 42754
rect 47794 42702 47796 42754
rect 47740 42700 47796 42702
rect 47852 41580 47908 41636
rect 48076 41468 48132 41524
rect 47740 40796 47796 40852
rect 48076 39506 48132 39508
rect 48076 39454 48078 39506
rect 48078 39454 48130 39506
rect 48130 39454 48132 39506
rect 48076 39452 48132 39454
rect 47740 38834 47796 38836
rect 47740 38782 47742 38834
rect 47742 38782 47794 38834
rect 47794 38782 47796 38834
rect 47740 38780 47796 38782
rect 47292 37436 47348 37492
rect 48076 38220 48132 38276
rect 47852 37100 47908 37156
rect 46284 35084 46340 35140
rect 48020 36540 48076 36596
rect 46620 35532 46676 35588
rect 47404 35698 47460 35700
rect 47404 35646 47406 35698
rect 47406 35646 47458 35698
rect 47458 35646 47460 35698
rect 47404 35644 47460 35646
rect 47292 35308 47348 35364
rect 47180 35084 47236 35140
rect 46060 34914 46116 34916
rect 46060 34862 46062 34914
rect 46062 34862 46114 34914
rect 46114 34862 46116 34914
rect 46060 34860 46116 34862
rect 45276 33964 45332 34020
rect 45892 34018 45948 34020
rect 45892 33966 45894 34018
rect 45894 33966 45946 34018
rect 45946 33966 45948 34018
rect 45892 33964 45948 33966
rect 44716 33516 44772 33572
rect 44828 33852 44884 33908
rect 44716 31948 44772 32004
rect 44716 31164 44772 31220
rect 45052 33122 45108 33124
rect 45052 33070 45054 33122
rect 45054 33070 45106 33122
rect 45106 33070 45108 33122
rect 45052 33068 45108 33070
rect 46172 33180 46228 33236
rect 46844 33964 46900 34020
rect 47852 35586 47908 35588
rect 47852 35534 47854 35586
rect 47854 35534 47906 35586
rect 47906 35534 47908 35586
rect 47852 35532 47908 35534
rect 48132 35308 48188 35364
rect 47516 34018 47572 34020
rect 47516 33966 47518 34018
rect 47518 33966 47570 34018
rect 47570 33966 47572 34018
rect 47516 33964 47572 33966
rect 47180 33628 47236 33684
rect 45612 32956 45668 33012
rect 46488 32620 46544 32676
rect 45612 32562 45668 32564
rect 45612 32510 45614 32562
rect 45614 32510 45666 32562
rect 45666 32510 45668 32562
rect 45612 32508 45668 32510
rect 46284 32508 46340 32564
rect 47292 32620 47348 32676
rect 44492 30380 44548 30436
rect 43820 30156 43876 30212
rect 45164 30044 45220 30100
rect 45836 32060 45892 32116
rect 45668 30434 45724 30436
rect 45668 30382 45670 30434
rect 45670 30382 45722 30434
rect 45722 30382 45724 30434
rect 45668 30380 45724 30382
rect 45388 30156 45444 30212
rect 45052 29372 45108 29428
rect 44492 29260 44548 29316
rect 43372 28924 43428 28980
rect 43260 28642 43316 28644
rect 43260 28590 43262 28642
rect 43262 28590 43314 28642
rect 43314 28590 43316 28642
rect 43260 28588 43316 28590
rect 43708 28866 43764 28868
rect 43708 28814 43710 28866
rect 43710 28814 43762 28866
rect 43762 28814 43764 28866
rect 43708 28812 43764 28814
rect 44324 28754 44380 28756
rect 44324 28702 44326 28754
rect 44326 28702 44378 28754
rect 44378 28702 44380 28754
rect 44324 28700 44380 28702
rect 43036 27804 43092 27860
rect 42588 26684 42644 26740
rect 43036 27580 43092 27636
rect 42476 26290 42532 26292
rect 42476 26238 42478 26290
rect 42478 26238 42530 26290
rect 42530 26238 42532 26290
rect 42476 26236 42532 26238
rect 41692 25788 41748 25844
rect 41580 24444 41636 24500
rect 42252 24892 42308 24948
rect 42140 24610 42196 24612
rect 42140 24558 42142 24610
rect 42142 24558 42194 24610
rect 42194 24558 42196 24610
rect 42140 24556 42196 24558
rect 41356 23436 41412 23492
rect 40908 21756 40964 21812
rect 40684 21532 40740 21588
rect 40348 20018 40404 20020
rect 40348 19966 40350 20018
rect 40350 19966 40402 20018
rect 40402 19966 40404 20018
rect 40348 19964 40404 19966
rect 39676 18172 39732 18228
rect 39564 18060 39620 18116
rect 39844 18060 39900 18116
rect 39340 17948 39396 18004
rect 40236 18338 40292 18340
rect 40236 18286 40238 18338
rect 40238 18286 40290 18338
rect 40290 18286 40292 18338
rect 40236 18284 40292 18286
rect 40124 17612 40180 17668
rect 40236 17948 40292 18004
rect 39228 16828 39284 16884
rect 39228 16380 39284 16436
rect 39564 16940 39620 16996
rect 38332 14812 38388 14868
rect 37940 14364 37996 14420
rect 38332 14364 38388 14420
rect 37716 14028 37772 14084
rect 38556 14252 38612 14308
rect 37100 13020 37156 13076
rect 37212 12908 37268 12964
rect 37324 13132 37380 13188
rect 37772 13132 37828 13188
rect 37884 13244 37940 13300
rect 37660 13074 37716 13076
rect 37660 13022 37662 13074
rect 37662 13022 37714 13074
rect 37714 13022 37716 13074
rect 37660 13020 37716 13022
rect 38220 13356 38276 13412
rect 37156 12684 37212 12740
rect 36876 12124 36932 12180
rect 36988 12572 37044 12628
rect 37324 12348 37380 12404
rect 37436 12460 37492 12516
rect 37324 12178 37380 12180
rect 37324 12126 37326 12178
rect 37326 12126 37378 12178
rect 37378 12126 37380 12178
rect 37324 12124 37380 12126
rect 37996 12684 38052 12740
rect 36764 11788 36820 11844
rect 37436 11788 37492 11844
rect 37100 11564 37156 11620
rect 36988 10834 37044 10836
rect 36988 10782 36990 10834
rect 36990 10782 37042 10834
rect 37042 10782 37044 10834
rect 36988 10780 37044 10782
rect 37100 10556 37156 10612
rect 37212 11340 37268 11396
rect 36988 10444 37044 10500
rect 35980 9811 36036 9828
rect 35980 9772 35982 9811
rect 35982 9772 36034 9811
rect 36034 9772 36036 9811
rect 35868 9100 35924 9156
rect 35532 9042 35588 9044
rect 35532 8990 35534 9042
rect 35534 8990 35586 9042
rect 35586 8990 35588 9042
rect 35532 8988 35588 8990
rect 35308 8876 35364 8932
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 33740 8204 33796 8260
rect 33404 7756 33460 7812
rect 34188 8258 34244 8260
rect 34188 8206 34190 8258
rect 34190 8206 34242 8258
rect 34242 8206 34244 8258
rect 34188 8204 34244 8206
rect 31276 7084 31332 7140
rect 30772 5906 30828 5908
rect 30772 5854 30774 5906
rect 30774 5854 30826 5906
rect 30826 5854 30828 5906
rect 31612 6412 31668 6468
rect 30772 5852 30828 5854
rect 30268 5292 30324 5348
rect 31388 5404 31444 5460
rect 31724 5794 31780 5796
rect 31724 5742 31726 5794
rect 31726 5742 31778 5794
rect 31778 5742 31780 5794
rect 31724 5740 31780 5742
rect 31892 5404 31948 5460
rect 33404 7308 33460 7364
rect 33180 6524 33236 6580
rect 33516 6578 33572 6580
rect 33516 6526 33518 6578
rect 33518 6526 33570 6578
rect 33570 6526 33572 6578
rect 33516 6524 33572 6526
rect 32956 6076 33012 6132
rect 33338 6412 33394 6468
rect 32508 5964 32564 6020
rect 32172 5234 32228 5236
rect 32172 5182 32174 5234
rect 32174 5182 32226 5234
rect 32226 5182 32228 5234
rect 32172 5180 32228 5182
rect 32508 5180 32564 5236
rect 32060 5068 32116 5124
rect 33740 5852 33796 5908
rect 34020 8034 34076 8036
rect 34020 7982 34022 8034
rect 34022 7982 34074 8034
rect 34074 7982 34076 8034
rect 34020 7980 34076 7982
rect 34188 6748 34244 6804
rect 34076 6076 34132 6132
rect 33964 5852 34020 5908
rect 33908 5628 33964 5684
rect 33740 5516 33796 5572
rect 33348 5292 33404 5348
rect 33180 5068 33236 5124
rect 31724 4956 31780 5012
rect 32732 4844 32788 4900
rect 32396 4732 32452 4788
rect 30772 3724 30828 3780
rect 31500 3836 31556 3892
rect 32396 3836 32452 3892
rect 33628 4732 33684 4788
rect 32788 3724 32844 3780
rect 32340 3666 32396 3668
rect 32340 3614 32342 3666
rect 32342 3614 32394 3666
rect 32394 3614 32396 3666
rect 32340 3612 32396 3614
rect 33964 4508 34020 4564
rect 33236 3666 33292 3668
rect 33236 3614 33238 3666
rect 33238 3614 33290 3666
rect 33290 3614 33292 3666
rect 33236 3612 33292 3614
rect 33628 3521 33684 3556
rect 33628 3500 33630 3521
rect 33630 3500 33682 3521
rect 33682 3500 33684 3521
rect 34412 7980 34468 8036
rect 34692 8258 34748 8260
rect 34692 8206 34694 8258
rect 34694 8206 34746 8258
rect 34746 8206 34748 8258
rect 34692 8204 34748 8206
rect 35308 8370 35364 8372
rect 35308 8318 35310 8370
rect 35310 8318 35362 8370
rect 35362 8318 35364 8370
rect 35308 8316 35364 8318
rect 35980 8258 36036 8260
rect 35980 8206 35982 8258
rect 35982 8206 36034 8258
rect 36034 8206 36036 8258
rect 35980 8204 36036 8206
rect 36316 9884 36372 9940
rect 36652 10332 36708 10388
rect 39228 14812 39284 14868
rect 39452 14530 39508 14532
rect 39452 14478 39454 14530
rect 39454 14478 39506 14530
rect 39506 14478 39508 14530
rect 39452 14476 39508 14478
rect 38444 12684 38500 12740
rect 38892 13468 38948 13524
rect 40012 16828 40068 16884
rect 39676 14252 39732 14308
rect 39956 13970 40012 13972
rect 39956 13918 39958 13970
rect 39958 13918 40010 13970
rect 40010 13918 40012 13970
rect 39956 13916 40012 13918
rect 39284 13244 39340 13300
rect 38668 13074 38724 13076
rect 38668 13022 38670 13074
rect 38670 13022 38722 13074
rect 38722 13022 38724 13074
rect 38668 13020 38724 13022
rect 38556 12460 38612 12516
rect 39396 12684 39452 12740
rect 38556 12290 38612 12292
rect 38556 12238 38558 12290
rect 38558 12238 38610 12290
rect 38610 12238 38612 12290
rect 38556 12236 38612 12238
rect 38892 12178 38948 12180
rect 38556 12012 38612 12068
rect 38892 12126 38894 12178
rect 38894 12126 38946 12178
rect 38946 12126 38948 12178
rect 38892 12124 38948 12126
rect 38332 11676 38388 11732
rect 39956 12178 40012 12180
rect 39956 12126 39958 12178
rect 39958 12126 40010 12178
rect 40010 12126 40012 12178
rect 39956 12124 40012 12126
rect 39004 11676 39060 11732
rect 37548 11394 37604 11396
rect 37548 11342 37550 11394
rect 37550 11342 37602 11394
rect 37602 11342 37604 11394
rect 37548 11340 37604 11342
rect 37324 10610 37380 10612
rect 37324 10558 37326 10610
rect 37326 10558 37378 10610
rect 37378 10558 37380 10610
rect 37324 10556 37380 10558
rect 38556 10892 38612 10948
rect 37996 10610 38052 10612
rect 37996 10558 37998 10610
rect 37998 10558 38050 10610
rect 38050 10558 38052 10610
rect 37996 10556 38052 10558
rect 36484 9154 36540 9156
rect 36484 9102 36486 9154
rect 36486 9102 36538 9154
rect 36538 9102 36540 9154
rect 36484 9100 36540 9102
rect 36204 8204 36260 8260
rect 34916 7644 34972 7700
rect 35420 7474 35476 7476
rect 35420 7422 35422 7474
rect 35422 7422 35474 7474
rect 35474 7422 35476 7474
rect 35420 7420 35476 7422
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 36428 7980 36484 8036
rect 36204 7532 36260 7588
rect 37156 9100 37212 9156
rect 36988 7644 37044 7700
rect 36316 7420 36372 7476
rect 36204 6972 36260 7028
rect 37604 9938 37660 9940
rect 37604 9886 37606 9938
rect 37606 9886 37658 9938
rect 37658 9886 37660 9938
rect 37604 9884 37660 9886
rect 38668 10610 38724 10612
rect 38668 10558 38670 10610
rect 38670 10558 38722 10610
rect 38722 10558 38724 10610
rect 38668 10556 38724 10558
rect 38332 10386 38388 10388
rect 38332 10334 38334 10386
rect 38334 10334 38386 10386
rect 38386 10334 38388 10386
rect 38332 10332 38388 10334
rect 38892 11394 38948 11396
rect 38892 11342 38894 11394
rect 38894 11342 38946 11394
rect 38946 11342 38948 11394
rect 38892 11340 38948 11342
rect 38780 10332 38836 10388
rect 39228 11170 39284 11172
rect 39228 11118 39230 11170
rect 39230 11118 39282 11170
rect 39282 11118 39284 11170
rect 39228 11116 39284 11118
rect 40348 15986 40404 15988
rect 40348 15934 40350 15986
rect 40350 15934 40402 15986
rect 40402 15934 40404 15986
rect 40348 15932 40404 15934
rect 40292 14476 40348 14532
rect 40460 14252 40516 14308
rect 41468 21868 41524 21924
rect 42084 24050 42140 24052
rect 42084 23998 42086 24050
rect 42086 23998 42138 24050
rect 42138 23998 42140 24050
rect 42084 23996 42140 23998
rect 42084 23548 42140 23604
rect 41580 21756 41636 21812
rect 42476 24780 42532 24836
rect 42588 24668 42644 24724
rect 43148 26908 43204 26964
rect 43820 26796 43876 26852
rect 44380 26908 44436 26964
rect 43484 26236 43540 26292
rect 43260 25676 43316 25732
rect 44044 25730 44100 25732
rect 44044 25678 44046 25730
rect 44046 25678 44098 25730
rect 44098 25678 44100 25730
rect 44044 25676 44100 25678
rect 43260 24892 43316 24948
rect 42980 24498 43036 24500
rect 42980 24446 42982 24498
rect 42982 24446 43034 24498
rect 43034 24446 43036 24498
rect 42980 24444 43036 24446
rect 43372 24780 43428 24836
rect 43876 24722 43932 24724
rect 43876 24670 43878 24722
rect 43878 24670 43930 24722
rect 43930 24670 43932 24722
rect 43876 24668 43932 24670
rect 43148 24444 43204 24500
rect 42532 24050 42588 24052
rect 42532 23998 42534 24050
rect 42534 23998 42586 24050
rect 42586 23998 42588 24050
rect 42532 23996 42588 23998
rect 42476 23660 42532 23716
rect 42252 22428 42308 22484
rect 42364 23212 42420 23268
rect 42140 22316 42196 22372
rect 42364 21868 42420 21924
rect 42588 22988 42644 23044
rect 42476 22540 42532 22596
rect 42700 22316 42756 22372
rect 43036 23660 43092 23716
rect 43036 22428 43092 22484
rect 43932 22428 43988 22484
rect 44044 22370 44100 22372
rect 44044 22318 44046 22370
rect 44046 22318 44098 22370
rect 44098 22318 44100 22370
rect 44044 22316 44100 22318
rect 43260 22204 43316 22260
rect 41020 20860 41076 20916
rect 40796 20636 40852 20692
rect 41524 20914 41580 20916
rect 41524 20862 41526 20914
rect 41526 20862 41578 20914
rect 41578 20862 41580 20914
rect 41524 20860 41580 20862
rect 42252 20972 42308 21028
rect 40908 19964 40964 20020
rect 41020 18450 41076 18452
rect 41020 18398 41022 18450
rect 41022 18398 41074 18450
rect 41074 18398 41076 18450
rect 41020 18396 41076 18398
rect 40908 17948 40964 18004
rect 40908 17500 40964 17556
rect 40796 17164 40852 17220
rect 40908 16857 40910 16884
rect 40910 16857 40962 16884
rect 40962 16857 40964 16884
rect 40908 16828 40964 16857
rect 40908 16604 40964 16660
rect 40908 15484 40964 15540
rect 42786 19628 42842 19684
rect 41804 18620 41860 18676
rect 41300 18508 41356 18564
rect 41692 18284 41748 18340
rect 42364 18284 42420 18340
rect 42700 18396 42756 18452
rect 41132 17724 41188 17780
rect 41634 17724 41690 17780
rect 41356 17276 41412 17332
rect 41468 17666 41524 17668
rect 41468 17614 41470 17666
rect 41470 17614 41522 17666
rect 41522 17614 41524 17666
rect 41468 17612 41524 17614
rect 40684 13916 40740 13972
rect 41132 15932 41188 15988
rect 41356 15372 41412 15428
rect 41132 15260 41188 15316
rect 40236 12236 40292 12292
rect 40348 11900 40404 11956
rect 40348 11676 40404 11732
rect 40236 11340 40292 11396
rect 38108 9938 38164 9940
rect 38108 9886 38110 9938
rect 38110 9886 38162 9938
rect 38162 9886 38164 9938
rect 38108 9884 38164 9886
rect 38668 9996 38724 10052
rect 37548 8316 37604 8372
rect 39732 10050 39788 10052
rect 39732 9998 39734 10050
rect 39734 9998 39786 10050
rect 39786 9998 39788 10050
rect 39732 9996 39788 9998
rect 39004 9660 39060 9716
rect 39228 9826 39284 9828
rect 39228 9774 39230 9826
rect 39230 9774 39282 9826
rect 39282 9774 39284 9826
rect 39228 9772 39284 9774
rect 39452 9826 39508 9828
rect 39452 9774 39454 9826
rect 39454 9774 39506 9826
rect 39506 9774 39508 9826
rect 39452 9772 39508 9774
rect 39956 9772 40012 9828
rect 40236 9884 40292 9940
rect 39452 9100 39508 9156
rect 37884 8258 37940 8260
rect 37884 8206 37886 8258
rect 37886 8206 37938 8258
rect 37938 8206 37940 8258
rect 37884 8204 37940 8206
rect 38108 7980 38164 8036
rect 37996 7868 38052 7924
rect 35084 6076 35140 6132
rect 34076 3948 34132 4004
rect 34748 5906 34804 5908
rect 34748 5854 34750 5906
rect 34750 5854 34802 5906
rect 34802 5854 34804 5906
rect 34748 5852 34804 5854
rect 35196 5852 35252 5908
rect 36204 5906 36260 5908
rect 36204 5854 36206 5906
rect 36206 5854 36258 5906
rect 36258 5854 36260 5906
rect 36204 5852 36260 5854
rect 35868 5794 35924 5796
rect 35868 5742 35870 5794
rect 35870 5742 35922 5794
rect 35922 5742 35924 5794
rect 35868 5740 35924 5742
rect 34972 5628 35028 5684
rect 34636 5068 34692 5124
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35196 5292 35252 5348
rect 35532 5068 35588 5124
rect 36204 5628 36260 5684
rect 35756 5068 35812 5124
rect 34748 4508 34804 4564
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 37436 7644 37492 7700
rect 36764 6412 36820 6468
rect 36652 5794 36708 5796
rect 36652 5742 36654 5794
rect 36654 5742 36706 5794
rect 36706 5742 36708 5794
rect 36652 5740 36708 5742
rect 36484 5122 36540 5124
rect 36484 5070 36486 5122
rect 36486 5070 36538 5122
rect 36538 5070 36540 5122
rect 36484 5068 36540 5070
rect 35980 3724 36036 3780
rect 37268 6412 37324 6468
rect 36988 6300 37044 6356
rect 37268 6076 37324 6132
rect 37100 5852 37156 5908
rect 36764 5068 36820 5124
rect 36876 5740 36932 5796
rect 36372 3666 36428 3668
rect 36372 3614 36374 3666
rect 36374 3614 36426 3666
rect 36426 3614 36428 3666
rect 36372 3612 36428 3614
rect 36652 3612 36708 3668
rect 38444 7980 38500 8036
rect 38220 7308 38276 7364
rect 38332 6076 38388 6132
rect 38892 8428 38948 8484
rect 38892 7756 38948 7812
rect 38780 7532 38836 7588
rect 38556 7308 38612 7364
rect 38668 6972 38724 7028
rect 38556 5852 38612 5908
rect 37660 5516 37716 5572
rect 37996 5516 38052 5572
rect 37324 5292 37380 5348
rect 37660 5292 37716 5348
rect 37324 5068 37380 5124
rect 37436 5180 37492 5236
rect 37996 5180 38052 5236
rect 37828 5122 37884 5124
rect 37828 5070 37830 5122
rect 37830 5070 37882 5122
rect 37882 5070 37884 5122
rect 37828 5068 37884 5070
rect 38780 5404 38836 5460
rect 38668 5068 38724 5124
rect 36876 3836 36932 3892
rect 36764 3521 36820 3556
rect 36764 3500 36766 3521
rect 36766 3500 36818 3521
rect 36818 3500 36820 3521
rect 37100 3517 37156 3556
rect 37100 3500 37102 3517
rect 37102 3500 37154 3517
rect 37154 3500 37156 3517
rect 39170 7980 39226 8036
rect 39340 6636 39396 6692
rect 39900 9100 39956 9156
rect 40572 12572 40628 12628
rect 40684 12796 40740 12852
rect 40684 11788 40740 11844
rect 41244 15202 41300 15204
rect 41244 15150 41246 15202
rect 41246 15150 41298 15202
rect 41298 15150 41300 15202
rect 41244 15148 41300 15150
rect 42588 17666 42644 17668
rect 42588 17614 42590 17666
rect 42590 17614 42642 17666
rect 42642 17614 42644 17666
rect 42588 17612 42644 17614
rect 43148 17612 43204 17668
rect 42924 17500 42980 17556
rect 42476 17388 42532 17444
rect 43148 16940 43204 16996
rect 42812 16828 42868 16884
rect 41580 15820 41636 15876
rect 41468 15148 41524 15204
rect 41692 15596 41748 15652
rect 40964 14364 41020 14420
rect 41412 13970 41468 13972
rect 41412 13918 41414 13970
rect 41414 13918 41466 13970
rect 41466 13918 41468 13970
rect 41412 13916 41468 13918
rect 42252 15708 42308 15764
rect 41972 15596 42028 15652
rect 42140 15372 42196 15428
rect 41804 13692 41860 13748
rect 41916 13580 41972 13636
rect 42028 15036 42084 15092
rect 41298 12796 41354 12852
rect 41132 12460 41188 12516
rect 41804 12460 41860 12516
rect 41020 12348 41076 12404
rect 42532 16098 42588 16100
rect 42532 16046 42534 16098
rect 42534 16046 42586 16098
rect 42586 16046 42588 16098
rect 42532 16044 42588 16046
rect 42364 15148 42420 15204
rect 42476 15484 42532 15540
rect 43596 22092 43652 22148
rect 43372 21980 43428 22036
rect 43372 20802 43428 20804
rect 43372 20750 43374 20802
rect 43374 20750 43426 20802
rect 43426 20750 43428 20802
rect 43372 20748 43428 20750
rect 43484 21586 43540 21588
rect 43484 21534 43486 21586
rect 43486 21534 43538 21586
rect 43538 21534 43540 21586
rect 43484 21532 43540 21534
rect 43372 17724 43428 17780
rect 43484 18396 43540 18452
rect 43260 16380 43316 16436
rect 42924 16210 42980 16212
rect 42924 16158 42926 16210
rect 42926 16158 42978 16210
rect 42978 16158 42980 16210
rect 42924 16156 42980 16158
rect 43932 20972 43988 21028
rect 43820 20914 43876 20916
rect 43820 20862 43822 20914
rect 43822 20862 43874 20914
rect 43874 20862 43876 20914
rect 43820 20860 43876 20862
rect 43820 20636 43876 20692
rect 43932 20524 43988 20580
rect 44268 21586 44324 21588
rect 44268 21534 44270 21586
rect 44270 21534 44322 21586
rect 44322 21534 44324 21586
rect 44268 21532 44324 21534
rect 44268 21308 44324 21364
rect 44044 20188 44100 20244
rect 44044 19628 44100 19684
rect 44940 29036 44996 29092
rect 45948 30210 46004 30212
rect 45948 30158 45950 30210
rect 45950 30158 46002 30210
rect 46002 30158 46004 30210
rect 45948 30156 46004 30158
rect 46172 31052 46228 31108
rect 48020 32732 48076 32788
rect 47628 32562 47684 32564
rect 47628 32510 47630 32562
rect 47630 32510 47682 32562
rect 47682 32510 47684 32562
rect 47628 32508 47684 32510
rect 48188 32508 48244 32564
rect 47628 31052 47684 31108
rect 48300 32284 48356 32340
rect 47964 30156 48020 30212
rect 45948 29260 46004 29316
rect 45388 28700 45444 28756
rect 45052 27916 45108 27972
rect 44716 27746 44772 27748
rect 44716 27694 44718 27746
rect 44718 27694 44770 27746
rect 44770 27694 44772 27746
rect 44716 27692 44772 27694
rect 44604 26012 44660 26068
rect 45836 28588 45892 28644
rect 46172 29148 46228 29204
rect 47964 29202 48020 29204
rect 47964 29150 47966 29202
rect 47966 29150 48018 29202
rect 48018 29150 48020 29202
rect 47964 29148 48020 29150
rect 48300 29426 48356 29428
rect 48300 29374 48302 29426
rect 48302 29374 48354 29426
rect 48354 29374 48356 29426
rect 48300 29372 48356 29374
rect 48300 28642 48356 28644
rect 48300 28590 48302 28642
rect 48302 28590 48354 28642
rect 48354 28590 48356 28642
rect 48300 28588 48356 28590
rect 45388 27858 45444 27860
rect 45388 27806 45390 27858
rect 45390 27806 45442 27858
rect 45442 27806 45444 27858
rect 45388 27804 45444 27806
rect 46060 27804 46116 27860
rect 45612 27356 45668 27412
rect 44940 26796 44996 26852
rect 46844 27804 46900 27860
rect 46264 27356 46320 27412
rect 45164 26402 45220 26404
rect 45164 26350 45166 26402
rect 45166 26350 45218 26402
rect 45218 26350 45220 26402
rect 45164 26348 45220 26350
rect 46396 26348 46452 26404
rect 45500 26124 45556 26180
rect 45612 26236 45668 26292
rect 45220 25730 45276 25732
rect 45220 25678 45222 25730
rect 45222 25678 45274 25730
rect 45274 25678 45276 25730
rect 45220 25676 45276 25678
rect 44940 25564 44996 25620
rect 45724 25676 45780 25732
rect 46172 25900 46228 25956
rect 46060 25506 46116 25508
rect 46060 25454 46062 25506
rect 46062 25454 46114 25506
rect 46114 25454 46116 25506
rect 46060 25452 46116 25454
rect 44828 24780 44884 24836
rect 45388 24722 45444 24724
rect 45388 24670 45390 24722
rect 45390 24670 45442 24722
rect 45442 24670 45444 24722
rect 45388 24668 45444 24670
rect 45164 24610 45220 24612
rect 45164 24558 45166 24610
rect 45166 24558 45218 24610
rect 45218 24558 45220 24610
rect 45164 24556 45220 24558
rect 45836 24556 45892 24612
rect 45500 23938 45556 23940
rect 45500 23886 45502 23938
rect 45502 23886 45554 23938
rect 45554 23886 45556 23938
rect 45500 23884 45556 23886
rect 46620 27020 46676 27076
rect 46956 27356 47012 27412
rect 47068 26796 47124 26852
rect 47292 27858 47348 27860
rect 47292 27806 47294 27858
rect 47294 27806 47346 27858
rect 47346 27806 47348 27858
rect 47292 27804 47348 27806
rect 47964 27468 48020 27524
rect 48300 27580 48356 27636
rect 47292 27074 47348 27076
rect 47292 27022 47294 27074
rect 47294 27022 47346 27074
rect 47346 27022 47348 27074
rect 47292 27020 47348 27022
rect 47292 26796 47348 26852
rect 47292 26572 47348 26628
rect 46620 25900 46676 25956
rect 46396 25506 46452 25508
rect 46396 25454 46398 25506
rect 46398 25454 46450 25506
rect 46450 25454 46452 25506
rect 46396 25452 46452 25454
rect 47124 26066 47180 26068
rect 47124 26014 47126 26066
rect 47126 26014 47178 26066
rect 47178 26014 47180 26066
rect 47124 26012 47180 26014
rect 47404 26684 47460 26740
rect 47404 26266 47406 26292
rect 47406 26266 47458 26292
rect 47458 26266 47460 26292
rect 47404 26236 47460 26266
rect 46788 25564 46844 25620
rect 48412 26236 48468 26292
rect 47180 25340 47236 25396
rect 46620 25004 46676 25060
rect 45276 23324 45332 23380
rect 45612 23436 45668 23492
rect 45052 23212 45108 23268
rect 44940 23100 44996 23156
rect 45724 23324 45780 23380
rect 46284 23212 46340 23268
rect 45836 23100 45892 23156
rect 44828 22988 44884 23044
rect 45220 22764 45276 22820
rect 44604 21980 44660 22036
rect 44604 21756 44660 21812
rect 44716 20802 44772 20804
rect 44716 20750 44718 20802
rect 44718 20750 44770 20802
rect 44770 20750 44772 20802
rect 44716 20748 44772 20750
rect 44492 19852 44548 19908
rect 45612 21308 45668 21364
rect 45612 21084 45668 21140
rect 45500 20914 45556 20916
rect 45500 20862 45502 20914
rect 45502 20862 45554 20914
rect 45554 20862 45556 20914
rect 45500 20860 45556 20862
rect 45276 20748 45332 20804
rect 45500 20300 45556 20356
rect 44940 19852 44996 19908
rect 45052 19794 45108 19796
rect 45052 19742 45054 19794
rect 45054 19742 45106 19794
rect 45106 19742 45108 19794
rect 45052 19740 45108 19742
rect 43708 19234 43764 19236
rect 43708 19182 43710 19234
rect 43710 19182 43762 19234
rect 43762 19182 43764 19234
rect 43708 19180 43764 19182
rect 44690 18844 44746 18900
rect 43708 18620 43764 18676
rect 44268 18620 44324 18676
rect 43820 17724 43876 17780
rect 44044 17836 44100 17892
rect 43708 17500 43764 17556
rect 43932 17666 43988 17668
rect 43932 17614 43934 17666
rect 43934 17614 43986 17666
rect 43986 17614 43988 17666
rect 43932 17612 43988 17614
rect 43708 16828 43764 16884
rect 43708 16492 43764 16548
rect 43708 16098 43764 16100
rect 43708 16046 43710 16098
rect 43710 16046 43762 16098
rect 43762 16046 43764 16098
rect 43708 16044 43764 16046
rect 43820 16156 43876 16212
rect 43372 15372 43428 15428
rect 43260 15314 43316 15316
rect 43260 15262 43262 15314
rect 43262 15262 43314 15314
rect 43314 15262 43316 15314
rect 43260 15260 43316 15262
rect 42812 15148 42868 15204
rect 42700 14588 42756 14644
rect 42140 12572 42196 12628
rect 41244 12236 41300 12292
rect 41356 12066 41412 12068
rect 41356 12014 41358 12066
rect 41358 12014 41410 12066
rect 41410 12014 41412 12066
rect 41356 12012 41412 12014
rect 41020 11900 41076 11956
rect 40572 11228 40628 11284
rect 40684 10332 40740 10388
rect 40460 9324 40516 9380
rect 40292 9212 40348 9268
rect 40460 8988 40516 9044
rect 39564 7868 39620 7924
rect 39676 8092 39732 8148
rect 40124 7980 40180 8036
rect 40348 7474 40404 7476
rect 40348 7422 40350 7474
rect 40350 7422 40402 7474
rect 40402 7422 40404 7474
rect 40348 7420 40404 7422
rect 39228 6524 39284 6580
rect 40460 6972 40516 7028
rect 40236 6524 40292 6580
rect 40572 6466 40628 6468
rect 40572 6414 40574 6466
rect 40574 6414 40626 6466
rect 40626 6414 40628 6466
rect 40572 6412 40628 6414
rect 39116 6076 39172 6132
rect 41020 10556 41076 10612
rect 41020 9826 41076 9828
rect 41020 9774 41022 9826
rect 41022 9774 41074 9826
rect 41074 9774 41076 9826
rect 41020 9772 41076 9774
rect 42028 12178 42084 12180
rect 42028 12126 42030 12178
rect 42030 12126 42082 12178
rect 42082 12126 42084 12178
rect 42028 12124 42084 12126
rect 41804 12012 41860 12068
rect 43518 15148 43574 15204
rect 44828 18396 44884 18452
rect 44940 19234 44996 19236
rect 44940 19182 44942 19234
rect 44942 19182 44994 19234
rect 44994 19182 44996 19234
rect 44940 19180 44996 19182
rect 44716 18338 44772 18340
rect 44716 18286 44718 18338
rect 44718 18286 44770 18338
rect 44770 18286 44772 18338
rect 44716 18284 44772 18286
rect 44380 17500 44436 17556
rect 44268 16044 44324 16100
rect 44380 16380 44436 16436
rect 42812 14252 42868 14308
rect 43036 13858 43092 13860
rect 43036 13806 43038 13858
rect 43038 13806 43090 13858
rect 43090 13806 43092 13858
rect 43036 13804 43092 13806
rect 42700 12460 42756 12516
rect 42886 12348 42942 12404
rect 43484 13634 43540 13636
rect 43484 13582 43486 13634
rect 43486 13582 43538 13634
rect 43538 13582 43540 13634
rect 43484 13580 43540 13582
rect 43260 13468 43316 13524
rect 43391 13356 43447 13412
rect 44604 17612 44660 17668
rect 45220 19234 45276 19236
rect 45220 19182 45222 19234
rect 45222 19182 45274 19234
rect 45274 19182 45276 19234
rect 45220 19180 45276 19182
rect 46956 22204 47012 22260
rect 46116 21698 46172 21700
rect 46116 21646 46118 21698
rect 46118 21646 46170 21698
rect 46170 21646 46172 21698
rect 46116 21644 46172 21646
rect 46620 21549 46622 21588
rect 46622 21549 46674 21588
rect 46674 21549 46676 21588
rect 46620 21532 46676 21549
rect 48188 25340 48244 25396
rect 47740 24780 47796 24836
rect 48076 24834 48132 24836
rect 48076 24782 48078 24834
rect 48078 24782 48130 24834
rect 48130 24782 48132 24834
rect 48076 24780 48132 24782
rect 47180 23212 47236 23268
rect 48020 23266 48076 23268
rect 48020 23214 48022 23266
rect 48022 23214 48074 23266
rect 48074 23214 48076 23266
rect 48020 23212 48076 23214
rect 47740 22258 47796 22260
rect 47740 22206 47742 22258
rect 47742 22206 47794 22258
rect 47794 22206 47796 22258
rect 47740 22204 47796 22206
rect 47068 21644 47124 21700
rect 45836 21084 45892 21140
rect 46396 20524 46452 20580
rect 45612 19964 45668 20020
rect 45948 19740 46004 19796
rect 45500 18956 45556 19012
rect 45724 19234 45780 19236
rect 45724 19182 45726 19234
rect 45726 19182 45778 19234
rect 45778 19182 45780 19234
rect 45724 19180 45780 19182
rect 45612 18844 45668 18900
rect 45948 18732 46004 18788
rect 44940 17052 44996 17108
rect 44996 16322 45052 16324
rect 44996 16270 44998 16322
rect 44998 16270 45050 16322
rect 45050 16270 45052 16322
rect 44996 16268 45052 16270
rect 44716 16044 44772 16100
rect 44380 14924 44436 14980
rect 44044 13356 44100 13412
rect 42476 11788 42532 11844
rect 41580 11228 41636 11284
rect 41804 11394 41860 11396
rect 41804 11342 41806 11394
rect 41806 11342 41858 11394
rect 41858 11342 41860 11394
rect 41804 11340 41860 11342
rect 44492 14476 44548 14532
rect 44268 13244 44324 13300
rect 44380 14028 44436 14084
rect 45836 18338 45892 18340
rect 45836 18286 45838 18338
rect 45838 18286 45890 18338
rect 45890 18286 45892 18338
rect 45836 18284 45892 18286
rect 45276 17500 45332 17556
rect 47628 21644 47684 21700
rect 47292 20524 47348 20580
rect 47404 21308 47460 21364
rect 46844 19234 46900 19236
rect 46844 19182 46846 19234
rect 46846 19182 46898 19234
rect 46898 19182 46900 19234
rect 46844 19180 46900 19182
rect 47740 21586 47796 21588
rect 47740 21534 47742 21586
rect 47742 21534 47794 21586
rect 47794 21534 47796 21586
rect 47740 21532 47796 21534
rect 48076 21532 48132 21588
rect 47964 20300 48020 20356
rect 48244 21196 48300 21252
rect 48300 20802 48356 20804
rect 48300 20750 48302 20802
rect 48302 20750 48354 20802
rect 48354 20750 48356 20802
rect 48300 20748 48356 20750
rect 48748 22428 48804 22484
rect 48748 20748 48804 20804
rect 47628 19964 47684 20020
rect 47292 18732 47348 18788
rect 45500 16940 45556 16996
rect 45164 14924 45220 14980
rect 45276 15148 45332 15204
rect 45164 14642 45220 14644
rect 45164 14590 45166 14642
rect 45166 14590 45218 14642
rect 45218 14590 45220 14642
rect 45164 14588 45220 14590
rect 44940 14252 44996 14308
rect 45164 14028 45220 14084
rect 45388 14924 45444 14980
rect 45612 16380 45668 16436
rect 46060 16268 46116 16324
rect 46956 16882 47012 16884
rect 46956 16830 46958 16882
rect 46958 16830 47010 16882
rect 47010 16830 47012 16882
rect 46956 16828 47012 16830
rect 48076 20018 48132 20020
rect 48076 19966 48078 20018
rect 48078 19966 48130 20018
rect 48130 19966 48132 20018
rect 48076 19964 48132 19966
rect 47740 18338 47796 18340
rect 47740 18286 47742 18338
rect 47742 18286 47794 18338
rect 47794 18286 47796 18338
rect 47740 18284 47796 18286
rect 47684 16882 47740 16884
rect 47684 16830 47686 16882
rect 47686 16830 47738 16882
rect 47738 16830 47740 16882
rect 47684 16828 47740 16830
rect 45612 16044 45668 16100
rect 45612 15596 45668 15652
rect 45500 15260 45556 15316
rect 45724 15148 45780 15204
rect 44492 13746 44548 13748
rect 44492 13694 44494 13746
rect 44494 13694 44546 13746
rect 44546 13694 44548 13746
rect 44828 13746 44884 13748
rect 44492 13692 44548 13694
rect 44828 13694 44830 13746
rect 44830 13694 44882 13746
rect 44882 13694 44884 13746
rect 44828 13692 44884 13694
rect 44660 13580 44716 13636
rect 45612 14924 45668 14980
rect 44940 13356 44996 13412
rect 45276 13580 45332 13636
rect 44268 12684 44324 12740
rect 43596 12348 43652 12404
rect 44604 13244 44660 13300
rect 45276 13244 45332 13300
rect 44268 12236 44324 12292
rect 43260 12124 43316 12180
rect 43148 11676 43204 11732
rect 43484 11788 43540 11844
rect 42588 11394 42644 11396
rect 42588 11342 42590 11394
rect 42590 11342 42642 11394
rect 42642 11342 42644 11394
rect 42588 11340 42644 11342
rect 42924 11228 42980 11284
rect 41692 10668 41748 10724
rect 41580 10610 41636 10612
rect 41580 10558 41582 10610
rect 41582 10558 41634 10610
rect 41634 10558 41636 10610
rect 41580 10556 41636 10558
rect 41468 9772 41524 9828
rect 41580 10332 41636 10388
rect 41132 9154 41188 9156
rect 41132 9102 41134 9154
rect 41134 9102 41186 9154
rect 41186 9102 41188 9154
rect 41132 9100 41188 9102
rect 40796 8316 40852 8372
rect 42644 10220 42700 10276
rect 41692 9826 41748 9828
rect 41692 9774 41694 9826
rect 41694 9774 41746 9826
rect 41746 9774 41748 9826
rect 41692 9772 41748 9774
rect 41804 8876 41860 8932
rect 43820 11676 43876 11732
rect 43372 10556 43428 10612
rect 44044 10722 44100 10724
rect 44044 10670 44046 10722
rect 44046 10670 44098 10722
rect 44098 10670 44100 10722
rect 44044 10668 44100 10670
rect 43372 10332 43428 10388
rect 44100 10444 44156 10500
rect 44940 12178 44996 12180
rect 44940 12126 44942 12178
rect 44942 12126 44994 12178
rect 44994 12126 44996 12178
rect 44940 12124 44996 12126
rect 45500 13356 45556 13412
rect 45388 12236 45444 12292
rect 45164 12012 45220 12068
rect 44660 11954 44716 11956
rect 44660 11902 44662 11954
rect 44662 11902 44714 11954
rect 44714 11902 44716 11954
rect 44660 11900 44716 11902
rect 47068 16098 47124 16100
rect 47068 16046 47070 16098
rect 47070 16046 47122 16098
rect 47122 16046 47124 16098
rect 47068 16044 47124 16046
rect 47292 16098 47348 16100
rect 47292 16046 47294 16098
rect 47294 16046 47346 16098
rect 47346 16046 47348 16098
rect 47292 16044 47348 16046
rect 46620 15596 46676 15652
rect 47516 15596 47572 15652
rect 46396 15148 46452 15204
rect 46844 14924 46900 14980
rect 46172 14588 46228 14644
rect 45836 14530 45892 14532
rect 45836 14478 45838 14530
rect 45838 14478 45890 14530
rect 45890 14478 45892 14530
rect 45836 14476 45892 14478
rect 48076 16492 48132 16548
rect 48300 19852 48356 19908
rect 47964 16044 48020 16100
rect 45948 14252 46004 14308
rect 45724 13804 45780 13860
rect 46508 13804 46564 13860
rect 45948 13746 46004 13748
rect 45948 13694 45950 13746
rect 45950 13694 46002 13746
rect 46002 13694 46004 13746
rect 45948 13692 46004 13694
rect 48412 16156 48468 16212
rect 48300 15314 48356 15316
rect 48300 15262 48302 15314
rect 48302 15262 48354 15314
rect 48354 15262 48356 15314
rect 48300 15260 48356 15262
rect 45724 12684 45780 12740
rect 45612 12236 45668 12292
rect 46172 12684 46228 12740
rect 46482 12572 46538 12628
rect 47292 12572 47348 12628
rect 47516 12460 47572 12516
rect 47628 13468 47684 13524
rect 47068 12178 47124 12180
rect 47068 12126 47070 12178
rect 47070 12126 47122 12178
rect 47122 12126 47124 12178
rect 47068 12124 47124 12126
rect 47292 12178 47348 12180
rect 47292 12126 47294 12178
rect 47294 12126 47346 12178
rect 47346 12126 47348 12178
rect 47292 12124 47348 12126
rect 48076 13468 48132 13524
rect 48300 12572 48356 12628
rect 48132 12460 48188 12516
rect 44492 10892 44548 10948
rect 42924 9772 42980 9828
rect 42028 9212 42084 9268
rect 43708 9660 43764 9716
rect 43036 8930 43092 8932
rect 43036 8878 43038 8930
rect 43038 8878 43090 8930
rect 43090 8878 43092 8930
rect 43036 8876 43092 8878
rect 41580 8258 41636 8260
rect 41580 8206 41582 8258
rect 41582 8206 41634 8258
rect 41634 8206 41636 8258
rect 44996 10892 45052 10948
rect 44828 10780 44884 10836
rect 45388 10780 45444 10836
rect 45388 10220 45444 10276
rect 46172 11900 46228 11956
rect 45836 11788 45892 11844
rect 46956 11788 47012 11844
rect 45724 10220 45780 10276
rect 45836 11116 45892 11172
rect 44716 9660 44772 9716
rect 44940 9436 44996 9492
rect 42364 8316 42420 8372
rect 41580 8204 41636 8206
rect 41020 7196 41076 7252
rect 41300 6972 41356 7028
rect 41356 6636 41412 6692
rect 41020 6412 41076 6468
rect 39004 5964 39060 6020
rect 39116 5906 39172 5908
rect 39116 5854 39118 5906
rect 39118 5854 39170 5906
rect 39170 5854 39172 5906
rect 39452 5964 39508 6020
rect 39116 5852 39172 5854
rect 39004 5404 39060 5460
rect 38108 3948 38164 4004
rect 37746 3388 37802 3444
rect 38780 4284 38836 4340
rect 39284 5404 39340 5460
rect 40180 5740 40236 5796
rect 40572 5740 40628 5796
rect 39116 4956 39172 5012
rect 39452 5068 39508 5124
rect 39788 5122 39844 5124
rect 39788 5070 39790 5122
rect 39790 5070 39842 5122
rect 39842 5070 39844 5122
rect 39788 5068 39844 5070
rect 40236 5404 40292 5460
rect 40348 4956 40404 5012
rect 39900 4338 39956 4340
rect 39900 4286 39902 4338
rect 39902 4286 39954 4338
rect 39954 4286 39956 4338
rect 39900 4284 39956 4286
rect 40236 3724 40292 3780
rect 39956 3666 40012 3668
rect 39956 3614 39958 3666
rect 39958 3614 40010 3666
rect 40010 3614 40012 3666
rect 39956 3612 40012 3614
rect 40292 3554 40348 3556
rect 40292 3502 40294 3554
rect 40294 3502 40346 3554
rect 40346 3502 40348 3554
rect 40292 3500 40348 3502
rect 39788 3388 39844 3444
rect 40908 5628 40964 5684
rect 43820 8316 43876 8372
rect 43036 8092 43092 8148
rect 42252 7868 42308 7924
rect 41580 7420 41636 7476
rect 42252 7474 42308 7476
rect 42252 7422 42254 7474
rect 42254 7422 42306 7474
rect 42306 7422 42308 7474
rect 42252 7420 42308 7422
rect 41692 7362 41748 7364
rect 41692 7310 41694 7362
rect 41694 7310 41746 7362
rect 41746 7310 41748 7362
rect 41692 7308 41748 7310
rect 43428 7980 43484 8036
rect 42588 7308 42644 7364
rect 42924 7474 42980 7476
rect 42924 7422 42926 7474
rect 42926 7422 42978 7474
rect 42978 7422 42980 7474
rect 42924 7420 42980 7422
rect 44130 8540 44186 8596
rect 44716 8316 44772 8372
rect 44268 8204 44324 8260
rect 43148 7308 43204 7364
rect 43764 7980 43820 8036
rect 43932 8092 43988 8148
rect 41692 6524 41748 6580
rect 41804 5906 41860 5908
rect 41804 5854 41806 5906
rect 41806 5854 41858 5906
rect 41858 5854 41860 5906
rect 41804 5852 41860 5854
rect 41132 5404 41188 5460
rect 41580 5740 41636 5796
rect 40684 5292 40740 5348
rect 40796 5180 40852 5236
rect 42140 5906 42196 5908
rect 42140 5854 42142 5906
rect 42142 5854 42194 5906
rect 42194 5854 42196 5906
rect 42140 5852 42196 5854
rect 42364 6188 42420 6244
rect 43036 6636 43092 6692
rect 43148 6748 43204 6804
rect 42644 6524 42700 6580
rect 42476 6412 42532 6468
rect 42476 5964 42532 6020
rect 42812 5852 42868 5908
rect 42028 5516 42084 5572
rect 41020 5068 41076 5124
rect 40684 4396 40740 4452
rect 40852 3836 40908 3892
rect 40684 3500 40740 3556
rect 41692 5068 41748 5124
rect 41412 4396 41468 4452
rect 42364 5122 42420 5124
rect 42364 5070 42366 5122
rect 42366 5070 42418 5122
rect 42418 5070 42420 5122
rect 42364 5068 42420 5070
rect 42476 4956 42532 5012
rect 41356 4226 41412 4228
rect 41356 4174 41358 4226
rect 41358 4174 41410 4226
rect 41410 4174 41412 4226
rect 41356 4172 41412 4174
rect 41468 3836 41524 3892
rect 42700 5292 42756 5348
rect 45948 10610 46004 10612
rect 45948 10558 45950 10610
rect 45950 10558 46002 10610
rect 46002 10558 46004 10610
rect 45948 10556 46004 10558
rect 46844 11394 46900 11396
rect 46482 11228 46538 11284
rect 46844 11342 46846 11394
rect 46846 11342 46898 11394
rect 46898 11342 46900 11394
rect 46844 11340 46900 11342
rect 46732 10220 46788 10276
rect 46956 11228 47012 11284
rect 47068 10610 47124 10612
rect 47068 10558 47070 10610
rect 47070 10558 47122 10610
rect 47122 10558 47124 10610
rect 47068 10556 47124 10558
rect 46844 10108 46900 10164
rect 45276 9042 45332 9044
rect 45276 8990 45278 9042
rect 45278 8990 45330 9042
rect 45330 8990 45332 9042
rect 45276 8988 45332 8990
rect 45612 9042 45668 9044
rect 45612 8990 45614 9042
rect 45614 8990 45666 9042
rect 45666 8990 45668 9042
rect 45612 8988 45668 8990
rect 45108 8316 45164 8372
rect 45500 8258 45556 8260
rect 45500 8206 45502 8258
rect 45502 8206 45554 8258
rect 45554 8206 45556 8258
rect 45500 8204 45556 8206
rect 44940 8092 44996 8148
rect 47124 9266 47180 9268
rect 47124 9214 47126 9266
rect 47126 9214 47178 9266
rect 47178 9214 47180 9266
rect 47124 9212 47180 9214
rect 46172 8540 46228 8596
rect 46620 9042 46676 9044
rect 46620 8990 46622 9042
rect 46622 8990 46674 9042
rect 46674 8990 46676 9042
rect 46620 8988 46676 8990
rect 47964 12348 48020 12404
rect 47964 11506 48020 11508
rect 47964 11454 47966 11506
rect 47966 11454 48018 11506
rect 48018 11454 48020 11506
rect 47964 11452 48020 11454
rect 48300 11116 48356 11172
rect 48132 10610 48188 10612
rect 48132 10558 48134 10610
rect 48134 10558 48186 10610
rect 48186 10558 48188 10610
rect 48132 10556 48188 10558
rect 47628 10108 47684 10164
rect 47572 9772 47628 9828
rect 47292 8988 47348 9044
rect 43932 6748 43988 6804
rect 43372 6300 43428 6356
rect 43820 6636 43876 6692
rect 44044 6690 44100 6692
rect 44044 6638 44046 6690
rect 44046 6638 44098 6690
rect 44098 6638 44100 6690
rect 44044 6636 44100 6638
rect 45052 7362 45108 7364
rect 45052 7310 45054 7362
rect 45054 7310 45106 7362
rect 45106 7310 45108 7362
rect 45052 7308 45108 7310
rect 44940 7084 44996 7140
rect 44716 6748 44772 6804
rect 42924 5516 42980 5572
rect 43820 5234 43876 5236
rect 43820 5182 43822 5234
rect 43822 5182 43874 5234
rect 43874 5182 43876 5234
rect 43820 5180 43876 5182
rect 43372 5068 43428 5124
rect 43932 5107 43988 5124
rect 43932 5068 43934 5107
rect 43934 5068 43986 5107
rect 43986 5068 43988 5107
rect 44996 6466 45052 6468
rect 44996 6414 44998 6466
rect 44998 6414 45050 6466
rect 45050 6414 45052 6466
rect 44996 6412 45052 6414
rect 44716 5180 44772 5236
rect 43148 4956 43204 5012
rect 43708 4396 43764 4452
rect 42588 3836 42644 3892
rect 41692 3554 41748 3556
rect 41692 3502 41694 3554
rect 41694 3502 41746 3554
rect 41746 3502 41748 3554
rect 41692 3500 41748 3502
rect 42476 3554 42532 3556
rect 42476 3502 42478 3554
rect 42478 3502 42530 3554
rect 42530 3502 42532 3554
rect 42476 3500 42532 3502
rect 43484 4226 43540 4228
rect 43484 4174 43486 4226
rect 43486 4174 43538 4226
rect 43538 4174 43540 4226
rect 43484 4172 43540 4174
rect 42700 3612 42756 3668
rect 43092 3666 43148 3668
rect 43092 3614 43094 3666
rect 43094 3614 43146 3666
rect 43146 3614 43148 3666
rect 44044 3724 44100 3780
rect 43092 3612 43148 3614
rect 43708 3554 43764 3556
rect 43708 3502 43710 3554
rect 43710 3502 43762 3554
rect 43762 3502 43764 3554
rect 43708 3500 43764 3502
rect 45612 6690 45668 6692
rect 45612 6638 45614 6690
rect 45614 6638 45666 6690
rect 45666 6638 45668 6690
rect 45612 6636 45668 6638
rect 45500 6412 45556 6468
rect 45724 6412 45780 6468
rect 45892 6188 45948 6244
rect 45810 5887 45812 5908
rect 45812 5887 45864 5908
rect 45864 5887 45866 5908
rect 45810 5852 45866 5887
rect 45388 5516 45444 5572
rect 45388 5292 45444 5348
rect 44940 5068 44996 5124
rect 45948 5180 46004 5236
rect 46284 6972 46340 7028
rect 46396 6690 46452 6692
rect 46396 6638 46398 6690
rect 46398 6638 46450 6690
rect 46450 6638 46452 6690
rect 46396 6636 46452 6638
rect 46396 6412 46452 6468
rect 47068 7084 47124 7140
rect 47516 7362 47572 7364
rect 47516 7310 47518 7362
rect 47518 7310 47570 7362
rect 47570 7310 47572 7362
rect 47516 7308 47572 7310
rect 47404 6972 47460 7028
rect 47404 6188 47460 6244
rect 47292 5852 47348 5908
rect 45052 3836 45108 3892
rect 47516 5234 47572 5236
rect 47516 5182 47518 5234
rect 47518 5182 47570 5234
rect 47570 5182 47572 5234
rect 47516 5180 47572 5182
rect 48636 17500 48692 17556
rect 47964 6860 48020 6916
rect 48300 8092 48356 8148
rect 48300 7644 48356 7700
rect 45332 3666 45388 3668
rect 45332 3614 45334 3666
rect 45334 3614 45386 3666
rect 45386 3614 45388 3666
rect 45332 3612 45388 3614
rect 46060 3948 46116 4004
rect 47460 3724 47516 3780
rect 46676 3666 46732 3668
rect 46676 3614 46678 3666
rect 46678 3614 46730 3666
rect 46730 3614 46732 3666
rect 46676 3612 46732 3614
rect 47572 3666 47628 3668
rect 47572 3614 47574 3666
rect 47574 3614 47626 3666
rect 47626 3614 47628 3666
rect 47572 3612 47628 3614
rect 48020 3666 48076 3668
rect 48020 3614 48022 3666
rect 48022 3614 48074 3666
rect 48074 3614 48076 3666
rect 48020 3612 48076 3614
rect 48300 3612 48356 3668
rect 46228 3500 46284 3556
rect 28924 2716 28980 2772
<< metal3 >>
rect 49200 47124 50000 47152
rect 33628 47068 50000 47124
rect 33628 47012 33684 47068
rect 49200 47040 50000 47068
rect 30146 46956 30156 47012
rect 30212 46956 33684 47012
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 30258 46060 30268 46116
rect 30324 46060 33180 46116
rect 33236 46060 33246 46116
rect 33394 46060 33404 46116
rect 33460 46060 36988 46116
rect 37044 46060 37054 46116
rect 38098 46060 38108 46116
rect 38164 46060 40796 46116
rect 40852 46060 40862 46116
rect 6850 45836 6860 45892
rect 6916 45836 7308 45892
rect 7364 45836 7374 45892
rect 20066 45836 20076 45892
rect 20132 45836 24780 45892
rect 24836 45836 24846 45892
rect 29698 45836 29708 45892
rect 29764 45836 30268 45892
rect 30324 45836 30334 45892
rect 30930 45836 30940 45892
rect 30996 45836 32172 45892
rect 32228 45836 32238 45892
rect 35018 45836 35028 45892
rect 35084 45836 38668 45892
rect 38724 45836 38734 45892
rect 41122 45836 41132 45892
rect 41188 45836 46284 45892
rect 46340 45836 46350 45892
rect 11834 45724 11844 45780
rect 11900 45724 14588 45780
rect 14644 45724 14654 45780
rect 17490 45724 17500 45780
rect 17556 45724 24332 45780
rect 24388 45724 24398 45780
rect 27122 45724 27132 45780
rect 27188 45724 31444 45780
rect 31500 45724 31510 45780
rect 33618 45724 33628 45780
rect 33684 45724 39172 45780
rect 39228 45724 39238 45780
rect 40450 45724 40460 45780
rect 40516 45724 42980 45780
rect 43036 45724 43046 45780
rect 2370 45612 2380 45668
rect 2436 45612 3108 45668
rect 3164 45612 4564 45668
rect 4620 45612 4630 45668
rect 6682 45612 6692 45668
rect 6748 45612 9212 45668
rect 9268 45612 9828 45668
rect 9884 45612 9894 45668
rect 17154 45612 17164 45668
rect 17220 45612 18508 45668
rect 18564 45612 18574 45668
rect 26002 45612 26012 45668
rect 26068 45612 26796 45668
rect 26852 45612 26862 45668
rect 35298 45612 35308 45668
rect 35364 45612 36652 45668
rect 36708 45612 36718 45668
rect 6290 45500 6300 45556
rect 6356 45500 8260 45556
rect 8316 45500 12236 45556
rect 12292 45500 12302 45556
rect 27234 45500 27244 45556
rect 27300 45500 29204 45556
rect 29260 45500 29270 45556
rect 36390 45500 36428 45556
rect 36484 45500 37884 45556
rect 37940 45500 39788 45556
rect 39844 45500 39854 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 4554 45388 4564 45444
rect 4620 45388 6188 45444
rect 6244 45388 6254 45444
rect 9762 45388 9772 45444
rect 9828 45388 10556 45444
rect 10612 45388 10622 45444
rect 12674 45388 12684 45444
rect 12740 45388 13916 45444
rect 13972 45388 13982 45444
rect 28354 45388 28364 45444
rect 28420 45388 29988 45444
rect 30044 45388 30054 45444
rect 35074 45388 35084 45444
rect 35140 45388 35980 45444
rect 36036 45388 36046 45444
rect 37650 45388 37660 45444
rect 37716 45388 38892 45444
rect 38948 45388 38958 45444
rect 41346 45388 41356 45444
rect 41412 45388 43260 45444
rect 43316 45388 43326 45444
rect 46778 45388 46788 45444
rect 46844 45388 47516 45444
rect 47572 45388 47582 45444
rect 4442 45276 4452 45332
rect 4508 45276 5012 45332
rect 5068 45276 5078 45332
rect 36530 45276 36540 45332
rect 36596 45276 37996 45332
rect 38052 45276 38062 45332
rect 41234 45276 41244 45332
rect 41300 45276 44604 45332
rect 44660 45276 44670 45332
rect 2650 45164 2660 45220
rect 2716 45164 27580 45220
rect 27636 45164 46172 45220
rect 46228 45164 46238 45220
rect 9202 45052 9212 45108
rect 9268 45052 10332 45108
rect 10388 45052 10398 45108
rect 12338 45052 12348 45108
rect 12404 45052 15484 45108
rect 15540 45052 15550 45108
rect 16258 45052 16268 45108
rect 16324 45052 17500 45108
rect 17556 45052 17566 45108
rect 20738 45052 20748 45108
rect 20804 45052 21756 45108
rect 21812 45052 21822 45108
rect 25218 45052 25228 45108
rect 25284 45052 29708 45108
rect 29764 45052 32732 45108
rect 32788 45052 33068 45108
rect 33124 45052 33134 45108
rect 42242 45052 42252 45108
rect 42308 45052 42588 45108
rect 42644 45052 45388 45108
rect 45444 45052 45454 45108
rect 3714 44940 3724 44996
rect 3780 44940 4004 44996
rect 4060 44940 4900 44996
rect 4956 44940 13916 44996
rect 13972 44940 13982 44996
rect 16930 44940 16940 44996
rect 16996 44940 18060 44996
rect 18116 44940 18126 44996
rect 19618 44940 19628 44996
rect 19684 44940 19964 44996
rect 20020 44940 20030 44996
rect 27906 44940 27916 44996
rect 27972 44940 28252 44996
rect 28308 44940 29148 44996
rect 29204 44940 29214 44996
rect 36642 44940 36652 44996
rect 36708 44940 37324 44996
rect 37380 44940 37390 44996
rect 40338 44940 40348 44996
rect 40404 44940 40852 44996
rect 40908 44940 40918 44996
rect 3546 44828 3556 44884
rect 3612 44828 9380 44884
rect 12786 44828 12796 44884
rect 12852 44828 15596 44884
rect 15652 44828 15662 44884
rect 16594 44828 16604 44884
rect 16660 44828 21308 44884
rect 21364 44828 21374 44884
rect 37202 44828 37212 44884
rect 37268 44828 41244 44884
rect 41300 44828 42700 44884
rect 42756 44828 42766 44884
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 9324 44660 9380 44828
rect 39004 44772 39060 44828
rect 13458 44716 13468 44772
rect 13524 44716 16548 44772
rect 17658 44716 17668 44772
rect 17724 44716 26908 44772
rect 26964 44716 27804 44772
rect 27860 44716 27870 44772
rect 38994 44716 39004 44772
rect 39060 44716 39070 44772
rect 16492 44660 16548 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 9324 44604 15148 44660
rect 15204 44604 15214 44660
rect 16492 44604 17948 44660
rect 18004 44604 18014 44660
rect 26852 44604 27020 44660
rect 27076 44604 28868 44660
rect 28924 44604 28934 44660
rect 26852 44548 26908 44604
rect 20850 44492 20860 44548
rect 20916 44492 22316 44548
rect 22372 44492 22382 44548
rect 22530 44492 22540 44548
rect 22596 44492 25004 44548
rect 25060 44492 25070 44548
rect 26226 44492 26236 44548
rect 26292 44492 26908 44548
rect 30482 44492 30492 44548
rect 30548 44492 35756 44548
rect 35812 44492 35822 44548
rect 39666 44492 39676 44548
rect 39732 44492 40908 44548
rect 40964 44492 40974 44548
rect 42802 44492 42812 44548
rect 42868 44492 45612 44548
rect 45668 44492 45678 44548
rect 9090 44380 9100 44436
rect 9156 44380 9436 44436
rect 9492 44380 9502 44436
rect 25890 44380 25900 44436
rect 25956 44380 27244 44436
rect 27300 44380 27310 44436
rect 41458 44380 41468 44436
rect 41524 44380 41804 44436
rect 41860 44380 43260 44436
rect 43316 44380 46396 44436
rect 46452 44380 46462 44436
rect 8418 44268 8428 44324
rect 8484 44268 9660 44324
rect 9716 44268 9726 44324
rect 9986 44268 9996 44324
rect 10052 44268 11004 44324
rect 11060 44268 11070 44324
rect 13010 44268 13020 44324
rect 13076 44268 13580 44324
rect 13636 44268 13646 44324
rect 23090 44268 23100 44324
rect 23156 44268 24220 44324
rect 24276 44268 24286 44324
rect 25330 44268 25340 44324
rect 25396 44268 28196 44324
rect 28252 44268 28262 44324
rect 35541 44268 35551 44324
rect 35607 44268 36428 44324
rect 36484 44268 36494 44324
rect 43754 44268 43764 44324
rect 43820 44268 44268 44324
rect 44324 44268 44940 44324
rect 44996 44268 45006 44324
rect 20626 44156 20636 44212
rect 20692 44156 26908 44212
rect 27794 44156 27804 44212
rect 27860 44156 30735 44212
rect 30791 44156 31836 44212
rect 31892 44156 31902 44212
rect 35298 44156 35308 44212
rect 35364 44156 37436 44212
rect 37492 44156 37502 44212
rect 4722 44044 4732 44100
rect 4788 44044 5964 44100
rect 6020 44044 6030 44100
rect 7074 44044 7084 44100
rect 7140 44044 7980 44100
rect 8036 44044 8046 44100
rect 19394 44044 19404 44100
rect 19460 44044 25228 44100
rect 25284 44044 25294 44100
rect 26852 43988 26908 44156
rect 27906 44044 27916 44100
rect 27972 44044 28364 44100
rect 28420 44044 30716 44100
rect 30772 44044 30782 44100
rect 38789 44044 38799 44100
rect 38855 44044 39900 44100
rect 39956 44044 41020 44100
rect 41076 44044 41086 44100
rect 42130 44044 42140 44100
rect 42196 44044 44100 44100
rect 44156 44044 44166 44100
rect 4274 43932 4284 43988
rect 4340 43932 7812 43988
rect 9986 43932 9996 43988
rect 10052 43932 10780 43988
rect 10836 43932 10846 43988
rect 26852 43932 47852 43988
rect 47908 43932 47918 43988
rect 5842 43820 5852 43876
rect 5908 43820 5918 43876
rect 5852 43764 5908 43820
rect 4946 43708 4956 43764
rect 5012 43708 6412 43764
rect 6468 43708 6478 43764
rect 3042 43596 3052 43652
rect 3108 43596 4060 43652
rect 4116 43596 4126 43652
rect 4386 43596 4396 43652
rect 4452 43596 7084 43652
rect 7140 43596 7150 43652
rect 7756 43540 7812 43932
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 14886 43820 14924 43876
rect 14980 43820 14990 43876
rect 20402 43820 20412 43876
rect 20468 43820 21644 43876
rect 21700 43820 21710 43876
rect 27570 43820 27580 43876
rect 27636 43820 43036 43876
rect 43092 43820 43102 43876
rect 47170 43820 47180 43876
rect 47236 43820 47404 43876
rect 47460 43820 47470 43876
rect 8530 43708 8540 43764
rect 8596 43708 10668 43764
rect 10724 43708 10734 43764
rect 17826 43708 17836 43764
rect 17892 43708 19292 43764
rect 19348 43708 19358 43764
rect 20514 43708 20524 43764
rect 20580 43708 20590 43764
rect 30482 43708 30492 43764
rect 30548 43708 30558 43764
rect 30706 43708 30716 43764
rect 30772 43708 48020 43764
rect 48076 43708 48086 43764
rect 20524 43652 20580 43708
rect 30492 43652 30548 43708
rect 13570 43596 13580 43652
rect 13636 43596 14140 43652
rect 14196 43596 15932 43652
rect 15988 43596 15998 43652
rect 17658 43596 17668 43652
rect 17724 43596 20580 43652
rect 21084 43596 27804 43652
rect 27860 43596 27870 43652
rect 29922 43596 29932 43652
rect 29988 43596 30716 43652
rect 30772 43596 30782 43652
rect 34962 43596 34972 43652
rect 35028 43596 36204 43652
rect 36260 43596 36270 43652
rect 36418 43596 36428 43652
rect 36484 43596 38052 43652
rect 38108 43596 38118 43652
rect 45042 43596 45052 43652
rect 45108 43596 46396 43652
rect 46452 43596 48188 43652
rect 48244 43596 48254 43652
rect 5058 43484 5068 43540
rect 5124 43484 7420 43540
rect 7476 43484 7486 43540
rect 7746 43484 7756 43540
rect 7812 43484 8876 43540
rect 8932 43484 8942 43540
rect 10210 43484 10220 43540
rect 10276 43484 11004 43540
rect 11060 43484 11070 43540
rect 13438 43484 13448 43540
rect 13504 43484 14476 43540
rect 14532 43484 14542 43540
rect 15026 43484 15036 43540
rect 1866 43372 1876 43428
rect 1932 43372 14588 43428
rect 14644 43372 14654 43428
rect 15092 43316 15148 43540
rect 16370 43484 16380 43540
rect 16436 43484 16716 43540
rect 16772 43484 16884 43540
rect 16940 43484 16950 43540
rect 20514 43484 20524 43540
rect 20580 43484 20860 43540
rect 20916 43484 20926 43540
rect 21084 43316 21140 43596
rect 22978 43484 22988 43540
rect 23044 43484 25900 43540
rect 25956 43484 25966 43540
rect 26786 43484 26796 43540
rect 26852 43484 27356 43540
rect 27412 43484 27422 43540
rect 27682 43484 27692 43540
rect 27748 43484 28252 43540
rect 28308 43484 29260 43540
rect 29316 43484 29326 43540
rect 30146 43484 30156 43540
rect 30212 43484 31276 43540
rect 31332 43484 31612 43540
rect 31668 43484 31678 43540
rect 31972 43484 31982 43540
rect 32038 43484 33068 43540
rect 33124 43484 33134 43540
rect 36642 43484 36652 43540
rect 36708 43484 37884 43540
rect 37940 43484 37950 43540
rect 38546 43484 38556 43540
rect 38612 43484 42476 43540
rect 42532 43484 42542 43540
rect 43474 43484 43484 43540
rect 43540 43484 44940 43540
rect 44996 43484 48300 43540
rect 48356 43484 48366 43540
rect 23538 43372 23548 43428
rect 23604 43372 24612 43428
rect 29642 43372 29652 43428
rect 29708 43372 33740 43428
rect 33796 43372 33806 43428
rect 34066 43372 34076 43428
rect 34132 43372 42700 43428
rect 42756 43372 45052 43428
rect 45108 43372 45118 43428
rect 24556 43316 24612 43372
rect 3658 43260 3668 43316
rect 3724 43260 5180 43316
rect 5236 43260 10052 43316
rect 13906 43260 13916 43316
rect 13972 43260 14252 43316
rect 14308 43260 14318 43316
rect 15092 43260 21140 43316
rect 21970 43260 21980 43316
rect 22036 43260 22876 43316
rect 22932 43260 23436 43316
rect 23492 43260 23502 43316
rect 24546 43260 24556 43316
rect 24612 43260 24622 43316
rect 26852 43260 28232 43316
rect 28288 43260 28476 43316
rect 28532 43260 28542 43316
rect 30342 43260 30380 43316
rect 30436 43260 30446 43316
rect 32386 43260 32396 43316
rect 32452 43260 34412 43316
rect 34468 43260 34478 43316
rect 9996 43204 10052 43260
rect 26852 43204 26908 43260
rect 7074 43148 7084 43204
rect 7140 43148 7868 43204
rect 7924 43148 8764 43204
rect 8820 43148 8830 43204
rect 9986 43148 9996 43204
rect 10052 43148 10220 43204
rect 10276 43148 10286 43204
rect 13682 43148 13692 43204
rect 13748 43148 26908 43204
rect 27804 43148 28084 43204
rect 28140 43148 28150 43204
rect 29932 43148 30492 43204
rect 30548 43148 30558 43204
rect 33058 43148 33068 43204
rect 33124 43148 33852 43204
rect 33908 43148 33918 43204
rect 40226 43148 40236 43204
rect 40292 43148 42420 43204
rect 42476 43148 47180 43204
rect 47236 43148 47246 43204
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 4946 43036 4956 43092
rect 5012 43036 5684 43092
rect 5740 43036 5750 43092
rect 6374 43036 6412 43092
rect 6468 43036 6478 43092
rect 8978 43036 8988 43092
rect 9044 43036 9660 43092
rect 9716 43036 10556 43092
rect 10612 43036 14756 43092
rect 14812 43036 14822 43092
rect 14914 43036 14924 43092
rect 14980 43036 15036 43092
rect 15092 43036 15102 43092
rect 20234 43036 20244 43092
rect 20300 43036 21868 43092
rect 21924 43036 22652 43092
rect 22708 43036 23660 43092
rect 23716 43036 23726 43092
rect 27804 42980 27860 43148
rect 29932 42980 29988 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 30706 43036 30716 43092
rect 30772 43036 31948 43092
rect 32004 43036 32014 43092
rect 33282 43036 33292 43092
rect 33348 43036 34188 43092
rect 34244 43036 34254 43092
rect 42242 43036 42252 43092
rect 42308 43036 47740 43092
rect 47796 43036 47806 43092
rect 2594 42924 2604 42980
rect 2660 42924 2670 42980
rect 2762 42924 2772 42980
rect 2828 42924 19460 42980
rect 20066 42924 20076 42980
rect 20132 42924 21420 42980
rect 21476 42924 21756 42980
rect 21812 42924 22316 42980
rect 22372 42924 27860 42980
rect 28466 42924 28476 42980
rect 28532 42924 29988 42980
rect 30818 42924 30828 42980
rect 30884 42924 32452 42980
rect 32508 42924 32518 42980
rect 33730 42924 33740 42980
rect 33796 42924 34748 42980
rect 34804 42924 34814 42980
rect 44594 42924 44604 42980
rect 44660 42924 45836 42980
rect 45892 42924 45902 42980
rect 2604 42868 2660 42924
rect 2604 42812 5292 42868
rect 5348 42812 6524 42868
rect 6580 42812 11340 42868
rect 11396 42812 11676 42868
rect 11732 42812 11742 42868
rect 12450 42812 12460 42868
rect 12516 42812 13580 42868
rect 13636 42812 13646 42868
rect 14914 42812 14924 42868
rect 14980 42812 16156 42868
rect 16212 42812 17500 42868
rect 17556 42812 17566 42868
rect 12002 42700 12012 42756
rect 12068 42700 12572 42756
rect 12628 42700 12638 42756
rect 12898 42700 12908 42756
rect 12964 42700 13804 42756
rect 13860 42700 15036 42756
rect 15092 42700 15102 42756
rect 16370 42700 16380 42756
rect 16436 42700 17164 42756
rect 17220 42700 17230 42756
rect 17378 42700 17388 42756
rect 17444 42700 18004 42756
rect 18060 42700 18070 42756
rect 12572 42644 12628 42700
rect 12572 42588 13916 42644
rect 13972 42588 14700 42644
rect 14756 42588 14766 42644
rect 15418 42588 15428 42644
rect 15484 42588 15932 42644
rect 15988 42588 16268 42644
rect 16324 42588 17724 42644
rect 17780 42588 17790 42644
rect 19404 42532 19460 42924
rect 21522 42812 21532 42868
rect 21588 42812 21980 42868
rect 22036 42812 22046 42868
rect 29932 42756 29988 42924
rect 35410 42812 35420 42868
rect 35476 42812 35644 42868
rect 35700 42812 35710 42868
rect 41122 42812 41132 42868
rect 41188 42812 41580 42868
rect 41636 42812 41646 42868
rect 44146 42812 44156 42868
rect 44212 42812 48076 42868
rect 48132 42812 48142 42868
rect 19730 42700 19740 42756
rect 19796 42700 19964 42756
rect 20020 42700 20030 42756
rect 22138 42700 22148 42756
rect 22204 42700 23212 42756
rect 23268 42700 23278 42756
rect 25442 42700 25452 42756
rect 25508 42700 25900 42756
rect 25956 42700 25966 42756
rect 29922 42700 29932 42756
rect 29988 42700 29998 42756
rect 32162 42700 32172 42756
rect 32228 42700 32620 42756
rect 32676 42700 38668 42756
rect 38612 42644 38668 42700
rect 19562 42588 19572 42644
rect 19628 42588 20524 42644
rect 20580 42588 21756 42644
rect 21812 42588 21822 42644
rect 29026 42588 29036 42644
rect 29092 42588 31724 42644
rect 31780 42588 31790 42644
rect 31938 42588 31948 42644
rect 32004 42588 37548 42644
rect 37604 42588 37614 42644
rect 38612 42588 43708 42644
rect 43764 42588 43774 42644
rect 43932 42532 43988 42756
rect 44044 42700 44054 42756
rect 47394 42700 47404 42756
rect 47460 42700 47740 42756
rect 47796 42700 47806 42756
rect 1474 42476 1484 42532
rect 1540 42476 1932 42532
rect 1988 42476 1998 42532
rect 3938 42476 3948 42532
rect 4004 42476 4676 42532
rect 4732 42476 5964 42532
rect 6020 42476 6030 42532
rect 19404 42476 21364 42532
rect 21522 42476 21532 42532
rect 21588 42476 22484 42532
rect 22540 42476 22988 42532
rect 23044 42476 23054 42532
rect 29362 42476 29372 42532
rect 29428 42476 40908 42532
rect 40964 42476 40974 42532
rect 43474 42476 43484 42532
rect 43540 42476 43988 42532
rect 10098 42364 10108 42420
rect 10164 42364 10174 42420
rect 700 42140 1596 42196
rect 1652 42140 1662 42196
rect 3210 42140 3220 42196
rect 3276 42140 3388 42196
rect 700 41748 756 42140
rect 3332 42084 3388 42140
rect 10108 42084 10164 42364
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 21308 42308 21364 42476
rect 26852 42364 33740 42420
rect 33796 42364 38668 42420
rect 39218 42364 39228 42420
rect 39284 42364 40236 42420
rect 40292 42364 40302 42420
rect 26852 42308 26908 42364
rect 38612 42308 38668 42364
rect 21308 42252 24892 42308
rect 24948 42252 26908 42308
rect 28578 42252 28588 42308
rect 28644 42252 30808 42308
rect 30864 42252 32284 42308
rect 32340 42252 32350 42308
rect 34402 42252 34412 42308
rect 34468 42252 38108 42308
rect 38164 42252 38174 42308
rect 38612 42252 44492 42308
rect 44548 42252 44558 42308
rect 49200 42196 50000 42224
rect 28690 42140 28700 42196
rect 28756 42140 30156 42196
rect 30212 42140 31948 42196
rect 32004 42140 32014 42196
rect 34290 42140 34300 42196
rect 34356 42140 37380 42196
rect 37436 42140 37446 42196
rect 37538 42140 37548 42196
rect 37604 42140 50000 42196
rect 49200 42112 50000 42140
rect 3332 42028 6580 42084
rect 8922 42028 8932 42084
rect 8988 42028 10388 42084
rect 6524 41972 6580 42028
rect 10332 41972 10388 42028
rect 16492 42028 16716 42084
rect 16772 42028 16782 42084
rect 16874 42028 16884 42084
rect 16940 42028 17164 42084
rect 17220 42028 17230 42084
rect 26562 42028 26572 42084
rect 26628 42028 26796 42084
rect 26852 42028 26862 42084
rect 35942 42028 35980 42084
rect 36036 42028 36046 42084
rect 36642 42028 36652 42084
rect 36708 42028 36876 42084
rect 36932 42028 36942 42084
rect 37090 42028 37100 42084
rect 37156 42028 37996 42084
rect 38052 42028 38062 42084
rect 38546 42028 38556 42084
rect 38612 42028 39452 42084
rect 39508 42028 39518 42084
rect 40002 42028 40012 42084
rect 40068 42028 41804 42084
rect 41860 42028 41870 42084
rect 16492 41972 16548 42028
rect 36652 41972 36708 42028
rect 4274 41916 4284 41972
rect 4340 41916 5964 41972
rect 6020 41916 6300 41972
rect 6356 41916 6366 41972
rect 6524 41916 7700 41972
rect 7756 41916 7766 41972
rect 8194 41916 8204 41972
rect 8260 41916 8764 41972
rect 8820 41916 8830 41972
rect 10294 41916 10332 41972
rect 10388 41916 10398 41972
rect 11890 41916 11900 41972
rect 11956 41916 13076 41972
rect 14858 41916 14868 41972
rect 14924 41916 15894 41972
rect 15950 41916 15960 41972
rect 16482 41916 16492 41972
rect 16548 41916 16558 41972
rect 21858 41916 21868 41972
rect 21924 41916 22764 41972
rect 22820 41916 23324 41972
rect 23380 41916 23390 41972
rect 24434 41916 24444 41972
rect 24500 41916 26236 41972
rect 26292 41916 27188 41972
rect 27244 41916 27254 41972
rect 28802 41916 28812 41972
rect 28868 41916 29484 41972
rect 29540 41916 29550 41972
rect 35838 41916 35848 41972
rect 35904 41916 36652 41972
rect 36708 41916 36718 41972
rect 37286 41916 37324 41972
rect 37380 41916 37390 41972
rect 37538 41916 37548 41972
rect 37604 41916 40796 41972
rect 40852 41916 42700 41972
rect 42756 41916 42766 41972
rect 43474 41916 43484 41972
rect 43540 41916 47516 41972
rect 47572 41916 47582 41972
rect 2594 41804 2604 41860
rect 2660 41804 5087 41860
rect 5143 41804 5153 41860
rect 6178 41804 6188 41860
rect 6244 41804 7084 41860
rect 7140 41804 7150 41860
rect 10546 41804 10556 41860
rect 10612 41804 11340 41860
rect 11396 41804 12796 41860
rect 12852 41804 12862 41860
rect 5087 41748 5143 41804
rect 700 41692 980 41748
rect 5087 41692 6860 41748
rect 6916 41692 6926 41748
rect 11890 41692 11900 41748
rect 11956 41692 12292 41748
rect 12348 41692 12358 41748
rect 0 41524 800 41552
rect 924 41524 980 41692
rect 6178 41580 6188 41636
rect 6244 41580 7532 41636
rect 7588 41580 7598 41636
rect 10882 41580 10892 41636
rect 10948 41580 11508 41636
rect 11564 41580 12012 41636
rect 12068 41580 12078 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 12796 41524 12852 41804
rect 13020 41636 13076 41916
rect 26094 41804 26104 41860
rect 26160 41804 27468 41860
rect 27524 41804 27804 41860
rect 27860 41804 27870 41860
rect 36082 41804 36092 41860
rect 36148 41804 36316 41860
rect 36372 41804 38220 41860
rect 38276 41804 38286 41860
rect 39218 41804 39228 41860
rect 39284 41804 39844 41860
rect 39900 41804 39910 41860
rect 44482 41804 44492 41860
rect 44548 41804 45724 41860
rect 45780 41804 45790 41860
rect 46050 41804 46060 41860
rect 46116 41804 46732 41860
rect 46788 41804 46798 41860
rect 15250 41692 15260 41748
rect 15316 41692 23436 41748
rect 23492 41692 23502 41748
rect 29474 41692 29484 41748
rect 29540 41692 30492 41748
rect 30548 41692 30558 41748
rect 34738 41692 34748 41748
rect 34804 41692 35588 41748
rect 36978 41692 36988 41748
rect 37044 41692 38444 41748
rect 38500 41692 38510 41748
rect 45266 41692 45276 41748
rect 45332 41692 45388 41748
rect 45444 41692 45454 41748
rect 35532 41636 35588 41692
rect 13010 41580 13020 41636
rect 13076 41580 13086 41636
rect 15138 41580 15148 41636
rect 15204 41580 15242 41636
rect 15362 41580 15372 41636
rect 15428 41580 16100 41636
rect 21522 41580 21532 41636
rect 21588 41580 22932 41636
rect 24770 41580 24780 41636
rect 24836 41580 26124 41636
rect 26180 41580 26908 41636
rect 26964 41580 26974 41636
rect 35532 41580 35644 41636
rect 35700 41580 37436 41636
rect 37492 41580 37502 41636
rect 37818 41580 37828 41636
rect 37884 41580 39228 41636
rect 39284 41580 39294 41636
rect 43922 41580 43932 41636
rect 43988 41580 47852 41636
rect 47908 41580 47918 41636
rect 16044 41524 16100 41580
rect 22876 41524 22932 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 0 41468 980 41524
rect 12796 41468 13580 41524
rect 13636 41468 13646 41524
rect 16034 41468 16044 41524
rect 16100 41468 16110 41524
rect 19506 41468 19516 41524
rect 19572 41468 22708 41524
rect 22764 41468 22774 41524
rect 22876 41468 27636 41524
rect 27692 41468 27702 41524
rect 29670 41468 29708 41524
rect 29764 41468 29774 41524
rect 36166 41468 36204 41524
rect 36260 41468 36270 41524
rect 38322 41468 38332 41524
rect 38388 41468 39564 41524
rect 39620 41468 39630 41524
rect 44492 41468 48076 41524
rect 48132 41468 48142 41524
rect 0 41440 800 41468
rect 44492 41412 44548 41468
rect 8922 41356 8932 41412
rect 8988 41356 9940 41412
rect 11778 41356 11788 41412
rect 11844 41356 12740 41412
rect 19618 41356 19628 41412
rect 19684 41356 19740 41412
rect 19796 41356 19806 41412
rect 20402 41356 20412 41412
rect 20468 41356 21644 41412
rect 21700 41356 26628 41412
rect 35914 41356 35924 41412
rect 35980 41356 36764 41412
rect 36820 41356 36830 41412
rect 43586 41356 43596 41412
rect 43652 41356 44492 41412
rect 44548 41356 44558 41412
rect 1978 41244 1988 41300
rect 2044 41244 2604 41300
rect 2660 41244 2670 41300
rect 9884 41188 9940 41356
rect 12684 41300 12740 41356
rect 10658 41244 10668 41300
rect 10724 41244 12460 41300
rect 12516 41244 12526 41300
rect 12674 41244 12684 41300
rect 12740 41244 12750 41300
rect 23986 41244 23996 41300
rect 24052 41244 25452 41300
rect 25508 41244 25518 41300
rect 26572 41188 26628 41356
rect 35522 41244 35532 41300
rect 35588 41244 46060 41300
rect 46116 41244 46126 41300
rect 2706 41132 2716 41188
rect 2772 41132 3388 41188
rect 3444 41132 3454 41188
rect 6972 41132 7868 41188
rect 7924 41132 7934 41188
rect 8082 41132 8092 41188
rect 8148 41132 8158 41188
rect 9874 41132 9884 41188
rect 9940 41132 9950 41188
rect 10882 41132 10892 41188
rect 10948 41132 11564 41188
rect 11620 41132 11630 41188
rect 15586 41132 15596 41188
rect 15652 41132 16716 41188
rect 16772 41132 16782 41188
rect 17490 41132 17500 41188
rect 17556 41132 19404 41188
rect 19460 41132 22876 41188
rect 22932 41132 22942 41188
rect 23202 41132 23212 41188
rect 23268 41132 23828 41188
rect 23884 41132 23894 41188
rect 25106 41132 25116 41188
rect 25172 41132 26348 41188
rect 26404 41132 26414 41188
rect 26562 41132 26572 41188
rect 26628 41132 26638 41188
rect 29586 41132 29596 41188
rect 29652 41132 30696 41188
rect 30752 41132 30762 41188
rect 30930 41132 30940 41188
rect 30996 41132 32264 41188
rect 32320 41132 32330 41188
rect 36194 41132 36204 41188
rect 36260 41132 36988 41188
rect 37044 41132 37054 41188
rect 37202 41132 37212 41188
rect 37268 41132 37324 41188
rect 37380 41132 37390 41188
rect 37538 41132 37548 41188
rect 37604 41132 38108 41188
rect 38164 41132 38174 41188
rect 38742 41132 38780 41188
rect 38836 41132 38846 41188
rect 41458 41132 41468 41188
rect 41524 41132 42196 41188
rect 42252 41132 42262 41188
rect 42466 41132 42476 41188
rect 42532 41132 43932 41188
rect 43988 41132 43998 41188
rect 44790 41132 44828 41188
rect 44884 41132 44894 41188
rect 6972 40964 7028 41132
rect 8092 41076 8148 41132
rect 7746 41020 7756 41076
rect 7812 41020 8764 41076
rect 8820 41020 8830 41076
rect 11638 41020 11676 41076
rect 11732 41020 11742 41076
rect 11974 41020 12012 41076
rect 12068 41020 12078 41076
rect 13906 41020 13916 41076
rect 13972 41020 15800 41076
rect 15856 41020 15866 41076
rect 17836 40964 17892 41132
rect 21970 41020 21980 41076
rect 22036 41020 22428 41076
rect 22484 41020 23548 41076
rect 23604 41020 23614 41076
rect 37398 41020 37436 41076
rect 37492 41020 37502 41076
rect 41794 41020 41804 41076
rect 41860 41020 43372 41076
rect 43428 41020 43438 41076
rect 43596 41020 45724 41076
rect 45780 41020 47516 41076
rect 47572 41020 47582 41076
rect 43596 40964 43652 41020
rect 6962 40908 6972 40964
rect 7028 40908 7038 40964
rect 17826 40908 17836 40964
rect 17892 40908 17902 40964
rect 18060 40908 28140 40964
rect 28196 40908 28206 40964
rect 29362 40908 29372 40964
rect 29428 40908 31052 40964
rect 31108 40908 31118 40964
rect 32274 40908 32284 40964
rect 32340 40908 42364 40964
rect 42420 40908 42430 40964
rect 42578 40908 42588 40964
rect 42644 40908 43596 40964
rect 43652 40908 43662 40964
rect 45042 40908 45052 40964
rect 45108 40908 45388 40964
rect 45444 40908 45836 40964
rect 45892 40908 45902 40964
rect 46050 40908 46060 40964
rect 46116 40908 46154 40964
rect 18060 40852 18116 40908
rect 32284 40852 32340 40908
rect 10892 40796 12796 40852
rect 12852 40796 12862 40852
rect 14700 40796 18116 40852
rect 26852 40796 32340 40852
rect 32396 40796 42924 40852
rect 42980 40796 42990 40852
rect 43810 40796 43820 40852
rect 43876 40796 46396 40852
rect 46452 40796 47740 40852
rect 47796 40796 47806 40852
rect 2874 40684 2884 40740
rect 2940 40684 6412 40740
rect 6468 40684 6478 40740
rect 10892 40628 10948 40796
rect 14700 40740 14756 40796
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 26852 40740 26908 40796
rect 32396 40740 32452 40796
rect 11218 40684 11228 40740
rect 11284 40684 11676 40740
rect 11732 40684 12908 40740
rect 12964 40684 13132 40740
rect 13188 40684 13198 40740
rect 14130 40684 14140 40740
rect 14196 40684 14456 40740
rect 14512 40684 14522 40740
rect 14690 40684 14700 40740
rect 14756 40684 14766 40740
rect 23314 40684 23324 40740
rect 23380 40684 26908 40740
rect 27122 40684 27132 40740
rect 27188 40684 27448 40740
rect 27504 40684 27514 40740
rect 28130 40684 28140 40740
rect 28196 40684 28680 40740
rect 28736 40684 28746 40740
rect 29810 40684 29820 40740
rect 29876 40684 32452 40740
rect 33842 40684 33852 40740
rect 33908 40684 42756 40740
rect 42812 40684 42822 40740
rect 43642 40684 43652 40740
rect 43708 40684 45836 40740
rect 45892 40684 45902 40740
rect 46060 40684 47404 40740
rect 47460 40684 47470 40740
rect 46060 40628 46116 40684
rect 3826 40572 3836 40628
rect 3892 40572 3902 40628
rect 6850 40572 6860 40628
rect 6916 40572 8204 40628
rect 8260 40572 9716 40628
rect 9772 40572 10164 40628
rect 10220 40572 10892 40628
rect 10948 40572 10958 40628
rect 12338 40572 12348 40628
rect 12404 40572 15148 40628
rect 15204 40572 15820 40628
rect 15876 40572 15886 40628
rect 17602 40572 17612 40628
rect 17668 40572 18620 40628
rect 18676 40572 18686 40628
rect 20906 40572 20916 40628
rect 20972 40572 21532 40628
rect 21588 40572 21598 40628
rect 24714 40572 24724 40628
rect 24780 40572 25788 40628
rect 25844 40572 25854 40628
rect 28802 40572 28812 40628
rect 28868 40572 31500 40628
rect 31556 40572 31566 40628
rect 34962 40572 34972 40628
rect 35028 40572 35084 40628
rect 35140 40572 38108 40628
rect 38164 40572 38332 40628
rect 38388 40572 38398 40628
rect 42354 40572 42364 40628
rect 42420 40572 42532 40628
rect 43474 40572 43484 40628
rect 43540 40572 43596 40628
rect 43652 40572 43662 40628
rect 44930 40572 44940 40628
rect 44996 40572 45276 40628
rect 45332 40572 45342 40628
rect 45500 40572 46116 40628
rect 46246 40572 46284 40628
rect 46340 40572 46350 40628
rect 3836 40516 3892 40572
rect 42476 40516 42532 40572
rect 45500 40516 45556 40572
rect 1978 40460 1988 40516
rect 2044 40460 4396 40516
rect 4452 40460 4462 40516
rect 5170 40460 5180 40516
rect 5236 40460 6244 40516
rect 6300 40460 8092 40516
rect 8148 40460 8596 40516
rect 8866 40460 8876 40516
rect 8932 40460 12572 40516
rect 12628 40460 12638 40516
rect 16594 40460 16604 40516
rect 16660 40460 18228 40516
rect 18284 40460 18294 40516
rect 28914 40460 28924 40516
rect 28980 40460 29932 40516
rect 29988 40460 30156 40516
rect 30212 40460 30222 40516
rect 30650 40460 30660 40516
rect 30716 40460 31388 40516
rect 31444 40460 31454 40516
rect 35644 40460 36708 40516
rect 36764 40460 36774 40516
rect 37650 40460 37660 40516
rect 37716 40460 39452 40516
rect 39508 40460 39518 40516
rect 39666 40460 39676 40516
rect 39732 40460 42252 40516
rect 42308 40460 42318 40516
rect 42476 40460 43372 40516
rect 43428 40460 45556 40516
rect 45714 40460 45724 40516
rect 45780 40460 46172 40516
rect 46228 40460 46238 40516
rect 46386 40460 46396 40516
rect 46452 40460 46490 40516
rect 46610 40460 46620 40516
rect 46676 40460 46732 40516
rect 46788 40460 46798 40516
rect 8540 40404 8596 40460
rect 35644 40404 35700 40460
rect 39676 40404 39732 40460
rect 2594 40348 2604 40404
rect 2660 40348 5348 40404
rect 5404 40348 5414 40404
rect 7522 40348 7532 40404
rect 7588 40348 8316 40404
rect 8372 40348 8382 40404
rect 8540 40348 8988 40404
rect 9044 40348 11452 40404
rect 11508 40348 11518 40404
rect 12898 40348 12908 40404
rect 12964 40348 13580 40404
rect 13636 40348 13646 40404
rect 16482 40348 16492 40404
rect 16548 40348 17276 40404
rect 17332 40348 17342 40404
rect 20290 40348 20300 40404
rect 20356 40348 20524 40404
rect 20580 40348 21308 40404
rect 21364 40348 21374 40404
rect 21578 40348 21588 40404
rect 21644 40348 22092 40404
rect 22148 40348 22820 40404
rect 22876 40348 22886 40404
rect 27514 40348 27524 40404
rect 27580 40348 29036 40404
rect 29092 40348 29102 40404
rect 29698 40348 29708 40404
rect 29820 40348 29830 40404
rect 30482 40348 30492 40404
rect 30548 40348 31780 40404
rect 31836 40348 31846 40404
rect 34850 40348 34860 40404
rect 34916 40348 35644 40404
rect 35700 40348 35710 40404
rect 36530 40348 36540 40404
rect 36596 40348 37828 40404
rect 37884 40348 37894 40404
rect 38322 40348 38332 40404
rect 38388 40348 39228 40404
rect 39284 40348 39732 40404
rect 41906 40348 41916 40404
rect 41972 40348 42476 40404
rect 42532 40348 42542 40404
rect 43372 40348 43932 40404
rect 43988 40348 43998 40404
rect 44156 40348 44380 40404
rect 44436 40348 44446 40404
rect 44566 40348 44604 40404
rect 44660 40348 44670 40404
rect 45602 40348 45612 40404
rect 45668 40348 46508 40404
rect 46564 40348 47124 40404
rect 47180 40348 47190 40404
rect 1810 40236 1820 40292
rect 1876 40236 2436 40292
rect 2492 40236 2502 40292
rect 3378 40236 3388 40292
rect 3444 40236 4004 40292
rect 4060 40236 4070 40292
rect 4162 40236 4172 40292
rect 4228 40236 5852 40292
rect 5908 40236 5918 40292
rect 11330 40236 11340 40292
rect 11396 40236 12124 40292
rect 12180 40236 12190 40292
rect 21410 40236 21420 40292
rect 21476 40236 22204 40292
rect 22260 40236 22270 40292
rect 25666 40236 25676 40292
rect 25732 40236 26964 40292
rect 27020 40236 27030 40292
rect 36194 40236 36204 40292
rect 36260 40236 38780 40292
rect 38836 40236 38846 40292
rect 43372 40180 43428 40348
rect 44156 40180 44212 40348
rect 19282 40124 19292 40180
rect 19348 40124 22316 40180
rect 22372 40124 22382 40180
rect 25330 40124 25340 40180
rect 25396 40124 25788 40180
rect 25844 40124 26684 40180
rect 26740 40124 26750 40180
rect 35410 40124 35420 40180
rect 35476 40124 36652 40180
rect 36708 40124 38220 40180
rect 38276 40124 38286 40180
rect 43362 40124 43372 40180
rect 43428 40124 43438 40180
rect 43922 40124 43932 40180
rect 43988 40124 44212 40180
rect 27458 40012 27468 40068
rect 27524 40012 29148 40068
rect 29204 40012 31276 40068
rect 31332 40012 31342 40068
rect 37874 40012 37884 40068
rect 37940 40012 41412 40068
rect 41514 40012 41524 40068
rect 41580 40012 42364 40068
rect 42420 40012 42430 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 41356 39956 41412 40012
rect 14242 39900 14252 39956
rect 14308 39900 18396 39956
rect 18452 39900 18462 39956
rect 38994 39900 39004 39956
rect 39060 39900 40124 39956
rect 40180 39900 40190 39956
rect 41356 39900 43484 39956
rect 43540 39900 43550 39956
rect 44818 39900 44828 39956
rect 44884 39900 44940 39956
rect 44996 39900 45006 39956
rect 43484 39844 43540 39900
rect 5842 39788 5852 39844
rect 5908 39788 10332 39844
rect 10388 39788 10398 39844
rect 32498 39788 32508 39844
rect 32564 39788 36876 39844
rect 36932 39788 36942 39844
rect 37986 39788 37996 39844
rect 38052 39788 41356 39844
rect 41412 39788 41422 39844
rect 43484 39788 46396 39844
rect 46452 39788 46462 39844
rect 5058 39676 5068 39732
rect 5124 39676 6300 39732
rect 6356 39676 6366 39732
rect 13906 39676 13916 39732
rect 13972 39676 17556 39732
rect 17612 39676 17622 39732
rect 32610 39676 32620 39732
rect 32676 39676 37156 39732
rect 37212 39676 37222 39732
rect 4050 39564 4060 39620
rect 4116 39564 4844 39620
rect 4900 39564 6076 39620
rect 6132 39564 6142 39620
rect 12282 39564 12292 39620
rect 12348 39564 13524 39620
rect 13580 39564 14364 39620
rect 14420 39564 14430 39620
rect 20122 39564 20132 39620
rect 20188 39564 21308 39620
rect 21364 39564 21374 39620
rect 22174 39564 22184 39620
rect 22240 39564 26236 39620
rect 26292 39564 26302 39620
rect 27346 39564 27356 39620
rect 27412 39564 29036 39620
rect 29092 39564 29102 39620
rect 30818 39564 30828 39620
rect 30884 39564 31612 39620
rect 31668 39564 32396 39620
rect 32452 39564 33068 39620
rect 33124 39564 33134 39620
rect 33562 39564 33572 39620
rect 33628 39564 37324 39620
rect 37380 39564 37390 39620
rect 38210 39564 38220 39620
rect 38276 39564 40684 39620
rect 40740 39564 41356 39620
rect 41412 39564 45500 39620
rect 45556 39564 45566 39620
rect 45714 39564 45724 39620
rect 45780 39564 46172 39620
rect 46228 39564 46238 39620
rect 9986 39452 9996 39508
rect 10052 39452 11284 39508
rect 11340 39452 12012 39508
rect 12068 39452 12078 39508
rect 12450 39452 12460 39508
rect 12516 39452 13244 39508
rect 13300 39452 13310 39508
rect 14914 39452 14924 39508
rect 14980 39452 23660 39508
rect 23716 39452 23726 39508
rect 28130 39452 28140 39508
rect 28196 39452 29204 39508
rect 29260 39452 29270 39508
rect 31714 39452 31724 39508
rect 31780 39452 32732 39508
rect 32788 39452 33292 39508
rect 33348 39452 33358 39508
rect 33516 39452 36540 39508
rect 36596 39452 36606 39508
rect 38434 39452 38444 39508
rect 38500 39452 42140 39508
rect 42196 39452 42206 39508
rect 45602 39452 45612 39508
rect 45668 39452 48076 39508
rect 48132 39452 48142 39508
rect 33516 39396 33572 39452
rect 6458 39340 6468 39396
rect 6524 39340 10556 39396
rect 10612 39340 10622 39396
rect 15362 39340 15372 39396
rect 15428 39340 28252 39396
rect 28308 39340 28904 39396
rect 28960 39340 28970 39396
rect 29362 39340 29372 39396
rect 29428 39340 33572 39396
rect 34626 39340 34636 39396
rect 34692 39340 41692 39396
rect 41748 39340 41758 39396
rect 42690 39340 42700 39396
rect 42756 39340 44940 39396
rect 44996 39340 45006 39396
rect 11666 39228 11676 39284
rect 11732 39228 13916 39284
rect 13972 39228 13982 39284
rect 23650 39228 23660 39284
rect 23716 39228 23726 39284
rect 24434 39228 24444 39284
rect 24500 39228 25676 39284
rect 25732 39228 25742 39284
rect 29922 39228 29932 39284
rect 29988 39228 30584 39284
rect 30640 39228 30650 39284
rect 36530 39228 36540 39284
rect 36596 39228 41972 39284
rect 42130 39228 42140 39284
rect 42196 39228 44044 39284
rect 44100 39228 45052 39284
rect 45108 39228 45118 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 3490 39116 3500 39172
rect 3556 39116 3948 39172
rect 4004 39116 15596 39172
rect 15652 39116 15662 39172
rect 21084 39116 23492 39172
rect 23548 39116 23558 39172
rect 15596 39060 15652 39116
rect 21084 39060 21140 39116
rect 23660 39060 23716 39228
rect 25554 39116 25564 39172
rect 25620 39116 25630 39172
rect 26114 39116 26124 39172
rect 26180 39116 27112 39172
rect 27168 39116 27178 39172
rect 36194 39116 36204 39172
rect 36260 39116 36652 39172
rect 36708 39116 36764 39172
rect 36820 39116 36830 39172
rect 38882 39116 38892 39172
rect 38948 39116 39564 39172
rect 39620 39116 39630 39172
rect 1586 39004 1596 39060
rect 1652 39004 4676 39060
rect 4732 39004 4742 39060
rect 9202 39004 9212 39060
rect 9268 39004 9660 39060
rect 9716 39004 9726 39060
rect 10322 39004 10332 39060
rect 10388 39004 10780 39060
rect 10836 39004 10846 39060
rect 12114 39004 12124 39060
rect 12180 39004 12728 39060
rect 12784 39004 12794 39060
rect 15596 39004 21140 39060
rect 21298 39004 21308 39060
rect 21364 39004 22184 39060
rect 22240 39004 22250 39060
rect 23660 39004 25060 39060
rect 25004 38948 25060 39004
rect 5170 38892 5180 38948
rect 5236 38892 6972 38948
rect 7028 38892 7038 38948
rect 21074 38892 21084 38948
rect 21140 38892 22540 38948
rect 22596 38892 22606 38948
rect 24994 38892 25004 38948
rect 25060 38892 25070 38948
rect 7074 38780 7084 38836
rect 7140 38780 8764 38836
rect 8820 38780 8830 38836
rect 10434 38780 10444 38836
rect 10500 38780 10510 38836
rect 13570 38780 13580 38836
rect 13636 38780 14252 38836
rect 14308 38780 14318 38836
rect 15922 38780 15932 38836
rect 15988 38780 16940 38836
rect 16996 38780 17006 38836
rect 20850 38780 20860 38836
rect 20916 38780 22428 38836
rect 22484 38780 22494 38836
rect 10444 38724 10500 38780
rect 25564 38724 25620 39116
rect 41916 39060 41972 39228
rect 42802 39116 42812 39172
rect 42868 39116 44604 39172
rect 44660 39116 44940 39172
rect 44996 39116 45006 39172
rect 45154 39116 45164 39172
rect 45220 39116 46732 39172
rect 46788 39116 46798 39172
rect 30706 39004 30716 39060
rect 30772 39004 31220 39060
rect 31276 39004 31286 39060
rect 33954 39004 33964 39060
rect 34020 39004 34030 39060
rect 35074 39004 35084 39060
rect 35140 39004 35868 39060
rect 35924 39004 36428 39060
rect 36484 39004 36494 39060
rect 37594 39004 37604 39060
rect 37660 39004 38108 39060
rect 38164 39004 38174 39060
rect 38994 39004 39004 39060
rect 39060 39004 39900 39060
rect 39956 39004 39966 39060
rect 41916 39004 47460 39060
rect 47516 39004 47526 39060
rect 33964 38948 34020 39004
rect 30370 38892 30380 38948
rect 30436 38892 30492 38948
rect 30548 38892 30558 38948
rect 33964 38892 36988 38948
rect 37044 38892 37054 38948
rect 37846 38892 37884 38948
rect 37940 38892 37950 38948
rect 38322 38892 38332 38948
rect 38388 38892 39228 38948
rect 39284 38892 39294 38948
rect 42242 38892 42252 38948
rect 42308 38892 43036 38948
rect 43092 38892 43102 38948
rect 44706 38892 44716 38948
rect 44772 38892 45612 38948
rect 45668 38892 45678 38948
rect 46386 38892 46396 38948
rect 46452 38892 46508 38948
rect 46564 38892 46574 38948
rect 27234 38780 27244 38836
rect 27300 38780 28252 38836
rect 28308 38780 28318 38836
rect 29138 38780 29148 38836
rect 29204 38780 29708 38836
rect 29764 38780 30492 38836
rect 30548 38780 30558 38836
rect 32722 38780 32732 38836
rect 32788 38780 33068 38836
rect 33124 38780 33134 38836
rect 34794 38780 34804 38836
rect 34860 38780 36540 38836
rect 36596 38780 36606 38836
rect 36866 38780 36876 38836
rect 36932 38780 40796 38836
rect 40852 38780 40862 38836
rect 41682 38780 41692 38836
rect 41748 38780 42812 38836
rect 42868 38780 42878 38836
rect 43866 38780 43876 38836
rect 43932 38780 46562 38836
rect 46618 38780 46628 38836
rect 46946 38780 46956 38836
rect 47012 38780 47740 38836
rect 47796 38780 47806 38836
rect 4666 38668 4676 38724
rect 4732 38668 5516 38724
rect 5572 38668 5964 38724
rect 6020 38668 7868 38724
rect 7924 38668 8428 38724
rect 8484 38668 9436 38724
rect 9492 38668 11564 38724
rect 11620 38668 13804 38724
rect 13860 38668 13870 38724
rect 21186 38668 21196 38724
rect 21252 38668 21980 38724
rect 22036 38668 22046 38724
rect 22204 38668 22932 38724
rect 22988 38668 23996 38724
rect 24052 38668 24062 38724
rect 25564 38668 26684 38724
rect 26740 38668 27132 38724
rect 27188 38668 27198 38724
rect 28690 38668 28700 38724
rect 28756 38668 29932 38724
rect 29988 38668 29998 38724
rect 30342 38668 30380 38724
rect 30436 38668 30446 38724
rect 31938 38668 31948 38724
rect 32004 38668 33944 38724
rect 34000 38668 34010 38724
rect 37958 38668 37996 38724
rect 38052 38668 38062 38724
rect 40674 38668 40684 38724
rect 40740 38668 41132 38724
rect 41188 38668 41198 38724
rect 41906 38668 41916 38724
rect 41972 38668 42588 38724
rect 42644 38668 44380 38724
rect 44436 38668 45388 38724
rect 45444 38668 45454 38724
rect 45826 38668 45836 38724
rect 45892 38668 46284 38724
rect 46340 38668 46350 38724
rect 22204 38612 22260 38668
rect 14354 38556 14364 38612
rect 14420 38556 15800 38612
rect 15856 38556 15866 38612
rect 22082 38556 22092 38612
rect 22148 38556 22260 38612
rect 28802 38556 28812 38612
rect 28868 38556 29820 38612
rect 29876 38556 29886 38612
rect 30156 38556 32060 38612
rect 32116 38556 34972 38612
rect 35028 38556 35038 38612
rect 35970 38556 35980 38612
rect 36036 38556 39452 38612
rect 39508 38556 41244 38612
rect 41300 38556 41310 38612
rect 43334 38556 43372 38612
rect 43428 38556 43438 38612
rect 43586 38556 43596 38612
rect 43652 38556 43708 38612
rect 43764 38556 43774 38612
rect 43922 38556 43932 38612
rect 43988 38556 44604 38612
rect 44660 38556 44670 38612
rect 46386 38556 46396 38612
rect 46452 38556 46508 38612
rect 46564 38556 46574 38612
rect 30156 38500 30212 38556
rect 10210 38444 10220 38500
rect 10276 38444 10286 38500
rect 23538 38444 23548 38500
rect 23604 38444 24612 38500
rect 24668 38444 30212 38500
rect 30370 38444 30380 38500
rect 30436 38444 30492 38500
rect 30548 38444 30558 38500
rect 31014 38444 31052 38500
rect 31108 38444 31118 38500
rect 38098 38444 38108 38500
rect 38164 38444 38174 38500
rect 38546 38444 38556 38500
rect 38612 38444 49364 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 6738 38332 6748 38388
rect 6804 38332 6814 38388
rect 3434 38220 3444 38276
rect 3500 38220 3836 38276
rect 3892 38220 4228 38276
rect 2986 38108 2996 38164
rect 3052 38108 3948 38164
rect 4004 38108 4014 38164
rect 2594 37996 2604 38052
rect 2660 37996 3780 38052
rect 3836 37996 3846 38052
rect 4172 37940 4228 38220
rect 6748 38052 6804 38332
rect 10220 38052 10276 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 38108 38388 38164 38444
rect 20178 38332 20188 38388
rect 20244 38332 21084 38388
rect 21140 38332 21150 38388
rect 25442 38332 25452 38388
rect 25508 38332 26572 38388
rect 26628 38332 26638 38388
rect 35970 38332 35980 38388
rect 36036 38332 37884 38388
rect 37940 38332 37950 38388
rect 38108 38332 42084 38388
rect 42140 38332 42150 38388
rect 45938 38332 45948 38388
rect 46004 38332 46732 38388
rect 46788 38332 46798 38388
rect 18274 38220 18284 38276
rect 18340 38220 18620 38276
rect 18676 38220 18686 38276
rect 20402 38220 20412 38276
rect 20468 38220 20524 38276
rect 20580 38220 20590 38276
rect 22810 38220 22820 38276
rect 22876 38220 23324 38276
rect 23380 38220 23390 38276
rect 25330 38220 25340 38276
rect 25396 38220 26124 38276
rect 26180 38220 26190 38276
rect 34178 38220 34188 38276
rect 34244 38220 35644 38276
rect 35700 38220 35710 38276
rect 36978 38220 36988 38276
rect 37044 38220 38444 38276
rect 38500 38220 38510 38276
rect 40898 38220 40908 38276
rect 40964 38220 41692 38276
rect 41748 38220 42364 38276
rect 42420 38220 42430 38276
rect 43474 38220 43484 38276
rect 43540 38220 44156 38276
rect 44212 38220 48076 38276
rect 48132 38220 48142 38276
rect 13346 38108 13356 38164
rect 13412 38108 14364 38164
rect 14420 38108 14430 38164
rect 16930 38108 16940 38164
rect 16996 38108 23212 38164
rect 23268 38108 23660 38164
rect 23716 38108 23726 38164
rect 34850 38108 34860 38164
rect 34916 38108 43820 38164
rect 43876 38108 43886 38164
rect 6738 37996 6748 38052
rect 6804 37996 6814 38052
rect 10210 37996 10220 38052
rect 10276 37996 10286 38052
rect 11666 37996 11676 38052
rect 11732 37996 11742 38052
rect 12114 37996 12124 38052
rect 12180 37996 12572 38052
rect 12628 37996 14252 38052
rect 14308 37996 14318 38052
rect 14578 37996 14588 38052
rect 14644 37996 14924 38052
rect 14980 37996 14990 38052
rect 16034 37996 16044 38052
rect 16100 37996 28028 38052
rect 28084 37996 30024 38052
rect 30080 37996 30090 38052
rect 30258 37996 30268 38052
rect 30324 37996 30716 38052
rect 30772 37996 32172 38052
rect 32228 37996 32238 38052
rect 36978 37996 36988 38052
rect 37044 37996 37436 38052
rect 37492 37996 38556 38052
rect 38612 37996 38622 38052
rect 44202 37996 44212 38052
rect 44268 37996 45388 38052
rect 45444 37996 45454 38052
rect 11676 37940 11732 37996
rect 4172 37884 11732 37940
rect 12002 37884 12012 37940
rect 12068 37884 13692 37940
rect 13748 37884 13758 37940
rect 19674 37884 19684 37940
rect 19740 37884 22540 37940
rect 22596 37884 22606 37940
rect 24210 37884 24220 37940
rect 24276 37884 27076 37940
rect 27132 37884 27142 37940
rect 28466 37884 28476 37940
rect 28532 37884 31592 37940
rect 31648 37884 31658 37940
rect 37202 37884 37212 37940
rect 37268 37884 40852 37940
rect 40908 37884 40918 37940
rect 9660 37828 9716 37884
rect 9650 37772 9660 37828
rect 9716 37772 9726 37828
rect 10974 37772 10984 37828
rect 11040 37772 11452 37828
rect 11508 37772 11676 37828
rect 11732 37772 11742 37828
rect 18218 37772 18228 37828
rect 18284 37772 18396 37828
rect 18452 37772 26908 37828
rect 33842 37772 33852 37828
rect 33908 37772 36988 37828
rect 37044 37772 37054 37828
rect 37706 37772 37716 37828
rect 37772 37772 38220 37828
rect 38276 37772 38286 37828
rect 42690 37772 42700 37828
rect 42756 37772 43596 37828
rect 43652 37772 43662 37828
rect 44482 37772 44492 37828
rect 44548 37772 45388 37828
rect 45444 37772 45454 37828
rect 46694 37772 46732 37828
rect 46788 37772 46798 37828
rect 26852 37716 26908 37772
rect 6850 37660 6860 37716
rect 6916 37660 10332 37716
rect 10388 37660 16604 37716
rect 16660 37660 16670 37716
rect 20178 37660 20188 37716
rect 20244 37660 20282 37716
rect 20374 37660 20412 37716
rect 20468 37660 20478 37716
rect 20570 37660 20580 37716
rect 20636 37660 21308 37716
rect 21364 37660 21374 37716
rect 25946 37660 25956 37716
rect 26012 37660 26572 37716
rect 26628 37660 26638 37716
rect 26852 37660 29764 37716
rect 29820 37660 29830 37716
rect 31042 37660 31052 37716
rect 31108 37660 38668 37716
rect 41570 37660 41580 37716
rect 41636 37660 42140 37716
rect 42196 37660 43372 37716
rect 43428 37660 43438 37716
rect 44818 37660 44828 37716
rect 44884 37660 46956 37716
rect 47012 37660 47022 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 38612 37604 38668 37660
rect 5786 37548 5796 37604
rect 5852 37548 6524 37604
rect 6580 37548 7420 37604
rect 7476 37548 13356 37604
rect 13412 37548 13422 37604
rect 21074 37548 21084 37604
rect 21140 37548 21150 37604
rect 25610 37548 25620 37604
rect 25676 37548 26460 37604
rect 26516 37548 26526 37604
rect 32386 37548 32396 37604
rect 32452 37548 33460 37604
rect 33516 37548 33526 37604
rect 36754 37548 36764 37604
rect 36820 37548 37884 37604
rect 37940 37548 37950 37604
rect 38612 37548 46172 37604
rect 46228 37548 46238 37604
rect 8754 37436 8764 37492
rect 8820 37436 9044 37492
rect 9100 37436 9436 37492
rect 9492 37436 20188 37492
rect 20244 37436 20254 37492
rect 7186 37324 7196 37380
rect 7252 37324 7644 37380
rect 7700 37324 7710 37380
rect 8026 37324 8036 37380
rect 8092 37324 8428 37380
rect 8484 37324 8494 37380
rect 12450 37324 12460 37380
rect 12516 37324 13132 37380
rect 13188 37324 13198 37380
rect 13346 37324 13356 37380
rect 13412 37324 16380 37380
rect 16436 37324 16446 37380
rect 18498 37324 18508 37380
rect 18564 37324 19068 37380
rect 19124 37324 19134 37380
rect 4274 37212 4284 37268
rect 4340 37212 5964 37268
rect 6020 37212 6244 37268
rect 6300 37212 6310 37268
rect 12562 37212 12572 37268
rect 12628 37212 13804 37268
rect 13860 37212 13870 37268
rect 16706 37212 16716 37268
rect 16772 37212 17332 37268
rect 17388 37212 17398 37268
rect 18274 37212 18284 37268
rect 18340 37212 18620 37268
rect 18676 37212 19292 37268
rect 19348 37212 19358 37268
rect 20290 37212 20300 37268
rect 20356 37212 20748 37268
rect 20804 37212 20814 37268
rect 21084 37156 21140 37548
rect 49308 37492 49364 38444
rect 21502 37436 21512 37492
rect 21568 37436 22428 37492
rect 22484 37436 27244 37492
rect 27300 37436 27310 37492
rect 30370 37436 30380 37492
rect 30436 37436 30660 37492
rect 30716 37436 33348 37492
rect 35634 37436 35644 37492
rect 35700 37436 36652 37492
rect 36708 37436 37324 37492
rect 37380 37436 37390 37492
rect 38612 37436 38892 37492
rect 38948 37436 40012 37492
rect 40068 37436 40078 37492
rect 40226 37436 40236 37492
rect 40292 37436 40572 37492
rect 40628 37436 42924 37492
rect 42980 37436 42990 37492
rect 47282 37436 47292 37492
rect 47348 37436 47358 37492
rect 49084 37436 49364 37492
rect 33292 37380 33348 37436
rect 38612 37380 38668 37436
rect 21634 37324 21644 37380
rect 21700 37324 22316 37380
rect 22372 37324 22382 37380
rect 24770 37324 24780 37380
rect 24836 37324 25564 37380
rect 25620 37324 25630 37380
rect 28354 37324 28364 37380
rect 28420 37324 29148 37380
rect 29204 37324 29214 37380
rect 32722 37324 32732 37380
rect 32788 37324 33068 37380
rect 33124 37324 33134 37380
rect 33292 37324 38668 37380
rect 47292 37268 47348 37436
rect 21746 37212 21756 37268
rect 21812 37212 22652 37268
rect 22708 37212 22718 37268
rect 30202 37212 30212 37268
rect 30268 37212 30604 37268
rect 30660 37212 30670 37268
rect 32162 37212 32172 37268
rect 32228 37212 33944 37268
rect 34000 37212 34010 37268
rect 34178 37212 34188 37268
rect 34244 37212 35308 37268
rect 35364 37212 35374 37268
rect 37036 37212 37046 37268
rect 37102 37212 40348 37268
rect 40404 37212 40414 37268
rect 41570 37212 41580 37268
rect 41636 37212 43932 37268
rect 43988 37212 43998 37268
rect 46386 37212 46396 37268
rect 46452 37212 47348 37268
rect 49084 37268 49140 37436
rect 49200 37268 50000 37296
rect 49084 37212 50000 37268
rect 49200 37184 50000 37212
rect 4722 37100 4732 37156
rect 4788 37100 4956 37156
rect 5012 37100 6748 37156
rect 6804 37100 6814 37156
rect 10546 37100 10556 37156
rect 10612 37100 11284 37156
rect 11340 37100 11350 37156
rect 12338 37100 12348 37156
rect 12404 37100 13188 37156
rect 13244 37100 13254 37156
rect 13682 37100 13692 37156
rect 13748 37100 15204 37156
rect 15260 37100 15270 37156
rect 16482 37100 16492 37156
rect 16548 37100 18732 37156
rect 18788 37100 18798 37156
rect 18890 37100 18900 37156
rect 18956 37100 20076 37156
rect 20132 37100 20142 37156
rect 20402 37100 20412 37156
rect 20468 37100 21140 37156
rect 21298 37100 21308 37156
rect 21364 37100 21532 37156
rect 21588 37100 21598 37156
rect 22194 37100 22204 37156
rect 22260 37100 22876 37156
rect 22932 37100 22942 37156
rect 26450 37100 26460 37156
rect 26516 37100 27916 37156
rect 27972 37100 27982 37156
rect 29754 37100 29764 37156
rect 29820 37100 32396 37156
rect 32452 37100 32462 37156
rect 32834 37100 32844 37156
rect 32900 37100 36260 37156
rect 36316 37100 36326 37156
rect 36642 37100 36652 37156
rect 36708 37100 37996 37156
rect 38052 37100 38062 37156
rect 43810 37100 43820 37156
rect 43876 37100 44156 37156
rect 44212 37100 44222 37156
rect 45154 37100 45164 37156
rect 45220 37100 45836 37156
rect 45892 37100 47852 37156
rect 47908 37100 47918 37156
rect 8754 36988 8764 37044
rect 8820 36988 9716 37044
rect 9772 36988 9782 37044
rect 18508 36988 21756 37044
rect 21812 36988 23492 37044
rect 23548 36988 23558 37044
rect 37202 36988 37212 37044
rect 37268 36988 37996 37044
rect 38052 36988 38062 37044
rect 41346 36988 41356 37044
rect 41412 36988 42028 37044
rect 42084 36988 42588 37044
rect 42644 36988 42654 37044
rect 44930 36988 44940 37044
rect 44996 36988 46172 37044
rect 46228 36988 46238 37044
rect 18508 36932 18564 36988
rect 6234 36876 6244 36932
rect 6300 36876 8148 36932
rect 8204 36876 8316 36932
rect 8372 36876 8382 36932
rect 8586 36876 8596 36932
rect 8708 36876 8718 36932
rect 15586 36876 15596 36932
rect 15652 36876 17780 36932
rect 17836 36876 18564 36932
rect 26114 36876 26124 36932
rect 26180 36876 26190 36932
rect 26338 36876 26348 36932
rect 26404 36876 26414 36932
rect 35634 36876 35644 36932
rect 35700 36876 37436 36932
rect 37492 36876 37502 36932
rect 42242 36876 42252 36932
rect 42308 36876 43036 36932
rect 43092 36876 43102 36932
rect 45266 36876 45276 36932
rect 45332 36876 46284 36932
rect 46340 36876 46350 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 11442 36764 11452 36820
rect 11508 36764 12012 36820
rect 12068 36764 12078 36820
rect 20178 36764 20188 36820
rect 20244 36764 20748 36820
rect 20804 36764 20814 36820
rect 9538 36652 9548 36708
rect 9604 36652 10500 36708
rect 10556 36652 10566 36708
rect 19170 36652 19180 36708
rect 19236 36652 22484 36708
rect 22540 36652 22550 36708
rect 5786 36540 5796 36596
rect 5852 36540 6524 36596
rect 6580 36540 6590 36596
rect 19282 36540 19292 36596
rect 19348 36540 20412 36596
rect 20468 36540 20478 36596
rect 25554 36540 25564 36596
rect 25620 36540 25788 36596
rect 25844 36540 25854 36596
rect 26124 36484 26180 36876
rect 26348 36708 26404 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 26878 36764 26888 36820
rect 26944 36764 28120 36820
rect 28176 36764 28186 36820
rect 26348 36652 27020 36708
rect 27076 36652 27086 36708
rect 30370 36652 30380 36708
rect 30436 36652 30828 36708
rect 30884 36652 31500 36708
rect 31556 36652 31566 36708
rect 35186 36652 35196 36708
rect 35252 36652 41524 36708
rect 41580 36652 41590 36708
rect 27906 36540 27916 36596
rect 27972 36540 30136 36596
rect 30192 36540 30202 36596
rect 31994 36540 32004 36596
rect 32060 36540 32844 36596
rect 32900 36540 32910 36596
rect 34290 36540 34300 36596
rect 34356 36540 34636 36596
rect 34692 36540 35364 36596
rect 35420 36540 35430 36596
rect 37538 36540 37548 36596
rect 37604 36540 40124 36596
rect 40180 36540 42588 36596
rect 42644 36540 42868 36596
rect 42924 36540 42934 36596
rect 45266 36540 45276 36596
rect 45332 36540 48020 36596
rect 48076 36540 48086 36596
rect 2594 36428 2604 36484
rect 2660 36428 3892 36484
rect 3948 36428 3958 36484
rect 4218 36428 4228 36484
rect 4284 36428 5628 36484
rect 5684 36428 5694 36484
rect 8194 36428 8204 36484
rect 8260 36428 8316 36484
rect 8372 36428 8382 36484
rect 9538 36428 9548 36484
rect 9604 36428 13804 36484
rect 13860 36428 13870 36484
rect 21354 36428 21364 36484
rect 21420 36428 21980 36484
rect 22036 36428 22046 36484
rect 26114 36428 26124 36484
rect 26180 36428 26190 36484
rect 31826 36428 31836 36484
rect 31892 36428 33404 36484
rect 33460 36428 34188 36484
rect 34244 36428 34254 36484
rect 39554 36428 39564 36484
rect 39620 36428 41132 36484
rect 41188 36428 41804 36484
rect 41860 36428 41870 36484
rect 43362 36428 43372 36484
rect 43428 36428 44716 36484
rect 44772 36428 44782 36484
rect 45490 36428 45500 36484
rect 45556 36428 45668 36484
rect 45724 36428 45734 36484
rect 5058 36316 5068 36372
rect 5124 36316 5908 36372
rect 5964 36316 9304 36372
rect 9360 36316 9370 36372
rect 17826 36316 17836 36372
rect 17892 36316 20860 36372
rect 20916 36316 20926 36372
rect 32386 36316 32396 36372
rect 32452 36316 34916 36372
rect 34972 36316 36876 36372
rect 36932 36316 37324 36372
rect 37380 36316 37390 36372
rect 41010 36316 41020 36372
rect 41076 36316 41692 36372
rect 41748 36316 41758 36372
rect 6626 36204 6636 36260
rect 6692 36204 6972 36260
rect 7028 36204 7038 36260
rect 8194 36204 8204 36260
rect 8260 36204 11788 36260
rect 11844 36204 11854 36260
rect 19954 36204 19964 36260
rect 20020 36204 21028 36260
rect 21084 36204 21094 36260
rect 34570 36204 34580 36260
rect 34636 36204 34748 36260
rect 34804 36204 35532 36260
rect 35588 36204 35598 36260
rect 43698 36204 43708 36260
rect 43764 36204 44604 36260
rect 44660 36204 45052 36260
rect 45108 36204 45118 36260
rect 7634 36092 7644 36148
rect 7700 36092 8988 36148
rect 9044 36092 11452 36148
rect 11508 36092 11518 36148
rect 20738 36092 20748 36148
rect 20804 36092 29148 36148
rect 29204 36092 29214 36148
rect 32554 36092 32564 36148
rect 32620 36092 36988 36148
rect 37044 36092 37054 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 20850 35980 20860 36036
rect 20916 35980 21308 36036
rect 21364 35980 21374 36036
rect 21634 35980 21644 36036
rect 21700 35980 21710 36036
rect 21858 35980 21868 36036
rect 21924 35980 29820 36036
rect 29876 35980 29886 36036
rect 29978 35980 29988 36036
rect 30044 35980 31108 36036
rect 31164 35980 32452 36036
rect 37650 35980 37660 36036
rect 37716 35980 41804 36036
rect 41860 35980 41870 36036
rect 21644 35924 21700 35980
rect 32396 35924 32452 35980
rect 15474 35868 15484 35924
rect 15540 35868 18452 35924
rect 18508 35868 18518 35924
rect 19730 35868 19740 35924
rect 19796 35868 21700 35924
rect 26226 35868 26236 35924
rect 26292 35868 27916 35924
rect 27972 35868 27982 35924
rect 32396 35868 33068 35924
rect 33124 35868 33134 35924
rect 35914 35868 35924 35924
rect 35980 35868 39452 35924
rect 39508 35868 39518 35924
rect 42466 35868 42476 35924
rect 42532 35868 42812 35924
rect 42868 35868 42878 35924
rect 3602 35756 3612 35812
rect 3668 35756 5404 35812
rect 5460 35756 5470 35812
rect 8866 35756 8876 35812
rect 8932 35756 9492 35812
rect 9548 35756 9558 35812
rect 11078 35756 11116 35812
rect 11172 35756 11182 35812
rect 18274 35756 18284 35812
rect 18340 35756 18788 35812
rect 18844 35756 20860 35812
rect 20916 35756 20926 35812
rect 21084 35756 27804 35812
rect 27860 35756 27870 35812
rect 30258 35756 30268 35812
rect 30324 35756 30716 35812
rect 30772 35756 33180 35812
rect 33236 35756 33246 35812
rect 38602 35756 38612 35812
rect 38668 35756 40796 35812
rect 40852 35756 40862 35812
rect 43026 35756 43036 35812
rect 43092 35756 44436 35812
rect 44492 35756 44502 35812
rect 45350 35756 45388 35812
rect 45444 35756 45454 35812
rect 4834 35644 4844 35700
rect 4900 35644 4910 35700
rect 12114 35644 12124 35700
rect 12180 35644 12572 35700
rect 12628 35644 12638 35700
rect 20150 35644 20188 35700
rect 20244 35644 20254 35700
rect 2650 35308 2660 35364
rect 2716 35308 3500 35364
rect 3556 35308 3566 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 4844 35140 4900 35644
rect 21084 35588 21140 35756
rect 26114 35644 26124 35700
rect 26180 35644 27132 35700
rect 27188 35644 27198 35700
rect 28242 35644 28252 35700
rect 28308 35644 32564 35700
rect 32722 35644 32732 35700
rect 32788 35644 33516 35700
rect 33572 35644 34076 35700
rect 34132 35644 34142 35700
rect 37202 35644 37212 35700
rect 37268 35644 37436 35700
rect 37492 35644 37940 35700
rect 38098 35644 38108 35700
rect 38164 35644 38892 35700
rect 38948 35644 38958 35700
rect 39722 35644 39732 35700
rect 39788 35644 41468 35700
rect 41524 35644 41534 35700
rect 44818 35644 44828 35700
rect 44884 35644 47404 35700
rect 47460 35644 47470 35700
rect 13682 35532 13692 35588
rect 13748 35532 21140 35588
rect 21298 35532 21308 35588
rect 21364 35532 21588 35588
rect 21644 35532 22428 35588
rect 22484 35532 22494 35588
rect 24434 35532 24444 35588
rect 24500 35532 25844 35588
rect 25900 35532 25910 35588
rect 28914 35532 28924 35588
rect 28980 35532 29988 35588
rect 30044 35532 30054 35588
rect 32508 35476 32564 35644
rect 37884 35588 37940 35644
rect 35634 35532 35644 35588
rect 35700 35532 36092 35588
rect 36148 35532 37548 35588
rect 37604 35532 37614 35588
rect 37884 35532 43708 35588
rect 43764 35532 43774 35588
rect 45378 35532 45388 35588
rect 45444 35532 45500 35588
rect 45556 35532 45566 35588
rect 46610 35532 46620 35588
rect 46676 35532 47852 35588
rect 47908 35532 47918 35588
rect 6066 35420 6076 35476
rect 6132 35420 6412 35476
rect 6468 35420 12236 35476
rect 12292 35420 12302 35476
rect 17826 35420 17836 35476
rect 17892 35420 18284 35476
rect 18340 35420 18350 35476
rect 19282 35420 19292 35476
rect 19348 35420 19628 35476
rect 19684 35420 27692 35476
rect 27748 35420 28792 35476
rect 28848 35420 28858 35476
rect 30268 35420 31724 35476
rect 31780 35420 31790 35476
rect 32508 35420 39060 35476
rect 39218 35420 39228 35476
rect 39284 35420 41132 35476
rect 41188 35420 41198 35476
rect 41682 35420 41692 35476
rect 41748 35420 43036 35476
rect 43092 35420 43102 35476
rect 7970 35308 7980 35364
rect 8036 35308 8204 35364
rect 8260 35308 8270 35364
rect 9874 35308 9884 35364
rect 9940 35308 9950 35364
rect 9884 35252 9940 35308
rect 8418 35196 8428 35252
rect 8484 35196 9940 35252
rect 11078 35196 11116 35252
rect 11172 35196 11182 35252
rect 4722 35084 4732 35140
rect 4788 35084 4900 35140
rect 11788 35028 11844 35420
rect 30268 35364 30324 35420
rect 39004 35364 39060 35420
rect 12796 35308 13448 35364
rect 13504 35308 13514 35364
rect 15586 35308 15596 35364
rect 15652 35308 21868 35364
rect 21924 35308 21934 35364
rect 22418 35308 22428 35364
rect 22484 35308 22876 35364
rect 22932 35308 22942 35364
rect 25330 35308 25340 35364
rect 25396 35308 26236 35364
rect 26292 35308 26302 35364
rect 27570 35308 27580 35364
rect 27636 35308 27646 35364
rect 28588 35308 30324 35364
rect 30492 35308 31592 35364
rect 31648 35308 33852 35364
rect 33908 35308 33918 35364
rect 39004 35308 45668 35364
rect 47282 35308 47292 35364
rect 47348 35308 48132 35364
rect 48188 35308 48198 35364
rect 12796 35252 12852 35308
rect 27580 35252 27636 35308
rect 12786 35196 12796 35252
rect 12852 35196 12862 35252
rect 13878 35196 13916 35252
rect 13972 35196 13982 35252
rect 16230 35196 16268 35252
rect 16324 35196 16334 35252
rect 19506 35196 19516 35252
rect 19572 35196 20524 35252
rect 20580 35196 21980 35252
rect 22036 35196 23324 35252
rect 23380 35196 23390 35252
rect 25666 35196 25676 35252
rect 25732 35196 26908 35252
rect 26964 35196 26974 35252
rect 27580 35196 28364 35252
rect 28420 35196 28430 35252
rect 28588 35140 28644 35308
rect 28802 35196 28812 35252
rect 28868 35196 29148 35252
rect 29204 35196 29214 35252
rect 30492 35140 30548 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 35858 35196 35868 35252
rect 35924 35196 37100 35252
rect 37156 35196 37166 35252
rect 37706 35196 37716 35252
rect 37772 35196 42420 35252
rect 42476 35196 42486 35252
rect 45612 35140 45668 35308
rect 12338 35084 12348 35140
rect 12404 35084 13580 35140
rect 13636 35084 13646 35140
rect 15138 35084 15148 35140
rect 15204 35084 21028 35140
rect 22418 35084 22428 35140
rect 22484 35084 22764 35140
rect 22820 35084 22830 35140
rect 25442 35084 25452 35140
rect 25508 35084 25564 35140
rect 25620 35084 25630 35140
rect 28466 35084 28476 35140
rect 28532 35084 28644 35140
rect 30482 35084 30492 35140
rect 30548 35084 30558 35140
rect 32956 35084 36876 35140
rect 36932 35084 36942 35140
rect 45602 35084 45612 35140
rect 45668 35084 45678 35140
rect 46274 35084 46284 35140
rect 46340 35084 47180 35140
rect 47236 35084 47246 35140
rect 20972 35028 21028 35084
rect 11778 34972 11788 35028
rect 11844 34972 11854 35028
rect 16706 34972 16716 35028
rect 16772 34972 17220 35028
rect 17276 34972 17286 35028
rect 17388 34972 18172 35028
rect 18228 34972 18238 35028
rect 20972 34972 26908 35028
rect 17388 34916 17444 34972
rect 26852 34916 26908 34972
rect 3154 34860 3164 34916
rect 3220 34860 4508 34916
rect 4564 34860 5068 34916
rect 5124 34860 5134 34916
rect 7298 34860 7308 34916
rect 7364 34860 8652 34916
rect 8708 34860 9212 34916
rect 9268 34860 9278 34916
rect 9445 34860 9455 34916
rect 9511 34860 9660 34916
rect 9716 34860 12516 34916
rect 12572 34860 12582 34916
rect 17042 34860 17052 34916
rect 17108 34860 17444 34916
rect 19058 34860 19068 34916
rect 19124 34860 21084 34916
rect 21140 34860 21150 34916
rect 21522 34860 21532 34916
rect 21588 34860 21756 34916
rect 21812 34860 21822 34916
rect 22530 34860 22540 34916
rect 22596 34860 26292 34916
rect 26852 34860 28028 34916
rect 28084 34860 30024 34916
rect 30080 34860 30090 34916
rect 26236 34804 26292 34860
rect 4274 34748 4284 34804
rect 4340 34748 5180 34804
rect 5236 34748 5246 34804
rect 7522 34748 7532 34804
rect 7588 34748 8428 34804
rect 8484 34748 8494 34804
rect 9090 34748 9100 34804
rect 9156 34748 11284 34804
rect 11340 34748 11350 34804
rect 16762 34748 16772 34804
rect 16828 34748 17948 34804
rect 18004 34748 18014 34804
rect 18162 34748 18172 34804
rect 18228 34748 19180 34804
rect 19236 34748 19246 34804
rect 20066 34748 20076 34804
rect 20132 34748 20300 34804
rect 20356 34748 20366 34804
rect 26226 34748 26236 34804
rect 26292 34748 26302 34804
rect 26450 34748 26460 34804
rect 26516 34748 31556 34804
rect 31612 34748 31622 34804
rect 32274 34748 32284 34804
rect 32340 34748 32732 34804
rect 32788 34748 32798 34804
rect 5180 34692 5236 34748
rect 5180 34636 12684 34692
rect 12740 34636 12750 34692
rect 15092 34636 15708 34692
rect 15764 34636 15774 34692
rect 25666 34636 25676 34692
rect 25732 34636 26796 34692
rect 26852 34636 26862 34692
rect 31098 34636 31108 34692
rect 31164 34636 32060 34692
rect 32116 34636 32126 34692
rect 4050 34524 4060 34580
rect 4116 34524 5012 34580
rect 5068 34524 5078 34580
rect 5562 34524 5572 34580
rect 5628 34524 6916 34580
rect 6972 34524 8652 34580
rect 8708 34524 11228 34580
rect 11284 34524 11294 34580
rect 15092 34468 15148 34636
rect 32956 34580 33012 35084
rect 36502 34972 36540 35028
rect 36596 34972 36606 35028
rect 36754 34972 36764 35028
rect 36820 34972 37660 35028
rect 37716 34972 37726 35028
rect 41122 34972 41132 35028
rect 41188 34972 42140 35028
rect 42196 34972 42206 35028
rect 43138 34972 43148 35028
rect 43204 34972 44604 35028
rect 44660 34972 44670 35028
rect 44930 34972 44940 35028
rect 44996 34972 46284 35028
rect 46340 34972 46350 35028
rect 40898 34860 40908 34916
rect 40964 34860 41916 34916
rect 41972 34860 41982 34916
rect 43418 34860 43428 34916
rect 43484 34860 43708 34916
rect 43764 34860 43774 34916
rect 44034 34860 44044 34916
rect 44100 34860 46060 34916
rect 46116 34860 46126 34916
rect 43362 34636 43372 34692
rect 43428 34636 44044 34692
rect 44100 34636 44110 34692
rect 20290 34524 20300 34580
rect 20356 34524 20412 34580
rect 20468 34524 20478 34580
rect 21756 34524 33012 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 21756 34468 21812 34524
rect 2594 34412 2604 34468
rect 2660 34412 5684 34468
rect 5740 34412 5750 34468
rect 5964 34412 10948 34468
rect 11050 34412 11060 34468
rect 11116 34412 15148 34468
rect 17490 34412 17500 34468
rect 17556 34412 18284 34468
rect 18340 34412 18350 34468
rect 20514 34412 20524 34468
rect 20580 34412 21812 34468
rect 23650 34412 23660 34468
rect 23716 34412 23996 34468
rect 24052 34412 24062 34468
rect 25106 34412 25116 34468
rect 25172 34412 27244 34468
rect 27300 34412 27310 34468
rect 31546 34412 31556 34468
rect 31612 34412 36204 34468
rect 36260 34412 38668 34468
rect 38724 34412 42924 34468
rect 42980 34412 45164 34468
rect 45220 34412 45230 34468
rect 5964 34356 6020 34412
rect 10892 34356 10948 34412
rect 3490 34300 3500 34356
rect 3556 34300 4172 34356
rect 4228 34300 4238 34356
rect 5282 34300 5292 34356
rect 5348 34300 6020 34356
rect 6178 34300 6188 34356
rect 6244 34300 7140 34356
rect 7196 34300 7206 34356
rect 8978 34300 8988 34356
rect 9044 34300 9660 34356
rect 9716 34300 9726 34356
rect 10892 34300 12460 34356
rect 12516 34300 12526 34356
rect 12674 34300 12684 34356
rect 12740 34300 14644 34356
rect 19954 34300 19964 34356
rect 20020 34300 21308 34356
rect 21364 34300 21374 34356
rect 23734 34300 23772 34356
rect 23828 34300 23838 34356
rect 33842 34300 33852 34356
rect 33908 34300 36988 34356
rect 37044 34300 37054 34356
rect 37548 34300 37828 34356
rect 37884 34300 37894 34356
rect 38882 34300 38892 34356
rect 38948 34300 39004 34356
rect 39060 34300 39070 34356
rect 2930 34188 2940 34244
rect 2996 34188 4284 34244
rect 4340 34188 4350 34244
rect 6290 34188 6300 34244
rect 6356 34188 6860 34244
rect 6916 34188 6926 34244
rect 12954 34188 12964 34244
rect 13020 34188 14364 34244
rect 14420 34188 14430 34244
rect 4284 34020 4340 34188
rect 14588 34132 14644 34300
rect 18778 34188 18788 34244
rect 18844 34188 21868 34244
rect 21924 34188 21934 34244
rect 25442 34188 25452 34244
rect 25508 34188 26572 34244
rect 26628 34188 26638 34244
rect 28354 34188 28364 34244
rect 28420 34188 29148 34244
rect 29204 34188 29214 34244
rect 31938 34188 31948 34244
rect 32004 34188 33964 34244
rect 34020 34188 34030 34244
rect 37548 34132 37604 34300
rect 44818 34188 44828 34244
rect 44884 34188 45276 34244
rect 45332 34188 45342 34244
rect 6738 34076 6748 34132
rect 6804 34076 8092 34132
rect 8148 34076 8158 34132
rect 9986 34076 9996 34132
rect 10052 34076 12012 34132
rect 12068 34076 12078 34132
rect 13906 34076 13916 34132
rect 13972 34076 13982 34132
rect 14588 34076 14812 34132
rect 14868 34076 15148 34132
rect 15204 34076 15214 34132
rect 16930 34076 16940 34132
rect 16996 34076 18060 34132
rect 18116 34076 18126 34132
rect 20962 34076 20972 34132
rect 21028 34076 21644 34132
rect 21700 34076 21710 34132
rect 22418 34076 22428 34132
rect 22484 34076 23772 34132
rect 23828 34076 23838 34132
rect 29754 34076 29764 34132
rect 29820 34076 30716 34132
rect 30772 34076 30782 34132
rect 31826 34076 31836 34132
rect 31892 34076 33068 34132
rect 33124 34076 33134 34132
rect 34682 34076 34692 34132
rect 34748 34076 36652 34132
rect 36708 34076 36718 34132
rect 36978 34076 36988 34132
rect 37044 34076 37604 34132
rect 40058 34076 40068 34132
rect 40124 34076 40796 34132
rect 40852 34076 40862 34132
rect 13916 34020 13972 34076
rect 30716 34020 30772 34076
rect 4284 33964 4732 34020
rect 4788 33964 10108 34020
rect 10164 33964 10174 34020
rect 13916 33964 15036 34020
rect 15092 33964 15102 34020
rect 20290 33964 20300 34020
rect 20356 33964 22036 34020
rect 22092 33964 22102 34020
rect 23538 33964 23548 34020
rect 23604 33964 25396 34020
rect 25452 33964 25676 34020
rect 25732 33964 25742 34020
rect 30716 33964 32284 34020
rect 32340 33964 32350 34020
rect 34290 33964 34300 34020
rect 34356 33964 35663 34020
rect 35719 33964 35729 34020
rect 42410 33964 42420 34020
rect 42476 33964 45276 34020
rect 45332 33964 45342 34020
rect 45714 33964 45724 34020
rect 45780 33964 45892 34020
rect 45948 33964 45958 34020
rect 46834 33964 46844 34020
rect 46900 33964 47516 34020
rect 47572 33964 47582 34020
rect 3658 33852 3668 33908
rect 3724 33852 5572 33908
rect 5628 33852 5638 33908
rect 6514 33852 6524 33908
rect 6580 33852 7532 33908
rect 7588 33852 7598 33908
rect 7690 33852 7700 33908
rect 7756 33852 11060 33908
rect 11116 33852 11126 33908
rect 12450 33852 12460 33908
rect 12516 33852 14924 33908
rect 14980 33852 14990 33908
rect 21494 33852 21532 33908
rect 21588 33852 21598 33908
rect 21858 33852 21868 33908
rect 21924 33852 22204 33908
rect 22260 33852 22270 33908
rect 22530 33852 22540 33908
rect 22596 33852 23324 33908
rect 23380 33852 23390 33908
rect 23762 33852 23772 33908
rect 23828 33852 24276 33908
rect 24332 33852 24342 33908
rect 26898 33852 26908 33908
rect 26964 33852 27412 33908
rect 41458 33852 41468 33908
rect 41524 33852 42588 33908
rect 42644 33852 42654 33908
rect 44594 33852 44604 33908
rect 44660 33852 44828 33908
rect 44884 33852 44894 33908
rect 8418 33740 8428 33796
rect 8484 33740 10668 33796
rect 10724 33740 10780 33796
rect 10836 33740 10846 33796
rect 12338 33740 12348 33796
rect 12404 33740 13580 33796
rect 13636 33740 13646 33796
rect 17602 33740 17612 33796
rect 17668 33740 17678 33796
rect 18610 33740 18620 33796
rect 18676 33740 20748 33796
rect 20804 33740 20814 33796
rect 21354 33740 21364 33796
rect 21420 33740 22316 33796
rect 22372 33740 22382 33796
rect 25218 33740 25228 33796
rect 25284 33740 26012 33796
rect 26068 33740 26078 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 17612 33684 17668 33740
rect 27356 33684 27412 33852
rect 27906 33740 27916 33796
rect 27972 33740 28140 33796
rect 28196 33740 28206 33796
rect 30118 33740 30156 33796
rect 30212 33740 30222 33796
rect 32134 33740 32172 33796
rect 32228 33740 32238 33796
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 6738 33628 6748 33684
rect 6804 33628 7700 33684
rect 7756 33628 7766 33684
rect 10770 33628 10780 33684
rect 10836 33628 10846 33684
rect 13682 33628 13692 33684
rect 13748 33628 15032 33684
rect 15088 33628 15098 33684
rect 17042 33628 17052 33684
rect 17108 33628 17668 33684
rect 22194 33628 22204 33684
rect 22260 33628 22988 33684
rect 23044 33628 23054 33684
rect 23762 33628 23772 33684
rect 23828 33628 25116 33684
rect 25172 33628 25182 33684
rect 26450 33628 26460 33684
rect 26516 33628 26852 33684
rect 26908 33628 26918 33684
rect 27346 33628 27356 33684
rect 27412 33628 27422 33684
rect 28466 33628 28476 33684
rect 28532 33628 29708 33684
rect 29764 33628 29774 33684
rect 30034 33628 30044 33684
rect 30100 33628 30110 33684
rect 31014 33628 31052 33684
rect 31108 33628 31118 33684
rect 31826 33628 31836 33684
rect 31892 33628 32564 33684
rect 32620 33628 32630 33684
rect 36306 33628 36316 33684
rect 36372 33628 37100 33684
rect 37156 33628 37166 33684
rect 38882 33628 38892 33684
rect 38948 33628 41132 33684
rect 41188 33628 41198 33684
rect 44492 33628 47180 33684
rect 47236 33628 47246 33684
rect 10780 33572 10836 33628
rect 30044 33572 30100 33628
rect 44492 33572 44548 33628
rect 9314 33516 9324 33572
rect 9380 33516 10836 33572
rect 11890 33516 11900 33572
rect 11956 33516 12348 33572
rect 12404 33516 12414 33572
rect 12842 33516 12852 33572
rect 12908 33516 14084 33572
rect 14140 33516 14588 33572
rect 14644 33516 14654 33572
rect 15810 33516 15820 33572
rect 15876 33516 29988 33572
rect 30044 33516 31948 33572
rect 32004 33516 32014 33572
rect 35186 33516 35196 33572
rect 35252 33516 35532 33572
rect 35588 33516 36876 33572
rect 36932 33516 36942 33572
rect 41234 33516 41244 33572
rect 41300 33516 41804 33572
rect 41860 33516 41870 33572
rect 43922 33516 43932 33572
rect 43988 33516 44548 33572
rect 44706 33516 44716 33572
rect 44772 33516 44782 33572
rect 29932 33460 29988 33516
rect 9090 33404 9100 33460
rect 9156 33404 9996 33460
rect 10052 33404 10062 33460
rect 16258 33404 16268 33460
rect 16324 33404 18508 33460
rect 18564 33404 18574 33460
rect 20066 33404 20076 33460
rect 20132 33404 20300 33460
rect 20356 33404 20366 33460
rect 20524 33404 23772 33460
rect 23828 33404 23838 33460
rect 25330 33404 25340 33460
rect 25396 33404 28980 33460
rect 29036 33404 29046 33460
rect 29932 33404 30920 33460
rect 30976 33404 31724 33460
rect 31780 33404 31790 33460
rect 36530 33404 36540 33460
rect 36596 33404 38108 33460
rect 38164 33404 42700 33460
rect 42756 33404 42766 33460
rect 20524 33348 20580 33404
rect 44716 33348 44772 33516
rect 1586 33292 1596 33348
rect 1652 33292 2156 33348
rect 2212 33292 2222 33348
rect 4106 33292 4116 33348
rect 4172 33292 5124 33348
rect 5180 33292 6188 33348
rect 6244 33292 6254 33348
rect 6412 33292 12572 33348
rect 12628 33292 12638 33348
rect 13794 33292 13804 33348
rect 13860 33292 14364 33348
rect 14420 33292 15708 33348
rect 15764 33292 15774 33348
rect 18254 33292 18264 33348
rect 18320 33292 20580 33348
rect 21858 33292 21868 33348
rect 21924 33292 21934 33348
rect 25106 33292 25116 33348
rect 25172 33292 25452 33348
rect 25508 33292 25518 33348
rect 29474 33292 29484 33348
rect 29540 33292 30044 33348
rect 30100 33292 31164 33348
rect 31220 33292 31500 33348
rect 31556 33292 31566 33348
rect 32722 33292 32732 33348
rect 32788 33292 33068 33348
rect 33124 33292 33134 33348
rect 34962 33292 34972 33348
rect 35028 33292 36316 33348
rect 36372 33292 36382 33348
rect 41794 33292 41804 33348
rect 41860 33292 42812 33348
rect 42868 33292 42878 33348
rect 43474 33292 43484 33348
rect 43540 33292 44156 33348
rect 44212 33292 44772 33348
rect 6412 33236 6468 33292
rect 6066 33180 6076 33236
rect 6132 33180 6468 33236
rect 7084 33124 7140 33292
rect 21868 33236 21924 33292
rect 8306 33180 8316 33236
rect 8372 33180 8876 33236
rect 8932 33180 8942 33236
rect 11218 33180 11228 33236
rect 11284 33180 11900 33236
rect 11956 33180 11966 33236
rect 16482 33180 16492 33236
rect 16548 33180 17500 33236
rect 17556 33180 18060 33236
rect 18116 33180 18126 33236
rect 19404 33180 21924 33236
rect 33730 33180 33740 33236
rect 33796 33180 37100 33236
rect 37156 33180 37166 33236
rect 43586 33180 43596 33236
rect 43652 33180 46172 33236
rect 46228 33180 46238 33236
rect 19404 33124 19460 33180
rect 7074 33068 7084 33124
rect 7140 33068 7150 33124
rect 19394 33068 19404 33124
rect 19460 33068 19470 33124
rect 29810 33068 29820 33124
rect 29876 33068 30828 33124
rect 30884 33068 30894 33124
rect 35858 33068 35868 33124
rect 35924 33068 37772 33124
rect 37828 33068 37838 33124
rect 44146 33068 44156 33124
rect 44212 33068 45052 33124
rect 45108 33068 45118 33124
rect 20794 32956 20804 33012
rect 20860 32956 21644 33012
rect 21700 32956 21710 33012
rect 23090 32956 23100 33012
rect 23156 32956 23772 33012
rect 23828 32956 23838 33012
rect 33394 32956 33404 33012
rect 33460 32956 34524 33012
rect 34580 32956 34590 33012
rect 37650 32956 37660 33012
rect 37716 32956 39116 33012
rect 39172 32956 39182 33012
rect 43138 32956 43148 33012
rect 43204 32956 45612 33012
rect 45668 32956 45678 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 11330 32844 11340 32900
rect 11396 32844 15148 32900
rect 23762 32844 23772 32900
rect 23828 32844 32564 32900
rect 33170 32844 33180 32900
rect 33236 32844 35364 32900
rect 35420 32844 35430 32900
rect 38658 32844 38668 32900
rect 38724 32844 40012 32900
rect 40068 32844 40078 32900
rect 15092 32788 15148 32844
rect 1586 32732 1596 32788
rect 1652 32732 3220 32788
rect 3276 32732 4116 32788
rect 4172 32732 4182 32788
rect 9202 32732 9212 32788
rect 9268 32732 11004 32788
rect 11060 32732 11676 32788
rect 11732 32732 12796 32788
rect 12852 32732 12862 32788
rect 15092 32732 15596 32788
rect 15652 32732 15662 32788
rect 15941 32732 15951 32788
rect 16007 32732 18284 32788
rect 18340 32732 21196 32788
rect 21252 32732 29372 32788
rect 29428 32732 30136 32788
rect 30192 32732 30202 32788
rect 15596 32676 15652 32732
rect 32508 32676 32564 32844
rect 32834 32732 32844 32788
rect 32900 32732 33964 32788
rect 34020 32732 35868 32788
rect 35924 32732 37100 32788
rect 37156 32732 37436 32788
rect 37492 32732 38556 32788
rect 38612 32732 38622 32788
rect 39890 32732 39900 32788
rect 39956 32732 40236 32788
rect 40292 32732 40302 32788
rect 41010 32732 41020 32788
rect 41076 32732 41356 32788
rect 41412 32732 41692 32788
rect 41748 32732 41758 32788
rect 43362 32732 43372 32788
rect 43428 32732 48020 32788
rect 48076 32732 48086 32788
rect 12562 32620 12572 32676
rect 12628 32620 14364 32676
rect 14420 32620 14430 32676
rect 15596 32620 23044 32676
rect 23202 32620 23212 32676
rect 23268 32620 23548 32676
rect 23604 32620 25228 32676
rect 25284 32620 25294 32676
rect 27878 32620 27916 32676
rect 27972 32620 27982 32676
rect 30370 32620 30380 32676
rect 30436 32620 32284 32676
rect 32340 32620 32350 32676
rect 32508 32620 36204 32676
rect 36260 32620 36270 32676
rect 46478 32620 46488 32676
rect 46544 32620 47292 32676
rect 47348 32620 47358 32676
rect 22988 32564 23044 32620
rect 6066 32508 6076 32564
rect 6132 32508 6636 32564
rect 6692 32508 6702 32564
rect 10882 32508 10892 32564
rect 10948 32508 14028 32564
rect 14084 32508 14094 32564
rect 16818 32508 16828 32564
rect 16884 32508 18788 32564
rect 18844 32508 18854 32564
rect 19282 32508 19292 32564
rect 19348 32508 20748 32564
rect 20804 32508 20814 32564
rect 22988 32508 26292 32564
rect 26348 32508 26358 32564
rect 29250 32508 29260 32564
rect 29316 32508 29326 32564
rect 38854 32508 38892 32564
rect 38948 32508 38958 32564
rect 39162 32508 39172 32564
rect 39228 32508 41748 32564
rect 41804 32508 41814 32564
rect 45602 32508 45612 32564
rect 45668 32508 46284 32564
rect 46340 32508 47628 32564
rect 47684 32508 48188 32564
rect 48244 32508 48254 32564
rect 17770 32396 17780 32452
rect 17836 32396 18620 32452
rect 18676 32396 18686 32452
rect 4284 32284 5740 32340
rect 5796 32284 5806 32340
rect 4284 32228 4340 32284
rect 29260 32228 29316 32508
rect 35522 32396 35532 32452
rect 35588 32396 36092 32452
rect 36148 32396 39004 32452
rect 39060 32396 39070 32452
rect 39778 32396 39788 32452
rect 39844 32396 40460 32452
rect 40516 32396 43932 32452
rect 43988 32396 43998 32452
rect 43596 32228 43652 32396
rect 49200 32340 50000 32368
rect 48290 32284 48300 32340
rect 48356 32284 50000 32340
rect 49200 32256 50000 32284
rect 4274 32172 4284 32228
rect 4340 32172 4350 32228
rect 11666 32172 11676 32228
rect 11732 32172 13916 32228
rect 13972 32172 15148 32228
rect 17154 32172 17164 32228
rect 17220 32172 17612 32228
rect 17668 32172 25004 32228
rect 25060 32172 25070 32228
rect 29138 32172 29148 32228
rect 29204 32172 29316 32228
rect 38210 32172 38220 32228
rect 38276 32172 38556 32228
rect 38612 32172 38622 32228
rect 43586 32172 43596 32228
rect 43652 32172 43662 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 11676 32116 11732 32172
rect 11564 32060 11732 32116
rect 11564 32004 11620 32060
rect 4162 31948 4172 32004
rect 4228 31948 4238 32004
rect 4834 31948 4844 32004
rect 4900 31948 6076 32004
rect 6132 31948 6142 32004
rect 7746 31948 7756 32004
rect 7812 31948 8316 32004
rect 8372 31948 8382 32004
rect 11452 31948 11620 32004
rect 12226 31948 12236 32004
rect 12292 31948 12460 32004
rect 12516 31948 13580 32004
rect 13636 31948 14868 32004
rect 14924 31948 14934 32004
rect 4172 31892 4228 31948
rect 2930 31836 2940 31892
rect 2996 31836 3500 31892
rect 3556 31836 3566 31892
rect 4172 31836 5628 31892
rect 5684 31836 5694 31892
rect 11452 31780 11508 31948
rect 12086 31836 12124 31892
rect 12180 31836 12190 31892
rect 15092 31780 15148 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 16258 32060 16268 32116
rect 16324 32060 19404 32116
rect 19460 32060 19470 32116
rect 21970 32060 21980 32116
rect 22036 32060 22540 32116
rect 22596 32060 22606 32116
rect 45798 32060 45836 32116
rect 45892 32060 45902 32116
rect 18946 31948 18956 32004
rect 19012 31948 20412 32004
rect 20468 31948 20478 32004
rect 22978 31948 22988 32004
rect 23044 31948 23772 32004
rect 23828 31948 24556 32004
rect 24612 31948 25116 32004
rect 25172 31948 25182 32004
rect 26562 31948 26572 32004
rect 26628 31948 26684 32004
rect 26740 31948 26750 32004
rect 28018 31948 28028 32004
rect 28084 31948 28364 32004
rect 28420 31948 28430 32004
rect 29026 31948 29036 32004
rect 29092 31948 29540 32004
rect 29596 31948 29606 32004
rect 37314 31948 37324 32004
rect 37380 31948 37390 32004
rect 41234 31948 41244 32004
rect 41300 31948 41916 32004
rect 41972 31948 41982 32004
rect 43866 31948 43876 32004
rect 43932 31948 44716 32004
rect 44772 31948 44782 32004
rect 37324 31892 37380 31948
rect 15698 31836 15708 31892
rect 15764 31836 16828 31892
rect 16884 31836 17388 31892
rect 17444 31836 17454 31892
rect 21970 31836 21980 31892
rect 22036 31836 23884 31892
rect 23940 31836 23950 31892
rect 27010 31836 27020 31892
rect 27076 31836 28532 31892
rect 28588 31836 28598 31892
rect 36306 31836 36316 31892
rect 36372 31836 37380 31892
rect 39666 31836 39676 31892
rect 39732 31836 41692 31892
rect 41748 31836 41758 31892
rect 2594 31724 2604 31780
rect 2660 31724 3052 31780
rect 3108 31724 3118 31780
rect 5282 31724 5292 31780
rect 5348 31724 6076 31780
rect 6132 31724 6142 31780
rect 7970 31724 7980 31780
rect 8036 31724 8540 31780
rect 8596 31724 8606 31780
rect 9538 31724 9548 31780
rect 9604 31724 10220 31780
rect 10276 31724 10286 31780
rect 11442 31724 11452 31780
rect 11508 31724 11518 31780
rect 13458 31724 13468 31780
rect 13524 31724 14476 31780
rect 14532 31724 14542 31780
rect 15092 31724 15876 31780
rect 15932 31724 18620 31780
rect 18676 31724 19628 31780
rect 19684 31724 22428 31780
rect 22484 31724 22494 31780
rect 25834 31724 25844 31780
rect 25900 31724 27020 31780
rect 27076 31724 27086 31780
rect 27234 31724 27244 31780
rect 27300 31724 27916 31780
rect 27972 31724 27982 31780
rect 28110 31724 28120 31780
rect 28196 31724 28214 31780
rect 28354 31724 28364 31780
rect 28420 31724 29036 31780
rect 29092 31724 29102 31780
rect 30930 31724 30940 31780
rect 30996 31724 31836 31780
rect 31892 31724 31902 31780
rect 32890 31724 32900 31780
rect 32956 31724 35196 31780
rect 35252 31724 35262 31780
rect 42354 31724 42364 31780
rect 42420 31724 43036 31780
rect 43092 31724 44044 31780
rect 44100 31724 44110 31780
rect 3602 31612 3612 31668
rect 3668 31612 4452 31668
rect 4508 31612 5124 31668
rect 5180 31612 5190 31668
rect 8540 31556 8596 31724
rect 9762 31612 9772 31668
rect 9828 31612 9996 31668
rect 10052 31612 12460 31668
rect 12516 31612 12526 31668
rect 21298 31612 21308 31668
rect 21364 31612 22204 31668
rect 22260 31612 22270 31668
rect 27906 31612 27916 31668
rect 27972 31612 28476 31668
rect 28532 31612 29260 31668
rect 29316 31612 32508 31668
rect 32564 31612 32574 31668
rect 40226 31612 40236 31668
rect 40292 31612 40684 31668
rect 40740 31612 40750 31668
rect 8540 31500 10556 31556
rect 10612 31500 10622 31556
rect 12086 31500 12124 31556
rect 12180 31500 12190 31556
rect 13964 31500 13974 31556
rect 14030 31500 14252 31556
rect 14308 31500 14318 31556
rect 16706 31500 16716 31556
rect 16772 31500 17164 31556
rect 17220 31500 18060 31556
rect 18116 31500 23996 31556
rect 24052 31500 24062 31556
rect 24770 31500 24780 31556
rect 24836 31500 25284 31556
rect 25340 31500 30212 31556
rect 30268 31500 30278 31556
rect 30706 31500 30716 31556
rect 30772 31500 42756 31556
rect 10070 31388 10108 31444
rect 10164 31388 10174 31444
rect 23090 31388 23100 31444
rect 23156 31388 23604 31444
rect 23660 31388 23670 31444
rect 24882 31388 24892 31444
rect 24948 31388 25844 31444
rect 25900 31388 25910 31444
rect 27794 31388 27804 31444
rect 27860 31388 28812 31444
rect 28868 31388 28878 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 42700 31332 42756 31500
rect 14140 31276 14588 31332
rect 14644 31276 14654 31332
rect 20626 31276 20636 31332
rect 20692 31276 21028 31332
rect 23874 31276 23884 31332
rect 23940 31276 25116 31332
rect 25172 31276 29596 31332
rect 29652 31276 29662 31332
rect 30258 31276 30268 31332
rect 30324 31276 31612 31332
rect 31668 31276 31678 31332
rect 42690 31276 42700 31332
rect 42756 31276 42766 31332
rect 13206 31164 13244 31220
rect 13300 31164 13310 31220
rect 6402 31052 6412 31108
rect 6468 31052 7812 31108
rect 7868 31052 7878 31108
rect 14140 30996 14196 31276
rect 20972 31220 21028 31276
rect 16482 31164 16492 31220
rect 16548 31164 18284 31220
rect 18340 31164 20748 31220
rect 20804 31164 20814 31220
rect 20972 31164 26740 31220
rect 26796 31164 26806 31220
rect 27010 31164 27020 31220
rect 27076 31164 28700 31220
rect 28756 31164 28766 31220
rect 32106 31164 32116 31220
rect 32172 31164 33944 31220
rect 34000 31164 34010 31220
rect 39442 31164 39452 31220
rect 39508 31164 42252 31220
rect 42308 31164 42318 31220
rect 43586 31164 43596 31220
rect 43652 31164 44716 31220
rect 44772 31164 44782 31220
rect 16594 31052 16604 31108
rect 16660 31052 17948 31108
rect 18004 31052 18014 31108
rect 19394 31052 19404 31108
rect 19460 31052 20188 31108
rect 20244 31052 20254 31108
rect 20402 31052 20412 31108
rect 20468 31052 21756 31108
rect 21812 31052 21822 31108
rect 23538 31052 23548 31108
rect 23604 31052 24668 31108
rect 24724 31052 25228 31108
rect 25284 31052 25294 31108
rect 28242 31052 28252 31108
rect 28308 31052 30604 31108
rect 30660 31052 31164 31108
rect 31220 31052 31230 31108
rect 36828 31052 36838 31108
rect 36894 31052 40404 31108
rect 40460 31052 40470 31108
rect 46162 31052 46172 31108
rect 46228 31052 47628 31108
rect 47684 31052 47694 31108
rect 6178 30940 6188 30996
rect 6244 30940 6748 30996
rect 6804 30940 6814 30996
rect 6962 30940 6972 30996
rect 7028 30940 8204 30996
rect 8260 30940 8540 30996
rect 8596 30940 9884 30996
rect 9940 30940 9950 30996
rect 10098 30940 10108 30996
rect 10164 30940 14140 30996
rect 14196 30940 14206 30996
rect 17658 30940 17668 30996
rect 17724 30940 18620 30996
rect 18676 30940 20636 30996
rect 20692 30940 20702 30996
rect 23202 30940 23212 30996
rect 23268 30940 24276 30996
rect 24332 30940 24342 30996
rect 25638 30940 25676 30996
rect 25732 30940 25742 30996
rect 29362 30940 29372 30996
rect 29428 30940 30716 30996
rect 30772 30940 30782 30996
rect 32274 30940 32284 30996
rect 32340 30940 33068 30996
rect 33124 30940 33134 30996
rect 34178 30940 34188 30996
rect 34244 30940 35512 30996
rect 35568 30940 35578 30996
rect 36530 30940 36540 30996
rect 36596 30940 38892 30996
rect 38948 30940 38958 30996
rect 5898 30828 5908 30884
rect 5964 30828 8428 30884
rect 8484 30828 8494 30884
rect 18386 30828 18396 30884
rect 18452 30828 18732 30884
rect 18788 30828 18798 30884
rect 19506 30828 19516 30884
rect 19572 30828 20132 30884
rect 20188 30828 20972 30884
rect 21028 30828 21038 30884
rect 29194 30828 29204 30884
rect 29260 30828 32040 30884
rect 32096 30828 32106 30884
rect 36194 30828 36204 30884
rect 36260 30828 38332 30884
rect 38388 30828 38398 30884
rect 3052 30716 4844 30772
rect 4900 30716 4910 30772
rect 20514 30716 20524 30772
rect 20580 30716 21644 30772
rect 21700 30716 21710 30772
rect 27990 30716 28028 30772
rect 28084 30716 28094 30772
rect 30454 30716 30492 30772
rect 30548 30716 30558 30772
rect 3052 30660 3108 30716
rect 2482 30604 2492 30660
rect 2548 30604 3052 30660
rect 3108 30604 3118 30660
rect 7746 30604 7756 30660
rect 7812 30604 8316 30660
rect 8372 30604 8382 30660
rect 13794 30604 13804 30660
rect 13860 30604 13870 30660
rect 15474 30604 15484 30660
rect 15540 30604 20636 30660
rect 20692 30604 20702 30660
rect 20850 30604 20860 30660
rect 20916 30604 21420 30660
rect 21476 30604 21486 30660
rect 25750 30604 25788 30660
rect 25844 30604 25854 30660
rect 28130 30604 28140 30660
rect 28196 30604 29540 30660
rect 29596 30604 29606 30660
rect 36306 30604 36316 30660
rect 36372 30604 38332 30660
rect 38388 30604 38398 30660
rect 40562 30604 40572 30660
rect 40628 30604 42588 30660
rect 42644 30604 42654 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 7074 30492 7084 30548
rect 7140 30492 7150 30548
rect 10742 30492 10780 30548
rect 10836 30492 10846 30548
rect 7084 30436 7140 30492
rect 4366 30380 4376 30436
rect 4432 30380 7140 30436
rect 8530 30380 8540 30436
rect 8596 30380 9212 30436
rect 9268 30380 9278 30436
rect 10994 30380 11004 30436
rect 11060 30380 13524 30436
rect 6290 30268 6300 30324
rect 6356 30268 8764 30324
rect 8820 30268 8830 30324
rect 9314 30268 9324 30324
rect 9380 30268 9390 30324
rect 9324 30212 9380 30268
rect 13468 30212 13524 30380
rect 3490 30156 3500 30212
rect 3556 30156 4172 30212
rect 4228 30156 4238 30212
rect 8194 30156 8204 30212
rect 8260 30156 9380 30212
rect 10994 30156 11004 30212
rect 11060 30156 11070 30212
rect 13458 30156 13468 30212
rect 13524 30156 13534 30212
rect 11004 30100 11060 30156
rect 13804 30100 13860 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 18834 30492 18844 30548
rect 18900 30492 20076 30548
rect 20132 30492 21980 30548
rect 22036 30492 22046 30548
rect 23650 30492 23660 30548
rect 23716 30492 34748 30548
rect 34804 30492 34814 30548
rect 38938 30492 38948 30548
rect 39004 30492 39452 30548
rect 39508 30492 39518 30548
rect 43474 30492 43484 30548
rect 43540 30492 43932 30548
rect 43988 30492 43998 30548
rect 15250 30380 15260 30436
rect 15316 30380 28252 30436
rect 28308 30380 28318 30436
rect 29698 30380 29708 30436
rect 29764 30380 29802 30436
rect 32498 30380 32508 30436
rect 32564 30380 33516 30436
rect 33572 30380 33582 30436
rect 44482 30380 44492 30436
rect 44548 30380 45668 30436
rect 45724 30380 45734 30436
rect 17938 30268 17948 30324
rect 18004 30268 18508 30324
rect 18564 30268 19516 30324
rect 19572 30268 19582 30324
rect 20626 30268 20636 30324
rect 20692 30268 21812 30324
rect 30482 30268 30492 30324
rect 30548 30268 30940 30324
rect 30996 30268 31006 30324
rect 32386 30268 32396 30324
rect 32452 30268 33180 30324
rect 33236 30268 33246 30324
rect 38882 30268 38892 30324
rect 38948 30268 39340 30324
rect 39396 30268 39406 30324
rect 21756 30212 21812 30268
rect 2818 30044 2828 30100
rect 2884 30044 4620 30100
rect 4676 30044 4956 30100
rect 5012 30044 5022 30100
rect 8082 30044 8092 30100
rect 8148 30044 8820 30100
rect 8876 30044 9156 30100
rect 9212 30044 9222 30100
rect 9286 30044 9324 30100
rect 9380 30044 9390 30100
rect 11004 30044 13356 30100
rect 13412 30044 13860 30100
rect 13916 30156 14344 30212
rect 14400 30156 14410 30212
rect 15026 30156 15036 30212
rect 15092 30156 18340 30212
rect 18396 30156 18406 30212
rect 21756 30156 22540 30212
rect 22596 30156 22606 30212
rect 25442 30156 25452 30212
rect 25508 30156 26796 30212
rect 26852 30156 26862 30212
rect 28242 30156 28252 30212
rect 28308 30156 29148 30212
rect 29204 30156 29214 30212
rect 30594 30156 30604 30212
rect 30660 30156 32172 30212
rect 32228 30156 32238 30212
rect 33618 30156 33628 30212
rect 33684 30156 35312 30212
rect 35368 30156 35378 30212
rect 35802 30156 35812 30212
rect 35868 30156 36428 30212
rect 36484 30156 38500 30212
rect 38556 30156 38566 30212
rect 39218 30156 39228 30212
rect 39284 30156 41692 30212
rect 41748 30156 41758 30212
rect 43810 30156 43820 30212
rect 43876 30156 45388 30212
rect 45444 30156 45454 30212
rect 45938 30156 45948 30212
rect 46004 30156 47964 30212
rect 48020 30156 48030 30212
rect 13916 29988 13972 30156
rect 20402 30044 20412 30100
rect 20468 30044 21868 30100
rect 21924 30044 21934 30100
rect 24658 30044 24668 30100
rect 24724 30044 25228 30100
rect 25284 30044 25676 30100
rect 25732 30044 25742 30100
rect 27906 30044 27916 30100
rect 27972 30044 28924 30100
rect 28980 30044 29260 30100
rect 29316 30044 29326 30100
rect 30818 30044 30828 30100
rect 30884 30044 31276 30100
rect 31332 30044 32564 30100
rect 32620 30044 32630 30100
rect 36530 30044 36540 30100
rect 36596 30044 38220 30100
rect 38276 30044 38286 30100
rect 38444 30044 38780 30100
rect 38836 30044 38846 30100
rect 42690 30044 42700 30100
rect 42756 30044 45164 30100
rect 45220 30044 45724 30100
rect 45780 30044 45790 30100
rect 38444 29988 38500 30044
rect 7410 29932 7420 29988
rect 7476 29932 13972 29988
rect 14214 29932 14252 29988
rect 14308 29932 14318 29988
rect 16482 29932 16492 29988
rect 16548 29932 17500 29988
rect 17556 29932 17566 29988
rect 20738 29932 20748 29988
rect 20804 29932 21084 29988
rect 21140 29932 21150 29988
rect 23986 29932 23996 29988
rect 24052 29932 24892 29988
rect 24948 29932 24958 29988
rect 30146 29932 30156 29988
rect 30212 29932 33180 29988
rect 33236 29932 33246 29988
rect 37090 29932 37100 29988
rect 37156 29932 37772 29988
rect 37828 29932 38500 29988
rect 38612 29932 40236 29988
rect 40292 29932 40302 29988
rect 20188 29820 21756 29876
rect 21812 29820 21822 29876
rect 25778 29820 25788 29876
rect 25844 29820 26124 29876
rect 26180 29820 26190 29876
rect 26338 29820 26348 29876
rect 26404 29820 26442 29876
rect 33730 29820 33740 29876
rect 33796 29820 38388 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 3332 29708 5740 29764
rect 5796 29708 5806 29764
rect 18834 29708 18844 29764
rect 18900 29708 19628 29764
rect 19684 29708 19694 29764
rect 3332 29652 3388 29708
rect 20188 29652 20244 29820
rect 3042 29596 3052 29652
rect 3108 29596 3388 29652
rect 4946 29596 4956 29652
rect 5012 29596 5516 29652
rect 5572 29596 7476 29652
rect 7532 29596 13244 29652
rect 13300 29596 13310 29652
rect 15474 29596 15484 29652
rect 15540 29596 16380 29652
rect 16436 29596 16446 29652
rect 17938 29596 17948 29652
rect 18004 29596 19740 29652
rect 19796 29596 20244 29652
rect 20972 29708 30548 29764
rect 30604 29708 30828 29764
rect 30884 29708 30894 29764
rect 34038 29708 34076 29764
rect 34132 29708 34142 29764
rect 36642 29708 36652 29764
rect 36708 29708 36718 29764
rect 20972 29540 21028 29708
rect 22530 29596 22540 29652
rect 22596 29596 22764 29652
rect 22820 29596 23828 29652
rect 23884 29596 23894 29652
rect 23986 29596 23996 29652
rect 24052 29596 24220 29652
rect 24276 29596 26012 29652
rect 26068 29596 26078 29652
rect 27570 29596 27580 29652
rect 27636 29596 34524 29652
rect 34580 29596 34590 29652
rect 36652 29540 36708 29708
rect 38332 29652 38388 29820
rect 38546 29708 38556 29764
rect 38612 29708 38668 29932
rect 38332 29596 39060 29652
rect 39116 29596 39126 29652
rect 40226 29596 40236 29652
rect 40292 29596 42196 29652
rect 42252 29596 42262 29652
rect 3266 29484 3276 29540
rect 3332 29484 5348 29540
rect 5404 29484 5414 29540
rect 5618 29484 5628 29540
rect 5684 29484 5852 29540
rect 5908 29484 5918 29540
rect 10658 29484 10668 29540
rect 10724 29484 21028 29540
rect 21186 29484 21196 29540
rect 21252 29484 22316 29540
rect 22372 29484 23436 29540
rect 23492 29484 23502 29540
rect 24546 29484 24556 29540
rect 24612 29484 25340 29540
rect 25396 29484 25406 29540
rect 34850 29484 34860 29540
rect 34916 29484 37192 29540
rect 37248 29484 37548 29540
rect 37604 29484 37614 29540
rect 3332 29372 3724 29428
rect 3780 29372 3790 29428
rect 5058 29372 5068 29428
rect 5124 29372 6636 29428
rect 6692 29372 6702 29428
rect 8306 29372 8316 29428
rect 8372 29372 8988 29428
rect 9044 29372 9054 29428
rect 9650 29372 9660 29428
rect 9716 29372 9726 29428
rect 12338 29372 12348 29428
rect 12404 29372 12796 29428
rect 12852 29372 12862 29428
rect 14578 29372 14588 29428
rect 14644 29372 14924 29428
rect 14980 29372 15484 29428
rect 15540 29372 15550 29428
rect 20010 29372 20020 29428
rect 20076 29372 20188 29428
rect 20244 29372 20254 29428
rect 20514 29372 20524 29428
rect 20580 29372 20860 29428
rect 20916 29372 20926 29428
rect 21802 29372 21812 29428
rect 21868 29372 22204 29428
rect 22260 29372 22270 29428
rect 22978 29372 22988 29428
rect 23044 29372 23548 29428
rect 25554 29372 25564 29428
rect 25620 29372 25676 29428
rect 25732 29372 25742 29428
rect 26002 29372 26012 29428
rect 26068 29372 27188 29428
rect 27244 29372 27254 29428
rect 27906 29372 27916 29428
rect 27972 29372 29148 29428
rect 29204 29372 29214 29428
rect 31938 29372 31948 29428
rect 32004 29372 33740 29428
rect 33796 29372 33806 29428
rect 36082 29372 36092 29428
rect 36148 29372 37324 29428
rect 37380 29372 37390 29428
rect 40562 29372 40572 29428
rect 40628 29372 41804 29428
rect 41860 29372 41870 29428
rect 45042 29372 45052 29428
rect 45108 29372 48300 29428
rect 48356 29372 48366 29428
rect 3332 29316 3388 29372
rect 1810 29260 1820 29316
rect 1876 29260 2772 29316
rect 2828 29260 3388 29316
rect 4590 29260 4600 29316
rect 4656 29260 5516 29316
rect 5572 29260 5582 29316
rect 4060 29148 6076 29204
rect 6132 29148 6142 29204
rect 4060 28980 4116 29148
rect 9314 29036 9324 29092
rect 9380 29036 9390 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 9324 28980 9380 29036
rect 9660 28980 9716 29372
rect 23492 29316 23548 29372
rect 20402 29260 20412 29316
rect 20468 29260 22652 29316
rect 22708 29260 22718 29316
rect 23492 29260 24332 29316
rect 24388 29260 26460 29316
rect 26516 29260 31612 29316
rect 31668 29260 31678 29316
rect 34962 29260 34972 29316
rect 35028 29260 35476 29316
rect 35532 29260 35542 29316
rect 44482 29260 44492 29316
rect 44548 29260 45948 29316
rect 46004 29260 46014 29316
rect 44492 29204 44548 29260
rect 17546 29148 17556 29204
rect 17612 29148 18956 29204
rect 19012 29148 19404 29204
rect 19460 29148 19470 29204
rect 21074 29148 21084 29204
rect 21140 29148 21532 29204
rect 21588 29148 21598 29204
rect 25218 29148 25228 29204
rect 25284 29148 26348 29204
rect 26404 29148 26740 29204
rect 26796 29148 27748 29204
rect 27804 29148 32284 29204
rect 32340 29148 33460 29204
rect 33516 29148 37660 29204
rect 37716 29148 39620 29204
rect 39676 29148 40236 29204
rect 40292 29148 41244 29204
rect 41300 29148 41310 29204
rect 42588 29148 44548 29204
rect 46162 29148 46172 29204
rect 46228 29148 47964 29204
rect 48020 29148 48030 29204
rect 42588 29092 42644 29148
rect 11442 29036 11452 29092
rect 11508 29036 12684 29092
rect 12740 29036 14140 29092
rect 14196 29036 15036 29092
rect 15092 29036 15596 29092
rect 15652 29036 15662 29092
rect 23202 29036 23212 29092
rect 23268 29036 26908 29092
rect 30034 29036 30044 29092
rect 30100 29036 30110 29092
rect 30604 29036 31892 29092
rect 37146 29036 37156 29092
rect 37212 29036 42644 29092
rect 42802 29036 42812 29092
rect 42868 29036 44940 29092
rect 44996 29036 45006 29092
rect 26852 28980 26908 29036
rect 30044 28980 30100 29036
rect 30604 28980 30660 29036
rect 31836 28980 31892 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 4050 28924 4060 28980
rect 4116 28924 4126 28980
rect 5506 28924 5516 28980
rect 5572 28924 8260 28980
rect 8418 28924 8428 28980
rect 8484 28924 9380 28980
rect 9650 28924 9660 28980
rect 9716 28924 9726 28980
rect 18162 28924 18172 28980
rect 18228 28924 18620 28980
rect 18676 28924 21420 28980
rect 21476 28924 21486 28980
rect 26852 28924 29988 28980
rect 30044 28924 30660 28980
rect 31826 28924 31836 28980
rect 31892 28924 31902 28980
rect 37650 28924 37660 28980
rect 37716 28924 37996 28980
rect 38052 28924 38062 28980
rect 38322 28924 38332 28980
rect 38388 28924 38668 28980
rect 38724 28924 38734 28980
rect 41122 28924 41132 28980
rect 41188 28924 43372 28980
rect 43428 28924 43438 28980
rect 8204 28868 8260 28924
rect 4162 28812 4172 28868
rect 4228 28812 4844 28868
rect 4900 28812 5740 28868
rect 5796 28812 5806 28868
rect 8204 28812 9324 28868
rect 9380 28812 9864 28868
rect 9920 28812 9930 28868
rect 11330 28812 11340 28868
rect 11396 28812 12236 28868
rect 12292 28812 12302 28868
rect 19506 28812 19516 28868
rect 19572 28812 19852 28868
rect 19908 28812 19918 28868
rect 21690 28812 21700 28868
rect 21756 28812 22428 28868
rect 22484 28812 22494 28868
rect 23062 28812 23100 28868
rect 23156 28812 23166 28868
rect 29138 28812 29148 28868
rect 29204 28812 29708 28868
rect 29764 28812 29774 28868
rect 29932 28756 29988 28924
rect 30146 28812 30156 28868
rect 30212 28812 32844 28868
rect 32900 28812 33404 28868
rect 33460 28812 33470 28868
rect 34738 28812 34748 28868
rect 34804 28812 34814 28868
rect 36306 28812 36316 28868
rect 36372 28812 39228 28868
rect 39284 28812 40124 28868
rect 40180 28812 40190 28868
rect 42466 28812 42476 28868
rect 42532 28812 43708 28868
rect 43764 28812 43774 28868
rect 34748 28756 34804 28812
rect 3714 28700 3724 28756
rect 3780 28700 6300 28756
rect 6356 28700 6366 28756
rect 20402 28700 20412 28756
rect 20468 28700 21140 28756
rect 21410 28700 21420 28756
rect 21476 28700 23884 28756
rect 23940 28700 23950 28756
rect 26852 28700 29708 28756
rect 29764 28700 29774 28756
rect 29932 28700 32564 28756
rect 34748 28700 37156 28756
rect 37212 28700 37222 28756
rect 41234 28700 41244 28756
rect 41300 28700 44324 28756
rect 44380 28700 45388 28756
rect 45444 28700 45454 28756
rect 21084 28644 21140 28700
rect 1698 28588 1708 28644
rect 1764 28588 4508 28644
rect 4564 28588 4574 28644
rect 5618 28588 5628 28644
rect 5684 28588 7420 28644
rect 7476 28588 7486 28644
rect 8286 28588 8296 28644
rect 8352 28588 10612 28644
rect 10668 28588 10678 28644
rect 14354 28588 14364 28644
rect 14420 28588 15372 28644
rect 15428 28588 15438 28644
rect 19730 28588 19740 28644
rect 19796 28588 20300 28644
rect 20356 28588 20916 28644
rect 20972 28588 20982 28644
rect 21084 28588 22260 28644
rect 22316 28588 24220 28644
rect 24276 28588 24286 28644
rect 25526 28588 25564 28644
rect 25620 28588 25630 28644
rect 14018 28476 14028 28532
rect 14084 28476 15036 28532
rect 15092 28476 15484 28532
rect 15540 28476 15550 28532
rect 17710 28476 17720 28532
rect 17776 28476 17948 28532
rect 18004 28476 18014 28532
rect 18274 28476 18284 28532
rect 18340 28476 19180 28532
rect 19236 28476 19246 28532
rect 19506 28476 19516 28532
rect 19572 28476 20524 28532
rect 20580 28476 20590 28532
rect 26534 28476 26572 28532
rect 26628 28476 26638 28532
rect 26852 28420 26908 28700
rect 27290 28588 27300 28644
rect 27356 28588 30604 28644
rect 30660 28588 31724 28644
rect 31780 28588 31790 28644
rect 32508 28588 32564 28700
rect 32620 28588 33012 28644
rect 33068 28588 33236 28644
rect 33394 28588 33404 28644
rect 33460 28588 34504 28644
rect 34560 28588 34570 28644
rect 34738 28588 34748 28644
rect 34804 28588 36072 28644
rect 36128 28588 36138 28644
rect 41010 28588 41020 28644
rect 41076 28588 43260 28644
rect 43316 28588 45836 28644
rect 45892 28588 48300 28644
rect 48356 28588 48366 28644
rect 33180 28532 33236 28588
rect 28578 28476 28588 28532
rect 28644 28476 29484 28532
rect 29540 28476 29550 28532
rect 33180 28476 33628 28532
rect 33684 28476 33694 28532
rect 42028 28420 42084 28588
rect 5170 28364 5180 28420
rect 5236 28364 6076 28420
rect 6132 28364 6142 28420
rect 6402 28364 6412 28420
rect 6468 28364 6860 28420
rect 6916 28364 7140 28420
rect 7196 28364 7206 28420
rect 10994 28364 11004 28420
rect 11060 28364 12180 28420
rect 12236 28364 15148 28420
rect 15204 28364 15214 28420
rect 23426 28364 23436 28420
rect 23492 28364 26908 28420
rect 27570 28364 27580 28420
rect 27636 28364 28476 28420
rect 28532 28364 29036 28420
rect 29092 28364 29102 28420
rect 30044 28364 32732 28420
rect 32788 28364 32798 28420
rect 35858 28364 35868 28420
rect 35924 28364 37436 28420
rect 37492 28364 37502 28420
rect 42018 28364 42028 28420
rect 42084 28364 42094 28420
rect 30044 28308 30100 28364
rect 15250 28252 15260 28308
rect 15316 28252 15484 28308
rect 15540 28252 15550 28308
rect 24434 28252 24444 28308
rect 24500 28252 25452 28308
rect 25508 28252 26572 28308
rect 26628 28252 26638 28308
rect 28802 28252 28812 28308
rect 28868 28252 30044 28308
rect 30100 28252 30110 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 22866 28140 22876 28196
rect 22932 28140 25116 28196
rect 25172 28140 25182 28196
rect 25666 28140 25676 28196
rect 25732 28140 35756 28196
rect 35812 28140 35822 28196
rect 6962 28028 6972 28084
rect 7028 28028 7476 28084
rect 7532 28028 7542 28084
rect 10210 28028 10220 28084
rect 10276 28028 11340 28084
rect 11396 28028 11900 28084
rect 11956 28028 11966 28084
rect 19730 28028 19740 28084
rect 19796 28028 20188 28084
rect 20244 28028 20254 28084
rect 29362 28028 29372 28084
rect 29428 28028 29438 28084
rect 32554 28028 32564 28084
rect 32620 28028 33740 28084
rect 33796 28028 34972 28084
rect 35028 28028 35038 28084
rect 29372 27972 29428 28028
rect 4890 27916 4900 27972
rect 4956 27916 6188 27972
rect 6244 27916 6804 27972
rect 6860 27916 6870 27972
rect 8922 27916 8932 27972
rect 8988 27916 10892 27972
rect 10948 27916 10958 27972
rect 11218 27916 11228 27972
rect 11284 27916 13468 27972
rect 13524 27916 13534 27972
rect 13794 27916 13804 27972
rect 13860 27916 14476 27972
rect 14532 27916 14542 27972
rect 26842 27916 26852 27972
rect 26908 27916 28252 27972
rect 28308 27916 28812 27972
rect 28868 27916 29428 27972
rect 32106 27916 32116 27972
rect 32172 27916 45052 27972
rect 45108 27916 45118 27972
rect 11228 27860 11284 27916
rect 5954 27804 5964 27860
rect 6020 27804 6636 27860
rect 6692 27804 7756 27860
rect 7812 27804 7822 27860
rect 8026 27804 8036 27860
rect 8092 27804 9324 27860
rect 9380 27804 9390 27860
rect 10434 27804 10444 27860
rect 10500 27804 10780 27860
rect 10836 27804 11284 27860
rect 12002 27804 12012 27860
rect 12068 27804 12460 27860
rect 12516 27804 12526 27860
rect 12674 27804 12684 27860
rect 12740 27804 12908 27860
rect 12964 27804 13020 27860
rect 13076 27804 14028 27860
rect 14084 27804 14094 27860
rect 14700 27748 14756 27860
rect 14812 27804 14822 27860
rect 15362 27804 15372 27860
rect 15428 27804 15596 27860
rect 15652 27804 15662 27860
rect 16930 27804 16940 27860
rect 16996 27804 18284 27860
rect 18340 27804 18350 27860
rect 26002 27804 26012 27860
rect 26068 27804 26348 27860
rect 26404 27804 27020 27860
rect 27076 27804 27636 27860
rect 27692 27804 27702 27860
rect 27794 27804 27804 27860
rect 27860 27804 29036 27860
rect 29092 27804 29102 27860
rect 37314 27804 37324 27860
rect 37380 27804 38444 27860
rect 38500 27804 38510 27860
rect 41010 27804 41020 27860
rect 41076 27804 41804 27860
rect 41860 27804 43036 27860
rect 43092 27804 43102 27860
rect 45378 27804 45388 27860
rect 45444 27804 46060 27860
rect 46116 27804 46126 27860
rect 46834 27804 46844 27860
rect 46900 27804 47292 27860
rect 47348 27804 47358 27860
rect 46844 27748 46900 27804
rect 9090 27692 9100 27748
rect 9156 27692 14140 27748
rect 14196 27692 14756 27748
rect 15026 27692 15036 27748
rect 10546 27580 10556 27636
rect 10612 27580 12124 27636
rect 12180 27580 14140 27636
rect 14196 27580 14206 27636
rect 14354 27580 14364 27636
rect 14420 27580 14430 27636
rect 5282 27468 5292 27524
rect 5348 27468 5740 27524
rect 5796 27468 6524 27524
rect 6580 27468 7868 27524
rect 7924 27468 7934 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 14364 27412 14420 27580
rect 14700 27524 14756 27692
rect 15092 27636 15148 27748
rect 20626 27692 20636 27748
rect 20692 27692 22652 27748
rect 22708 27692 23100 27748
rect 23156 27692 23166 27748
rect 28186 27692 28196 27748
rect 28252 27692 30940 27748
rect 30996 27692 31006 27748
rect 33898 27692 33908 27748
rect 33964 27692 38332 27748
rect 38388 27692 38398 27748
rect 41122 27692 41132 27748
rect 41188 27692 41198 27748
rect 44706 27692 44716 27748
rect 44772 27692 46900 27748
rect 41132 27636 41188 27692
rect 15092 27580 15372 27636
rect 15428 27580 15438 27636
rect 28914 27580 28924 27636
rect 28980 27580 29596 27636
rect 29652 27580 29662 27636
rect 37538 27580 37548 27636
rect 37604 27580 37996 27636
rect 38052 27580 39956 27636
rect 40012 27580 41188 27636
rect 43026 27580 43036 27636
rect 43092 27580 48300 27636
rect 48356 27580 48366 27636
rect 14700 27468 15596 27524
rect 15652 27468 15662 27524
rect 20486 27468 20524 27524
rect 20580 27468 20590 27524
rect 28354 27468 28364 27524
rect 28420 27468 29820 27524
rect 29876 27468 30492 27524
rect 30548 27468 30558 27524
rect 33786 27468 33796 27524
rect 33852 27468 35028 27524
rect 35634 27468 35644 27524
rect 35700 27468 47964 27524
rect 48020 27468 48030 27524
rect 9762 27356 9772 27412
rect 9828 27356 10220 27412
rect 10276 27356 10286 27412
rect 12114 27356 12124 27412
rect 12180 27356 13020 27412
rect 13076 27356 13086 27412
rect 14364 27356 14980 27412
rect 15036 27356 15046 27412
rect 34514 27356 34524 27412
rect 34580 27356 34590 27412
rect 2818 27244 2828 27300
rect 2884 27244 6244 27300
rect 6300 27244 6310 27300
rect 13626 27244 13636 27300
rect 13692 27244 14420 27300
rect 20290 27244 20300 27300
rect 20356 27244 20972 27300
rect 21028 27244 21038 27300
rect 27794 27244 27804 27300
rect 27860 27244 29932 27300
rect 29988 27244 29998 27300
rect 7634 27132 7644 27188
rect 7700 27132 9996 27188
rect 10052 27132 10062 27188
rect 10322 27132 10332 27188
rect 10388 27132 11116 27188
rect 11172 27132 11182 27188
rect 11554 27132 11564 27188
rect 11620 27132 11630 27188
rect 14364 27132 14420 27244
rect 14476 27132 14486 27188
rect 18498 27132 18508 27188
rect 18564 27132 18956 27188
rect 19012 27132 19022 27188
rect 19180 27132 19740 27188
rect 19796 27132 19806 27188
rect 21690 27132 21700 27188
rect 21756 27132 23100 27188
rect 23156 27132 24108 27188
rect 24164 27132 24174 27188
rect 24882 27132 24892 27188
rect 24948 27132 25676 27188
rect 25732 27132 29708 27188
rect 29764 27132 29774 27188
rect 32722 27132 32732 27188
rect 32788 27132 34188 27188
rect 34244 27132 34254 27188
rect 11564 27076 11620 27132
rect 19180 27076 19236 27132
rect 3042 27020 3052 27076
rect 3108 27020 4508 27076
rect 4564 27020 4574 27076
rect 4834 27020 4844 27076
rect 4900 27020 5628 27076
rect 5684 27020 5694 27076
rect 6748 27020 7080 27076
rect 7136 27020 8540 27076
rect 8596 27020 8606 27076
rect 9538 27020 9548 27076
rect 9604 27020 12460 27076
rect 12516 27020 12526 27076
rect 13234 27020 13244 27076
rect 13300 27020 13468 27076
rect 13524 27020 13534 27076
rect 13850 27020 13860 27076
rect 13972 27020 13982 27076
rect 14130 27020 14140 27076
rect 14196 27020 14234 27076
rect 14774 27020 14812 27076
rect 14868 27020 14878 27076
rect 17602 27020 17612 27076
rect 17668 27020 19236 27076
rect 19394 27020 19404 27076
rect 19460 27020 20300 27076
rect 20356 27020 22260 27076
rect 22316 27020 22326 27076
rect 22866 27020 22876 27076
rect 22932 27020 23660 27076
rect 23716 27020 23726 27076
rect 25750 27020 25788 27076
rect 25844 27020 27804 27076
rect 27860 27020 27870 27076
rect 29250 27020 29260 27076
rect 29316 27020 30380 27076
rect 30436 27020 30446 27076
rect 31602 27020 31612 27076
rect 31668 27020 33796 27076
rect 33852 27020 33862 27076
rect 4844 26964 4900 27020
rect 3826 26908 3836 26964
rect 3892 26908 4900 26964
rect 6748 26852 6804 27020
rect 7980 26852 8036 27020
rect 18508 26964 18564 27020
rect 8726 26908 8764 26964
rect 8820 26908 8830 26964
rect 10210 26908 10220 26964
rect 10276 26908 11340 26964
rect 11396 26908 11676 26964
rect 11732 26908 11742 26964
rect 13010 26908 13020 26964
rect 13076 26908 14084 26964
rect 14242 26908 14252 26964
rect 14308 26908 15372 26964
rect 15428 26908 15438 26964
rect 18498 26908 18508 26964
rect 18564 26908 18574 26964
rect 18834 26908 18844 26964
rect 18900 26908 21308 26964
rect 21364 26908 21980 26964
rect 22036 26908 22540 26964
rect 22596 26908 22606 26964
rect 23202 26908 23212 26964
rect 23268 26908 24892 26964
rect 24948 26908 24958 26964
rect 5842 26796 5852 26852
rect 5908 26796 6804 26852
rect 7858 26796 7868 26852
rect 7924 26796 8036 26852
rect 14028 26852 14084 26908
rect 25788 26852 25844 27020
rect 34524 26964 34580 27356
rect 34972 27300 35028 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 48300 27412 48356 27580
rect 49200 27412 50000 27440
rect 45602 27356 45612 27412
rect 45668 27356 46264 27412
rect 46320 27356 46956 27412
rect 47012 27356 47022 27412
rect 48300 27356 50000 27412
rect 49200 27328 50000 27356
rect 34972 27244 35196 27300
rect 35252 27244 35262 27300
rect 35746 27244 35756 27300
rect 35812 27244 38892 27300
rect 38948 27244 39340 27300
rect 39396 27244 39406 27300
rect 38322 27132 38332 27188
rect 38444 27132 38780 27188
rect 38836 27132 39228 27188
rect 39284 27132 39294 27188
rect 35018 27020 35028 27076
rect 35084 27020 35756 27076
rect 35812 27020 35822 27076
rect 37874 27020 37884 27076
rect 37940 27020 38556 27076
rect 38612 27020 40348 27076
rect 40404 27020 40414 27076
rect 46610 27020 46620 27076
rect 46676 27020 47292 27076
rect 47348 27020 47358 27076
rect 32946 26908 32956 26964
rect 33012 26908 35196 26964
rect 35252 26908 35262 26964
rect 35522 26908 35532 26964
rect 35588 26908 43148 26964
rect 43204 26908 44380 26964
rect 44436 26908 44446 26964
rect 14028 26796 14812 26852
rect 14868 26796 14878 26852
rect 18722 26796 18732 26852
rect 18788 26796 19964 26852
rect 20020 26796 21196 26852
rect 21252 26796 21262 26852
rect 25340 26796 25844 26852
rect 29026 26796 29036 26852
rect 29092 26796 30156 26852
rect 30212 26796 30222 26852
rect 31826 26796 31836 26852
rect 31892 26796 37884 26852
rect 37940 26796 37950 26852
rect 39554 26796 39564 26852
rect 39620 26796 40964 26852
rect 41020 26796 41030 26852
rect 43810 26796 43820 26852
rect 43876 26796 44940 26852
rect 44996 26796 45006 26852
rect 47058 26796 47068 26852
rect 47124 26796 47292 26852
rect 47348 26796 47358 26852
rect 10994 26684 11004 26740
rect 11060 26684 11788 26740
rect 11844 26684 14140 26740
rect 14196 26684 14812 26740
rect 14868 26684 14878 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 25340 26628 25396 26796
rect 34038 26684 34076 26740
rect 34132 26684 34142 26740
rect 34514 26684 34524 26740
rect 34636 26684 35532 26740
rect 35588 26684 35598 26740
rect 36754 26684 36764 26740
rect 36820 26684 37660 26740
rect 37716 26684 37726 26740
rect 39218 26684 39228 26740
rect 39284 26684 40068 26740
rect 40124 26684 40134 26740
rect 42578 26684 42588 26740
rect 42644 26684 47404 26740
rect 47460 26684 47470 26740
rect 11666 26572 11676 26628
rect 11732 26572 12348 26628
rect 12404 26572 12414 26628
rect 18386 26572 18396 26628
rect 18452 26572 18956 26628
rect 19012 26572 19022 26628
rect 24658 26572 24668 26628
rect 24724 26572 25340 26628
rect 25396 26572 25406 26628
rect 29138 26572 29148 26628
rect 29204 26572 29484 26628
rect 29540 26572 29550 26628
rect 31042 26572 31052 26628
rect 31108 26572 31668 26628
rect 31724 26572 31734 26628
rect 32106 26572 32116 26628
rect 32228 26572 32238 26628
rect 32722 26572 32732 26628
rect 32788 26572 33180 26628
rect 33236 26572 47292 26628
rect 47348 26572 47358 26628
rect 7522 26460 7532 26516
rect 7588 26460 8092 26516
rect 8148 26460 8158 26516
rect 8530 26460 8540 26516
rect 8596 26460 8652 26516
rect 8708 26460 8718 26516
rect 8866 26460 8876 26516
rect 8932 26460 33516 26516
rect 33572 26460 33582 26516
rect 33730 26460 33740 26516
rect 33796 26460 35644 26516
rect 35700 26460 35710 26516
rect 36082 26460 36092 26516
rect 36148 26460 36158 26516
rect 37202 26460 37212 26516
rect 37268 26460 37828 26516
rect 19730 26348 19740 26404
rect 19796 26348 20412 26404
rect 20468 26348 20478 26404
rect 23482 26348 23492 26404
rect 23548 26348 25564 26404
rect 25620 26348 25630 26404
rect 26562 26348 26572 26404
rect 26628 26348 29988 26404
rect 30044 26348 30054 26404
rect 5170 26236 5180 26292
rect 5236 26236 8092 26292
rect 8148 26236 9436 26292
rect 9492 26236 9502 26292
rect 11330 26236 11340 26292
rect 11396 26236 12460 26292
rect 12516 26236 12840 26292
rect 12896 26236 12906 26292
rect 16930 26236 16940 26292
rect 16996 26236 17948 26292
rect 18004 26236 18014 26292
rect 25218 26236 25228 26292
rect 25284 26236 26460 26292
rect 26516 26236 26526 26292
rect 26898 26236 26908 26292
rect 26964 26236 28028 26292
rect 28084 26236 28094 26292
rect 29474 26236 29484 26292
rect 29540 26236 29820 26292
rect 29876 26236 29886 26292
rect 33002 26236 33012 26292
rect 33124 26236 33134 26292
rect 6524 26180 6580 26236
rect 28028 26180 28084 26236
rect 36092 26180 36148 26460
rect 1698 26124 1708 26180
rect 1764 26124 2548 26180
rect 2604 26124 2614 26180
rect 6514 26124 6524 26180
rect 6580 26124 6590 26180
rect 12114 26124 12124 26180
rect 12180 26124 13244 26180
rect 13300 26124 13310 26180
rect 15474 26124 15484 26180
rect 15540 26124 17556 26180
rect 17612 26124 17622 26180
rect 24546 26124 24556 26180
rect 24612 26124 24622 26180
rect 28028 26124 30492 26180
rect 30548 26124 30558 26180
rect 36092 26124 36988 26180
rect 37044 26124 37054 26180
rect 24556 26068 24612 26124
rect 37772 26068 37828 26460
rect 38882 26348 38892 26404
rect 38948 26348 39844 26404
rect 39900 26348 39910 26404
rect 45154 26348 45164 26404
rect 45220 26348 46396 26404
rect 46452 26348 46462 26404
rect 38770 26236 38780 26292
rect 38836 26236 39116 26292
rect 39172 26236 40348 26292
rect 40404 26236 40414 26292
rect 40674 26236 40684 26292
rect 40740 26236 42476 26292
rect 42532 26236 42542 26292
rect 43474 26236 43484 26292
rect 43540 26236 45612 26292
rect 45668 26236 45678 26292
rect 47394 26236 47404 26292
rect 47460 26236 48412 26292
rect 48468 26236 48478 26292
rect 39498 26124 39508 26180
rect 39564 26124 41244 26180
rect 41300 26124 41310 26180
rect 43652 26124 45500 26180
rect 45556 26124 45566 26180
rect 1922 26012 1932 26068
rect 1988 26012 15148 26068
rect 15362 26012 15372 26068
rect 15428 26012 16212 26068
rect 16268 26012 16278 26068
rect 24098 26012 24108 26068
rect 24164 26012 24612 26068
rect 25106 26012 25116 26068
rect 25172 26012 26796 26068
rect 26852 26012 30716 26068
rect 30772 26012 31836 26068
rect 31892 26012 31902 26068
rect 37762 26012 37772 26068
rect 37828 26012 37838 26068
rect 15092 25956 15148 26012
rect 15092 25900 16604 25956
rect 16660 25900 16670 25956
rect 26338 25900 26348 25956
rect 26404 25900 28700 25956
rect 28756 25900 30940 25956
rect 30996 25900 31006 25956
rect 33170 25900 33180 25956
rect 33236 25900 33246 25956
rect 33506 25900 33516 25956
rect 33572 25900 34748 25956
rect 34804 25900 34814 25956
rect 39554 25900 39564 25956
rect 39620 25900 40460 25956
rect 40516 25900 40526 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 33180 25844 33236 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 43652 25844 43708 26124
rect 44594 26012 44604 26068
rect 44660 26012 47124 26068
rect 47180 26012 47190 26068
rect 46162 25900 46172 25956
rect 46228 25900 46620 25956
rect 46676 25900 46686 25956
rect 13552 25788 13562 25844
rect 13618 25788 13916 25844
rect 13972 25788 13982 25844
rect 15092 25732 15148 25844
rect 15204 25788 15214 25844
rect 18722 25788 18732 25844
rect 18788 25788 19068 25844
rect 19124 25788 19134 25844
rect 30482 25788 30492 25844
rect 30548 25788 30828 25844
rect 30884 25788 33236 25844
rect 41346 25788 41356 25844
rect 41412 25788 41692 25844
rect 41748 25788 43708 25844
rect 2650 25676 2660 25732
rect 2716 25676 5964 25732
rect 6020 25676 6636 25732
rect 6692 25676 6702 25732
rect 7522 25676 7532 25732
rect 7588 25676 8540 25732
rect 8596 25676 8606 25732
rect 12002 25676 12012 25732
rect 12068 25676 13132 25732
rect 13188 25676 15148 25732
rect 18396 25676 18620 25732
rect 18676 25676 18686 25732
rect 28802 25676 28812 25732
rect 28868 25676 38668 25732
rect 43250 25676 43260 25732
rect 43316 25676 44044 25732
rect 44100 25676 44110 25732
rect 45210 25676 45220 25732
rect 45276 25676 45724 25732
rect 45780 25676 45790 25732
rect 18396 25620 18452 25676
rect 6962 25564 6972 25620
rect 7028 25564 8428 25620
rect 8484 25564 8494 25620
rect 9874 25564 9884 25620
rect 9940 25564 9950 25620
rect 10098 25564 10108 25620
rect 10164 25564 10174 25620
rect 12226 25564 12236 25620
rect 12292 25564 13804 25620
rect 13860 25564 13870 25620
rect 18386 25564 18396 25620
rect 18452 25564 18462 25620
rect 31042 25564 31052 25620
rect 31108 25564 34076 25620
rect 34132 25564 34142 25620
rect 9884 25508 9940 25564
rect 6066 25452 6076 25508
rect 6132 25452 7084 25508
rect 7140 25452 7150 25508
rect 9090 25452 9100 25508
rect 9156 25452 9940 25508
rect 10108 25508 10164 25564
rect 10108 25452 10332 25508
rect 10388 25452 10398 25508
rect 12674 25452 12684 25508
rect 12740 25452 13580 25508
rect 13636 25452 14308 25508
rect 14364 25452 14924 25508
rect 14980 25452 14990 25508
rect 15474 25452 15484 25508
rect 15540 25452 15708 25508
rect 15764 25452 15774 25508
rect 18498 25452 18508 25508
rect 18564 25452 18956 25508
rect 19012 25452 19022 25508
rect 21186 25452 21196 25508
rect 21252 25452 23884 25508
rect 23940 25452 23950 25508
rect 28354 25452 28364 25508
rect 28420 25452 29260 25508
rect 29316 25452 29708 25508
rect 29764 25452 29774 25508
rect 29978 25452 29988 25508
rect 30044 25452 30604 25508
rect 30660 25452 31052 25508
rect 31108 25452 31118 25508
rect 34850 25452 34860 25508
rect 34916 25452 35644 25508
rect 35700 25452 35710 25508
rect 38612 25396 38668 25676
rect 44930 25564 44940 25620
rect 44996 25564 46788 25620
rect 46844 25564 46854 25620
rect 46050 25452 46060 25508
rect 46116 25452 46396 25508
rect 46452 25452 46462 25508
rect 2146 25340 2156 25396
rect 2212 25340 3164 25396
rect 3220 25340 6300 25396
rect 6356 25340 7756 25396
rect 7812 25340 7822 25396
rect 8418 25340 8428 25396
rect 8484 25340 9324 25396
rect 9380 25340 9390 25396
rect 10882 25340 10892 25396
rect 10948 25340 14476 25396
rect 14532 25340 15036 25396
rect 15092 25340 15102 25396
rect 19282 25340 19292 25396
rect 19348 25340 20804 25396
rect 20860 25340 21532 25396
rect 21588 25340 22428 25396
rect 22484 25340 22494 25396
rect 30454 25340 30492 25396
rect 30548 25340 30558 25396
rect 31154 25340 31164 25396
rect 31220 25340 32172 25396
rect 32228 25340 32238 25396
rect 38612 25340 38836 25396
rect 47170 25340 47180 25396
rect 47236 25340 48188 25396
rect 48244 25340 48254 25396
rect 38780 25284 38836 25340
rect 18 25228 28 25284
rect 84 25228 24836 25284
rect 24892 25228 25116 25284
rect 25172 25228 25182 25284
rect 30156 25228 31052 25284
rect 31108 25228 31118 25284
rect 31322 25228 31332 25284
rect 31388 25228 33944 25284
rect 34000 25228 34010 25284
rect 37202 25228 37212 25284
rect 37268 25228 37548 25284
rect 37604 25228 37614 25284
rect 38770 25228 38780 25284
rect 38836 25228 38846 25284
rect 30156 25172 30212 25228
rect 3378 25116 3388 25172
rect 3444 25116 4844 25172
rect 4900 25116 4910 25172
rect 7970 25116 7980 25172
rect 8036 25116 8540 25172
rect 8596 25116 9212 25172
rect 9268 25116 9278 25172
rect 10210 25116 10220 25172
rect 10276 25116 10780 25172
rect 10836 25116 11676 25172
rect 11732 25116 14028 25172
rect 14084 25116 14094 25172
rect 25778 25116 25788 25172
rect 25844 25116 26236 25172
rect 26292 25116 27804 25172
rect 27860 25116 28252 25172
rect 28308 25116 28318 25172
rect 30146 25116 30156 25172
rect 30212 25116 30222 25172
rect 33030 25116 33068 25172
rect 33124 25116 33134 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 33068 25060 33124 25116
rect 13122 25004 13132 25060
rect 13188 25004 16716 25060
rect 16772 25004 16782 25060
rect 25666 25004 25676 25060
rect 25732 25004 27916 25060
rect 27972 25004 27982 25060
rect 33068 25004 35644 25060
rect 35700 25004 35710 25060
rect 35868 25004 46620 25060
rect 46676 25004 46686 25060
rect 0 24948 800 24976
rect 0 24892 1708 24948
rect 1764 24892 1774 24948
rect 11106 24892 11116 24948
rect 11172 24892 11788 24948
rect 11844 24892 12684 24948
rect 12740 24892 12750 24948
rect 16482 24892 16492 24948
rect 16548 24892 17500 24948
rect 17556 24892 17566 24948
rect 22306 24892 22316 24948
rect 22372 24892 22652 24948
rect 22708 24892 22718 24948
rect 23762 24892 23772 24948
rect 23828 24892 25788 24948
rect 25844 24892 25854 24948
rect 26506 24892 26516 24948
rect 26572 24892 27132 24948
rect 27188 24892 27198 24948
rect 30482 24892 30492 24948
rect 30548 24892 32060 24948
rect 32116 24892 32126 24948
rect 0 24864 800 24892
rect 3154 24780 3164 24836
rect 3220 24780 5516 24836
rect 5572 24780 5582 24836
rect 8082 24780 8092 24836
rect 8148 24780 8540 24836
rect 8596 24780 8606 24836
rect 12086 24780 12124 24836
rect 12180 24780 12190 24836
rect 16258 24780 16268 24836
rect 16324 24780 22204 24836
rect 22260 24780 22270 24836
rect 25890 24780 25900 24836
rect 25956 24780 26740 24836
rect 26898 24780 26908 24836
rect 26964 24780 29036 24836
rect 29092 24780 29102 24836
rect 30258 24780 30268 24836
rect 30324 24780 31948 24836
rect 32004 24780 32014 24836
rect 26684 24724 26740 24780
rect 2482 24668 2492 24724
rect 2548 24668 3556 24724
rect 3612 24668 3622 24724
rect 6178 24668 6188 24724
rect 6244 24668 6972 24724
rect 7028 24668 7038 24724
rect 7746 24668 7756 24724
rect 7812 24668 8316 24724
rect 8372 24668 8382 24724
rect 8698 24668 8708 24724
rect 8764 24668 8988 24724
rect 9044 24668 9054 24724
rect 11554 24668 11564 24724
rect 11620 24668 12236 24724
rect 12292 24668 12302 24724
rect 22082 24668 22092 24724
rect 22148 24668 22316 24724
rect 22372 24668 22382 24724
rect 24714 24668 24724 24724
rect 24780 24668 26516 24724
rect 26572 24668 26582 24724
rect 26684 24668 27020 24724
rect 27076 24668 27086 24724
rect 27458 24668 27468 24724
rect 27524 24668 28476 24724
rect 28532 24668 29484 24724
rect 29540 24668 29550 24724
rect 31714 24668 31724 24724
rect 31780 24668 32396 24724
rect 32452 24668 33180 24724
rect 33236 24668 33246 24724
rect 4292 24556 4302 24612
rect 4358 24556 7644 24612
rect 7700 24556 9436 24612
rect 9492 24556 9502 24612
rect 24434 24556 24444 24612
rect 24500 24556 25284 24612
rect 25340 24556 27580 24612
rect 27636 24556 29148 24612
rect 29204 24556 29214 24612
rect 30454 24556 30492 24612
rect 30548 24556 30558 24612
rect 35868 24500 35924 25004
rect 38658 24892 38668 24948
rect 38724 24892 38892 24948
rect 38948 24892 38958 24948
rect 42242 24892 42252 24948
rect 42308 24892 43260 24948
rect 43316 24892 43326 24948
rect 42466 24780 42476 24836
rect 42532 24780 43372 24836
rect 43428 24780 43438 24836
rect 44818 24780 44828 24836
rect 44884 24780 47740 24836
rect 47796 24780 48076 24836
rect 48132 24780 48142 24836
rect 37650 24668 37660 24724
rect 37716 24668 38332 24724
rect 38388 24668 38398 24724
rect 40338 24668 40348 24724
rect 40404 24668 40908 24724
rect 40964 24668 40974 24724
rect 42578 24668 42588 24724
rect 42644 24668 43876 24724
rect 43932 24668 45388 24724
rect 45444 24668 45454 24724
rect 41346 24556 41356 24612
rect 41412 24556 42140 24612
rect 42196 24556 42206 24612
rect 45154 24556 45164 24612
rect 45220 24556 45836 24612
rect 45892 24556 45902 24612
rect 2818 24444 2828 24500
rect 2884 24444 3948 24500
rect 4004 24444 4014 24500
rect 16370 24444 16380 24500
rect 16436 24444 17052 24500
rect 17108 24444 17118 24500
rect 24098 24444 24108 24500
rect 24164 24444 24892 24500
rect 24948 24444 24958 24500
rect 26114 24444 26124 24500
rect 26180 24444 35924 24500
rect 41234 24444 41244 24500
rect 41300 24444 41580 24500
rect 41636 24444 42980 24500
rect 43036 24444 43046 24500
rect 43138 24444 43148 24500
rect 43204 24444 43260 24500
rect 43316 24444 43326 24500
rect 5506 24332 5516 24388
rect 5572 24332 6860 24388
rect 6916 24332 6926 24388
rect 16594 24332 16604 24388
rect 16660 24332 20188 24388
rect 20244 24332 20254 24388
rect 24994 24332 25004 24388
rect 25060 24332 28868 24388
rect 28924 24332 28934 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 19394 24220 19404 24276
rect 19460 24220 19470 24276
rect 24210 24220 24220 24276
rect 24276 24220 24286 24276
rect 27682 24220 27692 24276
rect 27748 24220 30156 24276
rect 30212 24220 30222 24276
rect 30594 24220 30604 24276
rect 30660 24220 31724 24276
rect 31780 24220 33068 24276
rect 33124 24220 33134 24276
rect 19404 24052 19460 24220
rect 24220 24164 24276 24220
rect 23650 24108 23660 24164
rect 23716 24108 26120 24164
rect 26176 24108 26684 24164
rect 26740 24108 26750 24164
rect 30370 24108 30380 24164
rect 30436 24108 30940 24164
rect 30996 24108 31006 24164
rect 38098 24108 38108 24164
rect 38164 24108 38220 24164
rect 38276 24108 39340 24164
rect 39396 24108 39406 24164
rect 4386 23996 4396 24052
rect 4452 23996 5628 24052
rect 5684 23996 5694 24052
rect 19404 23996 20636 24052
rect 20692 23996 20702 24052
rect 36082 23996 36092 24052
rect 36148 23996 36988 24052
rect 37044 23996 37054 24052
rect 42074 23996 42084 24052
rect 42140 23996 42532 24052
rect 42588 23996 42598 24052
rect 4162 23884 4172 23940
rect 4228 23884 6636 23940
rect 6692 23884 6702 23940
rect 6962 23884 6972 23940
rect 7028 23884 7756 23940
rect 7812 23884 7822 23940
rect 8024 23884 8034 23940
rect 8090 23884 9212 23940
rect 9268 23884 9278 23940
rect 12870 23884 12908 23940
rect 12964 23884 12974 23940
rect 14130 23884 14140 23940
rect 14196 23884 14364 23940
rect 14420 23884 15148 23940
rect 15204 23884 15214 23940
rect 7756 23828 7812 23884
rect 3826 23772 3836 23828
rect 3892 23772 4564 23828
rect 4620 23772 5292 23828
rect 5348 23772 5358 23828
rect 7756 23772 8876 23828
rect 8932 23772 8942 23828
rect 18834 23660 18844 23716
rect 18900 23660 19180 23716
rect 19236 23660 19246 23716
rect 19404 23604 19460 23996
rect 20178 23884 20188 23940
rect 20244 23884 21532 23940
rect 21588 23884 21598 23940
rect 21914 23884 21924 23940
rect 21980 23884 22876 23940
rect 22932 23884 22942 23940
rect 26786 23884 26796 23940
rect 21532 23716 21588 23884
rect 26852 23828 26908 23940
rect 29362 23884 29372 23940
rect 29428 23884 31836 23940
rect 31892 23884 31902 23940
rect 37090 23884 37100 23940
rect 37156 23884 40124 23940
rect 40180 23884 40908 23940
rect 40964 23884 40974 23940
rect 43652 23884 45500 23940
rect 45556 23884 45566 23940
rect 26852 23772 27692 23828
rect 27748 23772 28700 23828
rect 28756 23772 29260 23828
rect 29316 23772 29326 23828
rect 31042 23772 31052 23828
rect 31108 23772 32284 23828
rect 32340 23772 32350 23828
rect 36866 23772 36876 23828
rect 36932 23772 37436 23828
rect 37492 23772 40348 23828
rect 40404 23772 40684 23828
rect 40740 23772 40750 23828
rect 21532 23660 26908 23716
rect 28354 23660 28364 23716
rect 28420 23660 30000 23716
rect 30056 23660 30828 23716
rect 30884 23660 30894 23716
rect 31388 23660 37884 23716
rect 37940 23660 37950 23716
rect 42466 23660 42476 23716
rect 42532 23660 43036 23716
rect 43092 23660 43102 23716
rect 26852 23604 26908 23660
rect 31388 23604 31444 23660
rect 2590 23548 2600 23604
rect 2656 23548 4284 23604
rect 4340 23548 4350 23604
rect 11666 23548 11676 23604
rect 11732 23548 13468 23604
rect 13524 23548 13534 23604
rect 17938 23548 17948 23604
rect 18004 23548 18732 23604
rect 18788 23548 18798 23604
rect 19282 23548 19292 23604
rect 19348 23548 19460 23604
rect 22866 23548 22876 23604
rect 22932 23548 23548 23604
rect 23604 23548 23614 23604
rect 26852 23548 31444 23604
rect 31602 23548 31612 23604
rect 31668 23548 31948 23604
rect 32004 23548 33012 23604
rect 33068 23548 33404 23604
rect 33460 23548 33470 23604
rect 34290 23548 34300 23604
rect 34356 23548 35084 23604
rect 35140 23548 38332 23604
rect 38388 23548 38780 23604
rect 38836 23548 40292 23604
rect 40348 23548 42084 23604
rect 42140 23548 42150 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 43652 23492 43708 23884
rect 2034 23436 2044 23492
rect 2100 23436 3052 23492
rect 3108 23436 5740 23492
rect 5796 23436 5806 23492
rect 24770 23436 24780 23492
rect 24836 23436 28252 23492
rect 28308 23436 28318 23492
rect 32834 23436 32844 23492
rect 32900 23436 33516 23492
rect 33572 23436 33582 23492
rect 34626 23436 34636 23492
rect 34692 23436 37772 23492
rect 37828 23436 37838 23492
rect 40674 23436 40684 23492
rect 40740 23436 41356 23492
rect 41412 23436 45612 23492
rect 45668 23436 45678 23492
rect 3154 23324 3164 23380
rect 3220 23324 3230 23380
rect 5170 23324 5180 23380
rect 5236 23324 6076 23380
rect 6132 23324 7196 23380
rect 7252 23324 7532 23380
rect 7588 23324 7598 23380
rect 12562 23324 12572 23380
rect 12628 23324 13020 23380
rect 13076 23324 13916 23380
rect 13972 23324 13982 23380
rect 18246 23324 18284 23380
rect 18340 23324 18350 23380
rect 30930 23324 30940 23380
rect 30996 23324 31612 23380
rect 31668 23324 31678 23380
rect 32022 23324 32060 23380
rect 32116 23324 32126 23380
rect 34962 23324 34972 23380
rect 35028 23324 35756 23380
rect 35812 23324 35822 23380
rect 45266 23324 45276 23380
rect 45332 23324 45724 23380
rect 45780 23324 45790 23380
rect 3164 22820 3220 23324
rect 5618 23212 5628 23268
rect 5684 23212 5852 23268
rect 5908 23212 6524 23268
rect 6580 23212 7308 23268
rect 7364 23212 7374 23268
rect 23874 23212 23884 23268
rect 23940 23212 25452 23268
rect 25508 23212 25788 23268
rect 25844 23212 25854 23268
rect 27010 23212 27020 23268
rect 27076 23212 27692 23268
rect 27748 23212 27758 23268
rect 29362 23212 29372 23268
rect 29428 23212 32172 23268
rect 32228 23212 32238 23268
rect 32386 23212 32396 23268
rect 32452 23212 32732 23268
rect 32788 23212 33180 23268
rect 33236 23212 33246 23268
rect 34524 23212 42364 23268
rect 42420 23212 42430 23268
rect 45042 23212 45052 23268
rect 45108 23212 46284 23268
rect 46340 23212 47180 23268
rect 47236 23212 48020 23268
rect 48076 23212 48086 23268
rect 3882 23100 3892 23156
rect 3948 23100 4844 23156
rect 4900 23100 4910 23156
rect 5954 23100 5964 23156
rect 6020 23100 7756 23156
rect 7812 23100 7822 23156
rect 8082 23100 8092 23156
rect 8148 23100 8158 23156
rect 9762 23100 9772 23156
rect 9828 23100 10220 23156
rect 10276 23100 10286 23156
rect 18274 23100 18284 23156
rect 18340 23100 18620 23156
rect 18676 23100 18686 23156
rect 20402 23100 20412 23156
rect 20468 23100 21084 23156
rect 21140 23100 21150 23156
rect 21522 23100 21532 23156
rect 21588 23100 23626 23156
rect 23682 23100 23692 23156
rect 23762 23100 23772 23156
rect 23828 23100 25004 23156
rect 25060 23100 25070 23156
rect 25554 23100 25564 23156
rect 25620 23100 26124 23156
rect 26180 23100 27960 23156
rect 28016 23100 28026 23156
rect 28242 23100 28252 23156
rect 28308 23100 29932 23156
rect 29988 23100 29998 23156
rect 32246 23100 32284 23156
rect 32340 23100 32350 23156
rect 4844 23044 4900 23100
rect 8092 23044 8148 23100
rect 4844 22988 6860 23044
rect 6916 22988 8148 23044
rect 17490 22988 17500 23044
rect 17556 22988 32564 23044
rect 32620 22988 34300 23044
rect 34356 22988 34366 23044
rect 3332 22876 4788 22932
rect 4844 22876 5516 22932
rect 5572 22876 5582 22932
rect 7186 22876 7196 22932
rect 7252 22876 8204 22932
rect 8260 22876 8270 22932
rect 13804 22876 14196 22932
rect 14252 22876 20076 22932
rect 20132 22876 22540 22932
rect 22596 22876 22606 22932
rect 26562 22876 26572 22932
rect 26628 22876 27244 22932
rect 27300 22876 27310 22932
rect 28690 22876 28700 22932
rect 28756 22876 33964 22932
rect 34020 22876 34030 22932
rect 3332 22820 3388 22876
rect 3154 22764 3164 22820
rect 3220 22764 3230 22820
rect 3322 22764 3332 22820
rect 3388 22764 3398 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 11218 22652 11228 22708
rect 11284 22652 11676 22708
rect 11732 22652 11742 22708
rect 13738 22652 13748 22708
rect 13804 22652 13860 22876
rect 34524 22820 34580 23212
rect 38658 23100 38668 23156
rect 38724 23100 39676 23156
rect 39732 23100 39742 23156
rect 44930 23100 44940 23156
rect 44996 23100 45836 23156
rect 45892 23100 45902 23156
rect 42578 22988 42588 23044
rect 42644 22988 44828 23044
rect 44884 22988 44894 23044
rect 22194 22764 22204 22820
rect 22260 22764 22270 22820
rect 22754 22764 22764 22820
rect 22820 22764 23548 22820
rect 23604 22764 23614 22820
rect 24882 22764 24892 22820
rect 24948 22764 26796 22820
rect 26852 22764 28588 22820
rect 28644 22764 28654 22820
rect 29922 22764 29932 22820
rect 29988 22764 31052 22820
rect 31108 22764 31118 22820
rect 31276 22764 34580 22820
rect 40562 22764 40572 22820
rect 40628 22764 45220 22820
rect 45276 22764 45286 22820
rect 22204 22596 22260 22764
rect 22642 22652 22652 22708
rect 22708 22652 23212 22708
rect 23268 22652 23278 22708
rect 26226 22652 26236 22708
rect 26292 22652 26908 22708
rect 26964 22652 26974 22708
rect 31276 22596 31332 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 31714 22652 31724 22708
rect 31780 22652 32732 22708
rect 32788 22652 32798 22708
rect 7914 22540 7924 22596
rect 7980 22540 9212 22596
rect 9268 22540 9660 22596
rect 9716 22540 9726 22596
rect 10098 22540 10108 22596
rect 10164 22540 14700 22596
rect 14756 22540 14766 22596
rect 16986 22540 16996 22596
rect 17052 22540 21532 22596
rect 21588 22540 21598 22596
rect 22204 22540 31332 22596
rect 31434 22540 31444 22596
rect 31500 22540 33460 22596
rect 33516 22540 33526 22596
rect 42466 22540 42476 22596
rect 42532 22540 43708 22596
rect 43652 22484 43708 22540
rect 49200 22484 50000 22512
rect 2818 22428 2828 22484
rect 2884 22428 3500 22484
rect 3556 22428 4620 22484
rect 4676 22428 4686 22484
rect 15362 22428 15372 22484
rect 15428 22428 17780 22484
rect 17836 22428 23156 22484
rect 42242 22428 42252 22484
rect 42308 22428 43036 22484
rect 43092 22428 43102 22484
rect 43652 22428 43932 22484
rect 43988 22428 43998 22484
rect 48738 22428 48748 22484
rect 48804 22428 50000 22484
rect 23100 22372 23156 22428
rect 49200 22400 50000 22428
rect 4722 22316 4732 22372
rect 4788 22316 5404 22372
rect 5460 22316 6300 22372
rect 6356 22316 6366 22372
rect 6570 22316 6580 22372
rect 6636 22316 7196 22372
rect 7252 22316 9436 22372
rect 9492 22316 9884 22372
rect 9940 22316 9950 22372
rect 12450 22316 12460 22372
rect 12516 22316 13356 22372
rect 13412 22316 13422 22372
rect 14130 22316 14140 22372
rect 14196 22316 15092 22372
rect 15148 22316 15158 22372
rect 15978 22316 15988 22372
rect 16044 22316 16996 22372
rect 17052 22316 17062 22372
rect 18050 22316 18060 22372
rect 18116 22316 18396 22372
rect 18452 22316 18844 22372
rect 18900 22316 18910 22372
rect 23090 22316 23100 22372
rect 23156 22316 25340 22372
rect 25396 22316 25406 22372
rect 27682 22316 27692 22372
rect 27748 22316 29640 22372
rect 29696 22316 29706 22372
rect 32022 22316 32060 22372
rect 32116 22316 32126 22372
rect 32246 22316 32284 22372
rect 32340 22316 32350 22372
rect 34906 22316 34916 22372
rect 34972 22316 35644 22372
rect 35700 22316 35710 22372
rect 35858 22316 35868 22372
rect 35924 22316 37940 22372
rect 37996 22316 38668 22372
rect 42130 22316 42140 22372
rect 42196 22316 42700 22372
rect 42756 22316 44044 22372
rect 44100 22316 44110 22372
rect 3714 22204 3724 22260
rect 3780 22204 4508 22260
rect 4564 22204 6412 22260
rect 6468 22204 6478 22260
rect 15810 22204 15820 22260
rect 15876 22204 19628 22260
rect 19684 22204 19694 22260
rect 22754 22204 22764 22260
rect 22820 22204 22988 22260
rect 23044 22204 23054 22260
rect 11330 22092 11340 22148
rect 11396 22092 11788 22148
rect 11844 22092 11854 22148
rect 14690 22092 14700 22148
rect 14756 22092 15372 22148
rect 15428 22092 15438 22148
rect 17378 22092 17388 22148
rect 17444 22092 20076 22148
rect 20132 22092 21308 22148
rect 21364 22092 21374 22148
rect 21690 22092 21700 22148
rect 21756 22092 22652 22148
rect 22708 22092 24892 22148
rect 24948 22092 27356 22148
rect 27412 22092 27422 22148
rect 34626 22092 34636 22148
rect 34692 22092 35980 22148
rect 36036 22092 36876 22148
rect 36932 22092 36942 22148
rect 38612 22092 38668 22316
rect 38882 22204 38892 22260
rect 38948 22204 43092 22260
rect 43222 22204 43260 22260
rect 43316 22204 43326 22260
rect 46946 22204 46956 22260
rect 47012 22204 47740 22260
rect 47796 22204 47806 22260
rect 43036 22148 43092 22204
rect 38724 22092 39116 22148
rect 39172 22092 39182 22148
rect 43036 22092 43596 22148
rect 43652 22092 43662 22148
rect 4498 21980 4508 22036
rect 4564 21980 4732 22036
rect 4788 21980 4798 22036
rect 14018 21980 14028 22036
rect 14084 21980 14094 22036
rect 21522 21980 21532 22036
rect 21588 21980 26460 22036
rect 26516 21980 26526 22036
rect 43362 21980 43372 22036
rect 43428 21980 44604 22036
rect 44660 21980 44670 22036
rect 14028 21924 14084 21980
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 4610 21868 4620 21924
rect 4676 21868 5404 21924
rect 5460 21868 5470 21924
rect 5730 21868 5740 21924
rect 5796 21868 6524 21924
rect 6580 21868 6590 21924
rect 13682 21868 13692 21924
rect 13748 21868 15820 21924
rect 15876 21868 15886 21924
rect 17826 21868 17836 21924
rect 17892 21868 18284 21924
rect 18340 21868 19068 21924
rect 19124 21868 19134 21924
rect 23034 21868 23044 21924
rect 23100 21868 23660 21924
rect 23716 21868 24500 21924
rect 24556 21868 25060 21924
rect 25116 21812 25172 21924
rect 39330 21868 39340 21924
rect 39396 21868 40572 21924
rect 40628 21868 40638 21924
rect 41458 21868 41468 21924
rect 41524 21868 42364 21924
rect 42420 21868 42430 21924
rect 2146 21756 2156 21812
rect 2212 21756 3276 21812
rect 3332 21756 3500 21812
rect 3556 21756 4056 21812
rect 4112 21756 4122 21812
rect 10882 21756 10892 21812
rect 10948 21756 14812 21812
rect 14868 21756 14878 21812
rect 16146 21756 16156 21812
rect 16212 21756 17276 21812
rect 17332 21756 18172 21812
rect 18228 21756 20692 21812
rect 20748 21756 21868 21812
rect 21924 21756 21934 21812
rect 25116 21756 27198 21812
rect 27254 21756 27972 21812
rect 28028 21756 29820 21812
rect 29876 21756 29886 21812
rect 33506 21756 33516 21812
rect 33572 21756 34412 21812
rect 34468 21756 36092 21812
rect 36148 21756 36540 21812
rect 36596 21756 36606 21812
rect 38434 21756 38444 21812
rect 38500 21756 39788 21812
rect 39844 21756 39854 21812
rect 40898 21756 40908 21812
rect 40964 21756 41580 21812
rect 41636 21756 44604 21812
rect 44660 21756 44670 21812
rect 3602 21644 3612 21700
rect 3668 21644 4172 21700
rect 4228 21644 4238 21700
rect 8540 21644 9044 21700
rect 14578 21644 14588 21700
rect 14644 21644 15186 21700
rect 15242 21644 15252 21700
rect 17602 21644 17612 21700
rect 17668 21644 17678 21700
rect 17826 21644 17836 21700
rect 17892 21644 22204 21700
rect 24266 21644 24276 21700
rect 24332 21644 25116 21700
rect 25172 21644 26124 21700
rect 26180 21644 26190 21700
rect 33730 21644 33740 21700
rect 33796 21644 37436 21700
rect 37492 21644 37502 21700
rect 38154 21644 38164 21700
rect 38220 21644 40292 21700
rect 40348 21644 40358 21700
rect 46106 21644 46116 21700
rect 46172 21644 47068 21700
rect 47124 21644 47628 21700
rect 47684 21644 47694 21700
rect 2594 21532 2604 21588
rect 2660 21532 5852 21588
rect 5908 21532 5918 21588
rect 8540 21476 8596 21644
rect 8988 21588 9044 21644
rect 17612 21588 17668 21644
rect 22148 21588 22204 21644
rect 8754 21532 8764 21588
rect 8820 21532 8830 21588
rect 8988 21532 16884 21588
rect 16940 21532 16950 21588
rect 17154 21532 17164 21588
rect 17220 21532 17948 21588
rect 18004 21532 18014 21588
rect 21410 21532 21420 21588
rect 21476 21532 21980 21588
rect 22036 21532 22046 21588
rect 22148 21532 24724 21588
rect 24780 21532 25452 21588
rect 25508 21532 25518 21588
rect 26002 21532 26012 21588
rect 26068 21532 29148 21588
rect 29204 21532 29708 21588
rect 29764 21532 29774 21588
rect 32050 21532 32060 21588
rect 32116 21532 33236 21588
rect 33292 21532 38668 21588
rect 39666 21532 39676 21588
rect 39732 21532 40684 21588
rect 40740 21532 40750 21588
rect 43474 21532 43484 21588
rect 43540 21532 44268 21588
rect 44324 21532 44334 21588
rect 46610 21532 46620 21588
rect 46676 21532 47740 21588
rect 47796 21532 48076 21588
rect 48132 21532 48142 21588
rect 1474 21420 1484 21476
rect 1540 21420 8596 21476
rect 8764 21364 8820 21532
rect 38612 21476 38668 21532
rect 16426 21420 16436 21476
rect 16492 21420 26908 21476
rect 29362 21420 29372 21476
rect 29428 21420 34076 21476
rect 34132 21420 37212 21476
rect 37268 21420 37278 21476
rect 38612 21420 40124 21476
rect 40180 21420 40190 21476
rect 26852 21364 26908 21420
rect 8764 21308 10556 21364
rect 10612 21308 10622 21364
rect 15474 21308 15484 21364
rect 15540 21308 15988 21364
rect 16044 21308 17836 21364
rect 17892 21308 17902 21364
rect 18274 21308 18284 21364
rect 18396 21308 18406 21364
rect 26852 21308 32060 21364
rect 32116 21308 32126 21364
rect 37314 21308 37324 21364
rect 37380 21308 38556 21364
rect 38612 21308 38622 21364
rect 44258 21308 44268 21364
rect 44324 21308 45612 21364
rect 45668 21308 47404 21364
rect 47460 21308 47470 21364
rect 26114 21196 26124 21252
rect 26180 21196 26796 21252
rect 26852 21196 26862 21252
rect 36754 21196 36764 21252
rect 36820 21196 39004 21252
rect 39060 21196 39070 21252
rect 39890 21196 39900 21252
rect 39956 21196 48244 21252
rect 48300 21196 48310 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 16706 21084 16716 21140
rect 16772 21084 18900 21140
rect 18956 21084 23436 21140
rect 23492 21084 23502 21140
rect 45602 21084 45612 21140
rect 45668 21084 45836 21140
rect 45892 21084 45902 21140
rect 11218 20972 11228 21028
rect 11284 20972 11564 21028
rect 11620 20972 13580 21028
rect 13636 20972 13646 21028
rect 15138 20972 15148 21028
rect 15204 20972 15540 21028
rect 15596 20972 17668 21028
rect 17724 20972 18116 21028
rect 18172 20972 26796 21028
rect 26852 20972 26862 21028
rect 42242 20972 42252 21028
rect 42308 20972 43932 21028
rect 43988 20972 43998 21028
rect 9314 20860 9324 20916
rect 9380 20860 14364 20916
rect 14420 20860 14430 20916
rect 22418 20860 22428 20916
rect 22484 20860 23100 20916
rect 23156 20860 24892 20916
rect 24948 20860 24958 20916
rect 31714 20860 31724 20916
rect 31780 20860 32396 20916
rect 32452 20860 32462 20916
rect 41010 20860 41020 20916
rect 41076 20860 41524 20916
rect 41580 20860 41590 20916
rect 43810 20860 43820 20916
rect 43876 20860 45500 20916
rect 45556 20860 45566 20916
rect 5170 20748 5180 20804
rect 5236 20748 5516 20804
rect 5572 20748 7644 20804
rect 7700 20748 7710 20804
rect 14242 20748 14252 20804
rect 14308 20748 14756 20804
rect 14812 20748 14822 20804
rect 16594 20748 16604 20804
rect 16660 20748 16670 20804
rect 17154 20748 17164 20804
rect 17220 20748 17612 20804
rect 17668 20748 18732 20804
rect 18788 20748 18798 20804
rect 20178 20748 20188 20804
rect 20244 20748 21420 20804
rect 21476 20748 21486 20804
rect 23314 20748 23324 20804
rect 23380 20748 25676 20804
rect 25732 20748 25742 20804
rect 30930 20748 30940 20804
rect 30996 20748 31276 20804
rect 31332 20748 31342 20804
rect 38882 20748 38892 20804
rect 38948 20748 43372 20804
rect 43428 20748 43438 20804
rect 43820 20748 44716 20804
rect 44772 20748 45276 20804
rect 45332 20748 45342 20804
rect 48290 20748 48300 20804
rect 48356 20748 48748 20804
rect 48804 20748 48814 20804
rect 16604 20692 16660 20748
rect 43820 20692 43876 20748
rect 14914 20636 14924 20692
rect 14980 20636 21868 20692
rect 21924 20636 21934 20692
rect 39778 20636 39788 20692
rect 39844 20636 40124 20692
rect 40180 20636 40796 20692
rect 40852 20636 43820 20692
rect 43876 20636 43886 20692
rect 6598 20524 6636 20580
rect 6692 20524 6702 20580
rect 13962 20524 13972 20580
rect 14028 20524 15036 20580
rect 15092 20524 15102 20580
rect 16482 20524 16492 20580
rect 16548 20524 17500 20580
rect 17556 20524 17566 20580
rect 17770 20524 17780 20580
rect 17836 20524 25564 20580
rect 25620 20524 25630 20580
rect 34122 20524 34132 20580
rect 34188 20524 36540 20580
rect 36596 20524 36606 20580
rect 36764 20524 39340 20580
rect 39396 20524 39900 20580
rect 39956 20524 39966 20580
rect 40226 20524 40236 20580
rect 40292 20524 43932 20580
rect 43988 20524 43998 20580
rect 46386 20524 46396 20580
rect 46452 20524 47292 20580
rect 47348 20524 47358 20580
rect 36764 20468 36820 20524
rect 6236 20412 6246 20468
rect 6302 20412 11676 20468
rect 11732 20412 11742 20468
rect 16034 20412 16044 20468
rect 16100 20412 16604 20468
rect 16660 20412 16670 20468
rect 19058 20412 19068 20468
rect 19124 20412 19134 20468
rect 35074 20412 35084 20468
rect 35140 20412 36820 20468
rect 38098 20412 38108 20468
rect 38164 20412 39004 20468
rect 39060 20412 39070 20468
rect 16258 20300 16268 20356
rect 16324 20300 16716 20356
rect 16772 20300 16782 20356
rect 15026 20188 15036 20244
rect 15092 20188 17780 20244
rect 17836 20188 17846 20244
rect 19068 20132 19124 20412
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 23426 20300 23436 20356
rect 23492 20300 24780 20356
rect 24836 20300 24846 20356
rect 25414 20300 25452 20356
rect 25508 20300 25518 20356
rect 31210 20300 31220 20356
rect 31276 20300 32060 20356
rect 32116 20300 32126 20356
rect 45490 20300 45500 20356
rect 45556 20300 47964 20356
rect 48020 20300 48030 20356
rect 22530 20188 22540 20244
rect 22596 20188 23548 20244
rect 23604 20188 23614 20244
rect 25554 20188 25564 20244
rect 25620 20188 27020 20244
rect 27076 20188 27086 20244
rect 28018 20188 28028 20244
rect 28084 20188 28420 20244
rect 28476 20188 28868 20244
rect 28924 20188 33628 20244
rect 33684 20188 33694 20244
rect 37762 20188 37772 20244
rect 37828 20188 38444 20244
rect 38500 20188 38510 20244
rect 39116 20188 44044 20244
rect 44100 20188 44110 20244
rect 39116 20132 39172 20188
rect 6626 20076 6636 20132
rect 6692 20076 6972 20132
rect 7028 20076 7038 20132
rect 7308 20076 8708 20132
rect 10098 20076 10108 20132
rect 10164 20076 13412 20132
rect 13468 20076 13478 20132
rect 13682 20076 13692 20132
rect 13748 20076 14364 20132
rect 14420 20076 14812 20132
rect 14868 20076 15708 20132
rect 15764 20076 15774 20132
rect 19068 20076 19236 20132
rect 19562 20076 19572 20132
rect 19628 20076 20188 20132
rect 20244 20076 20254 20132
rect 24098 20076 24108 20132
rect 24164 20076 25116 20132
rect 25172 20076 25182 20132
rect 26562 20076 26572 20132
rect 26628 20076 27132 20132
rect 27188 20076 27198 20132
rect 32050 20076 32060 20132
rect 32116 20076 32732 20132
rect 32788 20076 32798 20132
rect 36866 20076 36876 20132
rect 36932 20076 39060 20132
rect 39116 20076 39452 20132
rect 39508 20076 39518 20132
rect 7308 20020 7364 20076
rect 8652 20020 8708 20076
rect 19180 20020 19236 20076
rect 39004 20020 39060 20076
rect 1586 19964 1596 20020
rect 1652 19964 2268 20020
rect 2324 19964 2334 20020
rect 6514 19964 6524 20020
rect 6580 19964 7364 20020
rect 7522 19964 7532 20020
rect 7588 19964 8428 20020
rect 8484 19964 8494 20020
rect 8652 19964 10500 20020
rect 13794 19964 13804 20020
rect 13860 19964 14924 20020
rect 14980 19964 15932 20020
rect 15988 19964 15998 20020
rect 16370 19964 16380 20020
rect 16436 19964 16828 20020
rect 16884 19964 17500 20020
rect 17556 19964 17566 20020
rect 19180 19964 19740 20020
rect 19796 19964 23492 20020
rect 23548 19964 23558 20020
rect 25442 19964 25452 20020
rect 25508 19964 28028 20020
rect 28084 19964 28094 20020
rect 31826 19964 31836 20020
rect 31892 19964 33012 20020
rect 33068 19964 33078 20020
rect 35522 19964 35532 20020
rect 35588 19964 36316 20020
rect 36372 19964 36382 20020
rect 37202 19964 37212 20020
rect 37268 19964 37996 20020
rect 38052 19964 38780 20020
rect 38836 19964 38846 20020
rect 39004 19964 40348 20020
rect 40404 19964 40908 20020
rect 40964 19964 40974 20020
rect 45602 19964 45612 20020
rect 45668 19964 47628 20020
rect 47684 19964 48076 20020
rect 48132 19964 48142 20020
rect 10444 19908 10500 19964
rect 3042 19852 3052 19908
rect 3108 19852 7196 19908
rect 7252 19852 7262 19908
rect 7858 19852 7868 19908
rect 7924 19852 9996 19908
rect 10052 19852 10062 19908
rect 10444 19852 14532 19908
rect 14588 19852 14598 19908
rect 16930 19852 16940 19908
rect 16996 19852 19068 19908
rect 19124 19852 19134 19908
rect 20738 19852 20748 19908
rect 20804 19852 21644 19908
rect 21700 19852 24108 19908
rect 24164 19852 24174 19908
rect 30370 19852 30380 19908
rect 30436 19852 32284 19908
rect 32340 19852 37548 19908
rect 37604 19852 37884 19908
rect 37940 19852 37950 19908
rect 38266 19852 38276 19908
rect 38332 19852 39900 19908
rect 39956 19852 39966 19908
rect 44482 19852 44492 19908
rect 44548 19852 44940 19908
rect 44996 19852 48300 19908
rect 48356 19852 48366 19908
rect 7868 19796 7924 19852
rect 2146 19740 2156 19796
rect 2212 19740 6076 19796
rect 6132 19740 6142 19796
rect 6598 19740 6636 19796
rect 6692 19740 6702 19796
rect 6962 19740 6972 19796
rect 7028 19740 7924 19796
rect 9034 19740 9044 19796
rect 9100 19740 9212 19796
rect 9268 19740 13020 19796
rect 13076 19740 13086 19796
rect 15810 19740 15820 19796
rect 15876 19740 16268 19796
rect 16324 19740 16334 19796
rect 19170 19740 19180 19796
rect 19236 19740 22820 19796
rect 23090 19740 23100 19796
rect 23156 19740 23772 19796
rect 23828 19740 24332 19796
rect 24388 19740 24398 19796
rect 26852 19740 39116 19796
rect 39172 19740 39182 19796
rect 45042 19740 45052 19796
rect 45108 19740 45948 19796
rect 46004 19740 46014 19796
rect 22764 19684 22820 19740
rect 26852 19684 26908 19740
rect 8026 19628 8036 19684
rect 8092 19628 15428 19684
rect 15484 19628 15494 19684
rect 18330 19628 18340 19684
rect 18396 19628 19628 19684
rect 19684 19628 19694 19684
rect 20514 19628 20524 19684
rect 20580 19628 22092 19684
rect 22148 19628 22540 19684
rect 22596 19628 22606 19684
rect 22764 19628 26908 19684
rect 38882 19628 38892 19684
rect 38948 19628 39452 19684
rect 39508 19628 39518 19684
rect 42776 19628 42786 19684
rect 42842 19628 44044 19684
rect 44100 19628 44110 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 14690 19516 14700 19572
rect 14756 19516 15036 19572
rect 15092 19516 15102 19572
rect 19282 19516 19292 19572
rect 19348 19516 20412 19572
rect 20468 19516 20478 19572
rect 22250 19516 22260 19572
rect 22316 19516 23156 19572
rect 23212 19516 23660 19572
rect 23716 19516 24052 19572
rect 24108 19516 24118 19572
rect 30706 19516 30716 19572
rect 30772 19516 31052 19572
rect 31108 19516 31118 19572
rect 6962 19404 6972 19460
rect 7028 19404 7756 19460
rect 7812 19404 7822 19460
rect 8978 19404 8988 19460
rect 9044 19404 10444 19460
rect 10500 19404 10510 19460
rect 15092 19404 15260 19460
rect 15316 19404 16156 19460
rect 16212 19404 16222 19460
rect 16762 19404 16772 19460
rect 16828 19404 19068 19460
rect 19124 19404 19516 19460
rect 19572 19404 20188 19460
rect 20244 19404 20254 19460
rect 38042 19404 38052 19460
rect 38108 19404 40012 19460
rect 40068 19404 40078 19460
rect 14130 19292 14140 19348
rect 14196 19292 15036 19348
rect 15092 19292 15148 19404
rect 17154 19292 17164 19348
rect 17220 19292 19292 19348
rect 19348 19292 20300 19348
rect 20356 19292 20366 19348
rect 22698 19292 22708 19348
rect 22764 19292 25004 19348
rect 25060 19292 25676 19348
rect 25732 19292 27860 19348
rect 27916 19292 27926 19348
rect 31714 19292 31724 19348
rect 31780 19292 32060 19348
rect 32116 19292 32126 19348
rect 32386 19292 32396 19348
rect 32452 19292 33180 19348
rect 33236 19292 33246 19348
rect 4946 19180 4956 19236
rect 5012 19180 6636 19236
rect 6692 19180 6702 19236
rect 14018 19180 14028 19236
rect 14084 19180 15820 19236
rect 15876 19180 15886 19236
rect 17042 19180 17052 19236
rect 17108 19180 18060 19236
rect 18116 19180 18126 19236
rect 20178 19180 20188 19236
rect 20244 19180 21028 19236
rect 21084 19180 21532 19236
rect 21588 19180 21598 19236
rect 23874 19180 23884 19236
rect 23940 19180 24836 19236
rect 24892 19180 25564 19236
rect 25620 19180 26124 19236
rect 26180 19180 27692 19236
rect 27748 19180 27758 19236
rect 28130 19180 28140 19236
rect 28196 19180 29820 19236
rect 29876 19180 29886 19236
rect 43698 19180 43708 19236
rect 43764 19180 44940 19236
rect 44996 19180 45006 19236
rect 45210 19180 45220 19236
rect 45276 19180 45724 19236
rect 45780 19180 45790 19236
rect 46806 19180 46844 19236
rect 46900 19180 46910 19236
rect 46844 19124 46900 19180
rect 11666 19068 11676 19124
rect 11732 19068 14308 19124
rect 14364 19068 14374 19124
rect 15138 19068 15148 19124
rect 15204 19068 15708 19124
rect 15764 19068 17780 19124
rect 17836 19068 17846 19124
rect 17948 19068 25284 19124
rect 25340 19068 25350 19124
rect 37762 19068 37772 19124
rect 37828 19068 38668 19124
rect 38724 19068 38734 19124
rect 39106 19068 39116 19124
rect 39172 19068 46900 19124
rect 17948 19012 18004 19068
rect 4274 18956 4284 19012
rect 4340 18956 5404 19012
rect 5460 18956 6524 19012
rect 6580 18956 7532 19012
rect 7588 18956 7598 19012
rect 9986 18956 9996 19012
rect 10052 18956 15596 19012
rect 15652 18956 15662 19012
rect 15922 18956 15932 19012
rect 15988 18956 18004 19012
rect 19628 18956 22764 19012
rect 22820 18956 22830 19012
rect 24210 18956 24220 19012
rect 24276 18956 24556 19012
rect 24612 18956 24622 19012
rect 24770 18956 24780 19012
rect 24836 18956 24874 19012
rect 27850 18956 27860 19012
rect 27916 18956 28308 19012
rect 28364 18956 45500 19012
rect 45556 18956 45566 19012
rect 19628 18900 19684 18956
rect 15810 18844 15820 18900
rect 15876 18844 16380 18900
rect 16436 18844 16446 18900
rect 16594 18844 16604 18900
rect 16660 18844 19684 18900
rect 23762 18844 23772 18900
rect 23828 18844 25340 18900
rect 25396 18844 25406 18900
rect 44680 18844 44690 18900
rect 44746 18844 45612 18900
rect 45668 18844 45678 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 3994 18732 4004 18788
rect 4060 18732 6412 18788
rect 6468 18732 19068 18788
rect 19124 18732 19180 18788
rect 19236 18732 19246 18788
rect 26422 18732 26460 18788
rect 26516 18732 26526 18788
rect 45938 18732 45948 18788
rect 46004 18732 47292 18788
rect 47348 18732 47358 18788
rect 12226 18620 12236 18676
rect 12292 18620 32340 18676
rect 32396 18620 32406 18676
rect 41794 18620 41804 18676
rect 41860 18620 43708 18676
rect 43764 18620 44268 18676
rect 44324 18620 44334 18676
rect 16930 18508 16940 18564
rect 16996 18508 17612 18564
rect 17668 18508 17678 18564
rect 20402 18508 20412 18564
rect 20468 18508 22428 18564
rect 22484 18508 24556 18564
rect 24612 18508 24622 18564
rect 26012 18508 26796 18564
rect 26852 18508 26862 18564
rect 37426 18508 37436 18564
rect 37492 18508 41300 18564
rect 41356 18508 41366 18564
rect 26012 18452 26068 18508
rect 2258 18396 2268 18452
rect 2324 18396 3052 18452
rect 3108 18396 5292 18452
rect 5348 18396 5358 18452
rect 5506 18396 5516 18452
rect 5572 18396 5740 18452
rect 5796 18396 5806 18452
rect 7914 18396 7924 18452
rect 7980 18396 13132 18452
rect 13188 18396 15148 18452
rect 15250 18396 15260 18452
rect 15316 18396 15932 18452
rect 15988 18396 17276 18452
rect 17332 18396 18732 18452
rect 18788 18396 18798 18452
rect 20066 18396 20076 18452
rect 20132 18396 21196 18452
rect 21252 18396 21262 18452
rect 21410 18396 21420 18452
rect 21476 18396 21868 18452
rect 21924 18396 21934 18452
rect 22082 18396 22092 18452
rect 22148 18396 22988 18452
rect 23044 18396 23660 18452
rect 23716 18396 23726 18452
rect 24434 18396 24444 18452
rect 24500 18396 26068 18452
rect 26226 18396 26236 18452
rect 26292 18396 27020 18452
rect 27076 18396 27086 18452
rect 35298 18396 35308 18452
rect 35364 18396 36316 18452
rect 36372 18396 38220 18452
rect 38276 18396 38286 18452
rect 38546 18396 38556 18452
rect 38612 18396 41020 18452
rect 41076 18396 41086 18452
rect 42690 18396 42700 18452
rect 42756 18396 43484 18452
rect 43540 18396 44828 18452
rect 44884 18396 47796 18452
rect 15092 18340 15148 18396
rect 47740 18340 47796 18396
rect 3826 18284 3836 18340
rect 3892 18284 6300 18340
rect 6356 18284 6366 18340
rect 8530 18284 8540 18340
rect 8596 18284 13916 18340
rect 13972 18284 13982 18340
rect 15092 18284 17388 18340
rect 17444 18284 17454 18340
rect 18834 18284 18844 18340
rect 18900 18284 21980 18340
rect 22036 18284 22316 18340
rect 22372 18284 22382 18340
rect 26618 18284 26628 18340
rect 26684 18284 27468 18340
rect 27524 18284 27534 18340
rect 29250 18284 29260 18340
rect 29316 18284 29820 18340
rect 29876 18284 29886 18340
rect 34850 18284 34860 18340
rect 34916 18284 36092 18340
rect 36148 18284 36158 18340
rect 39106 18284 39116 18340
rect 39172 18284 40236 18340
rect 40292 18284 41692 18340
rect 41748 18284 42364 18340
rect 42420 18284 42430 18340
rect 44706 18284 44716 18340
rect 44772 18284 45836 18340
rect 45892 18284 45902 18340
rect 47730 18284 47740 18340
rect 47796 18284 47806 18340
rect 7466 18172 7476 18228
rect 7532 18172 10052 18228
rect 9996 18116 10052 18172
rect 13916 18116 13972 18284
rect 16034 18172 16044 18228
rect 16100 18172 23212 18228
rect 23268 18172 23278 18228
rect 26226 18172 26236 18228
rect 26292 18172 26460 18228
rect 26516 18172 26526 18228
rect 28018 18172 28028 18228
rect 28084 18172 28588 18228
rect 28644 18172 28654 18228
rect 28802 18172 28812 18228
rect 28868 18172 32228 18228
rect 32284 18172 33404 18228
rect 33460 18172 33470 18228
rect 39638 18172 39676 18228
rect 39732 18172 39742 18228
rect 9986 18060 9996 18116
rect 10052 18060 10062 18116
rect 13916 18060 16492 18116
rect 16548 18060 16558 18116
rect 21858 18060 21868 18116
rect 21924 18060 22652 18116
rect 22708 18060 22718 18116
rect 25218 18060 25228 18116
rect 25284 18060 26796 18116
rect 26852 18060 26862 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 28588 18004 28644 18172
rect 29474 18060 29484 18116
rect 29540 18060 31612 18116
rect 31668 18060 33012 18116
rect 33068 18060 33078 18116
rect 36082 18060 36092 18116
rect 36148 18060 37996 18116
rect 38052 18060 39564 18116
rect 39620 18060 39630 18116
rect 39834 18060 39844 18116
rect 39900 18060 40964 18116
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 40908 18004 40964 18060
rect 10210 17948 10220 18004
rect 10276 17948 12460 18004
rect 12516 17948 12526 18004
rect 22754 17948 22764 18004
rect 22820 17948 24388 18004
rect 24444 17948 24454 18004
rect 26422 17948 26460 18004
rect 26516 17948 26526 18004
rect 26618 17948 26628 18004
rect 26684 17948 26908 18004
rect 26964 17948 26974 18004
rect 28588 17948 29708 18004
rect 29764 17948 29774 18004
rect 32620 17948 33292 18004
rect 33348 17948 33358 18004
rect 39330 17948 39340 18004
rect 39396 17948 40236 18004
rect 40292 17948 40302 18004
rect 40898 17948 40908 18004
rect 40964 17948 43596 18004
rect 43652 17948 43662 18004
rect 32620 17892 32676 17948
rect 8306 17836 8316 17892
rect 8372 17836 8652 17892
rect 8708 17836 9212 17892
rect 9268 17836 12236 17892
rect 12292 17836 12302 17892
rect 14188 17836 14198 17892
rect 14254 17836 26068 17892
rect 26124 17836 26134 17892
rect 29026 17836 29036 17892
rect 29092 17836 30716 17892
rect 30772 17836 32172 17892
rect 32228 17836 32620 17892
rect 32676 17836 32686 17892
rect 43372 17836 44044 17892
rect 44100 17836 44110 17892
rect 43372 17780 43428 17836
rect 5114 17724 5124 17780
rect 5180 17724 8540 17780
rect 8596 17724 8606 17780
rect 16604 17724 19292 17780
rect 19348 17724 20076 17780
rect 20132 17724 22764 17780
rect 22820 17724 23436 17780
rect 23492 17724 23502 17780
rect 28130 17724 28140 17780
rect 28196 17724 28588 17780
rect 28644 17724 30044 17780
rect 30100 17724 30110 17780
rect 37202 17724 37212 17780
rect 37268 17724 39004 17780
rect 39060 17724 39070 17780
rect 41122 17724 41132 17780
rect 41188 17724 41634 17780
rect 41690 17724 43372 17780
rect 43428 17724 43438 17780
rect 43586 17724 43596 17780
rect 43652 17724 43820 17780
rect 43876 17724 43886 17780
rect 5282 17612 5292 17668
rect 5348 17612 6412 17668
rect 6468 17612 10108 17668
rect 10164 17612 10174 17668
rect 12786 17612 12796 17668
rect 12852 17612 13020 17668
rect 13076 17612 14476 17668
rect 14532 17612 14542 17668
rect 4218 17500 4228 17556
rect 4284 17500 4676 17556
rect 4732 17500 5740 17556
rect 5796 17500 6860 17556
rect 6916 17500 6926 17556
rect 16604 17444 16660 17724
rect 17938 17612 17948 17668
rect 18004 17612 18172 17668
rect 18228 17612 18844 17668
rect 18900 17612 18910 17668
rect 19002 17612 19012 17668
rect 19068 17612 19628 17668
rect 19684 17612 19694 17668
rect 20290 17612 20300 17668
rect 20356 17612 21196 17668
rect 21252 17612 21262 17668
rect 23538 17612 23548 17668
rect 23604 17612 25228 17668
rect 25284 17612 25294 17668
rect 27178 17612 27188 17668
rect 27244 17612 35812 17668
rect 35868 17612 35878 17668
rect 37762 17612 37772 17668
rect 37828 17612 38220 17668
rect 38276 17612 38780 17668
rect 38836 17612 40124 17668
rect 40180 17612 40190 17668
rect 41458 17612 41468 17668
rect 41524 17612 42588 17668
rect 42644 17612 42654 17668
rect 43138 17612 43148 17668
rect 43204 17612 43932 17668
rect 43988 17612 44604 17668
rect 44660 17612 44670 17668
rect 49200 17556 50000 17584
rect 19170 17500 19180 17556
rect 19236 17500 20188 17556
rect 20244 17500 20254 17556
rect 21354 17500 21364 17556
rect 21420 17500 22092 17556
rect 22148 17500 22158 17556
rect 25890 17500 25900 17556
rect 25956 17500 26628 17556
rect 26684 17500 26694 17556
rect 38546 17500 38556 17556
rect 38612 17500 40908 17556
rect 40964 17500 40974 17556
rect 42914 17500 42924 17556
rect 42980 17500 43708 17556
rect 43764 17500 44380 17556
rect 44436 17500 44446 17556
rect 45266 17500 45276 17556
rect 45332 17500 48636 17556
rect 48692 17500 50000 17556
rect 49200 17472 50000 17500
rect 16594 17388 16604 17444
rect 16660 17388 16670 17444
rect 17938 17388 17948 17444
rect 18004 17388 19964 17444
rect 20020 17388 20030 17444
rect 25302 17388 25340 17444
rect 25396 17388 25406 17444
rect 26898 17388 26908 17444
rect 26964 17388 27244 17444
rect 27300 17388 28140 17444
rect 28196 17388 28206 17444
rect 34402 17388 34412 17444
rect 34468 17388 34860 17444
rect 34916 17388 42476 17444
rect 42532 17388 42542 17444
rect 22418 17276 22428 17332
rect 22484 17276 23324 17332
rect 23380 17276 23390 17332
rect 23706 17276 23716 17332
rect 23772 17276 28308 17332
rect 28364 17276 28700 17332
rect 28756 17276 28766 17332
rect 28924 17276 31164 17332
rect 31220 17276 31230 17332
rect 37202 17276 37212 17332
rect 37268 17276 37660 17332
rect 37716 17276 41356 17332
rect 41412 17276 41422 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 28924 17220 28980 17276
rect 20178 17164 20188 17220
rect 20244 17164 23212 17220
rect 23268 17164 24332 17220
rect 24388 17164 25452 17220
rect 25508 17164 25518 17220
rect 25722 17164 25732 17220
rect 25788 17164 26348 17220
rect 26404 17164 27580 17220
rect 27636 17164 27646 17220
rect 28130 17164 28140 17220
rect 28196 17164 28980 17220
rect 31042 17164 31052 17220
rect 31108 17164 33628 17220
rect 33684 17164 35980 17220
rect 36036 17164 36876 17220
rect 36932 17164 36942 17220
rect 38210 17164 38220 17220
rect 38276 17164 40796 17220
rect 40852 17164 40862 17220
rect 4330 17052 4340 17108
rect 4396 17052 5628 17108
rect 5684 17052 8316 17108
rect 8372 17052 8382 17108
rect 8754 17052 8764 17108
rect 8820 17052 9436 17108
rect 9492 17052 13356 17108
rect 13412 17052 15092 17108
rect 15148 17052 15158 17108
rect 19618 17052 19628 17108
rect 19684 17052 21196 17108
rect 21252 17052 21756 17108
rect 21812 17052 21822 17108
rect 23370 17052 23380 17108
rect 23436 17052 25116 17108
rect 25172 17052 26124 17108
rect 26180 17052 26190 17108
rect 26674 17052 26684 17108
rect 26740 17052 28476 17108
rect 28532 17052 28542 17108
rect 26124 16996 26180 17052
rect 29372 16996 29428 17108
rect 29484 17052 44940 17108
rect 44996 17052 45006 17108
rect 9986 16940 9996 16996
rect 10052 16940 12124 16996
rect 12180 16940 16268 16996
rect 16324 16940 16334 16996
rect 18050 16940 18060 16996
rect 18116 16940 23996 16996
rect 24052 16940 24062 16996
rect 26124 16940 29428 16996
rect 38612 16940 39564 16996
rect 39620 16940 43148 16996
rect 43204 16940 45500 16996
rect 45556 16940 45566 16996
rect 38612 16884 38668 16940
rect 9314 16828 9324 16884
rect 9380 16828 10108 16884
rect 10164 16828 11788 16884
rect 11844 16828 11854 16884
rect 16146 16828 16156 16884
rect 16212 16828 18732 16884
rect 18788 16828 18798 16884
rect 19058 16828 19068 16884
rect 19124 16828 21868 16884
rect 21924 16828 21934 16884
rect 22306 16828 22316 16884
rect 22372 16828 23660 16884
rect 23716 16828 23726 16884
rect 23874 16828 23884 16884
rect 23940 16828 25676 16884
rect 25732 16828 25742 16884
rect 26338 16828 26348 16884
rect 26404 16828 26908 16884
rect 26964 16828 26974 16884
rect 29698 16828 29708 16884
rect 29764 16828 33012 16884
rect 33068 16828 33078 16884
rect 33618 16828 33628 16884
rect 33684 16828 34244 16884
rect 34962 16828 34972 16884
rect 35028 16828 37548 16884
rect 37604 16828 38108 16884
rect 38164 16828 38668 16884
rect 39218 16828 39228 16884
rect 39284 16828 40012 16884
rect 40068 16828 40908 16884
rect 40964 16828 40974 16884
rect 42802 16828 42812 16884
rect 42868 16828 43708 16884
rect 43764 16828 43774 16884
rect 46946 16828 46956 16884
rect 47012 16828 47684 16884
rect 47740 16828 47750 16884
rect 34188 16772 34244 16828
rect 4722 16716 4732 16772
rect 4788 16716 5964 16772
rect 6020 16716 6030 16772
rect 16482 16716 16492 16772
rect 16548 16716 19180 16772
rect 19236 16716 19246 16772
rect 20962 16716 20972 16772
rect 21028 16716 21756 16772
rect 21812 16716 21822 16772
rect 22530 16716 22540 16772
rect 22596 16716 23436 16772
rect 23492 16716 23502 16772
rect 31826 16716 31836 16772
rect 31892 16716 33740 16772
rect 33796 16716 33806 16772
rect 34178 16716 34188 16772
rect 34244 16716 34254 16772
rect 34850 16716 34860 16772
rect 34916 16716 35644 16772
rect 35700 16716 35710 16772
rect 11554 16604 11564 16660
rect 11620 16604 12628 16660
rect 12684 16604 12694 16660
rect 19030 16604 19068 16660
rect 19124 16604 19134 16660
rect 26338 16604 26348 16660
rect 26404 16604 26460 16660
rect 26516 16604 26526 16660
rect 39666 16604 39676 16660
rect 39732 16604 40908 16660
rect 40964 16604 40974 16660
rect 19506 16492 19516 16548
rect 19572 16492 20636 16548
rect 20692 16492 20702 16548
rect 25442 16492 25452 16548
rect 25508 16492 29652 16548
rect 29708 16492 29718 16548
rect 37874 16492 37884 16548
rect 37940 16492 38892 16548
rect 38948 16492 38958 16548
rect 43698 16492 43708 16548
rect 43764 16492 48076 16548
rect 48132 16492 48142 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 14354 16380 14364 16436
rect 14420 16380 28028 16436
rect 28084 16380 28094 16436
rect 38612 16380 39228 16436
rect 39284 16380 39294 16436
rect 43250 16380 43260 16436
rect 43316 16380 43326 16436
rect 44370 16380 44380 16436
rect 44436 16380 45612 16436
rect 45668 16380 45678 16436
rect 16258 16268 16268 16324
rect 16324 16268 17052 16324
rect 17108 16268 17612 16324
rect 17668 16268 17678 16324
rect 20290 16268 20300 16324
rect 20356 16268 20366 16324
rect 22306 16268 22316 16324
rect 22372 16268 22876 16324
rect 22932 16268 22942 16324
rect 24994 16268 25004 16324
rect 25060 16268 25956 16324
rect 26012 16268 26684 16324
rect 26740 16268 26750 16324
rect 28354 16268 28364 16324
rect 28420 16268 34524 16324
rect 34580 16268 34590 16324
rect 20300 16212 20356 16268
rect 38612 16212 38668 16380
rect 43260 16324 43316 16380
rect 43260 16268 44884 16324
rect 44986 16268 44996 16324
rect 45052 16268 46060 16324
rect 46116 16268 46126 16324
rect 44828 16212 44884 16268
rect 6402 16156 6412 16212
rect 6468 16156 7196 16212
rect 7252 16156 7262 16212
rect 14924 16156 21252 16212
rect 22026 16156 22036 16212
rect 22092 16156 23884 16212
rect 23940 16156 23950 16212
rect 30594 16156 30604 16212
rect 30660 16156 30940 16212
rect 30996 16156 31164 16212
rect 31220 16156 36484 16212
rect 36540 16156 38668 16212
rect 42914 16156 42924 16212
rect 42980 16156 43820 16212
rect 43876 16156 44772 16212
rect 44828 16156 48412 16212
rect 48468 16156 48478 16212
rect 12898 16044 12908 16100
rect 12964 16044 13580 16100
rect 13636 16044 13646 16100
rect 14924 15988 14980 16156
rect 15810 16044 15820 16100
rect 15876 16044 16604 16100
rect 16660 16044 16670 16100
rect 17378 16044 17388 16100
rect 17444 16044 19740 16100
rect 19796 16044 19806 16100
rect 4274 15932 4284 15988
rect 4340 15932 4956 15988
rect 5012 15932 6188 15988
rect 6244 15932 6254 15988
rect 12002 15932 12012 15988
rect 12068 15932 12796 15988
rect 12852 15932 12862 15988
rect 14914 15932 14924 15988
rect 14980 15932 14990 15988
rect 17266 15932 17276 15988
rect 17332 15932 17948 15988
rect 18004 15932 20300 15988
rect 20356 15932 20366 15988
rect 4498 15820 4508 15876
rect 4564 15820 6972 15876
rect 7028 15820 7308 15876
rect 7364 15820 7374 15876
rect 13402 15820 13412 15876
rect 13468 15820 14756 15876
rect 14812 15820 14822 15876
rect 19170 15820 19180 15876
rect 19236 15820 20468 15876
rect 20524 15820 20534 15876
rect 21196 15764 21252 16156
rect 44716 16100 44772 16156
rect 22418 16044 22428 16100
rect 22484 16044 23212 16100
rect 23268 16044 23278 16100
rect 25414 16044 25452 16100
rect 25508 16044 25518 16100
rect 26226 16044 26236 16100
rect 26292 16044 26796 16100
rect 26852 16044 26862 16100
rect 29138 16044 29148 16100
rect 29204 16044 29820 16100
rect 29876 16044 29886 16100
rect 30202 16044 30212 16100
rect 30268 16044 33572 16100
rect 33628 16044 33638 16100
rect 38098 16044 38108 16100
rect 38164 16044 38444 16100
rect 38500 16044 38510 16100
rect 42522 16044 42532 16100
rect 42588 16044 43708 16100
rect 43764 16044 43774 16100
rect 44230 16044 44268 16100
rect 44324 16044 44334 16100
rect 44706 16044 44716 16100
rect 44772 16044 44782 16100
rect 45602 16044 45612 16100
rect 45668 16044 47068 16100
rect 47124 16044 47134 16100
rect 47282 16044 47292 16100
rect 47348 16044 47964 16100
rect 48020 16044 48030 16100
rect 21522 15932 21532 15988
rect 21588 15932 25004 15988
rect 25060 15932 25070 15988
rect 28522 15932 28532 15988
rect 28588 15932 33964 15988
rect 34020 15932 34030 15988
rect 40338 15932 40348 15988
rect 40404 15932 41132 15988
rect 41188 15932 41198 15988
rect 26058 15820 26068 15876
rect 26124 15820 26684 15876
rect 26740 15820 27468 15876
rect 27524 15820 27534 15876
rect 27906 15820 27916 15876
rect 27972 15820 29932 15876
rect 29988 15820 29998 15876
rect 35634 15820 35644 15876
rect 35700 15820 41580 15876
rect 41636 15820 41646 15876
rect 21196 15708 28532 15764
rect 28690 15708 28700 15764
rect 28756 15708 30044 15764
rect 30100 15708 42252 15764
rect 42308 15708 42318 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 28476 15652 28532 15708
rect 7130 15596 7140 15652
rect 7196 15596 8204 15652
rect 8260 15596 8270 15652
rect 21354 15596 21364 15652
rect 21420 15596 21868 15652
rect 21924 15596 21934 15652
rect 26338 15596 26348 15652
rect 26404 15596 26572 15652
rect 26628 15596 28420 15652
rect 28476 15596 33292 15652
rect 33348 15596 33358 15652
rect 41682 15596 41692 15652
rect 41748 15596 41972 15652
rect 42028 15596 45612 15652
rect 45668 15596 45678 15652
rect 46610 15596 46620 15652
rect 46676 15596 47516 15652
rect 47572 15596 47582 15652
rect 28364 15540 28420 15596
rect 3042 15484 3052 15540
rect 3108 15484 3500 15540
rect 3556 15484 3566 15540
rect 7420 15484 8316 15540
rect 8372 15484 8382 15540
rect 11330 15484 11340 15540
rect 11396 15484 13580 15540
rect 13636 15484 13646 15540
rect 19394 15484 19404 15540
rect 19460 15484 19740 15540
rect 19796 15484 19806 15540
rect 19964 15484 23324 15540
rect 23380 15484 28140 15540
rect 28196 15484 28206 15540
rect 28364 15484 29148 15540
rect 29204 15484 29214 15540
rect 40898 15484 40908 15540
rect 40964 15484 42476 15540
rect 42532 15484 42542 15540
rect 4946 15372 4956 15428
rect 5012 15372 5404 15428
rect 5460 15372 5964 15428
rect 6020 15372 6030 15428
rect 7420 15316 7476 15484
rect 19964 15428 20020 15484
rect 10322 15372 10332 15428
rect 10388 15372 15148 15428
rect 16202 15372 16212 15428
rect 16268 15372 18956 15428
rect 19012 15372 20020 15428
rect 20962 15372 20972 15428
rect 21028 15372 22540 15428
rect 22596 15372 22606 15428
rect 23426 15372 23436 15428
rect 23492 15372 30044 15428
rect 30100 15372 30110 15428
rect 41346 15372 41356 15428
rect 41412 15372 42140 15428
rect 42196 15372 43372 15428
rect 43428 15372 43438 15428
rect 3826 15260 3836 15316
rect 3892 15260 5068 15316
rect 5124 15260 5134 15316
rect 7410 15260 7420 15316
rect 7476 15260 7486 15316
rect 7746 15260 7756 15316
rect 7812 15260 8316 15316
rect 8372 15260 8382 15316
rect 8866 15260 8876 15316
rect 8932 15260 9492 15316
rect 9548 15260 9558 15316
rect 12562 15260 12572 15316
rect 12628 15260 14196 15316
rect 14252 15260 14262 15316
rect 7420 15204 7476 15260
rect 15092 15204 15148 15372
rect 17378 15260 17388 15316
rect 17444 15260 18620 15316
rect 18676 15260 22204 15316
rect 25218 15260 25228 15316
rect 25284 15260 26572 15316
rect 26628 15260 26638 15316
rect 28130 15260 28140 15316
rect 28196 15260 28532 15316
rect 28588 15260 28598 15316
rect 29362 15260 29372 15316
rect 29428 15260 29932 15316
rect 29988 15260 31836 15316
rect 31892 15260 31902 15316
rect 33730 15260 33740 15316
rect 33796 15260 34860 15316
rect 34916 15260 34926 15316
rect 41122 15260 41132 15316
rect 41188 15260 43260 15316
rect 43316 15260 43326 15316
rect 45490 15260 45500 15316
rect 45556 15260 48300 15316
rect 48356 15260 48366 15316
rect 4610 15148 4620 15204
rect 4676 15148 5292 15204
rect 5348 15148 5358 15204
rect 7420 15148 8092 15204
rect 8148 15148 8158 15204
rect 9650 15148 9660 15204
rect 9716 15148 10220 15204
rect 10276 15148 10286 15204
rect 13458 15148 13468 15204
rect 13524 15148 14924 15204
rect 14980 15148 14990 15204
rect 15092 15148 16212 15204
rect 16268 15148 16278 15204
rect 16594 15148 16604 15204
rect 16660 15148 21756 15204
rect 21812 15148 21822 15204
rect 22148 15092 22204 15260
rect 22306 15148 22316 15204
rect 22372 15148 22988 15204
rect 23044 15148 23212 15204
rect 23268 15148 23278 15204
rect 25722 15148 25732 15204
rect 25788 15148 25900 15204
rect 25956 15148 25966 15204
rect 29642 15148 29652 15204
rect 29764 15148 29774 15204
rect 32162 15148 32172 15204
rect 32228 15148 36036 15204
rect 36092 15148 36102 15204
rect 41234 15148 41244 15204
rect 41300 15148 41468 15204
rect 41524 15148 42364 15204
rect 42420 15148 42812 15204
rect 42868 15148 42878 15204
rect 43484 15148 43518 15204
rect 43574 15148 43584 15204
rect 45266 15148 45276 15204
rect 45332 15148 45724 15204
rect 45780 15148 45790 15204
rect 46386 15148 46396 15204
rect 46452 15148 46900 15204
rect 43484 15092 43540 15148
rect 9426 15036 9436 15092
rect 9492 15036 10332 15092
rect 10388 15036 12628 15092
rect 12572 14980 12628 15036
rect 15092 15036 15484 15092
rect 15540 15036 15550 15092
rect 22138 15036 22148 15092
rect 22204 15036 22214 15092
rect 24210 15036 24220 15092
rect 24276 15036 25900 15092
rect 25956 15036 25966 15092
rect 28914 15036 28924 15092
rect 28980 15036 29820 15092
rect 29876 15036 30492 15092
rect 30548 15036 30558 15092
rect 42018 15036 42028 15092
rect 42084 15036 43540 15092
rect 5842 14924 5852 14980
rect 5908 14924 6524 14980
rect 6580 14924 9548 14980
rect 9604 14924 10108 14980
rect 10164 14924 10174 14980
rect 12310 14924 12348 14980
rect 12404 14924 12414 14980
rect 12572 14924 12852 14980
rect 12908 14924 12918 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 15092 14868 15148 15036
rect 46844 14980 46900 15148
rect 20626 14924 20636 14980
rect 20692 14924 21196 14980
rect 21252 14924 24556 14980
rect 24612 14924 24622 14980
rect 25554 14924 25564 14980
rect 25620 14924 25788 14980
rect 25844 14924 25854 14980
rect 26114 14924 26124 14980
rect 26180 14924 26348 14980
rect 26404 14924 26414 14980
rect 27122 14924 27132 14980
rect 27188 14924 27692 14980
rect 27748 14924 27758 14980
rect 28802 14924 28812 14980
rect 28868 14924 29316 14980
rect 29372 14924 29382 14980
rect 44370 14924 44380 14980
rect 44436 14924 45164 14980
rect 45220 14924 45230 14980
rect 45378 14924 45388 14980
rect 45444 14924 45612 14980
rect 45668 14924 45678 14980
rect 46834 14924 46844 14980
rect 46900 14924 46910 14980
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 8530 14812 8540 14868
rect 8596 14812 8764 14868
rect 8820 14812 10614 14868
rect 10670 14812 15148 14868
rect 23314 14812 23324 14868
rect 23380 14812 29372 14868
rect 29428 14812 29438 14868
rect 38322 14812 38332 14868
rect 38388 14812 39228 14868
rect 39284 14812 39294 14868
rect 22418 14700 22428 14756
rect 22484 14700 23996 14756
rect 24052 14700 27244 14756
rect 27300 14700 27310 14756
rect 16034 14588 16044 14644
rect 16100 14588 18396 14644
rect 18452 14588 18462 14644
rect 27458 14588 27468 14644
rect 27524 14588 28364 14644
rect 28420 14588 28430 14644
rect 36306 14588 36316 14644
rect 36372 14588 37212 14644
rect 37268 14588 42700 14644
rect 42756 14588 42766 14644
rect 45126 14588 45164 14644
rect 45220 14588 46172 14644
rect 46228 14588 46238 14644
rect 4722 14476 4732 14532
rect 4788 14476 6076 14532
rect 6132 14476 6524 14532
rect 6580 14476 6590 14532
rect 10322 14476 10332 14532
rect 10388 14476 12348 14532
rect 12404 14476 12460 14532
rect 12516 14476 12526 14532
rect 14018 14476 14028 14532
rect 14084 14476 14476 14532
rect 14532 14476 14542 14532
rect 19338 14476 19348 14532
rect 19404 14476 19628 14532
rect 19684 14476 19694 14532
rect 24658 14476 24668 14532
rect 24724 14476 25228 14532
rect 25284 14476 26684 14532
rect 26740 14476 27804 14532
rect 27860 14476 29148 14532
rect 29204 14476 29214 14532
rect 30370 14476 30380 14532
rect 30436 14476 33180 14532
rect 33236 14476 33628 14532
rect 33684 14476 33964 14532
rect 34020 14476 35868 14532
rect 35924 14476 35934 14532
rect 39442 14476 39452 14532
rect 39508 14476 40292 14532
rect 40348 14476 40358 14532
rect 44482 14476 44492 14532
rect 44548 14476 45836 14532
rect 45892 14476 45902 14532
rect 8306 14364 8316 14420
rect 8372 14364 10444 14420
rect 10500 14364 10892 14420
rect 10948 14364 10958 14420
rect 12338 14364 12348 14420
rect 12404 14364 14924 14420
rect 14980 14364 14990 14420
rect 15082 14364 15092 14420
rect 15148 14364 20412 14420
rect 20468 14364 20478 14420
rect 26226 14364 26236 14420
rect 26292 14364 28140 14420
rect 28196 14364 28206 14420
rect 29306 14364 29316 14420
rect 29428 14364 29438 14420
rect 29866 14364 29876 14420
rect 29932 14364 37940 14420
rect 37996 14364 38006 14420
rect 38322 14364 38332 14420
rect 38388 14364 40964 14420
rect 41020 14364 41030 14420
rect 5058 14252 5068 14308
rect 5124 14252 8428 14308
rect 8484 14252 10108 14308
rect 10164 14252 10174 14308
rect 19338 14252 19348 14308
rect 19404 14252 28868 14308
rect 28924 14252 30940 14308
rect 30996 14252 31006 14308
rect 36642 14252 36652 14308
rect 36708 14252 38556 14308
rect 38612 14252 39676 14308
rect 39732 14252 39742 14308
rect 40450 14252 40460 14308
rect 40516 14252 42812 14308
rect 42868 14252 42878 14308
rect 44930 14252 44940 14308
rect 44996 14252 45948 14308
rect 46004 14252 46014 14308
rect 6962 14140 6972 14196
rect 7028 14140 11900 14196
rect 11956 14140 11966 14196
rect 19628 14084 19684 14252
rect 20962 14140 20972 14196
rect 21028 14140 21420 14196
rect 21476 14140 21486 14196
rect 22642 14140 22652 14196
rect 22708 14140 26908 14196
rect 27010 14140 27020 14196
rect 27076 14140 28140 14196
rect 28196 14140 29484 14196
rect 29540 14140 30604 14196
rect 30660 14140 30670 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 13794 14028 13804 14084
rect 13860 14028 14364 14084
rect 14420 14028 19404 14084
rect 19460 14028 19470 14084
rect 19618 14028 19628 14084
rect 19684 14028 19694 14084
rect 25414 14028 25452 14084
rect 25508 14028 25518 14084
rect 25722 14028 25732 14084
rect 25844 14028 25854 14084
rect 26646 14028 26684 14084
rect 26740 14028 26750 14084
rect 26852 14028 26908 14140
rect 26964 14028 26974 14084
rect 28242 14028 28252 14084
rect 28308 14028 29596 14084
rect 29652 14028 30716 14084
rect 30772 14028 30782 14084
rect 36306 14028 36316 14084
rect 36372 14028 37716 14084
rect 37772 14028 44380 14084
rect 44436 14028 44446 14084
rect 45154 14028 45164 14084
rect 45220 14028 45230 14084
rect 26908 13972 26964 14028
rect 2034 13916 2044 13972
rect 2100 13916 3388 13972
rect 3444 13916 4900 13972
rect 4956 13916 4966 13972
rect 14466 13916 14476 13972
rect 14532 13916 14700 13972
rect 14756 13916 22932 13972
rect 22988 13916 24108 13972
rect 24164 13916 24174 13972
rect 24770 13916 24780 13972
rect 24836 13916 25340 13972
rect 25396 13916 25900 13972
rect 25956 13916 26572 13972
rect 26628 13916 26638 13972
rect 26908 13916 30156 13972
rect 30212 13916 30222 13972
rect 30426 13916 30436 13972
rect 30492 13916 31276 13972
rect 31332 13916 31342 13972
rect 34402 13916 34412 13972
rect 34468 13916 36204 13972
rect 36260 13916 36270 13972
rect 39946 13916 39956 13972
rect 40012 13916 40684 13972
rect 40740 13916 41412 13972
rect 41468 13916 41478 13972
rect 45164 13860 45220 14028
rect 19842 13804 19852 13860
rect 19908 13804 21756 13860
rect 21812 13804 26684 13860
rect 26740 13804 27020 13860
rect 27076 13804 27086 13860
rect 27402 13804 27412 13860
rect 27468 13804 36036 13860
rect 36092 13804 36102 13860
rect 43026 13804 43036 13860
rect 43092 13804 45724 13860
rect 45780 13804 46508 13860
rect 46564 13804 46574 13860
rect 44828 13748 44884 13804
rect 3490 13692 3500 13748
rect 3556 13692 5964 13748
rect 6020 13692 6030 13748
rect 8530 13692 8540 13748
rect 8596 13692 10220 13748
rect 10276 13692 10286 13748
rect 14242 13692 14252 13748
rect 14308 13692 14476 13748
rect 14532 13692 15372 13748
rect 15428 13692 15438 13748
rect 15754 13692 15764 13748
rect 15820 13692 16380 13748
rect 16436 13692 17612 13748
rect 17668 13692 17948 13748
rect 18004 13692 18014 13748
rect 18106 13692 18116 13748
rect 18172 13692 18620 13748
rect 18676 13692 18686 13748
rect 19506 13692 19516 13748
rect 19572 13692 20300 13748
rect 20356 13692 20860 13748
rect 20916 13692 21980 13748
rect 22036 13692 22046 13748
rect 26338 13692 26348 13748
rect 26404 13692 26572 13748
rect 26628 13692 26638 13748
rect 26852 13692 30100 13748
rect 30258 13692 30268 13748
rect 30324 13692 31388 13748
rect 31444 13692 31454 13748
rect 31724 13692 32732 13748
rect 32788 13692 32798 13748
rect 33058 13692 33068 13748
rect 33124 13692 35532 13748
rect 35588 13692 36652 13748
rect 36708 13692 36718 13748
rect 41794 13692 41804 13748
rect 41860 13692 44492 13748
rect 44548 13692 44558 13748
rect 44818 13692 44828 13748
rect 44884 13692 44894 13748
rect 45938 13692 45948 13748
rect 46004 13692 46014 13748
rect 8866 13580 8876 13636
rect 8932 13580 9548 13636
rect 9604 13580 9614 13636
rect 14914 13580 14924 13636
rect 14980 13580 15596 13636
rect 15652 13580 15662 13636
rect 16874 13580 16884 13636
rect 16940 13580 18508 13636
rect 18564 13580 18574 13636
rect 21298 13580 21308 13636
rect 21364 13580 22428 13636
rect 22484 13580 22494 13636
rect 26786 13580 26796 13636
rect 26852 13580 26908 13692
rect 30044 13636 30100 13692
rect 31724 13636 31780 13692
rect 45948 13636 46004 13692
rect 27346 13580 27356 13636
rect 27412 13580 28252 13636
rect 28308 13580 28318 13636
rect 30044 13580 31164 13636
rect 31220 13580 31780 13636
rect 31938 13580 31948 13636
rect 32004 13580 33740 13636
rect 33796 13580 33806 13636
rect 41906 13580 41916 13636
rect 41972 13580 43484 13636
rect 43540 13580 43550 13636
rect 44650 13580 44660 13636
rect 44716 13580 45276 13636
rect 45332 13580 46004 13636
rect 6738 13468 6748 13524
rect 6804 13468 7420 13524
rect 7476 13468 7980 13524
rect 8036 13468 9100 13524
rect 9156 13468 9166 13524
rect 15138 13468 15148 13524
rect 15204 13468 16156 13524
rect 16212 13468 16222 13524
rect 22306 13468 22316 13524
rect 22372 13468 22540 13524
rect 22596 13468 25396 13524
rect 25452 13468 26908 13524
rect 28354 13468 28364 13524
rect 28420 13468 30436 13524
rect 30492 13468 30502 13524
rect 30986 13468 30996 13524
rect 31052 13468 38892 13524
rect 38948 13468 38958 13524
rect 43250 13468 43260 13524
rect 43316 13468 47628 13524
rect 47684 13468 48076 13524
rect 48132 13468 48142 13524
rect 26852 13412 26908 13468
rect 6290 13356 6300 13412
rect 6356 13356 6860 13412
rect 6916 13356 6926 13412
rect 8082 13356 8092 13412
rect 8148 13356 8652 13412
rect 8708 13356 8718 13412
rect 12954 13356 12964 13412
rect 13020 13356 16492 13412
rect 16548 13356 16558 13412
rect 20962 13356 20972 13412
rect 21028 13356 22092 13412
rect 22148 13356 22158 13412
rect 23062 13356 23100 13412
rect 23156 13356 23166 13412
rect 25442 13356 25452 13412
rect 25508 13356 25564 13412
rect 25620 13356 25630 13412
rect 26852 13356 27692 13412
rect 27748 13356 28700 13412
rect 28756 13356 28766 13412
rect 29810 13356 29820 13412
rect 29876 13356 30156 13412
rect 30212 13356 30222 13412
rect 36194 13356 36204 13412
rect 36260 13356 36876 13412
rect 36932 13356 38220 13412
rect 38276 13356 38286 13412
rect 43381 13356 43391 13412
rect 43447 13356 44044 13412
rect 44100 13356 44940 13412
rect 44996 13356 45500 13412
rect 45556 13356 45566 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 11890 13244 11900 13300
rect 11956 13244 34692 13300
rect 34748 13244 34758 13300
rect 37874 13244 37884 13300
rect 37940 13244 39284 13300
rect 14802 13132 14812 13188
rect 14868 13132 21700 13188
rect 21756 13132 21766 13188
rect 22306 13132 22316 13188
rect 22372 13132 23436 13188
rect 23492 13132 27076 13188
rect 27132 13132 27804 13188
rect 27860 13132 27870 13188
rect 30258 13132 30268 13188
rect 30324 13132 31724 13188
rect 31780 13132 31790 13188
rect 37314 13132 37324 13188
rect 37380 13132 37772 13188
rect 37828 13132 37838 13188
rect 6290 13020 6300 13076
rect 6356 13020 8092 13076
rect 8148 13020 8158 13076
rect 15474 13020 15484 13076
rect 15540 13020 17500 13076
rect 17556 13020 18788 13076
rect 18844 13020 18854 13076
rect 20738 13020 20748 13076
rect 20804 13020 22876 13076
rect 22932 13020 24892 13076
rect 24948 13020 25676 13076
rect 25732 13020 25742 13076
rect 25946 13020 25956 13076
rect 26012 13020 30548 13076
rect 30604 13020 30614 13076
rect 35802 13020 35812 13076
rect 35868 13020 37100 13076
rect 37156 13020 37166 13076
rect 37650 13020 37660 13076
rect 37716 13020 38668 13076
rect 38724 13020 38734 13076
rect 13682 12908 13692 12964
rect 13748 12908 13758 12964
rect 20626 12908 20636 12964
rect 20692 12908 21756 12964
rect 21812 12908 22764 12964
rect 22820 12908 22830 12964
rect 23314 12908 23324 12964
rect 23380 12908 23390 12964
rect 23538 12908 23548 12964
rect 23604 12908 24444 12964
rect 24500 12908 24510 12964
rect 25162 12908 25172 12964
rect 25228 12908 31668 12964
rect 31724 12908 31734 12964
rect 32050 12908 32060 12964
rect 32116 12908 33572 12964
rect 33628 12908 33638 12964
rect 34850 12908 34860 12964
rect 34916 12908 35196 12964
rect 35252 12908 36204 12964
rect 36260 12908 36270 12964
rect 37174 12908 37212 12964
rect 37268 12908 37278 12964
rect 6962 12796 6972 12852
rect 7028 12796 8652 12852
rect 8708 12796 8718 12852
rect 13692 12740 13748 12908
rect 23324 12852 23380 12908
rect 23034 12796 23044 12852
rect 23100 12796 24332 12852
rect 24388 12796 24398 12852
rect 24602 12796 24612 12852
rect 24668 12796 29596 12852
rect 29652 12796 29662 12852
rect 30706 12796 30716 12852
rect 30772 12796 31388 12852
rect 31444 12796 31454 12852
rect 8418 12684 8428 12740
rect 8484 12684 8764 12740
rect 8820 12684 8830 12740
rect 10770 12684 10780 12740
rect 10836 12684 11564 12740
rect 11620 12684 12124 12740
rect 12180 12684 12190 12740
rect 12506 12684 12516 12740
rect 12572 12684 13356 12740
rect 13412 12684 13422 12740
rect 13692 12684 13804 12740
rect 13860 12684 13870 12740
rect 23762 12684 23772 12740
rect 23828 12684 29036 12740
rect 29092 12684 29102 12740
rect 33730 12684 33740 12740
rect 33796 12684 35644 12740
rect 35700 12684 37156 12740
rect 37212 12684 37222 12740
rect 37986 12684 37996 12740
rect 38052 12684 38444 12740
rect 38500 12684 38510 12740
rect 39340 12684 39396 13300
rect 44258 13244 44268 13300
rect 44324 13244 44604 13300
rect 44660 13244 44670 13300
rect 45154 13244 45164 13300
rect 45220 13244 45276 13300
rect 45332 13244 45342 13300
rect 40674 12796 40684 12852
rect 40740 12796 41298 12852
rect 41354 12796 41364 12852
rect 39452 12684 39462 12740
rect 44258 12684 44268 12740
rect 44324 12684 45724 12740
rect 45780 12684 46172 12740
rect 46228 12684 46238 12740
rect 49200 12628 50000 12656
rect 14438 12572 14476 12628
rect 14532 12572 14542 12628
rect 25442 12572 25452 12628
rect 25508 12572 26012 12628
rect 26068 12572 30268 12628
rect 30324 12572 30334 12628
rect 30930 12572 30940 12628
rect 30996 12572 32340 12628
rect 32396 12572 32406 12628
rect 33282 12572 33292 12628
rect 33348 12572 36204 12628
rect 36260 12572 36484 12628
rect 36540 12572 36550 12628
rect 36978 12572 36988 12628
rect 37044 12572 40572 12628
rect 40628 12572 42140 12628
rect 42196 12572 42206 12628
rect 46472 12572 46482 12628
rect 46538 12572 47292 12628
rect 47348 12572 47358 12628
rect 48290 12572 48300 12628
rect 48356 12572 50000 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 49200 12544 50000 12572
rect 6402 12460 6412 12516
rect 6468 12460 16156 12516
rect 16212 12460 16222 12516
rect 23986 12460 23996 12516
rect 24052 12460 31612 12516
rect 31668 12460 31678 12516
rect 37426 12460 37436 12516
rect 37492 12460 38556 12516
rect 38612 12460 41132 12516
rect 41188 12460 41804 12516
rect 41860 12460 42700 12516
rect 42756 12460 42766 12516
rect 47506 12460 47516 12516
rect 47572 12460 48132 12516
rect 48188 12460 48198 12516
rect 18050 12348 18060 12404
rect 18116 12348 18564 12404
rect 18620 12348 18956 12404
rect 19012 12348 19022 12404
rect 19674 12348 19684 12404
rect 19740 12348 22484 12404
rect 22540 12348 22550 12404
rect 29978 12348 29988 12404
rect 30044 12348 31500 12404
rect 31556 12348 31566 12404
rect 33450 12348 33460 12404
rect 33516 12348 35756 12404
rect 35812 12348 35822 12404
rect 37314 12348 37324 12404
rect 37380 12348 37390 12404
rect 37538 12348 37548 12404
rect 37604 12348 41020 12404
rect 41076 12348 41086 12404
rect 42876 12348 42886 12404
rect 42942 12348 43596 12404
rect 43652 12348 47964 12404
rect 48020 12348 48030 12404
rect 37324 12292 37380 12348
rect 6626 12236 6636 12292
rect 6692 12236 7196 12292
rect 7252 12236 7262 12292
rect 13626 12236 13636 12292
rect 13692 12236 13916 12292
rect 13972 12236 13982 12292
rect 21634 12236 21644 12292
rect 21700 12236 22092 12292
rect 22148 12236 22158 12292
rect 23370 12236 23380 12292
rect 23436 12236 28364 12292
rect 28420 12236 28430 12292
rect 37324 12236 38556 12292
rect 38612 12236 38622 12292
rect 40226 12236 40236 12292
rect 40292 12236 41244 12292
rect 41300 12236 41310 12292
rect 44230 12236 44268 12292
rect 44324 12236 44334 12292
rect 45378 12236 45388 12292
rect 45444 12236 45612 12292
rect 45668 12236 45678 12292
rect 8978 12124 8988 12180
rect 9044 12124 9436 12180
rect 9492 12124 9502 12180
rect 17490 12124 17500 12180
rect 17556 12124 17836 12180
rect 17892 12124 17902 12180
rect 19394 12124 19404 12180
rect 19460 12124 19852 12180
rect 19908 12124 19918 12180
rect 21746 12124 21756 12180
rect 21812 12124 21980 12180
rect 22036 12124 23100 12180
rect 23156 12124 23166 12180
rect 24770 12124 24780 12180
rect 24836 12124 25676 12180
rect 25732 12124 25742 12180
rect 28466 12124 28476 12180
rect 28532 12124 29820 12180
rect 29876 12124 29886 12180
rect 30146 12124 30156 12180
rect 30212 12124 31106 12180
rect 31162 12124 31612 12180
rect 31668 12124 31678 12180
rect 34514 12124 34524 12180
rect 34580 12124 35644 12180
rect 35700 12124 35710 12180
rect 36866 12124 36876 12180
rect 36932 12124 37324 12180
rect 37380 12124 37390 12180
rect 37548 12124 38892 12180
rect 38948 12124 38958 12180
rect 39946 12124 39956 12180
rect 40012 12124 42028 12180
rect 42084 12124 42094 12180
rect 43250 12124 43260 12180
rect 43316 12124 44940 12180
rect 44996 12124 47068 12180
rect 47124 12124 47134 12180
rect 47282 12124 47292 12180
rect 47348 12124 47358 12180
rect 37548 12068 37604 12124
rect 47292 12068 47348 12124
rect 11554 12012 11564 12068
rect 11620 12012 14588 12068
rect 14644 12012 14654 12068
rect 18162 12012 18172 12068
rect 18228 12012 20804 12068
rect 20860 12012 21700 12068
rect 22418 12012 22428 12068
rect 22484 12012 23548 12068
rect 23604 12012 23614 12068
rect 30370 12012 30380 12068
rect 30436 12012 34692 12068
rect 34748 12012 34758 12068
rect 36194 12012 36204 12068
rect 36260 12012 37604 12068
rect 38546 12012 38556 12068
rect 38612 12012 41356 12068
rect 41412 12012 41804 12068
rect 41860 12012 41870 12068
rect 45154 12012 45164 12068
rect 45220 12012 47348 12068
rect 21644 11956 21700 12012
rect 30604 11956 30660 12012
rect 19058 11900 19068 11956
rect 19124 11900 20188 11956
rect 20244 11900 21420 11956
rect 21476 11900 21486 11956
rect 21644 11900 23772 11956
rect 23828 11900 23838 11956
rect 30594 11900 30604 11956
rect 30660 11900 30670 11956
rect 32498 11900 32508 11956
rect 32564 11900 37548 11956
rect 37604 11900 37614 11956
rect 40338 11900 40348 11956
rect 40404 11900 41020 11956
rect 41076 11900 44660 11956
rect 44716 11900 46172 11956
rect 46228 11900 46238 11956
rect 33404 11844 33460 11900
rect 6748 11788 7252 11844
rect 7308 11788 10108 11844
rect 10164 11788 10780 11844
rect 10836 11788 10846 11844
rect 17602 11788 17612 11844
rect 17668 11788 20300 11844
rect 20356 11788 21252 11844
rect 21308 11788 21924 11844
rect 22586 11788 22596 11844
rect 22652 11788 23380 11844
rect 23436 11788 23446 11844
rect 33394 11788 33404 11844
rect 33460 11788 33470 11844
rect 36754 11788 36764 11844
rect 36820 11788 37436 11844
rect 37492 11788 37502 11844
rect 40348 11788 40684 11844
rect 40740 11788 42476 11844
rect 42532 11788 43484 11844
rect 43540 11788 43550 11844
rect 45826 11788 45836 11844
rect 45892 11788 46956 11844
rect 47012 11788 47022 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 6748 11732 6804 11788
rect 21868 11732 21924 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 40348 11732 40404 11788
rect 3332 11508 3388 11732
rect 3444 11676 3948 11732
rect 4004 11676 4014 11732
rect 6188 11676 6804 11732
rect 16370 11676 16380 11732
rect 16436 11676 16716 11732
rect 16772 11676 16782 11732
rect 18722 11676 18732 11732
rect 18788 11676 19404 11732
rect 19460 11676 19470 11732
rect 21858 11676 21868 11732
rect 21924 11676 21934 11732
rect 22418 11676 22428 11732
rect 22484 11676 23156 11732
rect 23212 11676 25900 11732
rect 25956 11676 26124 11732
rect 26180 11676 26190 11732
rect 26348 11676 33292 11732
rect 33348 11676 34300 11732
rect 34356 11676 34366 11732
rect 36026 11676 36036 11732
rect 36092 11676 38332 11732
rect 38388 11676 39004 11732
rect 39060 11676 39070 11732
rect 40338 11676 40348 11732
rect 40404 11676 40414 11732
rect 43138 11676 43148 11732
rect 43204 11676 43820 11732
rect 43876 11676 43886 11732
rect 3948 11620 4004 11676
rect 6188 11620 6244 11676
rect 26348 11620 26404 11676
rect 3948 11564 5124 11620
rect 5180 11564 6188 11620
rect 6244 11564 6254 11620
rect 16156 11564 26404 11620
rect 26674 11564 26684 11620
rect 26740 11564 26750 11620
rect 27010 11564 27020 11620
rect 27076 11564 27086 11620
rect 33842 11564 33852 11620
rect 33908 11564 35476 11620
rect 35532 11564 35542 11620
rect 35858 11564 35868 11620
rect 35924 11564 37100 11620
rect 37156 11564 37166 11620
rect 1810 11452 1820 11508
rect 1876 11452 3388 11508
rect 5506 11452 5516 11508
rect 5572 11452 6860 11508
rect 6916 11452 6926 11508
rect 4498 11340 4508 11396
rect 4564 11340 5628 11396
rect 5684 11340 6412 11396
rect 6468 11340 6478 11396
rect 7858 11340 7868 11396
rect 7924 11340 8316 11396
rect 8372 11340 9100 11396
rect 9156 11340 9166 11396
rect 14130 11340 14140 11396
rect 14196 11340 14812 11396
rect 14868 11340 14878 11396
rect 15112 11340 15122 11396
rect 15178 11340 15596 11396
rect 15652 11340 15662 11396
rect 4386 11228 4396 11284
rect 4452 11228 5964 11284
rect 6020 11228 6860 11284
rect 6916 11228 7756 11284
rect 7812 11228 7822 11284
rect 10882 11228 10892 11284
rect 10948 11228 15260 11284
rect 15316 11228 15326 11284
rect 16156 11172 16212 11564
rect 26684 11508 26740 11564
rect 17154 11452 17164 11508
rect 17220 11452 17724 11508
rect 17780 11452 17790 11508
rect 24490 11452 24500 11508
rect 24556 11452 25564 11508
rect 25620 11452 26348 11508
rect 26404 11452 26740 11508
rect 27020 11508 27076 11564
rect 27020 11452 27580 11508
rect 27636 11452 47964 11508
rect 48020 11452 48030 11508
rect 16370 11340 16380 11396
rect 16436 11340 17052 11396
rect 17108 11340 17118 11396
rect 19618 11340 19628 11396
rect 19684 11340 21700 11396
rect 21756 11340 21766 11396
rect 24042 11340 24052 11396
rect 24108 11340 24332 11396
rect 24388 11340 26236 11396
rect 26292 11340 26302 11396
rect 26562 11340 26572 11396
rect 26628 11340 26796 11396
rect 26852 11340 27020 11396
rect 27076 11340 27086 11396
rect 34178 11340 34188 11396
rect 34244 11340 34972 11396
rect 35028 11340 35038 11396
rect 35130 11340 35140 11396
rect 35196 11340 35756 11396
rect 35812 11340 35822 11396
rect 37174 11340 37212 11396
rect 37268 11340 37278 11396
rect 37538 11340 37548 11396
rect 37604 11340 38892 11396
rect 38948 11340 38958 11396
rect 40226 11340 40236 11396
rect 40292 11340 41804 11396
rect 41860 11340 41870 11396
rect 42578 11340 42588 11396
rect 42644 11340 42654 11396
rect 43932 11340 46844 11396
rect 46900 11340 46910 11396
rect 42588 11284 42644 11340
rect 23090 11228 23100 11284
rect 23156 11228 30100 11284
rect 30156 11228 30940 11284
rect 30996 11228 31006 11284
rect 34514 11228 34524 11284
rect 34580 11228 35532 11284
rect 35588 11228 35868 11284
rect 35924 11228 35934 11284
rect 40562 11228 40572 11284
rect 40628 11228 41580 11284
rect 41636 11228 41646 11284
rect 42588 11228 42924 11284
rect 42980 11228 42990 11284
rect 43932 11172 43988 11340
rect 46472 11228 46482 11284
rect 46538 11228 46956 11284
rect 47012 11228 47022 11284
rect 5282 11116 5292 11172
rect 5348 11116 7532 11172
rect 7588 11116 7598 11172
rect 14018 11116 14028 11172
rect 14084 11116 15596 11172
rect 15652 11116 16212 11172
rect 17602 11116 17612 11172
rect 17668 11116 18844 11172
rect 18900 11116 18910 11172
rect 26450 11116 26460 11172
rect 26516 11116 26908 11172
rect 28018 11116 28028 11172
rect 28084 11116 29652 11172
rect 29708 11116 30268 11172
rect 30324 11116 30716 11172
rect 30772 11116 30782 11172
rect 32610 11116 32620 11172
rect 32676 11116 39228 11172
rect 39284 11116 43988 11172
rect 45826 11116 45836 11172
rect 45892 11116 48300 11172
rect 48356 11116 48366 11172
rect 26852 11060 26908 11116
rect 26852 11004 27356 11060
rect 27412 11004 27636 11060
rect 27692 11004 28364 11060
rect 28420 11004 28430 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 13346 10892 13356 10948
rect 13412 10892 14364 10948
rect 14420 10892 14430 10948
rect 23762 10892 23772 10948
rect 23828 10892 38556 10948
rect 38612 10892 44492 10948
rect 44548 10892 44996 10948
rect 45052 10892 45062 10948
rect 3266 10780 3276 10836
rect 3332 10780 5068 10836
rect 5124 10780 5134 10836
rect 15362 10780 15372 10836
rect 15428 10780 15764 10836
rect 15820 10780 15830 10836
rect 21746 10780 21756 10836
rect 21812 10780 21980 10836
rect 22036 10780 22046 10836
rect 24770 10780 24780 10836
rect 24836 10780 25452 10836
rect 25508 10780 26684 10836
rect 26740 10780 26750 10836
rect 26852 10780 36988 10836
rect 37044 10780 37054 10836
rect 44818 10780 44828 10836
rect 44884 10780 45388 10836
rect 45444 10780 45454 10836
rect 26852 10724 26908 10780
rect 12786 10668 12796 10724
rect 12852 10668 13962 10724
rect 14018 10668 16380 10724
rect 16436 10668 16446 10724
rect 17500 10668 26908 10724
rect 30706 10668 30716 10724
rect 30772 10668 32956 10724
rect 33012 10668 34020 10724
rect 34076 10668 34086 10724
rect 41682 10668 41692 10724
rect 41748 10668 44044 10724
rect 44100 10668 44110 10724
rect 17500 10612 17556 10668
rect 13234 10556 13244 10612
rect 13300 10556 14364 10612
rect 14420 10556 14924 10612
rect 14980 10556 14990 10612
rect 16482 10556 16492 10612
rect 16548 10556 17500 10612
rect 17556 10556 17566 10612
rect 26506 10556 26516 10612
rect 26572 10556 27636 10612
rect 27692 10556 27702 10612
rect 35970 10556 35980 10612
rect 36036 10556 37100 10612
rect 37156 10556 37324 10612
rect 37380 10556 37390 10612
rect 37986 10556 37996 10612
rect 38052 10556 38668 10612
rect 38724 10556 38734 10612
rect 41010 10556 41020 10612
rect 41076 10556 41580 10612
rect 41636 10556 41646 10612
rect 43362 10556 43372 10612
rect 43428 10556 45948 10612
rect 46004 10556 46014 10612
rect 47058 10556 47068 10612
rect 47124 10556 48132 10612
rect 48188 10556 48198 10612
rect 4498 10444 4508 10500
rect 4564 10444 5180 10500
rect 5236 10444 5246 10500
rect 6962 10444 6972 10500
rect 7028 10444 8204 10500
rect 8260 10444 8270 10500
rect 15026 10444 15036 10500
rect 15092 10444 19852 10500
rect 19908 10444 20524 10500
rect 20580 10444 20590 10500
rect 30706 10444 30716 10500
rect 30772 10444 32508 10500
rect 32564 10444 32574 10500
rect 36978 10444 36988 10500
rect 37044 10444 44100 10500
rect 44156 10444 44166 10500
rect 13794 10332 13804 10388
rect 13860 10332 14588 10388
rect 14644 10332 15372 10388
rect 15428 10332 15438 10388
rect 24210 10332 24220 10388
rect 24276 10332 26908 10388
rect 27066 10332 27076 10388
rect 27132 10332 27580 10388
rect 27636 10332 27646 10388
rect 29978 10332 29988 10388
rect 30044 10332 31276 10388
rect 31332 10332 31342 10388
rect 34972 10332 36652 10388
rect 36708 10332 38332 10388
rect 38388 10332 38668 10388
rect 38770 10332 38780 10388
rect 38836 10332 38846 10388
rect 40674 10332 40684 10388
rect 40740 10332 41580 10388
rect 41636 10332 43372 10388
rect 43428 10332 43438 10388
rect 26852 10276 26908 10332
rect 26852 10220 32340 10276
rect 32498 10220 32508 10276
rect 32564 10220 34412 10276
rect 34468 10220 34478 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 32284 10164 32340 10220
rect 34972 10164 35028 10332
rect 38612 10276 38668 10332
rect 38780 10276 38836 10332
rect 38612 10220 42644 10276
rect 42700 10220 42710 10276
rect 45378 10220 45388 10276
rect 45444 10220 45724 10276
rect 45780 10220 46732 10276
rect 46788 10220 46798 10276
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 20794 10108 20804 10164
rect 20860 10108 22652 10164
rect 22708 10108 22718 10164
rect 23426 10108 23436 10164
rect 23492 10108 24220 10164
rect 24276 10108 26908 10164
rect 26964 10108 26974 10164
rect 30538 10108 30548 10164
rect 30604 10108 30940 10164
rect 30996 10108 31836 10164
rect 31892 10108 31902 10164
rect 32284 10108 34132 10164
rect 34188 10108 35028 10164
rect 46834 10108 46844 10164
rect 46900 10108 47628 10164
rect 47684 10108 47694 10164
rect 26852 10052 26908 10108
rect 2594 9996 2604 10052
rect 2660 9996 5740 10052
rect 5796 9996 5806 10052
rect 12114 9996 12124 10052
rect 12180 9996 13020 10052
rect 13076 9996 13524 10052
rect 13580 9996 14700 10052
rect 14756 9996 14766 10052
rect 22764 9996 23660 10052
rect 23716 9996 25676 10052
rect 25732 9996 25742 10052
rect 26852 9996 31892 10052
rect 38658 9996 38668 10052
rect 38724 9996 39732 10052
rect 39788 9996 39798 10052
rect 6290 9884 6300 9940
rect 6356 9884 7308 9940
rect 7364 9884 7374 9940
rect 19394 9884 19404 9940
rect 19460 9884 22540 9940
rect 22596 9884 22606 9940
rect 22698 9884 22708 9940
rect 22764 9884 22820 9996
rect 31836 9940 31892 9996
rect 23370 9884 23380 9940
rect 23436 9884 23884 9940
rect 23940 9884 23950 9940
rect 25106 9884 25116 9940
rect 25172 9884 25452 9940
rect 25508 9884 25518 9940
rect 28802 9884 28812 9940
rect 28868 9884 29820 9940
rect 29876 9884 29886 9940
rect 31826 9884 31836 9940
rect 31892 9884 31902 9940
rect 36306 9884 36316 9940
rect 36372 9884 37604 9940
rect 37660 9884 37670 9940
rect 38098 9884 38108 9940
rect 38164 9884 40236 9940
rect 40292 9884 40302 9940
rect 39452 9828 39508 9884
rect 4274 9772 4284 9828
rect 4340 9772 6860 9828
rect 6916 9772 6926 9828
rect 18834 9772 18844 9828
rect 18900 9772 20076 9828
rect 20132 9772 20142 9828
rect 22418 9772 22428 9828
rect 22484 9772 23660 9828
rect 23716 9772 25564 9828
rect 25620 9772 25630 9828
rect 26898 9772 26908 9828
rect 26964 9772 27356 9828
rect 27412 9772 27422 9828
rect 34682 9772 34692 9828
rect 34748 9772 35980 9828
rect 36036 9772 39228 9828
rect 39284 9772 39294 9828
rect 39442 9772 39452 9828
rect 39508 9772 39518 9828
rect 39946 9772 39956 9828
rect 40012 9772 41020 9828
rect 41076 9772 41086 9828
rect 41458 9772 41468 9828
rect 41524 9772 41692 9828
rect 41748 9772 41758 9828
rect 42914 9772 42924 9828
rect 42980 9772 47572 9828
rect 47628 9772 47638 9828
rect 4386 9660 4396 9716
rect 4452 9660 5964 9716
rect 6020 9660 6030 9716
rect 6738 9660 6748 9716
rect 6804 9660 8652 9716
rect 8708 9660 8988 9716
rect 9044 9660 9054 9716
rect 22530 9660 22540 9716
rect 22596 9660 23548 9716
rect 23604 9660 24444 9716
rect 24500 9660 24510 9716
rect 24668 9604 24724 9772
rect 41468 9716 41524 9772
rect 26506 9660 26516 9716
rect 26572 9660 32620 9716
rect 32676 9660 32686 9716
rect 38994 9660 39004 9716
rect 39060 9660 41524 9716
rect 43698 9660 43708 9716
rect 43764 9660 44716 9716
rect 44772 9660 44782 9716
rect 4834 9548 4844 9604
rect 4900 9548 5628 9604
rect 5684 9548 5694 9604
rect 15250 9548 15260 9604
rect 15316 9548 16044 9604
rect 16100 9548 16380 9604
rect 16436 9548 22316 9604
rect 22372 9548 22988 9604
rect 23044 9548 23054 9604
rect 24210 9548 24220 9604
rect 24276 9548 24724 9604
rect 25778 9548 25788 9604
rect 25844 9548 26012 9604
rect 26068 9548 26078 9604
rect 26236 9548 28252 9604
rect 28308 9548 33684 9604
rect 33740 9548 33750 9604
rect 26236 9492 26292 9548
rect 11834 9436 11844 9492
rect 11900 9436 13468 9492
rect 13524 9436 13534 9492
rect 17658 9436 17668 9492
rect 17724 9436 18172 9492
rect 18228 9436 18238 9492
rect 25218 9436 25228 9492
rect 25284 9436 26292 9492
rect 26954 9436 26964 9492
rect 27020 9436 44940 9492
rect 44996 9436 45006 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 13346 9324 13356 9380
rect 13412 9324 14476 9380
rect 14532 9324 14756 9380
rect 14812 9324 14822 9380
rect 27234 9324 27244 9380
rect 27300 9324 30492 9380
rect 30548 9324 30558 9380
rect 33842 9324 33852 9380
rect 33908 9324 40460 9380
rect 40516 9324 40526 9380
rect 12898 9212 12908 9268
rect 12964 9212 13468 9268
rect 13524 9212 15036 9268
rect 15092 9212 15102 9268
rect 24490 9212 24500 9268
rect 24556 9212 25340 9268
rect 25396 9212 25406 9268
rect 40282 9212 40292 9268
rect 40348 9212 42028 9268
rect 42084 9212 42094 9268
rect 46834 9212 46844 9268
rect 46900 9212 47124 9268
rect 47180 9212 47190 9268
rect 16258 9100 16268 9156
rect 16324 9100 16772 9156
rect 16828 9100 35868 9156
rect 35924 9100 36484 9156
rect 36540 9100 37156 9156
rect 37212 9100 37222 9156
rect 39442 9100 39452 9156
rect 39508 9100 39900 9156
rect 39956 9100 41132 9156
rect 41188 9100 41198 9156
rect 5282 8988 5292 9044
rect 5348 8988 5628 9044
rect 5684 8988 5694 9044
rect 11442 8988 11452 9044
rect 11508 8988 11676 9044
rect 11732 8988 11742 9044
rect 25666 8988 25676 9044
rect 25732 8988 26628 9044
rect 26684 8988 29932 9044
rect 29988 8988 29998 9044
rect 34962 8988 34972 9044
rect 35028 8988 35532 9044
rect 35588 8988 35598 9044
rect 40450 8988 40460 9044
rect 40516 8988 45276 9044
rect 45332 8988 45342 9044
rect 45602 8988 45612 9044
rect 45668 8988 46620 9044
rect 46676 8988 47292 9044
rect 47348 8988 47358 9044
rect 3546 8876 3556 8932
rect 3612 8876 4900 8932
rect 4956 8876 4966 8932
rect 5842 8876 5852 8932
rect 5908 8876 6860 8932
rect 6916 8876 6926 8932
rect 7298 8876 7308 8932
rect 7364 8876 8428 8932
rect 8484 8876 8494 8932
rect 22642 8876 22652 8932
rect 22708 8876 25228 8932
rect 25284 8876 25396 8932
rect 25452 8876 25462 8932
rect 32218 8876 32228 8932
rect 32284 8876 33628 8932
rect 33684 8876 33694 8932
rect 34626 8876 34636 8932
rect 34692 8876 35308 8932
rect 35364 8876 35374 8932
rect 41794 8876 41804 8932
rect 41860 8876 43036 8932
rect 43092 8876 43102 8932
rect 12562 8764 12572 8820
rect 12628 8764 13804 8820
rect 13860 8764 13870 8820
rect 21242 8764 21252 8820
rect 21308 8764 23940 8820
rect 23996 8764 24006 8820
rect 26002 8764 26012 8820
rect 26068 8764 26796 8820
rect 26852 8764 26862 8820
rect 31154 8764 31164 8820
rect 31220 8764 32396 8820
rect 32452 8764 32462 8820
rect 1586 8652 1596 8708
rect 1652 8652 3556 8708
rect 3612 8652 3622 8708
rect 4946 8652 4956 8708
rect 5012 8652 7084 8708
rect 7140 8652 7420 8708
rect 7476 8652 7486 8708
rect 25638 8652 25676 8708
rect 25732 8652 25742 8708
rect 28354 8652 28364 8708
rect 28420 8652 28924 8708
rect 28980 8652 28990 8708
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 14914 8540 14924 8596
rect 14980 8540 14990 8596
rect 23762 8540 23772 8596
rect 23828 8540 26908 8596
rect 30482 8540 30492 8596
rect 30548 8540 30558 8596
rect 44120 8540 44130 8596
rect 44186 8540 46172 8596
rect 46228 8540 46238 8596
rect 14924 8484 14980 8540
rect 3042 8428 3052 8484
rect 3108 8428 5740 8484
rect 5796 8428 5806 8484
rect 14578 8428 14588 8484
rect 14644 8428 15932 8484
rect 15988 8428 16380 8484
rect 16436 8428 16446 8484
rect 18050 8428 18060 8484
rect 18116 8428 19404 8484
rect 19460 8428 19470 8484
rect 20122 8428 20132 8484
rect 20188 8428 21980 8484
rect 22036 8428 22316 8484
rect 22372 8428 22382 8484
rect 24658 8428 24668 8484
rect 24724 8428 25452 8484
rect 25508 8428 26460 8484
rect 26516 8428 26526 8484
rect 0 8372 800 8400
rect 26852 8372 26908 8540
rect 30492 8484 30548 8540
rect 30492 8428 38892 8484
rect 38948 8428 38958 8484
rect 0 8316 980 8372
rect 4162 8316 4172 8372
rect 4228 8316 4238 8372
rect 6066 8316 6076 8372
rect 6132 8316 6860 8372
rect 6916 8316 6926 8372
rect 7298 8316 7308 8372
rect 7364 8316 9380 8372
rect 9762 8316 9772 8372
rect 9828 8316 11004 8372
rect 11060 8316 11070 8372
rect 12170 8316 12180 8372
rect 12236 8316 14700 8372
rect 14756 8316 14766 8372
rect 26674 8316 26684 8372
rect 26740 8316 30940 8372
rect 30996 8316 31006 8372
rect 35298 8316 35308 8372
rect 35364 8316 37548 8372
rect 37604 8316 37614 8372
rect 40786 8316 40796 8372
rect 40852 8316 42364 8372
rect 42420 8316 43820 8372
rect 43876 8316 44716 8372
rect 44772 8316 45108 8372
rect 45164 8316 45174 8372
rect 0 8288 800 8316
rect 924 8148 980 8316
rect 4172 8260 4228 8316
rect 7308 8260 7364 8316
rect 9324 8260 9380 8316
rect 3826 8204 3836 8260
rect 3892 8204 4620 8260
rect 4676 8204 4686 8260
rect 6738 8204 6748 8260
rect 6804 8204 7364 8260
rect 7746 8204 7756 8260
rect 7812 8204 8204 8260
rect 8260 8204 9100 8260
rect 9156 8204 9166 8260
rect 9324 8204 9884 8260
rect 9940 8204 10892 8260
rect 10948 8204 10958 8260
rect 12506 8204 12516 8260
rect 12572 8204 13580 8260
rect 13636 8204 13646 8260
rect 13804 8204 15260 8260
rect 15316 8204 15326 8260
rect 21858 8204 21868 8260
rect 21924 8204 23324 8260
rect 23380 8204 23390 8260
rect 25890 8204 25900 8260
rect 25956 8204 27020 8260
rect 27076 8204 27086 8260
rect 33730 8204 33740 8260
rect 33796 8204 34188 8260
rect 34244 8204 34254 8260
rect 34682 8204 34692 8260
rect 34748 8204 35980 8260
rect 36036 8204 36046 8260
rect 36194 8204 36204 8260
rect 36260 8204 36270 8260
rect 37874 8204 37884 8260
rect 37940 8204 41580 8260
rect 41636 8204 41646 8260
rect 44258 8204 44268 8260
rect 44324 8204 45500 8260
rect 45556 8204 45566 8260
rect 13804 8148 13860 8204
rect 36204 8148 36260 8204
rect 18 8092 28 8148
rect 84 8092 980 8148
rect 12058 8092 12068 8148
rect 12124 8092 13804 8148
rect 13860 8092 13870 8148
rect 14242 8092 14252 8148
rect 14308 8092 18732 8148
rect 18788 8092 20300 8148
rect 20356 8092 20366 8148
rect 26170 8092 26180 8148
rect 26236 8092 26460 8148
rect 26516 8092 26526 8148
rect 36204 8092 39676 8148
rect 39732 8092 39742 8148
rect 43026 8092 43036 8148
rect 43092 8092 43932 8148
rect 43988 8092 43998 8148
rect 44930 8092 44940 8148
rect 44996 8092 48300 8148
rect 48356 8092 48366 8148
rect 16146 7980 16156 8036
rect 16212 7980 18508 8036
rect 18564 7980 18574 8036
rect 26730 7980 26740 8036
rect 26796 7980 27972 8036
rect 28028 7980 28812 8036
rect 28868 7980 28878 8036
rect 29474 7980 29484 8036
rect 29540 7980 30044 8036
rect 30100 7980 30828 8036
rect 30884 7980 30894 8036
rect 32128 7980 32138 8036
rect 32194 7980 33628 8036
rect 33684 7980 34020 8036
rect 34076 7980 34086 8036
rect 34402 7980 34412 8036
rect 34468 7980 36428 8036
rect 36484 7980 36494 8036
rect 38098 7980 38108 8036
rect 38164 7980 38444 8036
rect 38500 7980 39170 8036
rect 39226 7980 40124 8036
rect 40180 7980 40190 8036
rect 43418 7980 43428 8036
rect 43484 7980 43764 8036
rect 43820 7980 43830 8036
rect 37986 7868 37996 7924
rect 38052 7868 39564 7924
rect 39620 7868 42252 7924
rect 42308 7868 42318 7924
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 23314 7756 23324 7812
rect 23380 7756 25340 7812
rect 25396 7756 25676 7812
rect 25732 7756 25742 7812
rect 33394 7756 33404 7812
rect 33460 7756 38892 7812
rect 38948 7756 38958 7812
rect 49200 7700 50000 7728
rect 5170 7644 5180 7700
rect 5236 7644 7532 7700
rect 7588 7644 7598 7700
rect 12786 7644 12796 7700
rect 12852 7644 13524 7700
rect 13850 7644 13860 7700
rect 13916 7644 14812 7700
rect 14868 7644 14878 7700
rect 23090 7644 23100 7700
rect 23156 7644 23772 7700
rect 23828 7644 23838 7700
rect 31350 7644 31388 7700
rect 31444 7644 31454 7700
rect 34906 7644 34916 7700
rect 34972 7644 36988 7700
rect 37044 7644 37436 7700
rect 37492 7644 37502 7700
rect 48290 7644 48300 7700
rect 48356 7644 50000 7700
rect 13468 7588 13524 7644
rect 49200 7616 50000 7644
rect 8306 7532 8316 7588
rect 8372 7532 9548 7588
rect 9604 7532 9614 7588
rect 13458 7532 13468 7588
rect 13524 7532 13580 7588
rect 13636 7532 13646 7588
rect 26898 7532 26908 7588
rect 26964 7532 27692 7588
rect 27748 7532 27758 7588
rect 36194 7532 36204 7588
rect 36260 7532 38780 7588
rect 38836 7532 38846 7588
rect 6962 7420 6972 7476
rect 7028 7420 7644 7476
rect 7700 7420 7710 7476
rect 9650 7420 9660 7476
rect 9716 7420 11116 7476
rect 11172 7420 11182 7476
rect 12786 7420 12796 7476
rect 12852 7420 13692 7476
rect 13748 7420 13758 7476
rect 14130 7420 14140 7476
rect 14196 7420 15036 7476
rect 15092 7420 15102 7476
rect 16930 7420 16940 7476
rect 16996 7420 17948 7476
rect 18004 7420 18014 7476
rect 19170 7420 19180 7476
rect 19236 7420 21980 7476
rect 22036 7420 22046 7476
rect 24098 7420 24108 7476
rect 24164 7420 25900 7476
rect 25956 7420 25966 7476
rect 28802 7420 28812 7476
rect 28868 7420 35420 7476
rect 35476 7420 36316 7476
rect 36372 7420 36382 7476
rect 40338 7420 40348 7476
rect 40404 7420 41580 7476
rect 41636 7420 41646 7476
rect 42242 7420 42252 7476
rect 42308 7420 42924 7476
rect 42980 7420 42990 7476
rect 12674 7308 12684 7364
rect 12740 7308 14028 7364
rect 14084 7308 14094 7364
rect 18050 7308 18060 7364
rect 18116 7308 18322 7364
rect 18378 7308 18388 7364
rect 33394 7308 33404 7364
rect 33460 7308 38220 7364
rect 38276 7308 38556 7364
rect 38612 7308 38622 7364
rect 41682 7308 41692 7364
rect 41748 7308 42588 7364
rect 42644 7308 43148 7364
rect 43204 7308 43214 7364
rect 45042 7308 45052 7364
rect 45108 7308 47516 7364
rect 47572 7308 47582 7364
rect 29586 7196 29596 7252
rect 29652 7196 41020 7252
rect 41076 7196 41086 7252
rect 25666 7084 25676 7140
rect 25732 7084 31276 7140
rect 31332 7084 31342 7140
rect 44930 7084 44940 7140
rect 44996 7084 47068 7140
rect 47124 7084 47134 7140
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 14690 6972 14700 7028
rect 14756 6972 15912 7028
rect 15968 6972 16772 7028
rect 16828 6972 16838 7028
rect 25778 6972 25788 7028
rect 25844 6972 32788 7028
rect 36194 6972 36204 7028
rect 36260 6972 38668 7028
rect 38724 6972 38734 7028
rect 40450 6972 40460 7028
rect 40516 6972 41300 7028
rect 41356 6972 46284 7028
rect 46340 6972 47404 7028
rect 47460 6972 47470 7028
rect 32732 6916 32788 6972
rect 4498 6860 4508 6916
rect 4564 6860 5740 6916
rect 5796 6860 5806 6916
rect 14242 6860 14252 6916
rect 14308 6860 15148 6916
rect 15204 6860 15214 6916
rect 25442 6860 25452 6916
rect 25508 6860 26908 6916
rect 32732 6860 47964 6916
rect 48020 6860 48030 6916
rect 26852 6804 26908 6860
rect 8978 6748 8988 6804
rect 9044 6748 9660 6804
rect 9716 6748 9726 6804
rect 26852 6748 34188 6804
rect 34244 6748 34254 6804
rect 43138 6748 43148 6804
rect 43204 6748 43932 6804
rect 43988 6748 44716 6804
rect 44772 6748 44782 6804
rect 3938 6636 3948 6692
rect 4004 6636 4956 6692
rect 5012 6636 5796 6692
rect 5852 6636 7084 6692
rect 7140 6636 8148 6692
rect 8204 6636 10108 6692
rect 10164 6636 10388 6692
rect 10444 6636 10454 6692
rect 12394 6636 12404 6692
rect 12460 6636 13132 6692
rect 13188 6636 13198 6692
rect 13794 6636 13804 6692
rect 13860 6636 15036 6692
rect 15092 6636 15102 6692
rect 16370 6636 16380 6692
rect 16436 6636 17052 6692
rect 17108 6636 17118 6692
rect 17378 6636 17388 6692
rect 17444 6636 18844 6692
rect 18900 6636 19292 6692
rect 19348 6636 19358 6692
rect 20010 6636 20020 6692
rect 20076 6636 20468 6692
rect 20524 6636 20534 6692
rect 21746 6636 21756 6692
rect 21812 6636 23324 6692
rect 23380 6636 23390 6692
rect 23538 6636 23548 6692
rect 23604 6636 24276 6692
rect 24332 6636 24342 6692
rect 27570 6636 27580 6692
rect 27636 6636 29204 6692
rect 29260 6636 29270 6692
rect 29754 6636 29764 6692
rect 29820 6636 30268 6692
rect 30324 6636 30334 6692
rect 39330 6636 39340 6692
rect 39396 6636 41356 6692
rect 41412 6636 41422 6692
rect 43026 6636 43036 6692
rect 43092 6636 43820 6692
rect 43876 6636 44044 6692
rect 44100 6636 44110 6692
rect 45602 6636 45612 6692
rect 45668 6636 46396 6692
rect 46452 6636 46462 6692
rect 13430 6524 13468 6580
rect 13524 6524 13534 6580
rect 14466 6524 14476 6580
rect 14532 6524 15260 6580
rect 15316 6524 15932 6580
rect 15988 6524 15998 6580
rect 18386 6524 18396 6580
rect 18452 6524 19628 6580
rect 19684 6524 24892 6580
rect 24948 6524 24958 6580
rect 25050 6524 25060 6580
rect 25116 6524 26012 6580
rect 26068 6524 33180 6580
rect 33236 6524 33516 6580
rect 33572 6524 33582 6580
rect 39218 6524 39228 6580
rect 39284 6524 40236 6580
rect 40292 6524 40302 6580
rect 41682 6524 41692 6580
rect 41748 6524 42644 6580
rect 42700 6524 45780 6580
rect 45724 6468 45780 6524
rect 4834 6412 4844 6468
rect 4900 6412 5628 6468
rect 5684 6412 5694 6468
rect 14914 6412 14924 6468
rect 14980 6412 17836 6468
rect 17892 6412 17902 6468
rect 18498 6412 18508 6468
rect 18564 6412 25900 6468
rect 25956 6412 25966 6468
rect 26338 6412 26348 6468
rect 26404 6412 26852 6468
rect 26908 6412 26918 6468
rect 31378 6412 31388 6468
rect 31444 6412 31612 6468
rect 31668 6412 33338 6468
rect 33394 6412 33404 6468
rect 36754 6412 36764 6468
rect 36820 6412 37268 6468
rect 37324 6412 37334 6468
rect 40562 6412 40572 6468
rect 40628 6412 41020 6468
rect 41076 6412 42476 6468
rect 42532 6412 42542 6468
rect 44986 6412 44996 6468
rect 45052 6412 45500 6468
rect 45556 6412 45566 6468
rect 45714 6412 45724 6468
rect 45780 6412 46396 6468
rect 46452 6412 46462 6468
rect 14690 6300 14700 6356
rect 14756 6300 15764 6356
rect 15820 6300 17612 6356
rect 17668 6300 17678 6356
rect 36978 6300 36988 6356
rect 37044 6300 43372 6356
rect 43428 6300 43438 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 28578 6188 28588 6244
rect 28644 6188 29148 6244
rect 29204 6188 42364 6244
rect 42420 6188 42430 6244
rect 45882 6188 45892 6244
rect 45948 6188 47404 6244
rect 47460 6188 47470 6244
rect 7858 6076 7868 6132
rect 7924 6076 9660 6132
rect 9716 6076 9726 6132
rect 10378 6076 10388 6132
rect 10444 6076 11900 6132
rect 11956 6076 12068 6132
rect 12124 6076 12134 6132
rect 25106 6076 25116 6132
rect 25172 6076 25452 6132
rect 25508 6076 25518 6132
rect 27906 6076 27916 6132
rect 27972 6076 27982 6132
rect 32946 6076 32956 6132
rect 33012 6076 33022 6132
rect 34066 6076 34076 6132
rect 34132 6076 35084 6132
rect 35140 6076 35150 6132
rect 37258 6076 37268 6132
rect 37324 6076 38332 6132
rect 38388 6076 38398 6132
rect 39106 6076 39116 6132
rect 39172 6076 39508 6132
rect 10882 5964 10892 6020
rect 10948 5964 12348 6020
rect 12404 5964 12414 6020
rect 12786 5964 12796 6020
rect 12852 5964 13916 6020
rect 13972 5964 13982 6020
rect 13346 5852 13356 5908
rect 13412 5852 13580 5908
rect 13636 5852 15148 5908
rect 15204 5852 15214 5908
rect 15698 5852 15708 5908
rect 15764 5852 16492 5908
rect 16548 5852 18732 5908
rect 18788 5852 18798 5908
rect 20850 5852 20860 5908
rect 20916 5852 22204 5908
rect 22260 5852 22270 5908
rect 22642 5852 22652 5908
rect 22708 5852 23772 5908
rect 23828 5852 23838 5908
rect 24546 5852 24556 5908
rect 24612 5852 25228 5908
rect 25284 5852 25294 5908
rect 25516 5852 25526 5908
rect 25582 5852 26124 5908
rect 26180 5852 26190 5908
rect 7970 5740 7980 5796
rect 8036 5740 8540 5796
rect 8596 5740 8606 5796
rect 16034 5740 16044 5796
rect 16100 5740 16828 5796
rect 16884 5740 18172 5796
rect 18228 5740 18238 5796
rect 24434 5628 24444 5684
rect 24500 5628 25900 5684
rect 25956 5628 25966 5684
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 27916 5460 27972 6076
rect 32956 6020 33012 6076
rect 39452 6020 39508 6076
rect 32498 5964 32508 6020
rect 32564 5964 39004 6020
rect 39060 5964 39070 6020
rect 39442 5964 39452 6020
rect 39508 5964 39518 6020
rect 42466 5964 42476 6020
rect 42532 5964 42542 6020
rect 42476 5908 42532 5964
rect 30762 5852 30772 5908
rect 30828 5852 33740 5908
rect 33796 5852 33806 5908
rect 33954 5852 33964 5908
rect 34020 5852 34030 5908
rect 34738 5852 34748 5908
rect 34804 5852 35196 5908
rect 35252 5852 35262 5908
rect 36194 5852 36204 5908
rect 36260 5852 37100 5908
rect 37156 5852 38556 5908
rect 38612 5852 39116 5908
rect 39172 5852 41804 5908
rect 41860 5852 41870 5908
rect 42130 5852 42140 5908
rect 42196 5852 42812 5908
rect 42868 5852 42878 5908
rect 45800 5852 45810 5908
rect 45866 5852 47292 5908
rect 47348 5852 47358 5908
rect 33964 5796 34020 5852
rect 29586 5740 29596 5796
rect 29652 5740 31724 5796
rect 31780 5740 31790 5796
rect 33740 5740 35868 5796
rect 35924 5740 35934 5796
rect 36642 5740 36652 5796
rect 36708 5740 36876 5796
rect 36932 5740 36942 5796
rect 40170 5740 40180 5796
rect 40236 5740 40572 5796
rect 40628 5740 41580 5796
rect 41636 5740 41646 5796
rect 33740 5572 33796 5740
rect 33898 5628 33908 5684
rect 33964 5628 34972 5684
rect 35028 5628 36204 5684
rect 36260 5628 40908 5684
rect 40964 5628 40974 5684
rect 33730 5516 33740 5572
rect 33796 5516 33806 5572
rect 37650 5516 37660 5572
rect 37716 5516 37726 5572
rect 37986 5516 37996 5572
rect 38052 5516 40292 5572
rect 42018 5516 42028 5572
rect 42084 5516 42924 5572
rect 42980 5516 45388 5572
rect 45444 5516 45454 5572
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 37660 5460 37716 5516
rect 40236 5460 40292 5516
rect 22866 5404 22876 5460
rect 22932 5404 25116 5460
rect 25172 5404 25182 5460
rect 27916 5404 29316 5460
rect 29372 5404 29382 5460
rect 31378 5404 31388 5460
rect 31444 5404 31892 5460
rect 31948 5404 31958 5460
rect 37660 5404 38780 5460
rect 38836 5404 39004 5460
rect 39060 5404 39070 5460
rect 39274 5404 39284 5460
rect 39340 5404 40068 5460
rect 40226 5404 40236 5460
rect 40292 5404 40302 5460
rect 40460 5404 41132 5460
rect 41188 5404 45444 5460
rect 27916 5348 27972 5404
rect 40012 5348 40068 5404
rect 40460 5348 40516 5404
rect 45388 5348 45444 5404
rect 14186 5292 14196 5348
rect 14252 5292 15148 5348
rect 18946 5292 18956 5348
rect 19012 5292 20300 5348
rect 20356 5292 21196 5348
rect 21252 5292 21262 5348
rect 27906 5292 27916 5348
rect 27972 5292 27982 5348
rect 28802 5292 28812 5348
rect 28868 5292 29484 5348
rect 29540 5292 30268 5348
rect 30324 5292 33348 5348
rect 33404 5292 33414 5348
rect 35186 5292 35196 5348
rect 35252 5292 37324 5348
rect 37380 5292 37390 5348
rect 37650 5292 37660 5348
rect 37716 5292 39844 5348
rect 40012 5292 40516 5348
rect 40674 5292 40684 5348
rect 40740 5292 42700 5348
rect 42756 5292 42766 5348
rect 45378 5292 45388 5348
rect 45444 5292 45454 5348
rect 15092 5236 15148 5292
rect 13458 5180 13468 5236
rect 13524 5180 13748 5236
rect 15092 5180 15260 5236
rect 15316 5180 17164 5236
rect 17220 5180 19516 5236
rect 19572 5180 20804 5236
rect 20860 5180 21644 5236
rect 21700 5180 23436 5236
rect 23492 5180 23502 5236
rect 32162 5180 32172 5236
rect 32228 5180 32508 5236
rect 32564 5180 37436 5236
rect 37492 5180 37502 5236
rect 37660 5180 37996 5236
rect 38052 5180 38062 5236
rect 13692 5012 13748 5180
rect 37660 5124 37716 5180
rect 39788 5124 39844 5292
rect 40786 5180 40796 5236
rect 40852 5180 43820 5236
rect 43876 5180 44716 5236
rect 44772 5180 44782 5236
rect 45938 5180 45948 5236
rect 46004 5180 47516 5236
rect 47572 5180 47582 5236
rect 17938 5068 17948 5124
rect 18004 5068 18900 5124
rect 18956 5068 18966 5124
rect 19058 5068 19068 5124
rect 19124 5068 19292 5124
rect 19348 5068 20188 5124
rect 20244 5068 20254 5124
rect 23090 5068 23100 5124
rect 23156 5068 24444 5124
rect 24500 5068 24510 5124
rect 26450 5068 26460 5124
rect 26516 5068 28812 5124
rect 28868 5068 28878 5124
rect 32050 5068 32060 5124
rect 32116 5068 32126 5124
rect 33170 5068 33180 5124
rect 33236 5068 33246 5124
rect 34626 5068 34636 5124
rect 34692 5068 35532 5124
rect 35588 5068 35598 5124
rect 35746 5068 35756 5124
rect 35812 5068 36484 5124
rect 36540 5068 36764 5124
rect 36820 5068 36830 5124
rect 37314 5068 37324 5124
rect 37380 5068 37716 5124
rect 37818 5068 37828 5124
rect 37884 5068 38668 5124
rect 38724 5068 39452 5124
rect 39508 5068 39518 5124
rect 39778 5068 39788 5124
rect 39844 5068 41020 5124
rect 41076 5068 41086 5124
rect 41682 5068 41692 5124
rect 41748 5068 42364 5124
rect 42420 5068 42430 5124
rect 43362 5068 43372 5124
rect 43428 5068 43932 5124
rect 43988 5068 44940 5124
rect 44996 5068 45006 5124
rect 32060 5012 32116 5068
rect 33180 5012 33236 5068
rect 12674 4956 12684 5012
rect 12740 4956 13468 5012
rect 13524 4956 13534 5012
rect 13692 4956 14588 5012
rect 14644 4956 15372 5012
rect 15428 4956 15438 5012
rect 18274 4956 18284 5012
rect 18340 4956 20020 5012
rect 20076 4956 21924 5012
rect 23202 4956 23212 5012
rect 23268 4956 26012 5012
rect 26068 4956 26078 5012
rect 31714 4956 31724 5012
rect 31780 4956 33236 5012
rect 39106 4956 39116 5012
rect 39172 4956 40348 5012
rect 40404 4956 40414 5012
rect 42466 4956 42476 5012
rect 42532 4956 43148 5012
rect 43204 4956 43214 5012
rect 21868 4900 21924 4956
rect 21858 4844 21868 4900
rect 21924 4844 21934 4900
rect 23986 4844 23996 4900
rect 24052 4844 25900 4900
rect 25956 4844 25966 4900
rect 26852 4844 28252 4900
rect 28308 4844 32732 4900
rect 32788 4844 32798 4900
rect 26852 4788 26908 4844
rect 13794 4732 13804 4788
rect 13860 4732 14476 4788
rect 14532 4732 14542 4788
rect 26226 4732 26236 4788
rect 26292 4732 26908 4788
rect 32386 4732 32396 4788
rect 32452 4732 33628 4788
rect 33684 4732 33694 4788
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 33954 4508 33964 4564
rect 34020 4508 34748 4564
rect 34804 4508 34814 4564
rect 16034 4396 16044 4452
rect 16100 4396 17444 4452
rect 17500 4396 17510 4452
rect 21970 4396 21980 4452
rect 22036 4396 23156 4452
rect 23212 4396 23222 4452
rect 24210 4396 24220 4452
rect 24276 4396 25228 4452
rect 25284 4396 25294 4452
rect 28690 4396 28700 4452
rect 28756 4396 29484 4452
rect 29540 4396 40684 4452
rect 40740 4396 40750 4452
rect 41402 4396 41412 4452
rect 41468 4396 43708 4452
rect 43764 4396 43774 4452
rect 15026 4284 15036 4340
rect 15092 4284 17276 4340
rect 17332 4284 17342 4340
rect 21858 4284 21868 4340
rect 21924 4284 22316 4340
rect 22372 4284 22652 4340
rect 22708 4284 22718 4340
rect 24322 4284 24332 4340
rect 24388 4284 25564 4340
rect 25620 4284 25630 4340
rect 38770 4284 38780 4340
rect 38836 4284 39900 4340
rect 39956 4284 39966 4340
rect 24332 4228 24388 4284
rect 19058 4172 19068 4228
rect 19124 4172 20300 4228
rect 20356 4172 24388 4228
rect 41346 4172 41356 4228
rect 41412 4172 43484 4228
rect 43540 4172 43550 4228
rect 21970 4060 21980 4116
rect 22036 4060 22764 4116
rect 22820 4060 26348 4116
rect 26404 4060 26414 4116
rect 34076 4060 38164 4116
rect 34076 4004 34132 4060
rect 38108 4004 38164 4060
rect 12562 3948 12572 4004
rect 12628 3948 13356 4004
rect 13412 3948 13422 4004
rect 22866 3948 22876 4004
rect 22932 3948 23772 4004
rect 23828 3948 34076 4004
rect 34132 3948 34142 4004
rect 38098 3948 38108 4004
rect 38164 3948 38174 4004
rect 38612 3948 46060 4004
rect 46116 3948 46126 4004
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 25452 3892 25508 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 38612 3892 38668 3948
rect 18722 3836 18732 3892
rect 18788 3836 23436 3892
rect 23492 3836 23996 3892
rect 24052 3836 24062 3892
rect 25442 3836 25452 3892
rect 25508 3836 25518 3892
rect 31490 3836 31500 3892
rect 31556 3836 32396 3892
rect 32452 3836 32462 3892
rect 36866 3836 36876 3892
rect 36932 3836 38668 3892
rect 40842 3836 40852 3892
rect 40908 3836 41468 3892
rect 41524 3836 42588 3892
rect 42644 3836 45052 3892
rect 45108 3836 45118 3892
rect 13346 3724 13356 3780
rect 13412 3724 16044 3780
rect 16100 3724 22428 3780
rect 22484 3724 22494 3780
rect 26338 3724 26348 3780
rect 26404 3724 30772 3780
rect 30828 3724 32228 3780
rect 32778 3724 32788 3780
rect 32844 3724 35980 3780
rect 36036 3724 40236 3780
rect 40292 3724 44044 3780
rect 44100 3724 47460 3780
rect 47516 3724 47526 3780
rect 14466 3612 14476 3668
rect 14532 3612 17836 3668
rect 17892 3612 18396 3668
rect 18452 3612 18462 3668
rect 19506 3612 19516 3668
rect 19572 3612 22540 3668
rect 22596 3612 22764 3668
rect 22820 3612 22830 3668
rect 24098 3612 24108 3668
rect 24164 3612 24836 3668
rect 24892 3612 26236 3668
rect 26292 3612 26302 3668
rect 32172 3556 32228 3724
rect 32330 3612 32340 3668
rect 32396 3612 33236 3668
rect 33292 3612 33302 3668
rect 36362 3612 36372 3668
rect 36428 3612 36652 3668
rect 36708 3612 39956 3668
rect 40012 3612 42700 3668
rect 42756 3612 43092 3668
rect 43148 3612 45332 3668
rect 45388 3612 46676 3668
rect 46732 3612 47572 3668
rect 47628 3612 48020 3668
rect 48076 3612 48300 3668
rect 48356 3612 48366 3668
rect 16258 3500 16268 3556
rect 16324 3500 17556 3556
rect 17612 3500 17622 3556
rect 17948 3500 18732 3556
rect 18788 3500 18798 3556
rect 19170 3500 19180 3556
rect 19236 3500 21532 3556
rect 21588 3500 21598 3556
rect 25162 3500 25172 3556
rect 25228 3500 26012 3556
rect 26068 3500 26078 3556
rect 32172 3500 33628 3556
rect 33684 3500 36764 3556
rect 36820 3500 36830 3556
rect 37090 3500 37100 3556
rect 37156 3500 40292 3556
rect 40348 3500 40358 3556
rect 40674 3500 40684 3556
rect 40740 3500 41692 3556
rect 41748 3500 42476 3556
rect 42532 3500 42542 3556
rect 43698 3500 43708 3556
rect 43764 3500 46228 3556
rect 46284 3500 46294 3556
rect 17948 3444 18004 3500
rect 12618 3388 12628 3444
rect 12684 3388 18004 3444
rect 18162 3388 18172 3444
rect 18228 3388 19628 3444
rect 19684 3388 21084 3444
rect 21140 3388 21150 3444
rect 37736 3388 37746 3444
rect 37802 3388 39788 3444
rect 39844 3388 39854 3444
rect 19618 3276 19628 3332
rect 19684 3276 19796 3332
rect 19852 3276 19862 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 49200 2772 50000 2800
rect 28914 2716 28924 2772
rect 28980 2716 50000 2772
rect 49200 2688 50000 2716
<< via3 >>
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 36428 45500 36484 45556
rect 37884 45500 37940 45556
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 19628 44940 19684 44996
rect 37324 44940 37380 44996
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 36428 44268 36484 44324
rect 37436 44156 37492 44212
rect 30716 44044 30772 44100
rect 6412 43708 6468 43764
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 14924 43820 14980 43876
rect 30716 43708 30772 43764
rect 30380 43260 30436 43316
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 6412 43036 6468 43092
rect 14924 43036 14980 43092
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 35644 42812 35700 42868
rect 31948 42588 32004 42644
rect 37548 42588 37604 42644
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 31948 42140 32004 42196
rect 37548 42140 37604 42196
rect 26572 42028 26628 42084
rect 35980 42028 36036 42084
rect 10332 41916 10388 41972
rect 36652 41916 36708 41972
rect 37324 41916 37380 41972
rect 6860 41692 6916 41748
rect 12012 41580 12068 41636
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 45388 41692 45444 41748
rect 15148 41580 15204 41636
rect 35644 41580 35700 41636
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 29708 41468 29764 41524
rect 36204 41468 36260 41524
rect 19628 41356 19684 41412
rect 46060 41244 46116 41300
rect 37324 41132 37380 41188
rect 38780 41132 38836 41188
rect 44828 41132 44884 41188
rect 11676 41020 11732 41076
rect 12012 41020 12068 41076
rect 37436 41020 37492 41076
rect 42364 40908 42420 40964
rect 45836 40908 45892 40964
rect 46060 40908 46116 40964
rect 46396 40796 46452 40852
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 11676 40684 11732 40740
rect 29820 40684 29876 40740
rect 6860 40572 6916 40628
rect 8204 40572 8260 40628
rect 15148 40572 15204 40628
rect 34972 40572 35028 40628
rect 42364 40572 42420 40628
rect 43596 40572 43652 40628
rect 44940 40572 44996 40628
rect 46284 40572 46340 40628
rect 43372 40460 43428 40516
rect 46396 40460 46452 40516
rect 46732 40460 46788 40516
rect 29708 40348 29764 40404
rect 39228 40348 39284 40404
rect 44604 40348 44660 40404
rect 38780 40236 38836 40292
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 44940 39900 44996 39956
rect 36876 39788 36932 39844
rect 37996 39788 38052 39844
rect 36540 39452 36596 39508
rect 10556 39340 10612 39396
rect 36540 39228 36596 39284
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 36764 39116 36820 39172
rect 21308 39004 21364 39060
rect 30492 38892 30548 38948
rect 37884 38892 37940 38948
rect 39228 38892 39284 38948
rect 46508 38892 46564 38948
rect 28252 38780 28308 38836
rect 36876 38780 36932 38836
rect 8428 38668 8484 38724
rect 26684 38668 26740 38724
rect 30380 38668 30436 38724
rect 37996 38668 38052 38724
rect 45836 38668 45892 38724
rect 29820 38556 29876 38612
rect 34972 38556 35028 38612
rect 35980 38556 36036 38612
rect 43372 38556 43428 38612
rect 43596 38556 43652 38612
rect 44604 38556 44660 38612
rect 46508 38556 46564 38612
rect 30492 38444 30548 38500
rect 31052 38444 31108 38500
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 26572 38332 26628 38388
rect 20524 38220 20580 38276
rect 36988 37996 37044 38052
rect 46732 37772 46788 37828
rect 10332 37660 10388 37716
rect 20188 37660 20244 37716
rect 20412 37660 20468 37716
rect 31052 37660 31108 37716
rect 44828 37660 44884 37716
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 13356 37548 13412 37604
rect 26460 37548 26516 37604
rect 36764 37548 36820 37604
rect 20188 37436 20244 37492
rect 13356 37324 13412 37380
rect 36652 37436 36708 37492
rect 10556 37100 10612 37156
rect 21308 37100 21364 37156
rect 45836 37100 45892 37156
rect 8764 36988 8820 37044
rect 37996 36988 38052 37044
rect 8316 36876 8372 36932
rect 8652 36876 8708 36932
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 20188 36764 20244 36820
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 8204 36428 8260 36484
rect 45500 36428 45556 36484
rect 36988 36092 37044 36148
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 11116 35756 11172 35812
rect 45388 35756 45444 35812
rect 20188 35644 20244 35700
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 28252 35644 28308 35700
rect 45500 35532 45556 35588
rect 11116 35196 11172 35252
rect 13916 35196 13972 35252
rect 16268 35196 16324 35252
rect 20524 35196 20580 35252
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 25564 35084 25620 35140
rect 21532 34860 21588 34916
rect 20300 34748 20356 34804
rect 26460 34748 26516 34804
rect 8652 34524 8708 34580
rect 36540 34972 36596 35028
rect 46284 34972 46340 35028
rect 20412 34524 20468 34580
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 20524 34412 20580 34468
rect 23996 34412 24052 34468
rect 36204 34412 36260 34468
rect 23772 34300 23828 34356
rect 38892 34300 38948 34356
rect 26572 34188 26628 34244
rect 10108 33964 10164 34020
rect 20300 33964 20356 34020
rect 45724 33964 45780 34020
rect 21532 33852 21588 33908
rect 10780 33740 10836 33796
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 30156 33740 30212 33796
rect 32172 33740 32228 33796
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 26460 33628 26516 33684
rect 29708 33628 29764 33684
rect 31052 33628 31108 33684
rect 20300 33404 20356 33460
rect 36540 33404 36596 33460
rect 38108 33404 38164 33460
rect 23100 32956 23156 33012
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 23772 32844 23828 32900
rect 27916 32620 27972 32676
rect 38892 32508 38948 32564
rect 38220 32172 38276 32228
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 12124 31836 12180 31892
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 45836 32060 45892 32116
rect 26684 31948 26740 32004
rect 28028 31948 28084 32004
rect 27020 31724 27076 31780
rect 28140 31724 28176 31780
rect 28176 31724 28196 31780
rect 27916 31612 27972 31668
rect 12124 31500 12180 31556
rect 14252 31500 14308 31556
rect 10108 31388 10164 31444
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 20636 31276 20692 31332
rect 13244 31164 13300 31220
rect 27020 31164 27076 31220
rect 28252 31052 28308 31108
rect 25676 30940 25732 30996
rect 38892 30940 38948 30996
rect 28028 30716 28084 30772
rect 30492 30716 30548 30772
rect 20636 30604 20692 30660
rect 25788 30604 25844 30660
rect 28140 30604 28196 30660
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 10780 30492 10836 30548
rect 8540 30380 8596 30436
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 28252 30380 28308 30436
rect 29708 30380 29764 30436
rect 38892 30268 38948 30324
rect 9324 30044 9380 30100
rect 38220 30044 38276 30100
rect 45724 30044 45780 30100
rect 14252 29932 14308 29988
rect 30156 29932 30212 29988
rect 25788 29820 25844 29876
rect 26348 29820 26404 29876
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 34076 29708 34132 29764
rect 23996 29596 24052 29652
rect 34524 29596 34580 29652
rect 20188 29372 20244 29428
rect 25676 29372 25732 29428
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 26348 29148 26404 29204
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 9324 28812 9380 28868
rect 23100 28812 23156 28868
rect 29708 28812 29764 28868
rect 30156 28812 30212 28868
rect 25564 28588 25620 28644
rect 26572 28476 26628 28532
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 25676 28140 25732 28196
rect 35756 28140 35812 28196
rect 20188 28028 20244 28084
rect 12908 27804 12964 27860
rect 12124 27580 12180 27636
rect 14140 27580 14196 27636
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 38332 27692 38388 27748
rect 20524 27468 20580 27524
rect 35644 27468 35700 27524
rect 13020 27356 13076 27412
rect 13916 27020 13972 27076
rect 14140 27020 14196 27076
rect 14812 27020 14868 27076
rect 8764 26908 8820 26964
rect 13020 26908 13076 26964
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 35756 27244 35812 27300
rect 38332 27132 38388 27188
rect 14812 26684 14868 26740
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 34076 26684 34132 26740
rect 34524 26684 34580 26740
rect 32172 26572 32228 26628
rect 8540 26460 8596 26516
rect 35644 26460 35700 26516
rect 33068 26236 33124 26292
rect 13244 26124 13300 26180
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 30492 25788 30548 25844
rect 31052 25564 31108 25620
rect 30492 25340 30548 25396
rect 31052 25228 31108 25284
rect 33068 25116 33124 25172
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 30492 24892 30548 24948
rect 12124 24780 12180 24836
rect 16268 24780 16324 24836
rect 30492 24556 30548 24612
rect 43260 24444 43316 24500
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 38108 24108 38164 24164
rect 12908 23884 12964 23940
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 18284 23324 18340 23380
rect 32060 23324 32116 23380
rect 29372 23212 29428 23268
rect 32284 23100 32340 23156
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 25340 22316 25396 22372
rect 32060 22316 32116 22372
rect 32284 22316 32340 22372
rect 43260 22204 43316 22260
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 17836 21644 17892 21700
rect 17836 21308 17892 21364
rect 18284 21308 18340 21364
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 6636 20524 6692 20580
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 24780 20300 24836 20356
rect 25452 20300 25508 20356
rect 6636 19740 6692 19796
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 46844 19180 46900 19236
rect 24780 18956 24836 19012
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 19068 18732 19124 18788
rect 26460 18732 26516 18788
rect 39676 18172 39732 18228
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 26460 17948 26516 18004
rect 43596 17948 43652 18004
rect 43596 17724 43652 17780
rect 25340 17388 25396 17444
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 29708 16828 29764 16884
rect 19068 16604 19124 16660
rect 26460 16604 26516 16660
rect 39676 16604 39732 16660
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 22316 16268 22372 16324
rect 25452 16044 25508 16100
rect 44268 16044 44324 16100
rect 26684 15820 26740 15876
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 26348 15596 26404 15652
rect 25900 15148 25956 15204
rect 29708 15148 29764 15204
rect 12348 14924 12404 14980
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 25788 14924 25844 14980
rect 26348 14924 26404 14980
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 29372 14812 29428 14868
rect 45164 14588 45220 14644
rect 12348 14476 12404 14532
rect 29372 14364 29428 14420
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 25452 14028 25508 14084
rect 25788 14028 25844 14084
rect 26684 14028 26740 14084
rect 26908 14028 26964 14084
rect 14476 13916 14532 13972
rect 23100 13356 23156 13412
rect 25452 13356 25508 13412
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 37212 12908 37268 12964
rect 45164 13244 45220 13300
rect 14476 12572 14532 12628
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 37548 12348 37604 12404
rect 44268 12236 44324 12292
rect 37548 11900 37604 11956
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 25900 11676 25956 11732
rect 37212 11340 37268 11396
rect 23100 11228 23156 11284
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 26908 10108 26964 10164
rect 22316 9548 22372 9604
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 13468 9212 13524 9268
rect 46844 9212 46900 9268
rect 25676 8652 25732 8708
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 25676 7756 25732 7812
rect 31388 7644 31444 7700
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 25788 6972 25844 7028
rect 13468 6524 13524 6580
rect 31388 6412 31444 6468
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19628 3388 19684 3444
rect 19628 3276 19684 3332
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 46284 4768 46316
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 19808 45500 20128 46316
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 19628 44996 19684 45006
rect 14924 43876 14980 43886
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 6412 43764 6468 43774
rect 6412 43092 6468 43708
rect 6412 43026 6468 43036
rect 14924 43092 14980 43820
rect 14924 43026 14980 43036
rect 10332 41972 10388 41982
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 6860 41748 6916 41758
rect 6860 40628 6916 41692
rect 6860 40562 6916 40572
rect 8204 40628 8260 40638
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 8204 36484 8260 40572
rect 8428 38724 8484 38734
rect 8428 37018 8484 38668
rect 10332 37716 10388 41916
rect 12012 41636 12068 41646
rect 11676 41076 11732 41086
rect 11676 40740 11732 41020
rect 12012 41076 12068 41580
rect 12012 41010 12068 41020
rect 15148 41636 15204 41646
rect 11676 40674 11732 40684
rect 15148 40628 15204 41580
rect 19628 41412 19684 44940
rect 19628 41346 19684 41356
rect 19808 43932 20128 45444
rect 35168 46284 35488 46316
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 30716 44100 30772 44110
rect 30716 43764 30772 44044
rect 30716 43698 30772 43708
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 15148 40562 15204 40572
rect 19808 40796 20128 42308
rect 30380 43316 30436 43326
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 10332 37650 10388 37660
rect 10556 39396 10612 39406
rect 10556 37156 10612 39340
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 26572 42084 26628 42094
rect 21308 39060 21364 39070
rect 20524 38276 20580 38286
rect 13356 37604 13412 37614
rect 13356 37380 13412 37548
rect 13356 37314 13412 37324
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 10556 37090 10612 37100
rect 8316 36962 8484 37018
rect 8764 37044 8820 37054
rect 8316 36932 8372 36962
rect 8316 36866 8372 36876
rect 8652 36932 8708 36942
rect 8204 36418 8260 36428
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 8652 34580 8708 36876
rect 8652 34514 8708 34524
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 8540 30436 8596 30446
rect 8540 26516 8596 30380
rect 8764 26964 8820 36988
rect 19808 36092 20128 37604
rect 20188 37716 20244 37726
rect 20188 37492 20244 37660
rect 20188 36820 20244 37436
rect 20188 36754 20244 36764
rect 20412 37716 20468 37726
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 11116 35812 11172 35822
rect 11116 35252 11172 35756
rect 11116 35186 11172 35196
rect 13916 35252 13972 35262
rect 10108 34020 10164 34030
rect 10108 31444 10164 33964
rect 10108 31378 10164 31388
rect 10780 33796 10836 33806
rect 10780 30548 10836 33740
rect 12124 31892 12180 31902
rect 12124 31556 12180 31836
rect 12124 31490 12180 31500
rect 10780 30482 10836 30492
rect 13244 31220 13300 31230
rect 9324 30100 9380 30110
rect 9324 28868 9380 30044
rect 9324 28802 9380 28812
rect 12908 27860 12964 27870
rect 8764 26898 8820 26908
rect 12124 27636 12180 27646
rect 8540 26450 8596 26460
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 12124 24836 12180 27580
rect 12124 24770 12180 24780
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 12908 23940 12964 27804
rect 13020 27412 13076 27422
rect 13020 26964 13076 27356
rect 13020 26898 13076 26908
rect 13244 26180 13300 31164
rect 13916 27076 13972 35196
rect 16268 35252 16324 35262
rect 14252 31556 14308 31566
rect 14252 29988 14308 31500
rect 14252 29922 14308 29932
rect 13916 27010 13972 27020
rect 14140 27636 14196 27646
rect 14140 27076 14196 27580
rect 14140 27010 14196 27020
rect 14812 27076 14868 27086
rect 14812 26740 14868 27020
rect 14812 26674 14868 26684
rect 13244 26114 13300 26124
rect 16268 24836 16324 35196
rect 16268 24770 16324 24780
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 20188 35700 20244 35710
rect 20188 29428 20244 35644
rect 20300 34804 20356 34814
rect 20300 34020 20356 34748
rect 20412 34580 20468 37660
rect 20524 35252 20580 38220
rect 21308 37156 21364 39004
rect 26572 38388 26628 42028
rect 29708 41524 29764 41534
rect 29708 40404 29764 41468
rect 29708 40338 29764 40348
rect 29820 40740 29876 40750
rect 28252 38836 28308 38846
rect 26572 38322 26628 38332
rect 26684 38724 26740 38734
rect 21308 37090 21364 37100
rect 26460 37604 26516 37614
rect 20524 35186 20580 35196
rect 25564 35140 25620 35150
rect 20412 34514 20468 34524
rect 21532 34916 21588 34926
rect 20300 33460 20356 33964
rect 20300 33394 20356 33404
rect 20524 34468 20580 34478
rect 20188 28084 20244 29372
rect 20188 28018 20244 28028
rect 20524 27524 20580 34412
rect 21532 33908 21588 34860
rect 23996 34468 24052 34478
rect 21532 33842 21588 33852
rect 23772 34356 23828 34366
rect 23100 33012 23156 33022
rect 20636 31332 20692 31342
rect 20636 30660 20692 31276
rect 20636 30594 20692 30604
rect 23100 28868 23156 32956
rect 23772 32900 23828 34300
rect 23772 32834 23828 32844
rect 23996 29652 24052 34412
rect 23996 29586 24052 29596
rect 23100 28802 23156 28812
rect 25564 28644 25620 35084
rect 26460 34804 26516 37548
rect 26460 33684 26516 34748
rect 26460 33618 26516 33628
rect 26572 34244 26628 34254
rect 25564 28578 25620 28588
rect 25676 30996 25732 31006
rect 25676 29428 25732 30940
rect 25788 30660 25844 30670
rect 25788 29876 25844 30604
rect 25788 29810 25844 29820
rect 26348 29876 26404 29886
rect 25676 28196 25732 29372
rect 26348 29204 26404 29820
rect 26348 29138 26404 29148
rect 26572 28532 26628 34188
rect 26684 32004 26740 38668
rect 28252 35700 28308 38780
rect 29820 38612 29876 40684
rect 30380 38724 30436 43260
rect 35168 43148 35488 44660
rect 36428 45556 36484 45566
rect 36428 44324 36484 45500
rect 37884 45556 37940 45566
rect 36428 44258 36484 44268
rect 37324 44996 37380 45006
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 31948 42644 32004 42654
rect 31948 42196 32004 42588
rect 31948 42130 32004 42140
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35644 42868 35700 42878
rect 35644 41636 35700 42812
rect 35644 41570 35700 41580
rect 35980 42084 36036 42094
rect 34972 40628 35028 40638
rect 30380 38658 30436 38668
rect 30492 38948 30548 38958
rect 29820 38546 29876 38556
rect 30492 38500 30548 38892
rect 34972 38612 35028 40572
rect 34972 38546 35028 38556
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 30492 38434 30548 38444
rect 31052 38500 31108 38510
rect 28252 35634 28308 35644
rect 31052 37716 31108 38444
rect 30156 33796 30212 33806
rect 29708 33684 29764 33694
rect 26684 31938 26740 31948
rect 27916 32676 27972 32686
rect 27020 31780 27076 31790
rect 27020 31220 27076 31724
rect 27916 31668 27972 32620
rect 27916 31602 27972 31612
rect 28028 32004 28084 32014
rect 27020 31154 27076 31164
rect 28028 30772 28084 31948
rect 28028 30706 28084 30716
rect 28140 31780 28196 31790
rect 28140 30660 28196 31724
rect 28140 30594 28196 30604
rect 28252 31108 28308 31118
rect 28252 30436 28308 31052
rect 28252 30370 28308 30380
rect 29708 30436 29764 33628
rect 29708 30370 29764 30380
rect 30156 29988 30212 33740
rect 31052 33684 31108 37660
rect 35168 38444 35488 39956
rect 35980 38612 36036 42028
rect 36652 41972 36708 41982
rect 35980 38546 36036 38556
rect 36204 41524 36260 41534
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 31052 33618 31108 33628
rect 32172 33796 32228 33806
rect 30156 29922 30212 29932
rect 30492 30772 30548 30782
rect 29708 28868 30212 28918
rect 29764 28862 30156 28868
rect 29708 28802 29764 28812
rect 30156 28802 30212 28812
rect 26572 28466 26628 28476
rect 25676 28130 25732 28140
rect 20524 27458 20580 27468
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 30492 25844 30548 30716
rect 32172 26628 32228 33740
rect 35168 33740 35488 35252
rect 36204 34468 36260 41468
rect 36540 39508 36596 39518
rect 36540 39284 36596 39452
rect 36540 39218 36596 39228
rect 36652 37492 36708 41916
rect 37324 41972 37380 44940
rect 37324 41188 37380 41916
rect 37324 41122 37380 41132
rect 37436 44212 37492 44222
rect 37436 41076 37492 44156
rect 37548 42644 37604 42654
rect 37548 42196 37604 42588
rect 37548 42130 37604 42140
rect 37436 41010 37492 41020
rect 36876 39844 36932 39854
rect 36764 39172 36820 39182
rect 36764 37604 36820 39116
rect 36876 38836 36932 39788
rect 37884 38948 37940 45500
rect 45388 41748 45444 41758
rect 38780 41188 38836 41198
rect 38780 40292 38836 41132
rect 44828 41188 44884 41198
rect 42364 40964 42420 40974
rect 42364 40628 42420 40908
rect 42364 40562 42420 40572
rect 43596 40628 43652 40638
rect 43372 40516 43428 40526
rect 38780 40226 38836 40236
rect 39228 40404 39284 40414
rect 37884 38882 37940 38892
rect 37996 39844 38052 39854
rect 36876 38770 36932 38780
rect 37996 38724 38052 39788
rect 39228 38948 39284 40348
rect 39228 38882 39284 38892
rect 36764 37538 36820 37548
rect 36988 38052 37044 38062
rect 36652 37426 36708 37436
rect 36988 36148 37044 37996
rect 37996 37044 38052 38668
rect 43372 38612 43428 40460
rect 43372 38546 43428 38556
rect 43596 38612 43652 40572
rect 43596 38546 43652 38556
rect 44604 40404 44660 40414
rect 44604 38612 44660 40348
rect 44604 38546 44660 38556
rect 44828 37716 44884 41132
rect 44940 40628 44996 40638
rect 44940 39956 44996 40572
rect 44940 39890 44996 39900
rect 44828 37650 44884 37660
rect 37996 36978 38052 36988
rect 36988 36082 37044 36092
rect 45388 35812 45444 41692
rect 46060 41300 46116 41310
rect 45836 40964 45892 40974
rect 45836 38724 45892 40908
rect 46060 40964 46116 41244
rect 46060 40898 46116 40908
rect 46396 40852 46452 40862
rect 45836 38658 45892 38668
rect 46284 40628 46340 40638
rect 45836 37156 45892 37166
rect 45388 35746 45444 35756
rect 45500 36484 45556 36494
rect 45500 35588 45556 36428
rect 45500 35522 45556 35532
rect 36204 34402 36260 34412
rect 36540 35028 36596 35038
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 36540 33460 36596 34972
rect 38892 34356 38948 34366
rect 36540 33394 36596 33404
rect 38108 33460 38164 33470
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 34076 29764 34132 29774
rect 34076 26740 34132 29708
rect 34076 26674 34132 26684
rect 34524 29652 34580 29662
rect 34524 26740 34580 29596
rect 34524 26674 34580 26684
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35756 28196 35812 28206
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 32172 26562 32228 26572
rect 30492 25778 30548 25788
rect 33068 26292 33124 26302
rect 31052 25620 31108 25630
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 12908 23874 12964 23884
rect 19808 23548 20128 25060
rect 30492 25396 30548 25406
rect 30492 24948 30548 25340
rect 31052 25284 31108 25564
rect 31052 25218 31108 25228
rect 33068 25172 33124 26236
rect 33068 25106 33124 25116
rect 35168 25900 35488 27412
rect 35644 27524 35700 27534
rect 35644 26516 35700 27468
rect 35756 27300 35812 28140
rect 35756 27234 35812 27244
rect 35644 26450 35700 26460
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 30492 24612 30548 24892
rect 30492 24546 30548 24556
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 18284 23380 18340 23390
rect 17836 21700 17892 21710
rect 17836 21364 17892 21644
rect 17836 21298 17892 21308
rect 18284 21364 18340 23324
rect 18284 21298 18340 21308
rect 19808 21980 20128 23492
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 32060 23380 32116 23390
rect 29372 23268 29428 23278
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 6636 20580 6692 20590
rect 6636 19796 6692 20524
rect 6636 19730 6692 19740
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 25340 22372 25396 22382
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 19808 18844 20128 20356
rect 24780 20356 24836 20366
rect 24780 19012 24836 20300
rect 24780 18946 24836 18956
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 19068 18788 19124 18798
rect 19068 16660 19124 18732
rect 19068 16594 19124 16604
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 25340 17444 25396 22316
rect 25340 17378 25396 17388
rect 25452 20356 25508 20366
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 12348 14980 12404 14990
rect 12348 14532 12404 14924
rect 12348 14466 12404 14476
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 14476 13972 14532 13982
rect 14476 12628 14532 13916
rect 14476 12562 14532 12572
rect 19808 12572 20128 14084
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 22316 16324 22372 16334
rect 22316 9604 22372 16268
rect 25452 16100 25508 20300
rect 26460 18788 26516 18798
rect 26460 18004 26516 18732
rect 26460 16660 26516 17948
rect 26460 16594 26516 16604
rect 25452 16034 25508 16044
rect 26684 15876 26740 15886
rect 26348 15652 26404 15662
rect 25900 15204 25956 15214
rect 25788 14980 25844 14990
rect 25452 14084 25508 14094
rect 23100 13412 23156 13422
rect 23100 11284 23156 13356
rect 25452 13412 25508 14028
rect 25452 13346 25508 13356
rect 25788 14084 25844 14924
rect 23100 11218 23156 11228
rect 22316 9538 22372 9548
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 13468 9268 13524 9278
rect 13468 6580 13524 9212
rect 13468 6514 13524 6524
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 6300 20128 7812
rect 25676 8708 25732 8718
rect 25676 7812 25732 8652
rect 25676 7746 25732 7756
rect 25788 7028 25844 14028
rect 25900 11732 25956 15148
rect 26348 14980 26404 15596
rect 26348 14914 26404 14924
rect 26684 14084 26740 15820
rect 29372 14868 29428 23212
rect 32060 22372 32116 23324
rect 32060 22306 32116 22316
rect 32284 23156 32340 23166
rect 32284 22372 32340 23100
rect 32284 22306 32340 22316
rect 35168 22764 35488 24276
rect 38108 24164 38164 33404
rect 38892 32564 38948 34300
rect 38220 32228 38276 32238
rect 38220 30100 38276 32172
rect 38892 30996 38948 32508
rect 38892 30324 38948 30940
rect 38892 30258 38948 30268
rect 45724 34020 45780 34030
rect 38220 30034 38276 30044
rect 45724 30100 45780 33964
rect 45836 32116 45892 37100
rect 46284 35028 46340 40572
rect 46396 40516 46452 40796
rect 46396 40450 46452 40460
rect 46732 40516 46788 40526
rect 46508 38948 46564 38958
rect 46508 38612 46564 38892
rect 46508 38546 46564 38556
rect 46732 37828 46788 40460
rect 46732 37762 46788 37772
rect 46284 34962 46340 34972
rect 45836 32050 45892 32060
rect 45724 30034 45780 30044
rect 38332 27748 38388 27758
rect 38332 27188 38388 27692
rect 38332 27122 38388 27132
rect 38108 24098 38164 24108
rect 43260 24500 43316 24510
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 43260 22260 43316 24444
rect 43260 22194 43316 22204
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 46844 19236 46900 19246
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 29708 16884 29764 16894
rect 29708 15204 29764 16828
rect 29708 15138 29764 15148
rect 35168 16492 35488 18004
rect 39676 18228 39732 18238
rect 39676 16660 39732 18172
rect 43596 18004 43652 18014
rect 43596 17780 43652 17948
rect 43596 17714 43652 17724
rect 39676 16594 39732 16604
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 29372 14420 29428 14812
rect 29372 14354 29428 14364
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 26684 14018 26740 14028
rect 26908 14084 26964 14094
rect 25900 11666 25956 11676
rect 26908 10164 26964 14028
rect 26908 10098 26964 10108
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 44268 16100 44324 16110
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 37212 12964 37268 12974
rect 37212 11396 37268 12908
rect 37548 12404 37604 12414
rect 37548 11956 37604 12348
rect 44268 12292 44324 16044
rect 45164 14644 45220 14654
rect 45164 13300 45220 14588
rect 45164 13234 45220 13244
rect 44268 12226 44324 12236
rect 37548 11890 37604 11900
rect 37212 11330 37268 11340
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 46844 9268 46900 19180
rect 46844 9202 46900 9212
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 25788 6962 25844 6972
rect 31388 7700 31444 7710
rect 31388 6468 31444 7644
rect 31388 6402 31444 6412
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19628 3444 19684 3454
rect 19628 3332 19684 3388
rect 19628 3266 19684 3276
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1446_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751534193
transform -1 0 26208 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _1447_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1752061876
transform -1 0 29568 0 -1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1448_
timestamp 1751534193
transform -1 0 26880 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1449_
timestamp 1751534193
transform -1 0 34384 0 1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _1450_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751905124
transform 1 0 25984 0 1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1451_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753371985
transform 1 0 25536 0 -1 25088
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1452_
timestamp 1751534193
transform -1 0 28784 0 1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1453_
timestamp 1751534193
transform 1 0 29008 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1454_
timestamp 1751534193
transform 1 0 37184 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _1455_
timestamp 1751905124
transform 1 0 29568 0 1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1456_
timestamp 1751534193
transform -1 0 30912 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _1457_
timestamp 1751905124
transform -1 0 30128 0 1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _1458_
timestamp 1751905124
transform 1 0 27888 0 -1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1459_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751531619
transform -1 0 29792 0 -1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1460_
timestamp 1751531619
transform -1 0 31024 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1461_
timestamp 1751531619
transform -1 0 32368 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1462_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751740063
transform -1 0 29456 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1463_
timestamp 1751534193
transform -1 0 23744 0 -1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1464_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753868718
transform 1 0 29008 0 1 26656
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1465_
timestamp 1751534193
transform -1 0 10080 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _1466_
timestamp 1751905124
transform 1 0 19488 0 1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1467_
timestamp 1751534193
transform 1 0 20944 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1468_
timestamp 1751534193
transform -1 0 22960 0 1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1469_
timestamp 1751534193
transform 1 0 18592 0 1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _1470_
timestamp 1751905124
transform 1 0 17584 0 1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1471_
timestamp 1751534193
transform 1 0 19152 0 -1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1472_
timestamp 1751740063
transform 1 0 17808 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1473_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532043
transform -1 0 21168 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1474_
timestamp 1751531619
transform -1 0 19936 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1475_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751889808
transform 1 0 18592 0 1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1476_
timestamp 1751532043
transform -1 0 19152 0 1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _1477_
timestamp 1751905124
transform -1 0 19152 0 -1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1478_
timestamp 1751531619
transform 1 0 17696 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1479_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753960525
transform 1 0 18480 0 -1 29792
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1480_
timestamp 1751889808
transform -1 0 16800 0 1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_4  _1481_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753864693
transform -1 0 22064 0 -1 32928
box -86 -86 2998 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1482_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753277515
transform 1 0 29120 0 -1 32928
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1483_
timestamp 1751532043
transform 1 0 32256 0 1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1484_
timestamp 1751534193
transform -1 0 11648 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1485_
timestamp 1751534193
transform 1 0 12432 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1486_
timestamp 1751534193
transform 1 0 13328 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _1487_
timestamp 1751905124
transform 1 0 12768 0 -1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1488_
timestamp 1751534193
transform -1 0 13104 0 1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _1489_
timestamp 1752061876
transform -1 0 13552 0 -1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _1490_
timestamp 1751905124
transform 1 0 11648 0 1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1491_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751914308
transform -1 0 13104 0 1 23520
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1492_
timestamp 1751534193
transform 1 0 12656 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _1493_
timestamp 1751905124
transform -1 0 14560 0 -1 25088
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1494_
timestamp 1751534193
transform -1 0 11648 0 1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _1495_
timestamp 1752061876
transform -1 0 12768 0 1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1496_
timestamp 1751531619
transform 1 0 10528 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1497_
timestamp 1751914308
transform -1 0 14672 0 1 25088
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1498_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753441877
transform -1 0 14448 0 1 31360
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1499_
timestamp 1751534193
transform -1 0 5264 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _1500_
timestamp 1752061876
transform -1 0 3024 0 1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1501_
timestamp 1751534193
transform -1 0 2576 0 -1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _1502_
timestamp 1752061876
transform -1 0 7952 0 -1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1503_
timestamp 1751534193
transform -1 0 3248 0 -1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1504_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751889408
transform 1 0 2128 0 1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_4  _1505_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1752051650
transform -1 0 6832 0 -1 21952
box -86 -86 1881 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1506_
timestamp 1751740063
transform 1 0 5488 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1507_
timestamp 1751534193
transform 1 0 5488 0 1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1508_
timestamp 1751534193
transform 1 0 3248 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _1509_
timestamp 1751905124
transform 1 0 2464 0 1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1510_
timestamp 1751914308
transform 1 0 3248 0 -1 25088
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _1511_
timestamp 1751905124
transform 1 0 6944 0 1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_2  _1512_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753579406
transform 1 0 6160 0 1 25088
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1513_
timestamp 1751534193
transform -1 0 7504 0 1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1514_
timestamp 1751534193
transform 1 0 11088 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_2  _1515_
timestamp 1753579406
transform -1 0 12880 0 -1 25088
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _1516_
timestamp 1752061876
transform 1 0 13328 0 1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1517_
timestamp 1753371985
transform 1 0 12656 0 -1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_4  _1518_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753432499
transform -1 0 13104 0 1 25088
box -86 -86 2214 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1519_
timestamp 1751532043
transform -1 0 10528 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1520_
timestamp 1753868718
transform -1 0 10752 0 -1 28224
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1521_
timestamp 1751532043
transform -1 0 9072 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1522_
timestamp 1751532043
transform 1 0 4592 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1523_
timestamp 1751534193
transform -1 0 7952 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1524_
timestamp 1753960525
transform 1 0 3024 0 1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _1525_
timestamp 1752061876
transform 1 0 4144 0 1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1526_
timestamp 1753371985
transform 1 0 3584 0 1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_4  _1527_
timestamp 1753432499
transform -1 0 7616 0 1 23520
box -86 -86 2214 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1528_
timestamp 1751534193
transform 1 0 5488 0 1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_4  _1529_
timestamp 1753864693
transform 1 0 4592 0 -1 25088
box -86 -86 2998 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _1530_
timestamp 1751905124
transform 1 0 3920 0 -1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1531_
timestamp 1753441877
transform 1 0 6160 0 1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _1532_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1752345181
transform 1 0 6384 0 -1 23520
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _1533_
timestamp 1751905124
transform 1 0 4032 0 1 25088
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1534_
timestamp 1751531619
transform 1 0 4704 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1535_
timestamp 1751531619
transform -1 0 13104 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1536_
timestamp 1751534193
transform -1 0 11200 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1537_
timestamp 1753371985
transform -1 0 11984 0 1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_2  _1538_
timestamp 1753579406
transform 1 0 9296 0 1 26656
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1539_
timestamp 1753441877
transform 1 0 7616 0 -1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__maj3_4  _1540_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753273081
transform 1 0 9072 0 1 29792
box -86 -86 1766 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1541_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753272495
transform 1 0 14112 0 -1 32928
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1542_
timestamp 1751534193
transform -1 0 2464 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1543_
timestamp 1753371985
transform 1 0 2912 0 1 25088
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1544_
timestamp 1751534193
transform 1 0 6608 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1545_
timestamp 1753371985
transform 1 0 4144 0 1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1546_
timestamp 1751914308
transform 1 0 3024 0 -1 26656
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1547_
timestamp 1751889808
transform 1 0 3696 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1548_
timestamp 1751532043
transform 1 0 14784 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1549_
timestamp 1751534193
transform 1 0 15120 0 -1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1550_
timestamp 1753371985
transform 1 0 13776 0 -1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1551_
timestamp 1751534193
transform 1 0 15008 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1552_
timestamp 1753441877
transform 1 0 13888 0 -1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1553_
timestamp 1751531619
transform -1 0 15456 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1554_
timestamp 1753441877
transform -1 0 15232 0 -1 29792
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1555_
timestamp 1751889408
transform 1 0 14896 0 -1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1556_
timestamp 1751889808
transform 1 0 12432 0 -1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _1557_
timestamp 1751905124
transform 1 0 14896 0 1 32928
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1558_
timestamp 1753277515
transform 1 0 29904 0 1 32928
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1559_
timestamp 1753277515
transform 1 0 30576 0 -1 34496
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1560_
timestamp 1751531619
transform 1 0 21504 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1561_
timestamp 1751889808
transform -1 0 20720 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1562_
timestamp 1751889408
transform 1 0 20720 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1563_
timestamp 1751534193
transform -1 0 18032 0 -1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _1564_
timestamp 1752061876
transform 1 0 18816 0 -1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1565_
timestamp 1751534193
transform 1 0 20272 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1566_
timestamp 1753371985
transform 1 0 19824 0 -1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _1567_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753891287
transform 1 0 19376 0 1 29792
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1568_
timestamp 1753441877
transform 1 0 21168 0 1 31360
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1569_
timestamp 1751532043
transform 1 0 25088 0 1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1570_
timestamp 1751532043
transform -1 0 25536 0 -1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _1571_
timestamp 1752061876
transform 1 0 27552 0 1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1572_
timestamp 1751531619
transform 1 0 29008 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1573_
timestamp 1751889408
transform 1 0 29456 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1574_
timestamp 1751534193
transform 1 0 30688 0 1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1575_
timestamp 1751531619
transform 1 0 27776 0 1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1576_
timestamp 1751889808
transform 1 0 29792 0 -1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1577_
timestamp 1751532043
transform 1 0 30912 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_4  _1578_
timestamp 1753864693
transform 1 0 30016 0 1 25088
box -86 -86 2998 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1579_
timestamp 1751531619
transform -1 0 11536 0 1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _1580_
timestamp 1752061876
transform 1 0 10192 0 -1 32928
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1581_
timestamp 1753277515
transform 1 0 13328 0 1 29792
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1582_
timestamp 1753277515
transform 1 0 14000 0 -1 31360
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1583_
timestamp 1753272495
transform 1 0 30128 0 1 31360
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1584_
timestamp 1753277515
transform 1 0 29456 0 -1 31360
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1585_
timestamp 1751532043
transform -1 0 29456 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1586_
timestamp 1753277515
transform 1 0 31024 0 -1 31360
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1587_
timestamp 1751534193
transform 1 0 21616 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1588_
timestamp 1751531619
transform 1 0 20048 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _1589_
timestamp 1752345181
transform 1 0 23408 0 1 28224
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1590_
timestamp 1751889808
transform 1 0 21168 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_4  _1591_
timestamp 1753864693
transform 1 0 21952 0 -1 28224
box -86 -86 2998 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1592_
timestamp 1751534193
transform 1 0 27104 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_2  _1593_
timestamp 1753579406
transform -1 0 28448 0 -1 25088
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1594_
timestamp 1753371985
transform 1 0 23744 0 -1 25088
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1595_
timestamp 1751889408
transform -1 0 28112 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1596_
timestamp 1753960525
transform 1 0 27328 0 -1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1597_
timestamp 1751534193
transform 1 0 30912 0 -1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1598_
timestamp 1751531619
transform 1 0 31360 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1599_
timestamp 1753277515
transform 1 0 8848 0 1 28224
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1600_
timestamp 1753277515
transform 1 0 9408 0 -1 29792
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1601_
timestamp 1753868718
transform 1 0 22400 0 1 26656
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1602_
timestamp 1753277515
transform 1 0 29792 0 1 28224
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1603_
timestamp 1751531619
transform -1 0 31584 0 1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1604_
timestamp 1751531619
transform 1 0 30016 0 1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1605_
timestamp 1751889408
transform 1 0 21168 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1606_
timestamp 1753441877
transform 1 0 19600 0 -1 29792
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1607_
timestamp 1753371985
transform -1 0 22288 0 1 29792
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1608_
timestamp 1751889408
transform 1 0 21280 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_4  _1609_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753960842
transform 1 0 22064 0 -1 29792
box -86 -86 1542 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1610_
timestamp 1751531619
transform -1 0 30464 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1611_
timestamp 1751531619
transform 1 0 24080 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1612_
timestamp 1751889408
transform 1 0 26320 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _1613_
timestamp 1752345181
transform -1 0 29680 0 -1 28224
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1614_
timestamp 1751531619
transform -1 0 29792 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1615_
timestamp 1751889408
transform -1 0 6048 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1616_
timestamp 1753868718
transform -1 0 11648 0 1 28224
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1617_
timestamp 1753277515
transform 1 0 7280 0 1 28224
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1618_
timestamp 1753272495
transform 1 0 33152 0 -1 28224
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1619_
timestamp 1753277515
transform 1 0 30688 0 -1 29792
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _1620_
timestamp 1752061876
transform -1 0 34384 0 1 29792
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1621_
timestamp 1753272495
transform 1 0 31920 0 1 29792
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1622_
timestamp 1753272495
transform 1 0 31696 0 1 34496
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1623_
timestamp 1751740063
transform 1 0 21168 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_4  _1624_
timestamp 1753960842
transform 1 0 21952 0 1 28224
box -86 -86 1542 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1625_
timestamp 1751889808
transform 1 0 29008 0 1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1626_
timestamp 1751889408
transform 1 0 29008 0 1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1627_
timestamp 1753277515
transform 1 0 27104 0 -1 34496
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1628_
timestamp 1751534193
transform 1 0 7280 0 1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1629_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753182340
transform -1 0 6384 0 -1 23520
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1630_
timestamp 1753960525
transform 1 0 7616 0 -1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1631_
timestamp 1751532043
transform -1 0 9184 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1632_
timestamp 1751889408
transform 1 0 11648 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao22_4  _1633_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753869255
transform 1 0 10752 0 -1 28224
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1634_
timestamp 1751532043
transform -1 0 6160 0 -1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1635_
timestamp 1753277515
transform 1 0 8288 0 1 36064
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1636_
timestamp 1751889808
transform 1 0 12320 0 1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1637_
timestamp 1753960525
transform 1 0 13776 0 -1 34496
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1638_
timestamp 1753277515
transform 1 0 13888 0 1 34496
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1639_
timestamp 1753277515
transform 1 0 29008 0 1 34496
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1640_
timestamp 1751531619
transform -1 0 31472 0 -1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1641_
timestamp 1751889808
transform 1 0 31472 0 1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1642_
timestamp 1751889408
transform 1 0 29120 0 1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1643_
timestamp 1753960525
transform 1 0 29456 0 -1 34496
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1644_
timestamp 1753277515
transform 1 0 30576 0 -1 36064
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1645_
timestamp 1751531619
transform 1 0 33712 0 1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1646_
timestamp 1751889808
transform 1 0 34048 0 -1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1647_
timestamp 1751889408
transform 1 0 34496 0 -1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1648_
timestamp 1751534193
transform 1 0 34944 0 1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _1649_
timestamp 1752061876
transform -1 0 34048 0 -1 36064
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1650_
timestamp 1753441877
transform -1 0 33712 0 1 36064
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1651_
timestamp 1751889408
transform -1 0 27104 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1652_
timestamp 1753277515
transform 1 0 25312 0 1 28224
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1653_
timestamp 1751534193
transform 1 0 22960 0 1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _1654_
timestamp 1752345181
transform -1 0 20272 0 1 32928
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1655_
timestamp 1753277515
transform -1 0 20944 0 1 34496
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1656_
timestamp 1753277515
transform 1 0 27776 0 -1 36064
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1657_
timestamp 1751531619
transform 1 0 8736 0 1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1658_
timestamp 1751889408
transform 1 0 9408 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1659_
timestamp 1753277515
transform 1 0 9072 0 1 25088
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1660_
timestamp 1751889408
transform 1 0 11200 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1661_
timestamp 1751531619
transform -1 0 15456 0 1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1662_
timestamp 1753277515
transform -1 0 13104 0 1 29792
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1663_
timestamp 1753277515
transform 1 0 10864 0 -1 36064
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1664_
timestamp 1751534193
transform 1 0 9408 0 -1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _1665_
timestamp 1753891287
transform -1 0 14896 0 1 32928
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1666_
timestamp 1753272495
transform 1 0 11760 0 1 34496
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1667_
timestamp 1753277515
transform 1 0 12432 0 -1 36064
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1668_
timestamp 1753277515
transform 1 0 29120 0 1 36064
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1669_
timestamp 1751531619
transform -1 0 28448 0 1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1670_
timestamp 1753272495
transform 1 0 27440 0 1 34496
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1671_
timestamp 1753277515
transform 1 0 30912 0 -1 37632
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1672_
timestamp 1753277515
transform 1 0 32928 0 -1 37632
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1673_
timestamp 1751534193
transform 1 0 35280 0 -1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1674_
timestamp 1753272495
transform 1 0 31248 0 1 36064
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1675_
timestamp 1751532043
transform 1 0 32592 0 1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1676_
timestamp 1751532043
transform -1 0 21616 0 1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1677_
timestamp 1751889408
transform -1 0 19376 0 1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1678_
timestamp 1753960525
transform 1 0 21728 0 -1 34496
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1679_
timestamp 1751531619
transform 1 0 27888 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_2  _1680_
timestamp 1753579406
transform 1 0 27328 0 -1 29792
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1681_
timestamp 1753277515
transform 1 0 27104 0 -1 37632
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1682_
timestamp 1753441877
transform 1 0 7616 0 1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1683_
timestamp 1751532043
transform 1 0 9408 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1684_
timestamp 1753371985
transform 1 0 7728 0 -1 25088
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1685_
timestamp 1753960525
transform 1 0 7952 0 1 25088
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1686_
timestamp 1751531619
transform -1 0 15680 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1687_
timestamp 1753371985
transform -1 0 14672 0 1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1688_
timestamp 1753960525
transform -1 0 14784 0 1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1689_
timestamp 1751531619
transform 1 0 11536 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1690_
timestamp 1751889808
transform -1 0 14112 0 1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1691_
timestamp 1751531619
transform 1 0 14000 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1692_
timestamp 1751531619
transform -1 0 14112 0 1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1693_
timestamp 1751534193
transform -1 0 8512 0 -1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1694_
timestamp 1751534193
transform -1 0 10080 0 -1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_2  _1695_
timestamp 1753579406
transform -1 0 12880 0 1 36064
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1696_
timestamp 1751740063
transform 1 0 11536 0 -1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1697_
timestamp 1753371985
transform -1 0 14224 0 -1 37632
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1698_
timestamp 1753277515
transform 1 0 14784 0 1 37632
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1699_
timestamp 1753277515
transform 1 0 29008 0 1 37632
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1700_
timestamp 1753272495
transform 1 0 27440 0 1 36064
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1701_
timestamp 1753277515
transform 1 0 30576 0 1 37632
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1702_
timestamp 1753277515
transform 1 0 32928 0 -1 39200
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1703_
timestamp 1751534193
transform 1 0 35616 0 1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1704_
timestamp 1751531619
transform -1 0 22288 0 1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1705_
timestamp 1753868718
transform 1 0 20496 0 -1 34496
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1706_
timestamp 1751531619
transform -1 0 27104 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1707_
timestamp 1751889408
transform -1 0 24080 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_2  _1708_
timestamp 1753579406
transform -1 0 26320 0 1 26656
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1709_
timestamp 1753277515
transform 1 0 26096 0 1 39200
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1710_
timestamp 1751532043
transform 1 0 29008 0 1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1711_
timestamp 1751889408
transform -1 0 8848 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_4  _1712_
timestamp 1753864693
transform -1 0 9184 0 -1 26656
box -86 -86 2998 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_4  _1713_
timestamp 1753864693
transform 1 0 11200 0 -1 29792
box -86 -86 2998 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1714_
timestamp 1751740063
transform 1 0 10752 0 -1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1715_
timestamp 1751531619
transform 1 0 12656 0 -1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _1716_
timestamp 1751905124
transform 1 0 12656 0 -1 39200
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1717_
timestamp 1751532043
transform 1 0 14448 0 -1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1718_
timestamp 1753371985
transform 1 0 14112 0 -1 39200
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1719_
timestamp 1753277515
transform 1 0 14112 0 1 39200
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1720_
timestamp 1753277515
transform 1 0 27888 0 -1 39200
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1721_
timestamp 1753868718
transform 1 0 28896 0 -1 29792
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1722_
timestamp 1753272495
transform 1 0 27440 0 1 37632
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1723_
timestamp 1753277515
transform 1 0 29568 0 1 39200
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1724_
timestamp 1751532043
transform 1 0 32144 0 1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1725_
timestamp 1753272495
transform -1 0 32480 0 -1 39200
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1726_
timestamp 1751531619
transform 1 0 32256 0 1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1727_
timestamp 1751889808
transform 1 0 33040 0 1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1728_
timestamp 1751889408
transform 1 0 37296 0 -1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1729_
timestamp 1751534193
transform -1 0 36624 0 1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _1730_
timestamp 1752061876
transform 1 0 29792 0 -1 39200
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1731_
timestamp 1753371985
transform -1 0 32256 0 1 39200
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1732_
timestamp 1751531619
transform 1 0 20160 0 1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1733_
timestamp 1751889408
transform -1 0 28672 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1734_
timestamp 1753277515
transform 1 0 26432 0 1 40768
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1735_
timestamp 1751889808
transform 1 0 12320 0 -1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1736_
timestamp 1751531619
transform 1 0 12320 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1737_
timestamp 1753960525
transform 1 0 11984 0 1 39200
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _1738_
timestamp 1752061876
transform 1 0 5488 0 1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1739_
timestamp 1751889408
transform 1 0 15232 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1740_
timestamp 1753277515
transform 1 0 12880 0 -1 42336
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1741_
timestamp 1753277515
transform 1 0 13440 0 -1 40768
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1742_
timestamp 1753277515
transform 1 0 27664 0 -1 40768
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1743_
timestamp 1753868718
transform 1 0 25088 0 -1 26656
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1744_
timestamp 1751531619
transform 1 0 26656 0 -1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1745_
timestamp 1751889808
transform 1 0 28000 0 1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1746_
timestamp 1751531619
transform 1 0 29008 0 -1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1747_
timestamp 1753277515
transform 1 0 29680 0 1 40768
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1748_
timestamp 1753277515
transform 1 0 31248 0 1 40768
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1749_
timestamp 1751534193
transform 1 0 40768 0 -1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1750_
timestamp 1751889408
transform 1 0 31248 0 -1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1751_
timestamp 1753272495
transform 1 0 29904 0 -1 40768
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1752_
timestamp 1751740063
transform 1 0 20048 0 -1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1753_
timestamp 1751532043
transform 1 0 22288 0 1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1754_
timestamp 1751740063
transform 1 0 25536 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1755_
timestamp 1753277515
transform 1 0 25760 0 -1 43904
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1756_
timestamp 1751740063
transform -1 0 9744 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1757_
timestamp 1751740063
transform -1 0 12768 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1758_
timestamp 1753277515
transform 1 0 10864 0 -1 43904
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1759_
timestamp 1753272495
transform 1 0 13328 0 1 40768
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1760_
timestamp 1753277515
transform 1 0 12432 0 -1 43904
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1761_
timestamp 1753277515
transform 1 0 27216 0 1 42336
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1762_
timestamp 1751889408
transform 1 0 20384 0 -1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1763_
timestamp 1753272495
transform 1 0 27552 0 -1 42336
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1764_
timestamp 1753277515
transform 1 0 29792 0 1 42336
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1765_
timestamp 1753277515
transform 1 0 30800 0 -1 42336
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1766_
timestamp 1751534193
transform -1 0 32704 0 -1 40768
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1767_
timestamp 1751532043
transform 1 0 32256 0 1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1768_
timestamp 1753272495
transform 1 0 30240 0 -1 43904
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1769_
timestamp 1751534193
transform 1 0 27328 0 -1 43904
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1770_
timestamp 1753272495
transform 1 0 28000 0 -1 43904
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1771_
timestamp 1751534193
transform 1 0 10192 0 -1 43904
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1772_
timestamp 1751534193
transform 1 0 11760 0 1 43904
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1773_
timestamp 1753272495
transform 1 0 14000 0 -1 43904
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1774_
timestamp 1753277515
transform -1 0 31808 0 1 43904
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1775_
timestamp 1751740063
transform 1 0 31472 0 1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1776_
timestamp 1751889408
transform -1 0 30240 0 -1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_4  _1777_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751882821
transform 1 0 32928 0 -1 43904
box -86 -86 1542 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1778_
timestamp 1753441877
transform 1 0 31584 0 -1 43904
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1779_
timestamp 1751534193
transform 1 0 34384 0 -1 43904
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1780_
timestamp 1751534193
transform 1 0 37856 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1781_
timestamp 1751534193
transform 1 0 39312 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1782_
timestamp 1751534193
transform 1 0 38640 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1783_
timestamp 1751889408
transform -1 0 46256 0 1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1784_
timestamp 1751740063
transform -1 0 44800 0 -1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1785_
timestamp 1751534193
transform -1 0 43792 0 -1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1786_
timestamp 1751534193
transform 1 0 44688 0 1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1787_
timestamp 1751889408
transform 1 0 42896 0 1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1788_
timestamp 1751534193
transform 1 0 43680 0 1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1789_
timestamp 1751534193
transform 1 0 37968 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1790_
timestamp 1751534193
transform 1 0 38528 0 -1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1791_
timestamp 1751531619
transform 1 0 42896 0 1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1792_
timestamp 1751531619
transform 1 0 43680 0 1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1793_
timestamp 1751740063
transform 1 0 47264 0 -1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1794_
timestamp 1751889408
transform 1 0 47600 0 1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1795_
timestamp 1753182340
transform 1 0 46032 0 -1 36064
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1796_
timestamp 1751534193
transform -1 0 45360 0 1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1797_
timestamp 1751740063
transform -1 0 48160 0 -1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1798_
timestamp 1751889408
transform -1 0 47600 0 1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1799_
timestamp 1753182340
transform -1 0 47376 0 -1 34496
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1800_
timestamp 1751534193
transform -1 0 45360 0 1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1801_
timestamp 1753277515
transform 1 0 45472 0 -1 32928
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1802_
timestamp 1751740063
transform -1 0 47040 0 1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1803_
timestamp 1753371985
transform 1 0 47040 0 -1 32928
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1804_
timestamp 1751740063
transform 1 0 47040 0 1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1805_
timestamp 1751532043
transform 1 0 23520 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1806_
timestamp 1751532043
transform -1 0 21616 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1807_
timestamp 1751740063
transform 1 0 17472 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1808_
timestamp 1751889408
transform 1 0 23968 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1809_
timestamp 1751534193
transform 1 0 25424 0 1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1810_
timestamp 1751534193
transform -1 0 28112 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1811_
timestamp 1751534193
transform 1 0 22736 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1812_
timestamp 1751740063
transform -1 0 25872 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1813_
timestamp 1751534193
transform 1 0 26208 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1814_
timestamp 1751531619
transform -1 0 26320 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1815_
timestamp 1751534193
transform 1 0 26320 0 -1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1816_
timestamp 1751534193
transform 1 0 25088 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1817_
timestamp 1751532043
transform -1 0 21616 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1818_
timestamp 1751534193
transform 1 0 20048 0 1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1819_
timestamp 1751534193
transform 1 0 21168 0 1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1820_
timestamp 1753960525
transform 1 0 24192 0 1 10976
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1821_
timestamp 1753441877
transform 1 0 25088 0 -1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1822_
timestamp 1751534193
transform -1 0 24192 0 -1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1823_
timestamp 1751532043
transform -1 0 24528 0 1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1824_
timestamp 1751532043
transform -1 0 23968 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1825_
timestamp 1751534193
transform -1 0 24416 0 -1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1826_
timestamp 1751534193
transform -1 0 24864 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1827_
timestamp 1751534193
transform 1 0 25648 0 -1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1828_
timestamp 1751534193
transform -1 0 17024 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1829_
timestamp 1751534193
transform 1 0 22288 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1830_
timestamp 1751534193
transform -1 0 23520 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1831_
timestamp 1753960525
transform 1 0 23072 0 1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1832_
timestamp 1753371985
transform 1 0 22960 0 1 6272
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1833_
timestamp 1751532043
transform 1 0 21168 0 1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1834_
timestamp 1751532043
transform 1 0 26880 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1835_
timestamp 1751534193
transform 1 0 23408 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1836_
timestamp 1753960525
transform -1 0 23072 0 1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1837_
timestamp 1753371985
transform 1 0 21392 0 1 6272
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1838_
timestamp 1751532043
transform 1 0 21952 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1839_
timestamp 1751532043
transform -1 0 26208 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1840_
timestamp 1751534193
transform 1 0 24976 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1841_
timestamp 1751534193
transform 1 0 24192 0 1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1842_
timestamp 1753960525
transform -1 0 24864 0 -1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1843_
timestamp 1753371985
transform -1 0 22288 0 1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1844_
timestamp 1751532043
transform 1 0 25648 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1845_
timestamp 1751889408
transform 1 0 26096 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1846_
timestamp 1751534193
transform 1 0 26320 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1847_
timestamp 1751531619
transform 1 0 26544 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1848_
timestamp 1753960525
transform 1 0 26208 0 -1 10976
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1849_
timestamp 1753441877
transform 1 0 27104 0 1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1850_
timestamp 1751534193
transform 1 0 28112 0 1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1851_
timestamp 1751532043
transform -1 0 29456 0 1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1852_
timestamp 1751534193
transform 1 0 26880 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1853_
timestamp 1753960525
transform 1 0 26432 0 1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1854_
timestamp 1753371985
transform -1 0 28224 0 1 6272
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1855_
timestamp 1751532043
transform -1 0 28672 0 1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1856_
timestamp 1753960525
transform 1 0 26320 0 -1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1857_
timestamp 1753371985
transform -1 0 27888 0 1 4704
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1858_
timestamp 1751532043
transform -1 0 28672 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1859_
timestamp 1753960525
transform 1 0 25312 0 1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1860_
timestamp 1753371985
transform -1 0 28000 0 1 3136
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1861_
timestamp 1751534193
transform 1 0 23968 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1862_
timestamp 1751889408
transform 1 0 25200 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1863_
timestamp 1751534193
transform -1 0 27664 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1864_
timestamp 1751531619
transform 1 0 30128 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1865_
timestamp 1751534193
transform -1 0 26544 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1866_
timestamp 1753960525
transform 1 0 26320 0 1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1867_
timestamp 1753441877
transform -1 0 36288 0 1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1868_
timestamp 1751534193
transform -1 0 35280 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1869_
timestamp 1751532043
transform -1 0 37296 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1870_
timestamp 1751534193
transform 1 0 27552 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1871_
timestamp 1751534193
transform 1 0 30128 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1872_
timestamp 1753960525
transform 1 0 31248 0 -1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1873_
timestamp 1753371985
transform -1 0 37072 0 -1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1874_
timestamp 1751532043
transform -1 0 34496 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1875_
timestamp 1753960525
transform 1 0 28784 0 -1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1876_
timestamp 1753371985
transform -1 0 34048 0 -1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1877_
timestamp 1751532043
transform -1 0 28784 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1878_
timestamp 1753960525
transform 1 0 29344 0 1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1879_
timestamp 1753371985
transform -1 0 34608 0 1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1880_
timestamp 1751534193
transform 1 0 31808 0 1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1881_
timestamp 1751534193
transform 1 0 39872 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1882_
timestamp 1751740063
transform -1 0 33040 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1883_
timestamp 1751889408
transform 1 0 32928 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1884_
timestamp 1753182340
transform -1 0 32256 0 1 20384
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1885_
timestamp 1751534193
transform -1 0 31024 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1886_
timestamp 1751889808
transform -1 0 32144 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1887_
timestamp 1751531619
transform -1 0 33712 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1888_
timestamp 1753371985
transform 1 0 30240 0 1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1889_
timestamp 1751534193
transform 1 0 23296 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1890_
timestamp 1751534193
transform -1 0 23856 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1891_
timestamp 1753960525
transform 1 0 31136 0 -1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1892_
timestamp 1751740063
transform 1 0 32144 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1893_
timestamp 1753868718
transform 1 0 30352 0 -1 25088
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1894_
timestamp 1753277515
transform 1 0 32928 0 1 25088
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1895_
timestamp 1753272495
transform 1 0 32928 0 -1 23520
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1896_
timestamp 1751889808
transform 1 0 34160 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1897_
timestamp 1751534193
transform -1 0 17920 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1898_
timestamp 1751534193
transform 1 0 16352 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1899_
timestamp 1751534193
transform 1 0 26880 0 -1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1900_
timestamp 1753371985
transform 1 0 34496 0 1 25088
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1901_
timestamp 1751889408
transform 1 0 35616 0 1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1902_
timestamp 1751534193
transform 1 0 36848 0 1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1903_
timestamp 1751532043
transform -1 0 31696 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1904_
timestamp 1753277515
transform 1 0 31696 0 1 26656
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1905_
timestamp 1753272495
transform 1 0 32928 0 -1 26656
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1906_
timestamp 1751889808
transform 1 0 34496 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1907_
timestamp 1753371985
transform 1 0 34608 0 1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1908_
timestamp 1751889408
transform 1 0 35728 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1909_
timestamp 1751534193
transform -1 0 35952 0 -1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1910_
timestamp 1753277515
transform 1 0 27104 0 1 31360
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1911_
timestamp 1753272495
transform -1 0 34608 0 1 26656
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1912_
timestamp 1751889808
transform 1 0 29008 0 1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1913_
timestamp 1753371985
transform -1 0 28672 0 -1 31360
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1914_
timestamp 1751889408
transform -1 0 29120 0 -1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1915_
timestamp 1751534193
transform -1 0 27104 0 1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1916_
timestamp 1753272495
transform -1 0 28448 0 1 32928
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1917_
timestamp 1751532043
transform -1 0 24416 0 1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1918_
timestamp 1753277515
transform 1 0 24416 0 1 34496
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1919_
timestamp 1751534193
transform -1 0 40768 0 1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_4  _1920_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751558652
transform 1 0 22624 0 -1 9408
box -86 -86 1094 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1921_
timestamp 1751889808
transform -1 0 27104 0 -1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1922_
timestamp 1751531619
transform 1 0 25536 0 -1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1923_
timestamp 1753371985
transform -1 0 27104 0 1 34496
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1924_
timestamp 1753277515
transform 1 0 25872 0 1 36064
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1925_
timestamp 1753272495
transform 1 0 25088 0 -1 36064
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1926_
timestamp 1751889808
transform -1 0 26544 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1927_
timestamp 1751534193
transform -1 0 16352 0 1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1928_
timestamp 1753371985
transform -1 0 27552 0 -1 36064
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1929_
timestamp 1751889408
transform 1 0 26544 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1930_
timestamp 1751534193
transform -1 0 24304 0 -1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1931_
timestamp 1751534193
transform 1 0 22960 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1932_
timestamp 1751534193
transform -1 0 23632 0 1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1933_
timestamp 1751534193
transform -1 0 16016 0 -1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1934_
timestamp 1753277515
transform 1 0 25088 0 -1 39200
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1935_
timestamp 1753272495
transform -1 0 26768 0 -1 37632
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1936_
timestamp 1751740063
transform -1 0 26096 0 1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1937_
timestamp 1751889408
transform 1 0 26432 0 -1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1938_
timestamp 1753182340
transform 1 0 23632 0 -1 39200
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1939_
timestamp 1751534193
transform -1 0 24304 0 -1 40768
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1940_
timestamp 1751532043
transform -1 0 25536 0 -1 43904
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1941_
timestamp 1753277515
transform 1 0 25088 0 -1 42336
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1942_
timestamp 1753441877
transform 1 0 25312 0 -1 40768
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1943_
timestamp 1751740063
transform -1 0 25312 0 1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1944_
timestamp 1751889408
transform 1 0 26656 0 -1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1945_
timestamp 1753182340
transform 1 0 23632 0 -1 42336
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1946_
timestamp 1751534193
transform 1 0 24192 0 -1 43904
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1947_
timestamp 1751889808
transform 1 0 29008 0 1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1948_
timestamp 1751531619
transform 1 0 28224 0 1 45472
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1949_
timestamp 1751889408
transform -1 0 29792 0 1 45472
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1950_
timestamp 1753441877
transform 1 0 25760 0 1 42336
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1951_
timestamp 1751889808
transform -1 0 27328 0 1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1952_
timestamp 1753371985
transform -1 0 26544 0 1 43904
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1953_
timestamp 1751889408
transform -1 0 26432 0 1 45472
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1954_
timestamp 1751534193
transform 1 0 26432 0 1 45472
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1955_
timestamp 1753441877
transform -1 0 29344 0 -1 45472
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1956_
timestamp 1751889408
transform -1 0 30576 0 1 45472
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1957_
timestamp 1751889408
transform -1 0 28784 0 1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1958_
timestamp 1751534193
transform -1 0 25424 0 1 43904
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1959_
timestamp 1751532043
transform 1 0 4704 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1960_
timestamp 1751740063
transform -1 0 6384 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1961_
timestamp 1753960525
transform -1 0 7168 0 -1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1962_
timestamp 1751740063
transform -1 0 3360 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1963_
timestamp 1753277515
transform 1 0 3584 0 -1 29792
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1964_
timestamp 1751889808
transform 1 0 4480 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1965_
timestamp 1751531619
transform -1 0 7168 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1966_
timestamp 1753371985
transform 1 0 5488 0 1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1967_
timestamp 1753277515
transform 1 0 3360 0 1 29792
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1968_
timestamp 1751532043
transform -1 0 5600 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1969_
timestamp 1753272495
transform -1 0 3584 0 -1 29792
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1970_
timestamp 1751740063
transform 1 0 2576 0 1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1971_
timestamp 1751889408
transform 1 0 4592 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1972_
timestamp 1753182340
transform 1 0 2800 0 1 31360
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1973_
timestamp 1751534193
transform -1 0 2688 0 1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1974_
timestamp 1753277515
transform 1 0 4256 0 -1 32928
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1975_
timestamp 1751532043
transform -1 0 6160 0 1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1976_
timestamp 1753441877
transform 1 0 4032 0 1 31360
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1977_
timestamp 1751889808
transform 1 0 6608 0 -1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1978_
timestamp 1753371985
transform -1 0 6608 0 -1 34496
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1979_
timestamp 1751889408
transform -1 0 6272 0 1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1980_
timestamp 1751534193
transform -1 0 2688 0 -1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1981_
timestamp 1751532043
transform 1 0 9856 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1982_
timestamp 1753277515
transform -1 0 10528 0 1 34496
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _1983_
timestamp 1752061876
transform 1 0 5488 0 1 31360
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1984_
timestamp 1753441877
transform 1 0 5824 0 -1 32928
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1985_
timestamp 1751889808
transform -1 0 8736 0 1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1986_
timestamp 1753371985
transform -1 0 7952 0 1 34496
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1987_
timestamp 1751889408
transform -1 0 7840 0 1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1988_
timestamp 1751534193
transform -1 0 7056 0 1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1989_
timestamp 1753272495
transform 1 0 9408 0 -1 36064
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1990_
timestamp 1751532043
transform -1 0 10080 0 1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1991_
timestamp 1753277515
transform 1 0 9968 0 1 37632
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_4  _1992_
timestamp 1751558652
transform 1 0 38528 0 1 23520
box -86 -86 1094 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1993_
timestamp 1751889808
transform -1 0 11088 0 1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1994_
timestamp 1751531619
transform 1 0 9184 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1995_
timestamp 1753371985
transform -1 0 10976 0 -1 37632
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1996_
timestamp 1751532043
transform -1 0 3472 0 -1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1997_
timestamp 1753277515
transform 1 0 2800 0 -1 39200
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1998_
timestamp 1753272495
transform -1 0 11424 0 1 39200
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1999_
timestamp 1751889808
transform 1 0 4368 0 1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2000_
timestamp 1751534193
transform -1 0 16128 0 1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2001_
timestamp 1753371985
transform 1 0 5488 0 1 39200
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2002_
timestamp 1751889408
transform 1 0 4816 0 -1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2003_
timestamp 1751534193
transform -1 0 2688 0 -1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2004_
timestamp 1753277515
transform -1 0 6160 0 -1 42336
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _2005_
timestamp 1753272495
transform -1 0 4816 0 -1 40768
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2006_
timestamp 1751740063
transform -1 0 4144 0 1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2007_
timestamp 1751889408
transform 1 0 4144 0 1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2008_
timestamp 1753182340
transform 1 0 3136 0 1 40768
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2009_
timestamp 1751534193
transform -1 0 2800 0 1 40768
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2010_
timestamp 1751534193
transform -1 0 17024 0 1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2011_
timestamp 1751532043
transform -1 0 5936 0 -1 45472
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2012_
timestamp 1753277515
transform 1 0 5264 0 -1 43904
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _2013_
timestamp 1752061876
transform 1 0 6160 0 -1 42336
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2014_
timestamp 1751889808
transform -1 0 6272 0 1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2015_
timestamp 1751740063
transform 1 0 4480 0 -1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2016_
timestamp 1751889408
transform 1 0 5824 0 1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2017_
timestamp 1753182340
transform -1 0 8064 0 -1 43904
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2018_
timestamp 1751534193
transform -1 0 4480 0 -1 43904
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2019_
timestamp 1751740063
transform 1 0 9408 0 -1 45472
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2020_
timestamp 1751889408
transform 1 0 9408 0 -1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2021_
timestamp 1751740063
transform -1 0 11312 0 1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2022_
timestamp 1753441877
transform 1 0 6272 0 1 42336
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2023_
timestamp 1751889808
transform -1 0 8176 0 1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2024_
timestamp 1753371985
transform -1 0 9184 0 -1 43904
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2025_
timestamp 1751889408
transform -1 0 7392 0 1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2026_
timestamp 1751534193
transform 1 0 7280 0 1 45472
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2027_
timestamp 1753371985
transform -1 0 9296 0 1 43904
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2028_
timestamp 1753182340
transform -1 0 10528 0 1 43904
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2029_
timestamp 1751534193
transform 1 0 10528 0 1 45472
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2030_
timestamp 1751740063
transform 1 0 7504 0 1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2031_
timestamp 1751889408
transform 1 0 8288 0 1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2032_
timestamp 1753182340
transform 1 0 7616 0 -1 32928
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2033_
timestamp 1751534193
transform -1 0 7616 0 -1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2034_
timestamp 1753277515
transform -1 0 9184 0 -1 29792
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2035_
timestamp 1751889808
transform -1 0 8400 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2036_
timestamp 1753371985
transform -1 0 7616 0 -1 31360
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2037_
timestamp 1751889408
transform -1 0 6496 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2038_
timestamp 1751534193
transform 1 0 8400 0 -1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2039_
timestamp 1753277515
transform 1 0 11200 0 1 31360
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _2040_
timestamp 1753272495
transform 1 0 9408 0 -1 31360
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2041_
timestamp 1751889808
transform -1 0 9856 0 1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2042_
timestamp 1753371985
transform 1 0 10080 0 -1 34496
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2043_
timestamp 1751889408
transform 1 0 10752 0 1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2044_
timestamp 1751534193
transform -1 0 9184 0 -1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2045_
timestamp 1753277515
transform 1 0 3248 0 1 34496
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _2046_
timestamp 1753272495
transform -1 0 11200 0 1 31360
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2047_
timestamp 1751889808
transform -1 0 3248 0 1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2048_
timestamp 1751534193
transform 1 0 16128 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2049_
timestamp 1751534193
transform -1 0 16800 0 -1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2050_
timestamp 1753371985
transform 1 0 4592 0 -1 36064
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2051_
timestamp 1751889408
transform 1 0 3360 0 1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2052_
timestamp 1751534193
transform -1 0 2688 0 1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2053_
timestamp 1753277515
transform -1 0 6160 0 -1 37632
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2054_
timestamp 1751532043
transform -1 0 5264 0 1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _2055_
timestamp 1753272495
transform 1 0 3808 0 -1 34496
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2056_
timestamp 1751889808
transform -1 0 5152 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2057_
timestamp 1753371985
transform -1 0 5264 0 1 36064
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2058_
timestamp 1751889408
transform -1 0 4368 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2059_
timestamp 1751534193
transform -1 0 2688 0 1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _2060_
timestamp 1753272495
transform 1 0 6160 0 -1 37632
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2061_
timestamp 1751532043
transform -1 0 7056 0 1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2062_
timestamp 1753277515
transform 1 0 6608 0 1 37632
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2063_
timestamp 1751889808
transform 1 0 7504 0 -1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2064_
timestamp 1751531619
transform -1 0 8960 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2065_
timestamp 1753371985
transform 1 0 7952 0 -1 39200
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2066_
timestamp 1751532043
transform 1 0 8736 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2067_
timestamp 1753277515
transform -1 0 10080 0 1 40768
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _2068_
timestamp 1753272495
transform 1 0 7056 0 1 39200
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2069_
timestamp 1751889808
transform -1 0 7840 0 -1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2070_
timestamp 1753371985
transform -1 0 8736 0 -1 42336
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2071_
timestamp 1751889408
transform 1 0 7616 0 1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2072_
timestamp 1751534193
transform -1 0 7056 0 -1 40768
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2073_
timestamp 1753277515
transform 1 0 10752 0 1 40768
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _2074_
timestamp 1753272495
transform 1 0 7840 0 -1 40768
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2075_
timestamp 1751740063
transform -1 0 13104 0 1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2076_
timestamp 1751889408
transform -1 0 12096 0 -1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2077_
timestamp 1753182340
transform 1 0 10080 0 -1 42336
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2078_
timestamp 1751534193
transform -1 0 10080 0 -1 42336
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_4  _2079_
timestamp 1751558652
transform -1 0 17024 0 -1 39200
box -86 -86 1094 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2080_
timestamp 1751532043
transform -1 0 15568 0 -1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2081_
timestamp 1753277515
transform 1 0 14784 0 1 40768
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2082_
timestamp 1751532043
transform -1 0 12544 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2083_
timestamp 1753441877
transform 1 0 11536 0 -1 40768
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2084_
timestamp 1751740063
transform 1 0 15680 0 1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2085_
timestamp 1751889408
transform -1 0 15456 0 -1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2086_
timestamp 1753182340
transform -1 0 16912 0 -1 40768
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2087_
timestamp 1751534193
transform 1 0 17248 0 -1 40768
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2088_
timestamp 1751740063
transform -1 0 13104 0 1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2089_
timestamp 1751889408
transform 1 0 13664 0 1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2090_
timestamp 1751740063
transform 1 0 13888 0 1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2091_
timestamp 1753441877
transform 1 0 15456 0 -1 42336
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2092_
timestamp 1751889808
transform 1 0 17472 0 1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2093_
timestamp 1753371985
transform 1 0 15568 0 1 42336
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2094_
timestamp 1751889408
transform -1 0 17472 0 1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2095_
timestamp 1751534193
transform -1 0 17248 0 1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2096_
timestamp 1753371985
transform 1 0 14448 0 1 42336
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2097_
timestamp 1753182340
transform -1 0 16576 0 -1 43904
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2098_
timestamp 1751534193
transform -1 0 12768 0 1 45472
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2099_
timestamp 1751531619
transform -1 0 28672 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2100_
timestamp 1751740063
transform 1 0 13776 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2101_
timestamp 1751532043
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2102_
timestamp 1751531619
transform 1 0 31808 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2103_
timestamp 1751532043
transform -1 0 32480 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2104_
timestamp 1751532043
transform -1 0 31808 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2105_
timestamp 1753371985
transform -1 0 34048 0 -1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2106_
timestamp 1751531619
transform 1 0 33040 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2107_
timestamp 1753371985
transform -1 0 34048 0 -1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2108_
timestamp 1753868718
transform -1 0 33376 0 1 18816
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2109_
timestamp 1751740063
transform -1 0 8960 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2110_
timestamp 1751534193
transform -1 0 7840 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2111_
timestamp 1751532043
transform -1 0 13104 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2112_
timestamp 1751889808
transform -1 0 9072 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2113_
timestamp 1751534193
transform 1 0 8400 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2114_
timestamp 1751889808
transform -1 0 15904 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2115_
timestamp 1751534193
transform -1 0 8848 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2116_
timestamp 1753441877
transform -1 0 10528 0 -1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2117_
timestamp 1753371985
transform 1 0 8848 0 1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2118_
timestamp 1751534193
transform 1 0 8512 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2119_
timestamp 1751532043
transform -1 0 7392 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2120_
timestamp 1751534193
transform 1 0 7392 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2121_
timestamp 1753441877
transform 1 0 8064 0 -1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2122_
timestamp 1753371985
transform -1 0 10528 0 -1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2123_
timestamp 1751534193
transform 1 0 5040 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2124_
timestamp 1751534193
transform -1 0 8176 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2125_
timestamp 1751740063
transform -1 0 7840 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2126_
timestamp 1751740063
transform 1 0 6048 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2127_
timestamp 1753182340
transform 1 0 5824 0 1 15680
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2128_
timestamp 1751534193
transform -1 0 5152 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2129_
timestamp 1751740063
transform 1 0 4032 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2130_
timestamp 1751740063
transform -1 0 6384 0 1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2131_
timestamp 1753182340
transform 1 0 4816 0 -1 15680
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2132_
timestamp 1751534193
transform -1 0 3920 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2133_
timestamp 1751534193
transform -1 0 8512 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2134_
timestamp 1751740063
transform -1 0 7504 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2135_
timestamp 1751740063
transform 1 0 6384 0 1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2136_
timestamp 1753182340
transform 1 0 5712 0 -1 14112
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2137_
timestamp 1751534193
transform -1 0 3584 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2138_
timestamp 1751534193
transform -1 0 8176 0 -1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2139_
timestamp 1751740063
transform 1 0 5488 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2140_
timestamp 1751740063
transform 1 0 7504 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2141_
timestamp 1753182340
transform 1 0 5488 0 1 12544
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2142_
timestamp 1751534193
transform -1 0 5264 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2143_
timestamp 1751534193
transform -1 0 5264 0 1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2144_
timestamp 1751740063
transform 1 0 3920 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2145_
timestamp 1751740063
transform 1 0 6272 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2146_
timestamp 1753182340
transform 1 0 4704 0 -1 10976
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2147_
timestamp 1751534193
transform -1 0 3360 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2148_
timestamp 1751740063
transform 1 0 3696 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2149_
timestamp 1751534193
transform -1 0 10192 0 1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2150_
timestamp 1751740063
transform 1 0 6720 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2151_
timestamp 1753182340
transform 1 0 5488 0 1 9408
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2152_
timestamp 1751534193
transform -1 0 2688 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2153_
timestamp 1751740063
transform 1 0 4480 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2154_
timestamp 1751740063
transform 1 0 6272 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2155_
timestamp 1753182340
transform 1 0 5040 0 -1 9408
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2156_
timestamp 1751534193
transform -1 0 3136 0 1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2157_
timestamp 1751740063
transform -1 0 7504 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2158_
timestamp 1751740063
transform 1 0 5936 0 1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2159_
timestamp 1753182340
transform 1 0 5488 0 1 7840
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2160_
timestamp 1751534193
transform -1 0 4592 0 1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2161_
timestamp 1751534193
transform 1 0 7504 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2162_
timestamp 1751740063
transform -1 0 9184 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2163_
timestamp 1751740063
transform -1 0 7280 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2164_
timestamp 1753182340
transform -1 0 8512 0 -1 7840
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2165_
timestamp 1751534193
transform -1 0 5264 0 1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2166_
timestamp 1751740063
transform 1 0 8064 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2167_
timestamp 1751740063
transform -1 0 11424 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2168_
timestamp 1753182340
transform 1 0 9408 0 -1 7840
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2169_
timestamp 1751534193
transform -1 0 10080 0 -1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2170_
timestamp 1751740063
transform -1 0 7952 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2171_
timestamp 1751740063
transform -1 0 9520 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2172_
timestamp 1753182340
transform 1 0 7952 0 -1 9408
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2173_
timestamp 1751534193
transform 1 0 9408 0 -1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2174_
timestamp 1751740063
transform 1 0 9408 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2175_
timestamp 1751740063
transform -1 0 9184 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2176_
timestamp 1753182340
transform -1 0 9408 0 1 10976
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2177_
timestamp 1751534193
transform -1 0 8624 0 1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2178_
timestamp 1751889408
transform -1 0 13216 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2179_
timestamp 1753277515
transform -1 0 12656 0 1 14112
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2180_
timestamp 1753441877
transform -1 0 11088 0 1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2181_
timestamp 1753441877
transform 1 0 9408 0 -1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2182_
timestamp 1751534193
transform 1 0 10528 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2183_
timestamp 1751889808
transform 1 0 45584 0 -1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2184_
timestamp 1753182340
transform -1 0 48048 0 1 23520
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2185_
timestamp 1753182340
transform -1 0 47040 0 1 26656
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2186_
timestamp 1751889808
transform 1 0 47040 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2187_
timestamp 1751889808
transform 1 0 47152 0 1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2188_
timestamp 1751532043
transform 1 0 40992 0 1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2189_
timestamp 1753868718
transform -1 0 48160 0 -1 26656
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2190_
timestamp 1751534193
transform -1 0 38976 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2191_
timestamp 1751534193
transform -1 0 37520 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2192_
timestamp 1751534193
transform 1 0 35952 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2193_
timestamp 1751740063
transform -1 0 44576 0 -1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2194_
timestamp 1751889408
transform -1 0 43680 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2195_
timestamp 1753182340
transform 1 0 41664 0 1 20384
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2196_
timestamp 1751534193
transform -1 0 42112 0 1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2197_
timestamp 1751740063
transform -1 0 43568 0 1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2198_
timestamp 1751889408
transform -1 0 44240 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2199_
timestamp 1753182340
transform 1 0 42224 0 1 21952
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2200_
timestamp 1751534193
transform 1 0 43568 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2201_
timestamp 1751534193
transform 1 0 23632 0 1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2202_
timestamp 1751740063
transform -1 0 42784 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2203_
timestamp 1751889408
transform -1 0 43568 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2204_
timestamp 1753182340
transform 1 0 40768 0 -1 25088
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2205_
timestamp 1751534193
transform 1 0 41552 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2206_
timestamp 1751740063
transform -1 0 41776 0 1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2207_
timestamp 1751889408
transform -1 0 41552 0 -1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2208_
timestamp 1753182340
transform -1 0 40992 0 1 23520
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2209_
timestamp 1751534193
transform -1 0 40208 0 -1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2210_
timestamp 1751740063
transform -1 0 37632 0 1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2211_
timestamp 1751889408
transform -1 0 37632 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2212_
timestamp 1753182340
transform -1 0 36624 0 1 23520
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2213_
timestamp 1751534193
transform -1 0 35392 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2214_
timestamp 1751531619
transform 1 0 36400 0 -1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2215_
timestamp 1751889808
transform 1 0 34384 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2216_
timestamp 1751889408
transform -1 0 35952 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2217_
timestamp 1751889408
transform -1 0 35728 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2218_
timestamp 1751534193
transform -1 0 34944 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2219_
timestamp 1753277515
transform 1 0 34272 0 -1 20384
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2220_
timestamp 1751889408
transform -1 0 36624 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2221_
timestamp 1751534193
transform -1 0 36400 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2222_
timestamp 1751531619
transform -1 0 39312 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2223_
timestamp 1751534193
transform 1 0 40544 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2224_
timestamp 1751889808
transform 1 0 38976 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2225_
timestamp 1751889408
transform -1 0 41552 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2226_
timestamp 1751889408
transform 1 0 39312 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2227_
timestamp 1751534193
transform -1 0 38976 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2228_
timestamp 1753277515
transform 1 0 25536 0 1 29792
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2229_
timestamp 1751889808
transform -1 0 25872 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2230_
timestamp 1751534193
transform -1 0 17920 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2231_
timestamp 1753371985
transform -1 0 26208 0 -1 29792
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2232_
timestamp 1751889408
transform -1 0 24864 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2233_
timestamp 1751534193
transform -1 0 23296 0 -1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2234_
timestamp 1753277515
transform -1 0 24864 0 -1 32928
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2235_
timestamp 1751531619
transform -1 0 24864 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2236_
timestamp 1751531619
transform -1 0 24080 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2237_
timestamp 1751889808
transform -1 0 23296 0 -1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2238_
timestamp 1753371985
transform -1 0 25872 0 1 32928
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2239_
timestamp 1751889408
transform 1 0 23744 0 -1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2240_
timestamp 1751534193
transform -1 0 23744 0 -1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2241_
timestamp 1751532043
transform 1 0 18592 0 -1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2242_
timestamp 1753277515
transform -1 0 17024 0 -1 32928
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _2243_
timestamp 1753272495
transform -1 0 25088 0 1 31360
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2244_
timestamp 1751889808
transform -1 0 17024 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2245_
timestamp 1753371985
transform 1 0 16800 0 1 31360
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2246_
timestamp 1751889408
transform -1 0 16800 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2247_
timestamp 1751534193
transform -1 0 16240 0 -1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2248_
timestamp 1751532043
transform 1 0 17248 0 -1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2249_
timestamp 1753277515
transform 1 0 17248 0 1 32928
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _2250_
timestamp 1753272495
transform -1 0 18592 0 -1 32928
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2251_
timestamp 1751889808
transform 1 0 16240 0 1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2252_
timestamp 1753371985
transform 1 0 16128 0 1 32928
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2253_
timestamp 1751889408
transform 1 0 17920 0 -1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2254_
timestamp 1751534193
transform -1 0 15568 0 1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _2255_
timestamp 1753272495
transform 1 0 17136 0 1 34496
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2256_
timestamp 1751532043
transform 1 0 20832 0 -1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2257_
timestamp 1753277515
transform -1 0 20160 0 1 36064
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2258_
timestamp 1751889808
transform 1 0 19040 0 -1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2259_
timestamp 1751531619
transform -1 0 20944 0 1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2260_
timestamp 1753371985
transform 1 0 17920 0 -1 37632
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2261_
timestamp 1751532043
transform -1 0 20496 0 -1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2262_
timestamp 1753277515
transform 1 0 20496 0 -1 37632
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _2263_
timestamp 1753272495
transform 1 0 18704 0 -1 36064
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2264_
timestamp 1751889808
transform -1 0 21952 0 1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2265_
timestamp 1751534193
transform -1 0 22960 0 1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2266_
timestamp 1753371985
transform 1 0 22064 0 -1 37632
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2267_
timestamp 1751889408
transform 1 0 21952 0 1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2268_
timestamp 1751534193
transform -1 0 19040 0 1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2269_
timestamp 1751532043
transform -1 0 20384 0 -1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2270_
timestamp 1753277515
transform 1 0 21168 0 1 39200
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _2271_
timestamp 1753272495
transform 1 0 21168 0 1 37632
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2272_
timestamp 1751740063
transform 1 0 20608 0 -1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2273_
timestamp 1751889408
transform 1 0 22288 0 -1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2274_
timestamp 1753182340
transform -1 0 22624 0 -1 39200
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2275_
timestamp 1751534193
transform -1 0 19376 0 -1 40768
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2276_
timestamp 1753277515
transform 1 0 20608 0 -1 42336
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2277_
timestamp 1753441877
transform 1 0 21168 0 -1 40768
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2278_
timestamp 1751889808
transform 1 0 23296 0 1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2279_
timestamp 1753371985
transform 1 0 22176 0 -1 42336
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2280_
timestamp 1751889408
transform -1 0 23296 0 1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2281_
timestamp 1751534193
transform -1 0 19264 0 1 42336
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2282_
timestamp 1751532043
transform -1 0 19824 0 1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2283_
timestamp 1753277515
transform 1 0 20720 0 -1 43904
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _2284_
timestamp 1753272495
transform 1 0 21168 0 1 40768
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2285_
timestamp 1751889808
transform 1 0 23408 0 -1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2286_
timestamp 1753371985
transform 1 0 22288 0 -1 43904
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2287_
timestamp 1751889408
transform 1 0 23968 0 1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2288_
timestamp 1751534193
transform -1 0 17584 0 1 45472
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2289_
timestamp 1753441877
transform 1 0 19824 0 1 42336
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2290_
timestamp 1753371985
transform 1 0 21168 0 1 42336
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2291_
timestamp 1751889408
transform 1 0 20944 0 -1 45472
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2292_
timestamp 1751534193
transform -1 0 20160 0 1 40768
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2293_
timestamp 1751534193
transform 1 0 37520 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2294_
timestamp 1751534193
transform 1 0 38640 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2295_
timestamp 1751889808
transform -1 0 38752 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2296_
timestamp 1751740063
transform -1 0 44016 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2297_
timestamp 1751740063
transform -1 0 44352 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2298_
timestamp 1751740063
transform 1 0 42000 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2299_
timestamp 1751740063
transform -1 0 44128 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _2300_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753172561
transform -1 0 43120 0 -1 15680
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2301_
timestamp 1753182340
transform 1 0 41552 0 1 14112
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2302_
timestamp 1753441877
transform 1 0 39424 0 -1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2303_
timestamp 1751534193
transform 1 0 34272 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2304_
timestamp 1753371985
transform -1 0 39424 0 -1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2305_
timestamp 1751889408
transform 1 0 40768 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2306_
timestamp 1751534193
transform -1 0 37520 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2307_
timestamp 1751534193
transform 1 0 37968 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2308_
timestamp 1751534193
transform 1 0 36624 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2309_
timestamp 1751534193
transform 1 0 40880 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2310_
timestamp 1753441877
transform 1 0 41216 0 1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2311_
timestamp 1751531619
transform 1 0 41552 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2312_
timestamp 1751889808
transform 1 0 42336 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2313_
timestamp 1751534193
transform 1 0 44576 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2314_
timestamp 1751534193
transform 1 0 38192 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2315_
timestamp 1751889808
transform 1 0 43456 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2316_
timestamp 1751531619
transform -1 0 44688 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _2317_
timestamp 1753891287
transform 1 0 41552 0 1 18816
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2318_
timestamp 1753441877
transform 1 0 42336 0 1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2319_
timestamp 1751531619
transform 1 0 43456 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2320_
timestamp 1751889808
transform 1 0 44352 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2321_
timestamp 1751534193
transform 1 0 44688 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2322_
timestamp 1751889808
transform 1 0 44688 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2323_
timestamp 1751531619
transform -1 0 46256 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _2324_
timestamp 1753891287
transform 1 0 43456 0 -1 18816
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2325_
timestamp 1751534193
transform 1 0 37296 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2326_
timestamp 1751534193
transform 1 0 44688 0 1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2327_
timestamp 1753441877
transform 1 0 42112 0 1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2328_
timestamp 1751531619
transform -1 0 44464 0 1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2329_
timestamp 1751740063
transform 1 0 44240 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2330_
timestamp 1751534193
transform 1 0 44688 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2331_
timestamp 1751532043
transform 1 0 44800 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2332_
timestamp 1751534193
transform 1 0 38864 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2333_
timestamp 1751534193
transform 1 0 46816 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2334_
timestamp 1751889808
transform -1 0 48272 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2335_
timestamp 1751531619
transform -1 0 47488 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _2336_
timestamp 1753891287
transform 1 0 45136 0 -1 17248
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2337_
timestamp 1751534193
transform 1 0 42784 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2338_
timestamp 1753371985
transform 1 0 42224 0 -1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2339_
timestamp 1751889808
transform 1 0 46256 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2340_
timestamp 1751531619
transform -1 0 46256 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2341_
timestamp 1751889808
transform 1 0 47600 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2342_
timestamp 1751531619
transform 1 0 47040 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _2343_
timestamp 1753891287
transform 1 0 45248 0 -1 12544
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2344_
timestamp 1751534193
transform -1 0 43792 0 1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2345_
timestamp 1753441877
transform 1 0 43120 0 -1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2346_
timestamp 1751532043
transform 1 0 44016 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2347_
timestamp 1753277515
transform -1 0 44464 0 1 12544
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2348_
timestamp 1751534193
transform 1 0 37744 0 1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2349_
timestamp 1751889808
transform 1 0 41552 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2350_
timestamp 1751531619
transform 1 0 42336 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2351_
timestamp 1753371985
transform -1 0 44240 0 1 10976
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2352_
timestamp 1753371985
transform 1 0 40992 0 1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2353_
timestamp 1753960525
transform 1 0 44352 0 -1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _2354_
timestamp 1753172561
transform 1 0 44688 0 1 14112
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2355_
timestamp 1751889808
transform 1 0 47040 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2356_
timestamp 1751531619
transform -1 0 47488 0 1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _2357_
timestamp 1753891287
transform 1 0 45248 0 1 15680
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2358_
timestamp 1751534193
transform -1 0 42224 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2359_
timestamp 1753441877
transform 1 0 42448 0 -1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2360_
timestamp 1751531619
transform -1 0 47600 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2361_
timestamp 1751889808
transform -1 0 45248 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2362_
timestamp 1751534193
transform 1 0 45248 0 -1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2363_
timestamp 1751889808
transform 1 0 47600 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2364_
timestamp 1751531619
transform -1 0 47600 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _2365_
timestamp 1753891287
transform 1 0 45248 0 1 10976
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2366_
timestamp 1753441877
transform 1 0 40880 0 1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2367_
timestamp 1751889408
transform -1 0 40544 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2368_
timestamp 1751740063
transform 1 0 40768 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2369_
timestamp 1751740063
transform -1 0 42336 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2370_
timestamp 1751534193
transform -1 0 37296 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2371_
timestamp 1751889808
transform -1 0 40544 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2372_
timestamp 1751531619
transform -1 0 41552 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2373_
timestamp 1753371985
transform 1 0 40208 0 1 10976
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2374_
timestamp 1751534193
transform -1 0 36176 0 -1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2375_
timestamp 1751534193
transform -1 0 36624 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2376_
timestamp 1753960525
transform 1 0 36848 0 -1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2377_
timestamp 1753371985
transform 1 0 37072 0 -1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2378_
timestamp 1751534193
transform -1 0 21168 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2379_
timestamp 1753960525
transform -1 0 39088 0 -1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2380_
timestamp 1751740063
transform 1 0 37072 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2381_
timestamp 1751889408
transform 1 0 38192 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2382_
timestamp 1751889808
transform 1 0 37520 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2383_
timestamp 1751531619
transform -1 0 40544 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2384_
timestamp 1753371985
transform 1 0 37296 0 -1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2385_
timestamp 1751889808
transform -1 0 38640 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2386_
timestamp 1751740063
transform -1 0 42224 0 1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2387_
timestamp 1751740063
transform -1 0 40656 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2388_
timestamp 1751740063
transform 1 0 35504 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2389_
timestamp 1751740063
transform 1 0 40768 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _2390_
timestamp 1753172561
transform -1 0 40544 0 -1 7840
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2391_
timestamp 1753182340
transform 1 0 38976 0 1 6272
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2392_
timestamp 1753441877
transform 1 0 38752 0 1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2393_
timestamp 1753371985
transform -1 0 38304 0 1 6272
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2394_
timestamp 1751889408
transform -1 0 37856 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2395_
timestamp 1751534193
transform 1 0 38304 0 1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2396_
timestamp 1751534193
transform -1 0 43456 0 -1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2397_
timestamp 1751534193
transform 1 0 40208 0 1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2398_
timestamp 1753441877
transform 1 0 40880 0 -1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2399_
timestamp 1751531619
transform 1 0 42112 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2400_
timestamp 1751889808
transform 1 0 42896 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2401_
timestamp 1751534193
transform -1 0 47152 0 -1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2402_
timestamp 1751889808
transform 1 0 46144 0 1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2403_
timestamp 1751531619
transform -1 0 46816 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _2404_
timestamp 1753891287
transform 1 0 42896 0 1 7840
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2405_
timestamp 1753441877
transform 1 0 42224 0 1 6272
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2406_
timestamp 1751531619
transform 1 0 43568 0 1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2407_
timestamp 1751889808
transform 1 0 43456 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2408_
timestamp 1751889808
transform 1 0 46368 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2409_
timestamp 1751531619
transform -1 0 47712 0 1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _2410_
timestamp 1753891287
transform 1 0 43792 0 -1 7840
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2411_
timestamp 1753441877
transform 1 0 42560 0 1 4704
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2412_
timestamp 1751531619
transform 1 0 44240 0 1 3136
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2413_
timestamp 1751740063
transform -1 0 44464 0 1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2414_
timestamp 1751534193
transform 1 0 44688 0 1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2415_
timestamp 1751532043
transform 1 0 44800 0 1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2416_
timestamp 1751889808
transform 1 0 45360 0 1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2417_
timestamp 1751531619
transform -1 0 47936 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _2418_
timestamp 1753891287
transform 1 0 44576 0 -1 6272
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2419_
timestamp 1751534193
transform -1 0 42224 0 -1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2420_
timestamp 1753371985
transform 1 0 38304 0 1 4704
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2421_
timestamp 1751889808
transform -1 0 42784 0 1 3136
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2422_
timestamp 1751531619
transform 1 0 41216 0 1 3136
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2423_
timestamp 1751534193
transform 1 0 27888 0 1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2424_
timestamp 1751889808
transform 1 0 45696 0 -1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2425_
timestamp 1751531619
transform -1 0 44240 0 1 3136
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _2426_
timestamp 1753891287
transform -1 0 42672 0 -1 4704
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2427_
timestamp 1753441877
transform 1 0 38864 0 -1 6272
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2428_
timestamp 1751532043
transform 1 0 39984 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2429_
timestamp 1753277515
transform -1 0 42560 0 1 4704
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2430_
timestamp 1751889808
transform 1 0 39760 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2431_
timestamp 1751531619
transform 1 0 41552 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2432_
timestamp 1753371985
transform 1 0 40992 0 1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2433_
timestamp 1751534193
transform -1 0 37072 0 -1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2434_
timestamp 1753371985
transform 1 0 36848 0 1 4704
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2435_
timestamp 1753960525
transform -1 0 41216 0 1 3136
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _2436_
timestamp 1753172561
transform -1 0 40992 0 1 4704
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2437_
timestamp 1751534193
transform 1 0 23408 0 -1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2438_
timestamp 1751889808
transform 1 0 38080 0 1 3136
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2439_
timestamp 1751531619
transform -1 0 40432 0 -1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _2440_
timestamp 1753891287
transform 1 0 36512 0 1 3136
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2441_
timestamp 1751534193
transform -1 0 36288 0 -1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2442_
timestamp 1753441877
transform 1 0 33488 0 1 4704
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2443_
timestamp 1751531619
transform -1 0 35392 0 1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2444_
timestamp 1751889808
transform -1 0 34832 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2445_
timestamp 1751889808
transform 1 0 34832 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2446_
timestamp 1751531619
transform -1 0 36176 0 1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _2447_
timestamp 1753891287
transform 1 0 33376 0 1 3136
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2448_
timestamp 1753441877
transform 1 0 34272 0 1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2449_
timestamp 1751889408
transform 1 0 35280 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2450_
timestamp 1751740063
transform 1 0 34496 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2451_
timestamp 1751740063
transform -1 0 35952 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2452_
timestamp 1751889808
transform 1 0 39200 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2453_
timestamp 1751531619
transform -1 0 39200 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2454_
timestamp 1753371985
transform 1 0 37296 0 1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2455_
timestamp 1753960525
transform 1 0 34384 0 -1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2456_
timestamp 1753371985
transform 1 0 34160 0 1 10976
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2457_
timestamp 1753960525
transform -1 0 36400 0 1 10976
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2458_
timestamp 1751740063
transform -1 0 34384 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2459_
timestamp 1751889408
transform -1 0 35280 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_4  _2460_
timestamp 1751558652
transform 1 0 38752 0 -1 20384
box -86 -86 1094 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2461_
timestamp 1751889808
transform 1 0 5488 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2462_
timestamp 1751531619
transform -1 0 6608 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2463_
timestamp 1753371985
transform -1 0 7168 0 -1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2464_
timestamp 1751889808
transform 1 0 33152 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2465_
timestamp 1751740063
transform 1 0 17808 0 -1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2466_
timestamp 1751740063
transform -1 0 26544 0 1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2467_
timestamp 1751740063
transform 1 0 16576 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2468_
timestamp 1751740063
transform 1 0 14336 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _2469_
timestamp 1753172561
transform -1 0 19040 0 1 6272
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2470_
timestamp 1753182340
transform 1 0 17472 0 -1 6272
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2471_
timestamp 1753441877
transform 1 0 24640 0 1 6272
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2472_
timestamp 1753371985
transform 1 0 33936 0 -1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2473_
timestamp 1751889408
transform 1 0 34160 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2474_
timestamp 1751534193
transform 1 0 35952 0 1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2475_
timestamp 1753441877
transform 1 0 25088 0 -1 6272
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2476_
timestamp 1751531619
transform 1 0 22624 0 1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2477_
timestamp 1751889808
transform -1 0 24864 0 -1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2478_
timestamp 1751889808
transform -1 0 25760 0 1 3136
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2479_
timestamp 1751531619
transform -1 0 26544 0 1 3136
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _2480_
timestamp 1753891287
transform -1 0 26656 0 -1 4704
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2481_
timestamp 1751534193
transform -1 0 19712 0 1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2482_
timestamp 1753441877
transform -1 0 20496 0 1 4704
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2483_
timestamp 1751531619
transform 1 0 18816 0 -1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2484_
timestamp 1751889808
transform -1 0 20384 0 1 3136
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2485_
timestamp 1751534193
transform -1 0 22848 0 1 3136
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2486_
timestamp 1751889808
transform 1 0 22624 0 -1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2487_
timestamp 1751531619
transform -1 0 22400 0 1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _2488_
timestamp 1753891287
transform -1 0 22176 0 1 3136
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2489_
timestamp 1751534193
transform 1 0 14672 0 -1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2490_
timestamp 1753441877
transform -1 0 19376 0 1 4704
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2491_
timestamp 1751531619
transform -1 0 16240 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2492_
timestamp 1751740063
transform -1 0 17024 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2493_
timestamp 1751534193
transform -1 0 15456 0 1 3136
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2494_
timestamp 1751532043
transform 1 0 17248 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2495_
timestamp 1751534193
transform -1 0 18816 0 1 3136
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2496_
timestamp 1751889808
transform -1 0 18144 0 1 3136
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2497_
timestamp 1751531619
transform 1 0 15792 0 1 3136
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _2498_
timestamp 1753891287
transform 1 0 15120 0 -1 4704
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2499_
timestamp 1751534193
transform -1 0 17472 0 1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2500_
timestamp 1753371985
transform -1 0 14896 0 -1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2501_
timestamp 1751889808
transform -1 0 12992 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2502_
timestamp 1751531619
transform 1 0 13328 0 1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2503_
timestamp 1751889808
transform -1 0 13776 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2504_
timestamp 1751531619
transform 1 0 12320 0 1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _2505_
timestamp 1753891287
transform -1 0 13776 0 -1 6272
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2506_
timestamp 1753441877
transform -1 0 18816 0 -1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2507_
timestamp 1751532043
transform -1 0 17024 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2508_
timestamp 1753277515
transform 1 0 14896 0 -1 7840
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2509_
timestamp 1751889808
transform -1 0 18480 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2510_
timestamp 1751531619
transform -1 0 18032 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2511_
timestamp 1753371985
transform 1 0 15904 0 -1 10976
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2512_
timestamp 1753371985
transform -1 0 16800 0 1 6272
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2513_
timestamp 1753960525
transform -1 0 15456 0 -1 6272
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _2514_
timestamp 1753172561
transform -1 0 15680 0 1 6272
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2515_
timestamp 1751889808
transform -1 0 14784 0 1 3136
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2516_
timestamp 1751531619
transform 1 0 13216 0 1 3136
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _2517_
timestamp 1753891287
transform -1 0 14896 0 1 4704
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2518_
timestamp 1753441877
transform -1 0 15232 0 1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2519_
timestamp 1751531619
transform -1 0 14448 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2520_
timestamp 1751889808
transform -1 0 14112 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2521_
timestamp 1751889808
transform -1 0 13104 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2522_
timestamp 1751531619
transform -1 0 14112 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _2523_
timestamp 1753891287
transform -1 0 13104 0 1 9408
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2524_
timestamp 1751534193
transform -1 0 16016 0 -1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2525_
timestamp 1753441877
transform 1 0 13552 0 -1 10976
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2526_
timestamp 1751531619
transform 1 0 12768 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2527_
timestamp 1751889808
transform 1 0 14672 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2528_
timestamp 1751889808
transform -1 0 16576 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2529_
timestamp 1751531619
transform -1 0 16240 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _2530_
timestamp 1753891287
transform 1 0 13888 0 1 10976
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2531_
timestamp 1753371985
transform 1 0 14784 0 -1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2532_
timestamp 1753277515
transform 1 0 13888 0 1 12544
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2533_
timestamp 1751889808
transform 1 0 17584 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2534_
timestamp 1751531619
transform -1 0 19152 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2535_
timestamp 1753371985
transform 1 0 15904 0 -1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2536_
timestamp 1753371985
transform -1 0 14448 0 1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2537_
timestamp 1753960525
transform -1 0 15120 0 -1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2538_
timestamp 1751740063
transform -1 0 13104 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2539_
timestamp 1751534193
transform 1 0 39312 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2540_
timestamp 1753277515
transform 1 0 33488 0 1 28224
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2541_
timestamp 1753277515
transform 1 0 35056 0 1 28224
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2542_
timestamp 1751740063
transform -1 0 42224 0 1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2543_
timestamp 1751889408
transform -1 0 40544 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2544_
timestamp 1753182340
transform -1 0 42000 0 -1 28224
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2545_
timestamp 1751534193
transform 1 0 43344 0 1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2546_
timestamp 1751532043
transform -1 0 36176 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2547_
timestamp 1753277515
transform 1 0 33600 0 -1 29792
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2548_
timestamp 1753277515
transform 1 0 36176 0 -1 29792
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2549_
timestamp 1751889808
transform 1 0 37744 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2550_
timestamp 1753371985
transform -1 0 38192 0 -1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2551_
timestamp 1751889408
transform 1 0 38192 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2552_
timestamp 1751534193
transform 1 0 38976 0 -1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2553_
timestamp 1751532043
transform -1 0 33152 0 1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _2554_
timestamp 1751905124
transform -1 0 35504 0 1 29792
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2555_
timestamp 1751889408
transform 1 0 31584 0 1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2556_
timestamp 1753277515
transform 1 0 32928 0 -1 31360
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2557_
timestamp 1753277515
transform 1 0 34496 0 -1 31360
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2558_
timestamp 1753277515
transform 1 0 35056 0 1 31360
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _2559_
timestamp 1753272495
transform -1 0 38192 0 1 29792
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2560_
timestamp 1751889808
transform 1 0 38528 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2561_
timestamp 1751534193
transform 1 0 35056 0 1 40768
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2562_
timestamp 1753371985
transform -1 0 37968 0 1 32928
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2563_
timestamp 1751889408
transform -1 0 33936 0 1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2564_
timestamp 1751534193
transform 1 0 34496 0 -1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2565_
timestamp 1751532043
transform 1 0 36064 0 1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2566_
timestamp 1753277515
transform 1 0 32928 0 -1 34496
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2567_
timestamp 1753277515
transform 1 0 32928 0 1 32928
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2568_
timestamp 1753277515
transform -1 0 36736 0 -1 34496
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _2569_
timestamp 1753272495
transform 1 0 35280 0 1 32928
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2570_
timestamp 1751889808
transform -1 0 35280 0 1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2571_
timestamp 1753371985
transform 1 0 36848 0 1 34496
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2572_
timestamp 1751889408
transform 1 0 36512 0 -1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2573_
timestamp 1751534193
transform -1 0 37408 0 -1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2574_
timestamp 1751532043
transform -1 0 34384 0 1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2575_
timestamp 1753277515
transform 1 0 34384 0 1 39200
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _2576_
timestamp 1753272495
transform -1 0 36512 0 -1 36064
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2577_
timestamp 1751889808
transform -1 0 35392 0 -1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2578_
timestamp 1753371985
transform 1 0 35392 0 -1 39200
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2579_
timestamp 1751889408
transform 1 0 36512 0 -1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2580_
timestamp 1751534193
transform -1 0 34160 0 1 40768
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2581_
timestamp 1751532043
transform -1 0 34832 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2582_
timestamp 1753277515
transform 1 0 34832 0 -1 42336
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _2583_
timestamp 1753272495
transform 1 0 35952 0 -1 40768
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2584_
timestamp 1751889808
transform -1 0 36512 0 1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2585_
timestamp 1753371985
transform -1 0 38864 0 -1 42336
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2586_
timestamp 1751889408
transform 1 0 36848 0 1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2587_
timestamp 1751534193
transform -1 0 34384 0 -1 42336
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2588_
timestamp 1751532043
transform 1 0 37856 0 -1 43904
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2589_
timestamp 1753277515
transform -1 0 36624 0 1 43904
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _2590_
timestamp 1753272495
transform 1 0 36400 0 -1 42336
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2591_
timestamp 1751889808
transform -1 0 35616 0 1 45472
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2592_
timestamp 1751534193
transform 1 0 39872 0 -1 43904
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2593_
timestamp 1753371985
transform 1 0 36848 0 1 40768
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2594_
timestamp 1751889408
transform 1 0 38640 0 1 45472
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2595_
timestamp 1751534193
transform -1 0 33488 0 1 40768
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2596_
timestamp 1751532043
transform -1 0 40432 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2597_
timestamp 1753277515
transform -1 0 39872 0 -1 43904
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _2598_
timestamp 1753272495
transform 1 0 36176 0 -1 45472
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2599_
timestamp 1751889808
transform 1 0 42448 0 1 45472
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2600_
timestamp 1753371985
transform 1 0 38864 0 -1 42336
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2601_
timestamp 1751889408
transform -1 0 40544 0 -1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2602_
timestamp 1751534193
transform -1 0 40320 0 1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2603_
timestamp 1751532043
transform -1 0 44352 0 1 43904
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2604_
timestamp 1753277515
transform -1 0 42336 0 -1 43904
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _2605_
timestamp 1753272495
transform 1 0 40768 0 -1 45472
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2606_
timestamp 1751889808
transform 1 0 46256 0 1 45472
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2607_
timestamp 1753371985
transform 1 0 41440 0 1 42336
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2608_
timestamp 1751889408
transform 1 0 47488 0 1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2609_
timestamp 1751534193
transform -1 0 28000 0 1 43904
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2610_
timestamp 1751531619
transform -1 0 43904 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2611_
timestamp 1751889808
transform 1 0 47488 0 1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _2612_
timestamp 1753272495
transform -1 0 43904 0 1 43904
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2613_
timestamp 1753371985
transform -1 0 44240 0 1 40768
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2614_
timestamp 1753960525
transform -1 0 43120 0 1 40768
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2615_
timestamp 1751740063
transform -1 0 42000 0 1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2616_
timestamp 1751531619
transform 1 0 42896 0 -1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2617_
timestamp 1753277515
transform 1 0 44352 0 -1 40768
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2618_
timestamp 1753371985
transform -1 0 48160 0 -1 40768
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2619_
timestamp 1751534193
transform 1 0 21168 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2620_
timestamp 1753960525
transform 1 0 45920 0 -1 40768
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2621_
timestamp 1751740063
transform -1 0 46704 0 -1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2622_
timestamp 1751532043
transform -1 0 44240 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2623_
timestamp 1753277515
transform 1 0 43792 0 -1 43904
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _2624_
timestamp 1753272495
transform -1 0 44128 0 1 42336
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _2625_
timestamp 1753272495
transform 1 0 42448 0 -1 43904
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2626_
timestamp 1751889808
transform 1 0 46704 0 -1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2627_
timestamp 1753371985
transform -1 0 48384 0 1 45472
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2628_
timestamp 1751889408
transform 1 0 47488 0 -1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2629_
timestamp 1751534193
transform -1 0 45360 0 1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _2630_
timestamp 1753272495
transform 1 0 44240 0 -1 42336
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2631_
timestamp 1751889408
transform 1 0 45136 0 -1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2632_
timestamp 1751534193
transform -1 0 28000 0 1 45472
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2633_
timestamp 1751534193
transform -1 0 45360 0 1 40768
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2634_
timestamp 1751534193
transform -1 0 41664 0 -1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2635_
timestamp 1751531619
transform -1 0 36512 0 1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _2636_
timestamp 1752061876
transform -1 0 44912 0 -1 31360
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2637_
timestamp 1751740063
transform -1 0 45472 0 1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2638_
timestamp 1753182340
transform 1 0 42896 0 1 29792
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2639_
timestamp 1751534193
transform 1 0 44688 0 1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2640_
timestamp 1751889408
transform -1 0 45024 0 -1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2641_
timestamp 1751534193
transform -1 0 43008 0 -1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2642_
timestamp 1751889408
transform -1 0 42896 0 1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2643_
timestamp 1751534193
transform 1 0 42112 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2644_
timestamp 1751889408
transform -1 0 42112 0 1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2645_
timestamp 1753960525
transform -1 0 39872 0 1 29792
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2646_
timestamp 1751534193
transform 1 0 42224 0 1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2647_
timestamp 1751534193
transform -1 0 40544 0 -1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2648_
timestamp 1751534193
transform -1 0 43456 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2649_
timestamp 1751534193
transform 1 0 41440 0 -1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2650_
timestamp 1753868718
transform -1 0 41440 0 1 31360
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2651_
timestamp 1753441877
transform 1 0 36400 0 -1 31360
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2652_
timestamp 1751889408
transform -1 0 39536 0 -1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2653_
timestamp 1751534193
transform -1 0 36624 0 1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2654_
timestamp 1753868718
transform 1 0 40768 0 -1 32928
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2655_
timestamp 1753441877
transform 1 0 38752 0 -1 32928
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2656_
timestamp 1751889408
transform 1 0 39536 0 -1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2657_
timestamp 1751534193
transform 1 0 40768 0 -1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2658_
timestamp 1751534193
transform -1 0 44128 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2659_
timestamp 1753868718
transform 1 0 41440 0 1 34496
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2660_
timestamp 1753441877
transform 1 0 37296 0 -1 36064
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2661_
timestamp 1751889408
transform -1 0 39200 0 -1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2662_
timestamp 1751534193
transform 1 0 40768 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2663_
timestamp 1751534193
transform 1 0 46032 0 1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2664_
timestamp 1753868718
transform -1 0 42560 0 1 36064
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2665_
timestamp 1753960525
transform 1 0 35056 0 1 36064
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2666_
timestamp 1751889408
transform 1 0 39200 0 -1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2667_
timestamp 1751534193
transform 1 0 41440 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2668_
timestamp 1751534193
transform 1 0 38864 0 -1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2669_
timestamp 1753868718
transform -1 0 41328 0 1 36064
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2670_
timestamp 1753441877
transform -1 0 37520 0 -1 37632
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2671_
timestamp 1751889408
transform -1 0 38304 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2672_
timestamp 1751534193
transform 1 0 38304 0 1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2673_
timestamp 1751534193
transform -1 0 34944 0 1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2674_
timestamp 1751534193
transform -1 0 42336 0 -1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2675_
timestamp 1753868718
transform -1 0 43120 0 1 37632
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2676_
timestamp 1753441877
transform 1 0 37744 0 -1 39200
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2677_
timestamp 1751889408
transform 1 0 38192 0 -1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2678_
timestamp 1751534193
transform 1 0 39536 0 -1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2679_
timestamp 1753868718
transform -1 0 41888 0 1 37632
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2680_
timestamp 1753960525
transform 1 0 36848 0 1 39200
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2681_
timestamp 1751889408
transform -1 0 39760 0 -1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2682_
timestamp 1751534193
transform 1 0 38976 0 1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2683_
timestamp 1753868718
transform 1 0 41440 0 -1 39200
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2684_
timestamp 1753441877
transform 1 0 41104 0 -1 40768
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2685_
timestamp 1751889408
transform 1 0 42224 0 -1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2686_
timestamp 1751534193
transform -1 0 34272 0 1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2687_
timestamp 1753868718
transform 1 0 44912 0 -1 39200
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2688_
timestamp 1753441877
transform 1 0 43232 0 -1 40768
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2689_
timestamp 1751889408
transform 1 0 45136 0 -1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2690_
timestamp 1751534193
transform 1 0 45360 0 1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2691_
timestamp 1753868718
transform -1 0 44912 0 -1 39200
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2692_
timestamp 1753441877
transform 1 0 46144 0 -1 39200
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2693_
timestamp 1751889408
transform -1 0 48048 0 -1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2694_
timestamp 1751534193
transform 1 0 29008 0 1 40768
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2695_
timestamp 1753868718
transform -1 0 44240 0 1 36064
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2696_
timestamp 1753868718
transform 1 0 42896 0 1 31360
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2697_
timestamp 1751534193
transform 1 0 44688 0 1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2698_
timestamp 1751740063
transform -1 0 8848 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2699_
timestamp 1751532043
transform -1 0 40544 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2700_
timestamp 1751532043
transform 1 0 20272 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2701_
timestamp 1751740063
transform -1 0 16688 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2702_
timestamp 1751534193
transform 1 0 23856 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2703_
timestamp 1751534193
transform -1 0 21616 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2704_
timestamp 1751534193
transform -1 0 17584 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2705_
timestamp 1753182340
transform -1 0 19936 0 1 18816
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2706_
timestamp 1751534193
transform -1 0 20272 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2707_
timestamp 1751531619
transform 1 0 26208 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2708_
timestamp 1751534193
transform 1 0 32704 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2709_
timestamp 1751532043
transform 1 0 22400 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2710_
timestamp 1751534193
transform 1 0 25872 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2711_
timestamp 1751534193
transform 1 0 26992 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2712_
timestamp 1753960525
transform 1 0 30128 0 -1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2713_
timestamp 1753371985
transform -1 0 40096 0 1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2714_
timestamp 1751532043
transform -1 0 41216 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2715_
timestamp 1751534193
transform 1 0 24304 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2716_
timestamp 1753960525
transform 1 0 29008 0 1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2717_
timestamp 1753371985
transform -1 0 38976 0 1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2718_
timestamp 1751532043
transform -1 0 34944 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2719_
timestamp 1753960525
transform 1 0 27664 0 1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2720_
timestamp 1753371985
transform -1 0 35728 0 1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2721_
timestamp 1751532043
transform -1 0 37296 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2722_
timestamp 1753960525
transform 1 0 26544 0 1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2723_
timestamp 1753371985
transform -1 0 37072 0 -1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2724_
timestamp 1751532043
transform -1 0 32592 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2725_
timestamp 1751534193
transform 1 0 26992 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2726_
timestamp 1751534193
transform 1 0 20160 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2727_
timestamp 1753960525
transform 1 0 25088 0 -1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2728_
timestamp 1753371985
transform -1 0 31584 0 1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2729_
timestamp 1751532043
transform -1 0 33824 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2730_
timestamp 1751532043
transform -1 0 25536 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2731_
timestamp 1751534193
transform -1 0 24976 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2732_
timestamp 1751534193
transform -1 0 24304 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2733_
timestamp 1753960525
transform 1 0 24304 0 1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2734_
timestamp 1753371985
transform -1 0 32704 0 1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2735_
timestamp 1751532043
transform 1 0 21168 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2736_
timestamp 1751534193
transform 1 0 20160 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2737_
timestamp 1751532043
transform 1 0 21168 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2738_
timestamp 1751740063
transform -1 0 17472 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2739_
timestamp 1751534193
transform -1 0 17024 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2740_
timestamp 1751531619
transform -1 0 23968 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2741_
timestamp 1753182340
transform 1 0 21616 0 -1 17248
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2742_
timestamp 1751534193
transform 1 0 29120 0 1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2743_
timestamp 1751532043
transform -1 0 33376 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2744_
timestamp 1751534193
transform 1 0 20048 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _2745_
timestamp 1753172561
transform 1 0 21616 0 1 17248
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2746_
timestamp 1751534193
transform 1 0 30800 0 -1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2747_
timestamp 1753441877
transform -1 0 32704 0 -1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2748_
timestamp 1753371985
transform 1 0 30688 0 1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2749_
timestamp 1751532043
transform -1 0 32592 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2750_
timestamp 1753441877
transform -1 0 32592 0 -1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2751_
timestamp 1753371985
transform 1 0 30352 0 -1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2752_
timestamp 1751532043
transform 1 0 32480 0 1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2753_
timestamp 1751534193
transform 1 0 29456 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2754_
timestamp 1753441877
transform 1 0 32928 0 -1 6272
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2755_
timestamp 1753371985
transform 1 0 29792 0 -1 6272
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2756_
timestamp 1751532043
transform -1 0 32480 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2757_
timestamp 1753441877
transform -1 0 32032 0 -1 4704
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2758_
timestamp 1753371985
transform 1 0 30912 0 -1 6272
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2759_
timestamp 1751532043
transform -1 0 32592 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2760_
timestamp 1753441877
transform -1 0 32144 0 -1 10976
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2761_
timestamp 1753371985
transform 1 0 29008 0 1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2762_
timestamp 1751532043
transform -1 0 30688 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2763_
timestamp 1753441877
transform 1 0 30688 0 -1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2764_
timestamp 1753371985
transform 1 0 29008 0 1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2765_
timestamp 1751532043
transform 1 0 20272 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2766_
timestamp 1751534193
transform 1 0 19488 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2767_
timestamp 1751531619
transform -1 0 20048 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2768_
timestamp 1751534193
transform 1 0 19824 0 -1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2769_
timestamp 1751534193
transform 1 0 20272 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2770_
timestamp 1753960525
transform -1 0 23744 0 -1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2771_
timestamp 1753371985
transform 1 0 19824 0 1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2772_
timestamp 1751532043
transform 1 0 18816 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2773_
timestamp 1753960525
transform -1 0 23408 0 1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2774_
timestamp 1753371985
transform 1 0 18704 0 -1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2775_
timestamp 1751532043
transform 1 0 18480 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2776_
timestamp 1751534193
transform -1 0 21840 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2777_
timestamp 1753960525
transform -1 0 22624 0 -1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2778_
timestamp 1753371985
transform 1 0 18592 0 1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2779_
timestamp 1751532043
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2780_
timestamp 1751534193
transform 1 0 23632 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2781_
timestamp 1753960525
transform 1 0 21168 0 1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2782_
timestamp 1753371985
transform 1 0 21168 0 1 10976
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2783_
timestamp 1751532043
transform 1 0 13440 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2784_
timestamp 1753960525
transform -1 0 22624 0 -1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2785_
timestamp 1753371985
transform 1 0 13776 0 -1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2786_
timestamp 1751532043
transform -1 0 14112 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2787_
timestamp 1753960525
transform -1 0 21504 0 -1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2788_
timestamp 1753371985
transform 1 0 14112 0 1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2789_
timestamp 1753960525
transform -1 0 24416 0 1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2790_
timestamp 1751534193
transform -1 0 19600 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2791_
timestamp 1753960525
transform -1 0 19376 0 1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2792_
timestamp 1751534193
transform -1 0 18928 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2793_
timestamp 1751531619
transform -1 0 19376 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2794_
timestamp 1751534193
transform 1 0 16800 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2795_
timestamp 1753960525
transform 1 0 17808 0 -1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2796_
timestamp 1753441877
transform 1 0 18704 0 1 25088
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2797_
timestamp 1751534193
transform 1 0 19824 0 1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2798_
timestamp 1751534193
transform -1 0 25760 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2799_
timestamp 1753960525
transform 1 0 17472 0 1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2800_
timestamp 1753441877
transform -1 0 19040 0 -1 25088
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2801_
timestamp 1751534193
transform -1 0 17920 0 -1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2802_
timestamp 1751534193
transform -1 0 27552 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2803_
timestamp 1753960525
transform 1 0 17472 0 1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2804_
timestamp 1753441877
transform -1 0 18816 0 -1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2805_
timestamp 1751534193
transform -1 0 17024 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2806_
timestamp 1751534193
transform -1 0 25200 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2807_
timestamp 1753960525
transform 1 0 18592 0 1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2808_
timestamp 1753441877
transform -1 0 19488 0 -1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2809_
timestamp 1751534193
transform -1 0 18368 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _2810_
timestamp 1752345181
transform -1 0 25424 0 1 20384
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _2811_
timestamp 1752345181
transform 1 0 21168 0 -1 18816
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2812_
timestamp 1751889808
transform 1 0 19040 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2813_
timestamp 1751534193
transform -1 0 21504 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_4  _2814_
timestamp 1753864693
transform -1 0 24192 0 1 20384
box -86 -86 2998 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2815_
timestamp 1753868718
transform -1 0 22736 0 -1 21952
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2816_
timestamp 1753441877
transform 1 0 24640 0 1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2817_
timestamp 1753441877
transform 1 0 25424 0 -1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2818_
timestamp 1751534193
transform 1 0 26880 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2819_
timestamp 1753441877
transform -1 0 24080 0 -1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2820_
timestamp 1753441877
transform 1 0 22960 0 1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2821_
timestamp 1751534193
transform 1 0 24080 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2822_
timestamp 1753441877
transform -1 0 27664 0 -1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2823_
timestamp 1753441877
transform 1 0 25648 0 -1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2824_
timestamp 1751534193
transform 1 0 26768 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2825_
timestamp 1751534193
transform -1 0 20496 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2826_
timestamp 1753441877
transform -1 0 22960 0 1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2827_
timestamp 1753441877
transform -1 0 22960 0 -1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2828_
timestamp 1751534193
transform 1 0 22288 0 -1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2829_
timestamp 1753960525
transform 1 0 24416 0 1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2830_
timestamp 1751534193
transform -1 0 14112 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2831_
timestamp 1753960525
transform -1 0 18704 0 1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2832_
timestamp 1751534193
transform -1 0 15232 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2833_
timestamp 1751531619
transform -1 0 16240 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2834_
timestamp 1751534193
transform -1 0 15904 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2835_
timestamp 1753960525
transform -1 0 15456 0 -1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2836_
timestamp 1753441877
transform -1 0 6944 0 -1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2837_
timestamp 1751534193
transform -1 0 2240 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2838_
timestamp 1753960525
transform -1 0 15232 0 1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2839_
timestamp 1753441877
transform -1 0 6720 0 1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2840_
timestamp 1751534193
transform -1 0 2688 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2841_
timestamp 1753960525
transform -1 0 14336 0 -1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2842_
timestamp 1753441877
transform 1 0 9744 0 1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2843_
timestamp 1751534193
transform -1 0 8848 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2844_
timestamp 1753960525
transform -1 0 16352 0 1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2845_
timestamp 1753441877
transform 1 0 7616 0 -1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2846_
timestamp 1751534193
transform -1 0 7616 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _2847_
timestamp 1752345181
transform -1 0 24640 0 -1 20384
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _2848_
timestamp 1752345181
transform -1 0 20944 0 1 17248
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_4  _2849_
timestamp 1753864693
transform -1 0 22736 0 -1 20384
box -86 -86 2998 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2850_
timestamp 1753868718
transform -1 0 20944 0 1 20384
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2851_
timestamp 1753441877
transform 1 0 13776 0 -1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2852_
timestamp 1753441877
transform -1 0 15680 0 -1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2853_
timestamp 1751534193
transform -1 0 10976 0 1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2854_
timestamp 1753441877
transform 1 0 13328 0 1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2855_
timestamp 1753441877
transform -1 0 15568 0 1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2856_
timestamp 1751534193
transform -1 0 10192 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2857_
timestamp 1753441877
transform 1 0 13440 0 -1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2858_
timestamp 1753441877
transform -1 0 15232 0 1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2859_
timestamp 1751534193
transform -1 0 9408 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2860_
timestamp 1753441877
transform 1 0 15568 0 1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2861_
timestamp 1753441877
transform -1 0 16912 0 -1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2862_
timestamp 1751534193
transform 1 0 16016 0 -1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2863_
timestamp 1751740063
transform -1 0 44464 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2864_
timestamp 1751889408
transform 1 0 47376 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2865_
timestamp 1751531619
transform 1 0 46592 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2866_
timestamp 1751740063
transform -1 0 47936 0 -1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2867_
timestamp 1751740063
transform -1 0 47152 0 -1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2868_
timestamp 1751889408
transform 1 0 47488 0 -1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2869_
timestamp 1753182340
transform 1 0 45472 0 -1 23520
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2870_
timestamp 1751534193
transform -1 0 45360 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2871_
timestamp 1751740063
transform 1 0 44576 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2872_
timestamp 1751889408
transform -1 0 47488 0 -1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2873_
timestamp 1753182340
transform 1 0 45360 0 1 23520
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2874_
timestamp 1751534193
transform 1 0 46256 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2875_
timestamp 1751740063
transform -1 0 46256 0 1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2876_
timestamp 1751889408
transform 1 0 46256 0 1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2877_
timestamp 1753182340
transform 1 0 43008 0 1 26656
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2878_
timestamp 1751534193
transform 1 0 43680 0 1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2879_
timestamp 1751531619
transform -1 0 47600 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2880_
timestamp 1751889808
transform 1 0 44688 0 1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2881_
timestamp 1751889408
transform 1 0 45472 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2882_
timestamp 1751889408
transform -1 0 45696 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2883_
timestamp 1751534193
transform -1 0 45360 0 1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2884_
timestamp 1753277515
transform 1 0 45248 0 -1 28224
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2885_
timestamp 1751889408
transform 1 0 45920 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2886_
timestamp 1751534193
transform 1 0 46704 0 -1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2887_
timestamp 1753441877
transform 1 0 22176 0 1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2888_
timestamp 1753371985
transform 1 0 22400 0 -1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2889_
timestamp 1753441877
transform 1 0 21728 0 -1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2890_
timestamp 1753371985
transform 1 0 19824 0 -1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2891_
timestamp 1753441877
transform -1 0 19376 0 -1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2892_
timestamp 1751740063
transform -1 0 19040 0 1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2893_
timestamp 1753960525
transform 1 0 27104 0 -1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2894_
timestamp 1753371985
transform -1 0 29008 0 -1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2895_
timestamp 1753960525
transform 1 0 28000 0 -1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2896_
timestamp 1753371985
transform -1 0 30128 0 1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2897_
timestamp 1753960525
transform -1 0 26992 0 -1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2898_
timestamp 1753441877
transform -1 0 14672 0 1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2899_
timestamp 1751534193
transform -1 0 14000 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2900_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751632746
transform 1 0 42560 0 -1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2901_
timestamp 1751632746
transform 1 0 45360 0 1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2902_
timestamp 1751632746
transform 1 0 45360 0 1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2903_
timestamp 1751632746
transform 1 0 45360 0 -1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2904_
timestamp 1751632746
transform 1 0 45360 0 1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2905_
timestamp 1751632746
transform 1 0 22288 0 1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2906_
timestamp 1751632746
transform 1 0 21840 0 -1 6272
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2907_
timestamp 1751632746
transform -1 0 21728 0 -1 6272
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2908_
timestamp 1751632746
transform -1 0 21952 0 -1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2909_
timestamp 1751632746
transform 1 0 27776 0 -1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2910_
timestamp 1751632746
transform 1 0 26880 0 -1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2911_
timestamp 1751632746
transform 1 0 26432 0 -1 6272
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2912_
timestamp 1751632746
transform 1 0 26768 0 -1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2913_
timestamp 1751632746
transform 1 0 35280 0 -1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2914_
timestamp 1751632746
transform 1 0 34944 0 -1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2915_
timestamp 1751632746
transform 1 0 32144 0 1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2916_
timestamp 1751632746
transform -1 0 32704 0 -1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2917_
timestamp 1751632746
transform 1 0 29680 0 -1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2918_
timestamp 1751632746
transform -1 0 34384 0 1 23520
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2919_
timestamp 1751632746
transform -1 0 38416 0 -1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2920_
timestamp 1751632746
transform -1 0 37856 0 -1 26656
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2921_
timestamp 1751632746
transform 1 0 25312 0 -1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2922_
timestamp 1751632746
transform 1 0 21728 0 -1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2923_
timestamp 1751632746
transform 1 0 22848 0 1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2924_
timestamp 1751632746
transform 1 0 22736 0 1 39200
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2925_
timestamp 1751632746
transform 1 0 22736 0 1 42336
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2926_
timestamp 1751632746
transform 1 0 25200 0 -1 45472
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2927_
timestamp 1751632746
transform 1 0 21728 0 -1 45472
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2928_
timestamp 1751632746
transform 1 0 1568 0 -1 28224
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2929_
timestamp 1751632746
transform -1 0 4592 0 1 28224
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2930_
timestamp 1751632746
transform 1 0 1568 0 -1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2931_
timestamp 1751632746
transform 1 0 1568 0 1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2932_
timestamp 1751632746
transform 1 0 6160 0 -1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2933_
timestamp 1751632746
transform 1 0 9408 0 -1 39200
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2934_
timestamp 1751632746
transform 1 0 1568 0 1 39200
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2935_
timestamp 1751632746
transform 1 0 1568 0 -1 42336
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2936_
timestamp 1751632746
transform 1 0 2240 0 1 43904
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2937_
timestamp 1751632746
transform 1 0 6160 0 -1 45472
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2938_
timestamp 1751632746
transform 1 0 10304 0 -1 45472
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2939_
timestamp 1751632746
transform 1 0 6160 0 1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2940_
timestamp 1751632746
transform 1 0 5488 0 1 29792
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2941_
timestamp 1751632746
transform 1 0 9184 0 1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2942_
timestamp 1751632746
transform 1 0 1568 0 -1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2943_
timestamp 1751632746
transform 1 0 1568 0 -1 37632
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2944_
timestamp 1751632746
transform -1 0 7952 0 -1 39200
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2945_
timestamp 1751632746
transform 1 0 5488 0 1 40768
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2946_
timestamp 1751632746
transform 1 0 9072 0 1 42336
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2947_
timestamp 1751632746
transform -1 0 19488 0 1 40768
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2948_
timestamp 1751632746
transform -1 0 17696 0 1 43904
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2949_
timestamp 1751632746
transform -1 0 16352 0 -1 45472
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2950_
timestamp 1751632746
transform 1 0 13328 0 -1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2951_
timestamp 1751632746
transform 1 0 9408 0 -1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2952_
timestamp 1751632746
transform 1 0 9296 0 1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2953_
timestamp 1751632746
transform 1 0 5152 0 -1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2954_
timestamp 1751632746
transform 1 0 2240 0 1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2955_
timestamp 1751632746
transform 1 0 2016 0 1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2956_
timestamp 1751632746
transform 1 0 3920 0 -1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2957_
timestamp 1751632746
transform 1 0 1792 0 1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2958_
timestamp 1751632746
transform 1 0 1568 0 1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2959_
timestamp 1751632746
transform 1 0 1568 0 -1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2960_
timestamp 1751632746
transform 1 0 3248 0 -1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2961_
timestamp 1751632746
transform 1 0 4816 0 -1 6272
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2962_
timestamp 1751632746
transform 1 0 7056 0 1 6272
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2963_
timestamp 1751632746
transform -1 0 11872 0 1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2964_
timestamp 1751632746
transform 1 0 6160 0 -1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2965_
timestamp 1751632746
transform -1 0 12208 0 1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2966_
timestamp 1751632746
transform 1 0 40768 0 -1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2967_
timestamp 1751632746
transform -1 0 44912 0 -1 23520
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2968_
timestamp 1751632746
transform 1 0 40656 0 1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2969_
timestamp 1751632746
transform 1 0 38416 0 1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2970_
timestamp 1751632746
transform 1 0 34944 0 -1 23520
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2971_
timestamp 1751632746
transform 1 0 33376 0 -1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2972_
timestamp 1751632746
transform -1 0 36624 0 1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2973_
timestamp 1751632746
transform 1 0 37632 0 1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2974_
timestamp 1751632746
transform 1 0 22512 0 1 29792
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2975_
timestamp 1751632746
transform 1 0 21728 0 1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2976_
timestamp 1751632746
transform 1 0 15008 0 1 29792
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2977_
timestamp 1751632746
transform 1 0 14000 0 -1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2978_
timestamp 1751632746
transform 1 0 15568 0 1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2979_
timestamp 1751632746
transform 1 0 17472 0 -1 39200
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2980_
timestamp 1751632746
transform 1 0 17808 0 1 39200
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2981_
timestamp 1751632746
transform 1 0 17584 0 -1 42336
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2982_
timestamp 1751632746
transform 1 0 17696 0 1 43904
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2983_
timestamp 1751632746
transform -1 0 20832 0 -1 45472
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2984_
timestamp 1751632746
transform 1 0 38192 0 1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2985_
timestamp 1751632746
transform -1 0 43904 0 -1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2986_
timestamp 1751632746
transform 1 0 45024 0 -1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2987_
timestamp 1751632746
transform 1 0 45360 0 1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2988_
timestamp 1751632746
transform 1 0 45360 0 1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2989_
timestamp 1751632746
transform -1 0 46816 0 -1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2990_
timestamp 1751632746
transform -1 0 48384 0 -1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2991_
timestamp 1751632746
transform 1 0 45360 0 1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2992_
timestamp 1751632746
transform 1 0 40768 0 -1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2993_
timestamp 1751632746
transform 1 0 37856 0 1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2994_
timestamp 1751632746
transform -1 0 39872 0 1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2995_
timestamp 1751632746
transform 1 0 35392 0 -1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2996_
timestamp 1751632746
transform 1 0 44688 0 1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2997_
timestamp 1751632746
transform -1 0 48384 0 -1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2998_
timestamp 1751632746
transform -1 0 48384 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2999_
timestamp 1751632746
transform 1 0 42672 0 -1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3000_
timestamp 1751632746
transform -1 0 43904 0 -1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3001_
timestamp 1751632746
transform 1 0 36624 0 -1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3002_
timestamp 1751632746
transform 1 0 33600 0 -1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3003_
timestamp 1751632746
transform 1 0 36624 0 -1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3004_
timestamp 1751632746
transform 1 0 32928 0 -1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3005_
timestamp 1751632746
transform 1 0 3024 0 -1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3006_
timestamp 1751632746
transform -1 0 36288 0 1 6272
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3007_
timestamp 1751632746
transform 1 0 23408 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3008_
timestamp 1751632746
transform 1 0 19600 0 -1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3009_
timestamp 1751632746
transform 1 0 15232 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3010_
timestamp 1751632746
transform 1 0 10080 0 1 6272
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3011_
timestamp 1751632746
transform 1 0 15568 0 1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3012_
timestamp 1751632746
transform 1 0 11872 0 -1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3013_
timestamp 1751632746
transform 1 0 10640 0 -1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3014_
timestamp 1751632746
transform 1 0 10080 0 1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3015_
timestamp 1751632746
transform 1 0 15456 0 1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3016_
timestamp 1751632746
transform 1 0 9408 0 1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3017_
timestamp 1751632746
transform -1 0 43344 0 1 28224
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3018_
timestamp 1751632746
transform -1 0 40320 0 1 28224
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3019_
timestamp 1751632746
transform -1 0 35952 0 -1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3020_
timestamp 1751632746
transform 1 0 33040 0 1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3021_
timestamp 1751632746
transform 1 0 32928 0 -1 40768
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3022_
timestamp 1751632746
transform 1 0 32704 0 1 42336
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3023_
timestamp 1751632746
transform 1 0 33040 0 -1 45472
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3024_
timestamp 1751632746
transform 1 0 37520 0 -1 45472
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3025_
timestamp 1751632746
transform 1 0 42224 0 -1 45472
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3026_
timestamp 1751632746
transform 1 0 40768 0 -1 42336
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3027_
timestamp 1751632746
transform 1 0 45360 0 1 40768
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3028_
timestamp 1751632746
transform 1 0 45360 0 -1 43904
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3029_
timestamp 1751632746
transform 1 0 45360 0 -1 45472
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3030_
timestamp 1751632746
transform 1 0 29680 0 -1 45472
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3031_
timestamp 1751632746
transform -1 0 45472 0 -1 29792
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3032_
timestamp 1751632746
transform -1 0 43792 0 -1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3033_
timestamp 1751632746
transform 1 0 37520 0 -1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3034_
timestamp 1751632746
transform 1 0 38080 0 1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3035_
timestamp 1751632746
transform 1 0 38416 0 1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3036_
timestamp 1751632746
transform 1 0 36848 0 1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3037_
timestamp 1751632746
transform 1 0 37520 0 -1 37632
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3038_
timestamp 1751632746
transform 1 0 38192 0 1 39200
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3039_
timestamp 1751632746
transform 1 0 38080 0 1 40768
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3040_
timestamp 1751632746
transform 1 0 41328 0 1 39200
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3041_
timestamp 1751632746
transform 1 0 45360 0 1 39200
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3042_
timestamp 1751632746
transform 1 0 45360 0 1 37632
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3043_
timestamp 1751632746
transform -1 0 45024 0 -1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3044_
timestamp 1751632746
transform -1 0 40880 0 1 42336
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3045_
timestamp 1751632746
transform 1 0 6384 0 1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3046_
timestamp 1751632746
transform 1 0 37520 0 -1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3047_
timestamp 1751632746
transform 1 0 37632 0 1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3048_
timestamp 1751632746
transform 1 0 32928 0 -1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3049_
timestamp 1751632746
transform 1 0 33600 0 1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3050_
timestamp 1751632746
transform 1 0 30688 0 1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3051_
timestamp 1751632746
transform 1 0 32928 0 -1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3052_
timestamp 1751632746
transform 1 0 30688 0 1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3053_
timestamp 1751632746
transform 1 0 30240 0 1 6272
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3054_
timestamp 1751632746
transform 1 0 29456 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3055_
timestamp 1751632746
transform 1 0 28784 0 1 3136
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3056_
timestamp 1751632746
transform 1 0 28000 0 -1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3057_
timestamp 1751632746
transform 1 0 27664 0 -1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3058_
timestamp 1751632746
transform -1 0 22064 0 -1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3059_
timestamp 1751632746
transform -1 0 20384 0 1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3060_
timestamp 1751632746
transform -1 0 18928 0 1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3061_
timestamp 1751632746
transform -1 0 22624 0 -1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3062_
timestamp 1751632746
transform 1 0 10752 0 -1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3063_
timestamp 1751632746
transform 1 0 11536 0 -1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3064_
timestamp 1751632746
transform 1 0 19264 0 -1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3065_
timestamp 1751632746
transform 1 0 15680 0 1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3066_
timestamp 1751632746
transform 1 0 15456 0 1 26656
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3067_
timestamp 1751632746
transform 1 0 17920 0 1 23520
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3068_
timestamp 1751632746
transform 1 0 25760 0 1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3069_
timestamp 1751632746
transform 1 0 22848 0 1 23520
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3070_
timestamp 1751632746
transform 1 0 25760 0 1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3071_
timestamp 1751632746
transform 1 0 21504 0 1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3072_
timestamp 1751632746
transform 1 0 1568 0 1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3073_
timestamp 1751632746
transform 1 0 1568 0 -1 23520
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3074_
timestamp 1751632746
transform -1 0 9744 0 1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3075_
timestamp 1751632746
transform 1 0 2240 0 -1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3076_
timestamp 1751632746
transform 1 0 9632 0 -1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3077_
timestamp 1751632746
transform 1 0 9408 0 -1 23520
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3078_
timestamp 1751632746
transform 1 0 9632 0 -1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3079_
timestamp 1751632746
transform -1 0 17920 0 1 23520
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3080_
timestamp 1751632746
transform 1 0 44688 0 1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3081_
timestamp 1751632746
transform 1 0 45360 0 -1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3082_
timestamp 1751632746
transform 1 0 45024 0 1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3083_
timestamp 1751632746
transform 1 0 45360 0 -1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3084_
timestamp 1751632746
transform 1 0 42448 0 -1 26656
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3085_
timestamp 1751632746
transform 1 0 42000 0 -1 28224
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3086_
timestamp 1751632746
transform -1 0 48384 0 1 28224
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3087_
timestamp 1751632746
transform 1 0 15232 0 1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3088_
timestamp 1751632746
transform 1 0 18704 0 -1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3089_
timestamp 1751632746
transform 1 0 15232 0 1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3090_
timestamp 1751632746
transform 1 0 29008 0 1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3091_
timestamp 1751632746
transform 1 0 29008 0 -1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _3092_
timestamp 1751632746
transform 1 0 10080 0 1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _3105_
timestamp 1751534193
transform -1 0 13104 0 1 43904
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _3106_
timestamp 1751534193
transform 1 0 13104 0 1 45472
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _3107_
timestamp 1751534193
transform 1 0 24416 0 1 45472
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _3108_
timestamp 1751534193
transform -1 0 17024 0 -1 45472
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _3109_
timestamp 1751534193
transform 1 0 20720 0 1 45472
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _3110_
timestamp 1751534193
transform 1 0 30576 0 1 45472
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _3111_
timestamp 1751534193
transform 1 0 32928 0 -1 42336
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _3112_
timestamp 1751534193
transform -1 0 34832 0 1 40768
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1465__A dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532392
transform -1 0 7616 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1466__B
timestamp 1751532392
transform 1 0 22176 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1470__B
timestamp 1751532392
transform 1 0 16912 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1474__B
timestamp 1751532392
transform 1 0 17360 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1477__B
timestamp 1751532392
transform 1 0 16800 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1479__C
timestamp 1751532392
transform -1 0 17696 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1564__A
timestamp 1751532392
transform 1 0 16128 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1603__A
timestamp 1751532392
transform 1 0 32480 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1618__A
timestamp 1751532392
transform 1 0 32928 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1618__C
timestamp 1751532392
transform -1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1619__A
timestamp 1751532392
transform 1 0 30464 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1689__A
timestamp 1751532392
transform 1 0 9632 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1689__B
timestamp 1751532392
transform 1 0 15120 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1690__A
timestamp 1751532392
transform 1 0 17472 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1690__B
timestamp 1751532392
transform 1 0 11760 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1714__A
timestamp 1751532392
transform 1 0 9632 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1715__A
timestamp 1751532392
transform 1 0 10080 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1740__A
timestamp 1751532392
transform 1 0 11536 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1758__A
timestamp 1751532392
transform -1 0 5488 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1758__B
timestamp 1751532392
transform -1 0 8400 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1759__B
timestamp 1751532392
transform 1 0 10528 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1771__A
timestamp 1751532392
transform -1 0 3808 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1772__A
timestamp 1751532392
transform -1 0 6384 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1780__A
timestamp 1751532392
transform -1 0 38304 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1781__A
timestamp 1751532392
transform 1 0 45136 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1782__A
timestamp 1751532392
transform 1 0 40096 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1787__A
timestamp 1751532392
transform 1 0 31472 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1789__A
timestamp 1751532392
transform 1 0 40208 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1805__A
timestamp 1751532392
transform -1 0 22400 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1806__A
timestamp 1751532392
transform 1 0 20944 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1807__A
timestamp 1751532392
transform 1 0 15680 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1810__A
timestamp 1751532392
transform 1 0 28784 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1811__A
timestamp 1751532392
transform -1 0 22848 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1815__A
timestamp 1751532392
transform -1 0 27440 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1817__A
timestamp 1751532392
transform 1 0 19824 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1820__A
timestamp 1751532392
transform 1 0 25536 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1820__D
timestamp 1751532392
transform 1 0 23968 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1824__A
timestamp 1751532392
transform -1 0 22176 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1834__A
timestamp 1751532392
transform 1 0 27552 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1839__A
timestamp 1751532392
transform 1 0 29344 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1844__A
timestamp 1751532392
transform -1 0 28000 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1848__A
timestamp 1751532392
transform 1 0 27552 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1848__D
timestamp 1751532392
transform 1 0 25984 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1862__A
timestamp 1751532392
transform -1 0 26768 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1865__A
timestamp 1751532392
transform 1 0 27552 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1866__A
timestamp 1751532392
transform 1 0 25648 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1866__D
timestamp 1751532392
transform 1 0 26096 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1881__A
timestamp 1751532392
transform 1 0 34384 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1884__A
timestamp 1751532392
transform -1 0 33376 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1891__D
timestamp 1751532392
transform 1 0 30912 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1899__A
timestamp 1751532392
transform 1 0 26656 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1900__C
timestamp 1751532392
transform -1 0 35392 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1907__C
timestamp 1751532392
transform 1 0 34496 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1913__C
timestamp 1751532392
transform 1 0 27328 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1919__A
timestamp 1751532392
transform -1 0 41328 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1920__A
timestamp 1751532392
transform 1 0 25312 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1922__A
timestamp 1751532392
transform -1 0 25536 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1927__A
timestamp 1751532392
transform 1 0 16352 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1928__C
timestamp 1751532392
transform 1 0 26208 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1932__A
timestamp 1751532392
transform 1 0 24528 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1938__A
timestamp 1751532392
transform 1 0 23408 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1945__A
timestamp 1751532392
transform 1 0 23408 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1952__C
timestamp 1751532392
transform 1 0 24640 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1956__A
timestamp 1751532392
transform 1 0 30576 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1961__D
timestamp 1751532392
transform -1 0 7616 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1965__A
timestamp 1751532392
transform 1 0 7056 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1972__A
timestamp 1751532392
transform 1 0 3584 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1978__C
timestamp 1751532392
transform -1 0 3808 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1986__C
timestamp 1751532392
transform 1 0 8512 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1994__A
timestamp 1751532392
transform 1 0 8960 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1997__B
timestamp 1751532392
transform 1 0 3360 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2000__A
timestamp 1751532392
transform -1 0 16128 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2001__C
timestamp 1751532392
transform -1 0 3024 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2004__B
timestamp 1751532392
transform -1 0 2128 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2005__B
timestamp 1751532392
transform -1 0 2128 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2008__A
timestamp 1751532392
transform 1 0 2912 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2012__B
timestamp 1751532392
transform -1 0 3248 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2013__B
timestamp 1751532392
transform -1 0 2912 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2017__A
timestamp 1751532392
transform -1 0 5152 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2022__B
timestamp 1751532392
transform -1 0 2464 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2024__C
timestamp 1751532392
transform -1 0 3360 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2028__A
timestamp 1751532392
transform -1 0 4592 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2032__A
timestamp 1751532392
transform 1 0 6608 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2036__C
timestamp 1751532392
transform 1 0 7616 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2042__C
timestamp 1751532392
transform 1 0 11200 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2049__A
timestamp 1751532392
transform -1 0 17920 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2050__C
timestamp 1751532392
transform 1 0 5712 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2057__C
timestamp 1751532392
transform 1 0 5712 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2064__A
timestamp 1751532392
transform -1 0 9184 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2067__B
timestamp 1751532392
transform 1 0 6160 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2070__C
timestamp 1751532392
transform -1 0 3360 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2074__B
timestamp 1751532392
transform -1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2077__A
timestamp 1751532392
transform 1 0 8848 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2086__A
timestamp 1751532392
transform 1 0 18144 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2093__C
timestamp 1751532392
transform 1 0 16800 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2097__A
timestamp 1751532392
transform -1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2100__A
timestamp 1751532392
transform -1 0 16576 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2109__B
timestamp 1751532392
transform -1 0 9856 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2111__A
timestamp 1751532392
transform -1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2112__B
timestamp 1751532392
transform -1 0 4480 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2186__A
timestamp 1751532392
transform 1 0 32480 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2187__A
timestamp 1751532392
transform 1 0 47712 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2189__D
timestamp 1751532392
transform 1 0 48048 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2192__A
timestamp 1751532392
transform 1 0 36400 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2193__B
timestamp 1751532392
transform 1 0 43792 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2195__A
timestamp 1751532392
transform -1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2199__A
timestamp 1751532392
transform -1 0 41552 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2204__A
timestamp 1751532392
transform 1 0 37408 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2208__A
timestamp 1751532392
transform 1 0 41440 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2212__A
timestamp 1751532392
transform 1 0 36176 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2216__A
timestamp 1751532392
transform 1 0 37856 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2220__A
timestamp 1751532392
transform 1 0 34048 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2222__B
timestamp 1751532392
transform 1 0 38304 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2223__A
timestamp 1751532392
transform 1 0 40320 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2224__B
timestamp 1751532392
transform 1 0 39984 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2230__A
timestamp 1751532392
transform -1 0 17472 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2259__A
timestamp 1751532392
transform 1 0 20048 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2265__A
timestamp 1751532392
transform 1 0 21504 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2274__A
timestamp 1751532392
transform -1 0 23072 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2303__A
timestamp 1751532392
transform 1 0 32480 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2304__A
timestamp 1751532392
transform 1 0 37632 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2304__C
timestamp 1751532392
transform 1 0 37296 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2308__A
timestamp 1751532392
transform 1 0 34048 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2315__B
timestamp 1751532392
transform 1 0 44912 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2316__A
timestamp 1751532392
transform 1 0 48048 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2317__A
timestamp 1751532392
transform 1 0 44240 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2322__B
timestamp 1751532392
transform -1 0 44688 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2324__A
timestamp 1751532392
transform 1 0 44016 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2325__A
timestamp 1751532392
transform -1 0 37296 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2333__A
timestamp 1751532392
transform 1 0 47824 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2350__A
timestamp 1751532392
transform 1 0 47488 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2362__A
timestamp 1751532392
transform 1 0 33600 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2374__A
timestamp 1751532392
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2377__A
timestamp 1751532392
transform 1 0 35728 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2379__A
timestamp 1751532392
transform 1 0 42560 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2379__D
timestamp 1751532392
transform -1 0 37744 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2393__A
timestamp 1751532392
transform -1 0 39312 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2393__C
timestamp 1751532392
transform -1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2401__A
timestamp 1751532392
transform 1 0 26432 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2423__A
timestamp 1751532392
transform 1 0 29232 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2425__A
timestamp 1751532392
transform -1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2437__A
timestamp 1751532392
transform -1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2439__A
timestamp 1751532392
transform 1 0 47376 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2440__A
timestamp 1751532392
transform 1 0 46144 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2446__A
timestamp 1751532392
transform -1 0 32928 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2447__A
timestamp 1751532392
transform 1 0 30688 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2456__A
timestamp 1751532392
transform 1 0 33376 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2457__D
timestamp 1751532392
transform 1 0 36400 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2461__B
timestamp 1751532392
transform -1 0 4368 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2462__A
timestamp 1751532392
transform -1 0 4144 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2463__B
timestamp 1751532392
transform 1 0 4592 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2472__A
timestamp 1751532392
transform 1 0 38640 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2472__C
timestamp 1751532392
transform 1 0 36400 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2479__A
timestamp 1751532392
transform -1 0 24976 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2480__A
timestamp 1751532392
transform -1 0 26992 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2485__A
timestamp 1751532392
transform -1 0 19600 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2488__A
timestamp 1751532392
transform -1 0 22960 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2489__A
timestamp 1751532392
transform -1 0 12320 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2495__A
timestamp 1751532392
transform -1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2509__B
timestamp 1751532392
transform -1 0 17808 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2510__A
timestamp 1751532392
transform -1 0 18256 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2511__A
timestamp 1751532392
transform -1 0 17696 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2522__A
timestamp 1751532392
transform -1 0 12208 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2528__B
timestamp 1751532392
transform 1 0 16688 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2529__A
timestamp 1751532392
transform 1 0 16240 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2530__A
timestamp 1751532392
transform -1 0 15680 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2533__B
timestamp 1751532392
transform 1 0 20720 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2534__A
timestamp 1751532392
transform 1 0 18480 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2535__A
timestamp 1751532392
transform -1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2536__A
timestamp 1751532392
transform 1 0 13664 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2537__B
timestamp 1751532392
transform 1 0 22848 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2537__D
timestamp 1751532392
transform -1 0 12656 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2539__A
timestamp 1751532392
transform 1 0 48160 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2540__A
timestamp 1751532392
transform 1 0 32480 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2541__A
timestamp 1751532392
transform 1 0 35392 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2550__C
timestamp 1751532392
transform -1 0 37072 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2561__A
timestamp 1751532392
transform 1 0 37520 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2592__A
timestamp 1751532392
transform 1 0 32032 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2609__A
timestamp 1751532392
transform -1 0 27888 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2610__B
timestamp 1751532392
transform 1 0 22736 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2611__B
timestamp 1751532392
transform -1 0 24752 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2614__D
timestamp 1751532392
transform 1 0 25760 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2620__D
timestamp 1751532392
transform 1 0 30128 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2623__B
timestamp 1751532392
transform -1 0 2912 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2630__B
timestamp 1751532392
transform 1 0 25088 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2631__A
timestamp 1751532392
transform 1 0 26880 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2632__A
timestamp 1751532392
transform -1 0 17808 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2635__A
timestamp 1751532392
transform -1 0 25760 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2637__A
timestamp 1751532392
transform 1 0 45808 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2642__A
timestamp 1751532392
transform -1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2668__A
timestamp 1751532392
transform 1 0 30352 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2688__A
timestamp 1751532392
transform 1 0 27104 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2689__A
timestamp 1751532392
transform -1 0 19824 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2693__A
timestamp 1751532392
transform 1 0 23520 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2694__A
timestamp 1751532392
transform -1 0 27664 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2695__A
timestamp 1751532392
transform 1 0 24640 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2698__A
timestamp 1751532392
transform -1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2698__B
timestamp 1751532392
transform -1 0 5824 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2701__B
timestamp 1751532392
transform -1 0 15904 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2705__C
timestamp 1751532392
transform -1 0 19824 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2709__A
timestamp 1751532392
transform -1 0 23296 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2730__A
timestamp 1751532392
transform 1 0 28336 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2736__A
timestamp 1751532392
transform -1 0 16912 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2738__B
timestamp 1751532392
transform 1 0 15232 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2746__A
timestamp 1751532392
transform -1 0 30688 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2747__C
timestamp 1751532392
transform 1 0 33600 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2750__C
timestamp 1751532392
transform 1 0 33936 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2753__A
timestamp 1751532392
transform 1 0 29232 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2760__B
timestamp 1751532392
transform 1 0 30464 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2763__B
timestamp 1751532392
transform 1 0 30016 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2789__A
timestamp 1751532392
transform 1 0 23072 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2795__A
timestamp 1751532392
transform -1 0 17808 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2798__A
timestamp 1751532392
transform 1 0 25648 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2802__A
timestamp 1751532392
transform 1 0 27664 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2806__A
timestamp 1751532392
transform -1 0 23520 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2810__A
timestamp 1751532392
transform 1 0 24192 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2812__A
timestamp 1751532392
transform 1 0 16800 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2816__C
timestamp 1751532392
transform 1 0 24416 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2817__A
timestamp 1751532392
transform -1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2819__C
timestamp 1751532392
transform -1 0 23184 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2822__C
timestamp 1751532392
transform -1 0 28112 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2829__C
timestamp 1751532392
transform -1 0 28448 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2835__A
timestamp 1751532392
transform 1 0 15456 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2850__A
timestamp 1751532392
transform 1 0 20160 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2852__A
timestamp 1751532392
transform -1 0 16128 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2860__C
timestamp 1751532392
transform 1 0 16912 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2863__B
timestamp 1751532392
transform 1 0 31136 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2865__A
timestamp 1751532392
transform 1 0 47040 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2877__A
timestamp 1751532392
transform 1 0 44240 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2885__A
timestamp 1751532392
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2891__C
timestamp 1751532392
transform 1 0 16128 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2895__D
timestamp 1751532392
transform 1 0 28448 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2897__A
timestamp 1751532392
transform -1 0 26208 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2897__D
timestamp 1751532392
transform -1 0 24528 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2900__CLK
timestamp 1751532392
transform 1 0 32480 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2901__CLK
timestamp 1751532392
transform 1 0 26208 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2902__CLK
timestamp 1751532392
transform 1 0 31024 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2903__CLK
timestamp 1751532392
transform 1 0 33376 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2904__CLK
timestamp 1751532392
transform 1 0 32032 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2905__CLK
timestamp 1751532392
transform 1 0 22288 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2906__CLK
timestamp 1751532392
transform 1 0 20720 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2907__CLK
timestamp 1751532392
transform 1 0 20384 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2908__CLK
timestamp 1751532392
transform 1 0 19936 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2909__CLK
timestamp 1751532392
transform 1 0 30016 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2910__CLK
timestamp 1751532392
transform 1 0 30128 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2911__CLK
timestamp 1751532392
transform 1 0 29680 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2912__CLK
timestamp 1751532392
transform 1 0 30016 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2914__CLK
timestamp 1751532392
transform 1 0 39312 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2918__CLK
timestamp 1751532392
transform 1 0 33936 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2919__CLK
timestamp 1751532392
transform 1 0 40208 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2920__CLK
timestamp 1751532392
transform 1 0 38080 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2921__CLK
timestamp 1751532392
transform 1 0 28896 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2922__CLK
timestamp 1751532392
transform -1 0 23632 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2926__CLK
timestamp 1751532392
transform 1 0 28896 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2928__CLK
timestamp 1751532392
transform 1 0 4816 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2929__CLK
timestamp 1751532392
transform 1 0 2016 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2930__CLK
timestamp 1751532392
transform 1 0 4032 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2931__CLK
timestamp 1751532392
transform 1 0 3136 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2932__CLK
timestamp 1751532392
transform 1 0 8064 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2933__CLK
timestamp 1751532392
transform 1 0 10528 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2934__CLK
timestamp 1751532392
transform 1 0 2352 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2935__CLK
timestamp 1751532392
transform 1 0 2016 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2936__CLK
timestamp 1751532392
transform -1 0 3248 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2937__CLK
timestamp 1751532392
transform -1 0 4704 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2938__CLK
timestamp 1751532392
transform -1 0 6832 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2939__CLK
timestamp 1751532392
transform 1 0 5040 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2940__CLK
timestamp 1751532392
transform 1 0 7392 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2941__CLK
timestamp 1751532392
transform -1 0 11200 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2942__CLK
timestamp 1751532392
transform 1 0 6160 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2943__CLK
timestamp 1751532392
transform 1 0 4592 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2944__CLK
timestamp 1751532392
transform 1 0 9408 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2945__CLK
timestamp 1751532392
transform 1 0 6384 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2946__CLK
timestamp 1751532392
transform -1 0 9968 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2950__CLK
timestamp 1751532392
transform 1 0 14896 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2951__CLK
timestamp 1751532392
transform -1 0 8736 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2954__CLK
timestamp 1751532392
transform 1 0 3808 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2955__CLK
timestamp 1751532392
transform 1 0 4816 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2956__CLK
timestamp 1751532392
transform 1 0 7168 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2957__CLK
timestamp 1751532392
transform 1 0 5040 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2958__CLK
timestamp 1751532392
transform 1 0 4816 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2959__CLK
timestamp 1751532392
transform 1 0 3472 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2960__CLK
timestamp 1751532392
transform 1 0 5712 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2961__CLK
timestamp 1751532392
transform 1 0 8064 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2962__CLK
timestamp 1751532392
transform 1 0 10304 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2963__CLK
timestamp 1751532392
transform 1 0 11312 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2964__CLK
timestamp 1751532392
transform 1 0 10416 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2965__CLK
timestamp 1751532392
transform 1 0 11200 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2967__CLK
timestamp 1751532392
transform 1 0 36400 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2968__CLK
timestamp 1751532392
transform 1 0 48160 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2970__CLK
timestamp 1751532392
transform 1 0 38528 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2973__CLK
timestamp 1751532392
transform 1 0 42448 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2974__CLK
timestamp 1751532392
transform 1 0 23744 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2975__CLK
timestamp 1751532392
transform 1 0 20720 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2976__CLK
timestamp 1751532392
transform 1 0 18256 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2977__CLK
timestamp 1751532392
transform 1 0 13776 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2978__CLK
timestamp 1751532392
transform -1 0 17920 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2988__CLK
timestamp 1751532392
transform 1 0 48160 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2989__CLK
timestamp 1751532392
transform -1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2990__CLK
timestamp 1751532392
transform 1 0 45024 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2991__CLK
timestamp 1751532392
transform -1 0 47712 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2992__CLK
timestamp 1751532392
transform -1 0 45472 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2993__CLK
timestamp 1751532392
transform 1 0 42336 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2995__CLK
timestamp 1751532392
transform -1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2996__CLK
timestamp 1751532392
transform 1 0 27888 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2997__CLK
timestamp 1751532392
transform -1 0 26880 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2998__CLK
timestamp 1751532392
transform 1 0 28560 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2999__CLK
timestamp 1751532392
transform 1 0 28560 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3000__CLK
timestamp 1751532392
transform -1 0 46816 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3001__CLK
timestamp 1751532392
transform -1 0 48160 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3002__CLK
timestamp 1751532392
transform -1 0 33376 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3003__CLK
timestamp 1751532392
transform 1 0 42448 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3004__CLK
timestamp 1751532392
transform 1 0 33152 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3006__CLK
timestamp 1751532392
transform -1 0 36512 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3007__CLK
timestamp 1751532392
transform -1 0 23408 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3008__CLK
timestamp 1751532392
transform -1 0 17360 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3009__CLK
timestamp 1751532392
transform -1 0 14336 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3010__CLK
timestamp 1751532392
transform 1 0 11984 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3011__CLK
timestamp 1751532392
transform 1 0 19152 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3012__CLK
timestamp 1751532392
transform 1 0 11648 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3013__CLK
timestamp 1751532392
transform 1 0 10416 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3014__CLK
timestamp 1751532392
transform 1 0 10752 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3015__CLK
timestamp 1751532392
transform 1 0 17472 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3017__CLK
timestamp 1751532392
transform 1 0 43792 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3018__CLK
timestamp 1751532392
transform 1 0 39536 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3019__CLK
timestamp 1751532392
transform 1 0 32480 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3020__CLK
timestamp 1751532392
transform 1 0 38192 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3021__CLK
timestamp 1751532392
transform 1 0 36176 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3022__CLK
timestamp 1751532392
transform 1 0 29904 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3023__CLK
timestamp 1751532392
transform -1 0 19936 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3024__CLK
timestamp 1751532392
transform 1 0 4816 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3025__CLK
timestamp 1751532392
transform 1 0 3920 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3026__CLK
timestamp 1751532392
transform -1 0 30912 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3027__CLK
timestamp 1751532392
transform 1 0 25312 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3028__CLK
timestamp 1751532392
transform -1 0 2016 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3029__CLK
timestamp 1751532392
transform -1 0 3696 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3029__D
timestamp 1751532392
transform -1 0 2800 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3030__CLK
timestamp 1751532392
transform 1 0 31024 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3031__CLK
timestamp 1751532392
transform 1 0 42336 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3032__CLK
timestamp 1751532392
transform 1 0 44128 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3033__CLK
timestamp 1751532392
transform 1 0 45136 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3034__CLK
timestamp 1751532392
transform 1 0 42784 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3035__CLK
timestamp 1751532392
transform 1 0 34832 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3036__CLK
timestamp 1751532392
transform 1 0 33376 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3037__CLK
timestamp 1751532392
transform 1 0 29680 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3038__CLK
timestamp 1751532392
transform 1 0 25088 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3039__CLK
timestamp 1751532392
transform 1 0 18144 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3040__CLK
timestamp 1751532392
transform 1 0 26656 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3041__CLK
timestamp 1751532392
transform 1 0 27216 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3042__CLK
timestamp 1751532392
transform 1 0 26208 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3042__D
timestamp 1751532392
transform -1 0 31808 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3043__CLK
timestamp 1751532392
transform 1 0 45248 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3044__CLK
timestamp 1751532392
transform 1 0 27664 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3046__CLK
timestamp 1751532392
transform 1 0 39536 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3049__CLK
timestamp 1751532392
transform 1 0 34048 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3050__CLK
timestamp 1751532392
transform 1 0 33936 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3052__CLK
timestamp 1751532392
transform 1 0 34048 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3053__CLK
timestamp 1751532392
transform 1 0 33264 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3054__CLK
timestamp 1751532392
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3055__CLK
timestamp 1751532392
transform -1 0 32480 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3056__CLK
timestamp 1751532392
transform 1 0 32704 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3057__CLK
timestamp 1751532392
transform 1 0 29568 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3058__CLK
timestamp 1751532392
transform 1 0 19600 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3059__CLK
timestamp 1751532392
transform 1 0 21168 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3060__CLK
timestamp 1751532392
transform 1 0 20048 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3061__CLK
timestamp 1751532392
transform 1 0 21392 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3062__CLK
timestamp 1751532392
transform 1 0 11648 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3063__CLK
timestamp 1751532392
transform 1 0 12096 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3064__CLK
timestamp 1751532392
transform -1 0 22512 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3065__CLK
timestamp 1751532392
transform 1 0 22512 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3066__CLK
timestamp 1751532392
transform 1 0 17472 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3067__CLK
timestamp 1751532392
transform 1 0 20608 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3069__CLK
timestamp 1751532392
transform 1 0 21840 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3071__CLK
timestamp 1751532392
transform 1 0 20720 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3079__CLK
timestamp 1751532392
transform 1 0 17472 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3083__CLK
timestamp 1751532392
transform -1 0 46704 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3084__CLK
timestamp 1751532392
transform 1 0 48048 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3085__CLK
timestamp 1751532392
transform 1 0 42000 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3086__CLK
timestamp 1751532392
transform 1 0 48048 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3087__CLK
timestamp 1751532392
transform 1 0 15008 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3088__CLK
timestamp 1751532392
transform 1 0 22064 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3089__CLK
timestamp 1751532392
transform -1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3109__A
timestamp 1751532392
transform -1 0 17808 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__3110__A
timestamp 1751532392
transform -1 0 30352 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_0_wb_clk_i_A
timestamp 1751532392
transform 1 0 24752 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_4_0_0_wb_clk_i_A
timestamp 1751532392
transform -1 0 8064 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_4_1_0_wb_clk_i_A
timestamp 1751532392
transform -1 0 12768 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_4_2_0_wb_clk_i_A
timestamp 1751532392
transform 1 0 19376 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_4_3_0_wb_clk_i_A
timestamp 1751532392
transform 1 0 19264 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_4_4_0_wb_clk_i_A
timestamp 1751532392
transform 1 0 15792 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_4_5_0_wb_clk_i_A
timestamp 1751532392
transform 1 0 13664 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_4_6_0_wb_clk_i_A
timestamp 1751532392
transform 1 0 22288 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_4_7_0_wb_clk_i_A
timestamp 1751532392
transform -1 0 20720 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_4_8_0_wb_clk_i_A
timestamp 1751532392
transform 1 0 28784 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_4_9_0_wb_clk_i_A
timestamp 1751532392
transform 1 0 30464 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_4_10_0_wb_clk_i_A
timestamp 1751532392
transform 1 0 39984 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_4_11_0_wb_clk_i_A
timestamp 1751532392
transform 1 0 36400 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_4_12_0_wb_clk_i_A
timestamp 1751532392
transform 1 0 35728 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_4_13_0_wb_clk_i_A
timestamp 1751532392
transform 1 0 38416 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_4_14_0_wb_clk_i_A
timestamp 1751532392
transform 1 0 42112 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_4_15_0_wb_clk_i_A
timestamp 1751532392
transform 1 0 37856 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkload1_A
timestamp 1751532392
transform 1 0 18704 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkload2_A
timestamp 1751532392
transform 1 0 15904 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkload3_A
timestamp 1751532392
transform 1 0 13552 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkload4_A
timestamp 1751532392
transform 1 0 14336 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkload5_A
timestamp 1751532392
transform 1 0 17584 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkload7_A
timestamp 1751532392
transform 1 0 35952 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkload9_A
timestamp 1751532392
transform 1 0 39200 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkload11_A
timestamp 1751532392
transform -1 0 37296 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkload12_A
timestamp 1751532392
transform 1 0 40208 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkload13_A
timestamp 1751532392
transform 1 0 45696 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkload14_A
timestamp 1751532392
transform 1 0 44240 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input1_A
timestamp 1751532392
transform -1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input2_A
timestamp 1751532392
transform -1 0 29904 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input3_A
timestamp 1751532392
transform -1 0 27104 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input4_A
timestamp 1751532392
transform -1 0 45920 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input5_A
timestamp 1751532392
transform -1 0 48272 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input6_A
timestamp 1751532392
transform -1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input7_A
timestamp 1751532392
transform -1 0 48384 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input8_A
timestamp 1751532392
transform -1 0 32256 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input9_A
timestamp 1751532392
transform -1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input10_A
timestamp 1751532392
transform 1 0 2128 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input11_A
timestamp 1751532392
transform 1 0 2464 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_output23_A
timestamp 1751532392
transform -1 0 3696 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_output25_A
timestamp 1751532392
transform -1 0 29008 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_0_wb_clk_i dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751661108
transform 1 0 24976 0 1 25088
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_4_0_0_wb_clk_i
timestamp 1751661108
transform -1 0 13664 0 -1 18816
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_4_1_0_wb_clk_i
timestamp 1751661108
transform -1 0 13328 0 -1 15680
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_4_2_0_wb_clk_i
timestamp 1751661108
transform -1 0 20272 0 1 15680
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_4_3_0_wb_clk_i
timestamp 1751661108
transform 1 0 17248 0 -1 18816
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_4_4_0_wb_clk_i
timestamp 1751661108
transform 1 0 11200 0 -1 31360
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_4_5_0_wb_clk_i
timestamp 1751661108
transform 1 0 11312 0 -1 32928
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_4_6_0_wb_clk_i
timestamp 1751661108
transform 1 0 18144 0 1 31360
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_4_7_0_wb_clk_i
timestamp 1751661108
transform -1 0 20496 0 -1 34496
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_4_8_0_wb_clk_i
timestamp 1751661108
transform 1 0 30800 0 1 14112
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_4_9_0_wb_clk_i
timestamp 1751661108
transform 1 0 30688 0 1 15680
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_4_10_0_wb_clk_i
timestamp 1751661108
transform 1 0 40768 0 -1 17248
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_4_11_0_wb_clk_i
timestamp 1751661108
transform 1 0 38752 0 1 18816
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_4_12_0_wb_clk_i
timestamp 1751661108
transform 1 0 35952 0 -1 32928
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_4_13_0_wb_clk_i
timestamp 1751661108
transform 1 0 37408 0 1 31360
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_4_14_0_wb_clk_i
timestamp 1751661108
transform 1 0 39872 0 1 29792
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_4_15_0_wb_clk_i
timestamp 1751661108
transform 1 0 40208 0 1 26656
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__inv_6  clkload0 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751896485
transform 1 0 9744 0 -1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_6  clkload1
timestamp 1751896485
transform 1 0 17472 0 -1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_6  clkload2
timestamp 1751896485
transform 1 0 15904 0 -1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_6  clkload3
timestamp 1751896485
transform 1 0 14448 0 1 31360
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_6  clkload4
timestamp 1751896485
transform 1 0 11312 0 -1 34496
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_6  clkload5
timestamp 1751896485
transform 1 0 18592 0 -1 31360
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_6  clkload6
timestamp 1751896485
transform -1 0 17024 0 -1 34496
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkload7
timestamp 1751661108
transform 1 0 29904 0 -1 15680
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__inv_6  clkload8
timestamp 1751896485
transform 1 0 30688 0 1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_4  clkload9
timestamp 1751558652
transform -1 0 38192 0 1 17248
box -86 -86 1094 870
use gf180mcu_as_sc_mcu7t3v3__inv_6  clkload10
timestamp 1751896485
transform 1 0 38752 0 -1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_6  clkload11
timestamp 1751896485
transform 1 0 33936 0 1 31360
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_6  clkload12
timestamp 1751896485
transform 1 0 37408 0 -1 34496
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_6  clkload13
timestamp 1751896485
transform 1 0 40768 0 -1 29792
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_4  clkload14 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751633659
transform 1 0 39760 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532351
transform 1 0 1568 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_18
timestamp 1751532351
transform 1 0 3360 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_36
timestamp 1751532351
transform 1 0 5376 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_52
timestamp 1751532351
transform 1 0 7168 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_70
timestamp 1751532351
transform 1 0 9184 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_0_86 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532312
transform 1 0 10976 0 1 3136
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_0_94 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532246
transform 1 0 11872 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_98 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532440
transform 1 0 12320 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_104
timestamp 1751532440
transform 1 0 12992 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_126
timestamp 1751532440
transform 1 0 15456 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_128 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532423
transform 1 0 15680 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_138
timestamp 1751532440
transform 1 0 16800 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_140
timestamp 1751532423
transform 1 0 17024 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_0_156
timestamp 1751532246
transform 1 0 18816 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_160
timestamp 1751532423
transform 1 0 19264 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_192
timestamp 1751532440
transform 1 0 22848 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_194
timestamp 1751532423
transform 1 0 23072 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_0_197
timestamp 1751532246
transform 1 0 23408 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_201
timestamp 1751532423
transform 1 0 23856 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_206
timestamp 1751532440
transform 1 0 24416 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_208
timestamp 1751532423
transform 1 0 24640 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_225
timestamp 1751532440
transform 1 0 26544 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_227
timestamp 1751532423
transform 1 0 26768 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_244
timestamp 1751532423
transform 1 0 28672 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_274
timestamp 1751532440
transform 1 0 32032 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_278
timestamp 1751532440
transform 1 0 32480 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_282
timestamp 1751532440
transform 1 0 32928 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_0_300
timestamp 1751532246
transform 1 0 34944 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_0_308
timestamp 1751532246
transform 1 0 35840 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_335
timestamp 1751532440
transform 1 0 38864 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_339
timestamp 1751532423
transform 1 0 39312 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_342
timestamp 1751532440
transform 1 0 39648 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_370
timestamp 1751532440
transform 1 0 42784 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_390
timestamp 1751532440
transform 1 0 45024 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_394
timestamp 1751532440
transform 1 0 45472 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_398
timestamp 1751532440
transform 1 0 45920 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_402
timestamp 1751532440
transform 1 0 46368 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_406
timestamp 1751532440
transform 1 0 46816 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_410
timestamp 1751532440
transform 1 0 47264 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_414
timestamp 1751532440
transform 1 0 47712 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_418
timestamp 1751532440
transform 1 0 48160 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_2
timestamp 1751532351
transform 1 0 1568 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_18
timestamp 1751532351
transform 1 0 3360 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_34
timestamp 1751532351
transform 1 0 5152 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_50
timestamp 1751532351
transform 1 0 6944 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_1_66
timestamp 1751532246
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_72
timestamp 1751532351
transform 1 0 9408 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_1_88
timestamp 1751532246
transform 1 0 11200 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_121
timestamp 1751532440
transform 1 0 14896 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_137
timestamp 1751532440
transform 1 0 16688 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_139
timestamp 1751532423
transform 1 0 16912 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_146
timestamp 1751532423
transform 1 0 17696 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_154
timestamp 1751532440
transform 1 0 18592 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_226
timestamp 1751532423
transform 1 0 26656 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_254
timestamp 1751532440
transform 1 0 29792 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_1_258
timestamp 1751532246
transform 1 0 30240 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_278
timestamp 1751532440
transform 1 0 32480 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_282
timestamp 1751532440
transform 1 0 32928 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_286
timestamp 1751532440
transform 1 0 33376 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_349
timestamp 1751532423
transform 1 0 40432 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_352
timestamp 1751532440
transform 1 0 40768 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_354
timestamp 1751532423
transform 1 0 40992 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_409
timestamp 1751532440
transform 1 0 47152 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_413
timestamp 1751532440
transform 1 0 47600 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_417
timestamp 1751532440
transform 1 0 48048 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_419
timestamp 1751532423
transform 1 0 48272 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_2_2
timestamp 1751532351
transform 1 0 1568 0 1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_2_18
timestamp 1751532351
transform 1 0 3360 0 1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_34
timestamp 1751532423
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_2_37
timestamp 1751532351
transform 1 0 5488 0 1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_2_53
timestamp 1751532351
transform 1 0 7280 0 1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_2_69
timestamp 1751532351
transform 1 0 9072 0 1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_2_85
timestamp 1751532312
transform 1 0 10864 0 1 4704
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_2_93
timestamp 1751532246
transform 1 0 11760 0 1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_97
timestamp 1751532423
transform 1 0 12208 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_121
timestamp 1751532440
transform 1 0 14896 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_123
timestamp 1751532423
transform 1 0 15120 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_171
timestamp 1751532440
transform 1 0 20496 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_188
timestamp 1751532440
transform 1 0 22400 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_224
timestamp 1751532440
transform 1 0 26432 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_226
timestamp 1751532423
transform 1 0 26656 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_243
timestamp 1751532440
transform 1 0 28560 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_247
timestamp 1751532440
transform 1 0 29008 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_282
timestamp 1751532440
transform 1 0 32928 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_284
timestamp 1751532423
transform 1 0 33152 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_311
timestamp 1751532440
transform 1 0 36176 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_327
timestamp 1751532440
transform 1 0 37968 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_329
timestamp 1751532423
transform 1 0 38192 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_2
timestamp 1751532351
transform 1 0 1568 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_3_18
timestamp 1751532312
transform 1 0 3360 0 -1 6272
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_26
timestamp 1751532246
transform 1 0 4256 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_30
timestamp 1751532423
transform 1 0 4704 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_58
timestamp 1751532440
transform 1 0 7840 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_62
timestamp 1751532423
transform 1 0 8288 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_78
timestamp 1751532440
transform 1 0 10080 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_3_82
timestamp 1751532312
transform 1 0 10528 0 -1 6272
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_90
timestamp 1751532246
transform 1 0 11424 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_94
timestamp 1751532423
transform 1 0 11872 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_111
timestamp 1751532440
transform 1 0 13776 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_113
timestamp 1751532423
transform 1 0 14000 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_142
timestamp 1751532440
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_182
timestamp 1751532423
transform 1 0 21728 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_222
timestamp 1751532440
transform 1 0 26208 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_251
timestamp 1751532440
transform 1 0 29456 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_253
timestamp 1751532423
transform 1 0 29680 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_274
timestamp 1751532423
transform 1 0 32032 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_279
timestamp 1751532423
transform 1 0 32592 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_312
timestamp 1751532423
transform 1 0 36288 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_333
timestamp 1751532440
transform 1 0 38640 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_349
timestamp 1751532423
transform 1 0 40432 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_365
timestamp 1751532440
transform 1 0 42224 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_369
timestamp 1751532423
transform 1 0 42672 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_383
timestamp 1751532440
transform 1 0 44240 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_385
timestamp 1751532423
transform 1 0 44464 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_400
timestamp 1751532440
transform 1 0 46144 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_416
timestamp 1751532440
transform 1 0 47936 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_2
timestamp 1751532351
transform 1 0 1568 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_4_18
timestamp 1751532246
transform 1 0 3360 0 1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_22
timestamp 1751532423
transform 1 0 3808 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_37
timestamp 1751532440
transform 1 0 5488 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_48
timestamp 1751532440
transform 1 0 6720 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_50
timestamp 1751532423
transform 1 0 6944 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_164
timestamp 1751532440
transform 1 0 19712 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_168
timestamp 1751532440
transform 1 0 20160 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_172
timestamp 1751532440
transform 1 0 20608 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_174
timestamp 1751532423
transform 1 0 20832 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_177
timestamp 1751532440
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_189
timestamp 1751532440
transform 1 0 22512 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_207
timestamp 1751532423
transform 1 0 24528 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_225
timestamp 1751532440
transform 1 0 26544 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_229
timestamp 1751532423
transform 1 0 26992 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_244
timestamp 1751532423
transform 1 0 28672 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_251
timestamp 1751532440
transform 1 0 29456 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_255
timestamp 1751532440
transform 1 0 29904 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_257
timestamp 1751532423
transform 1 0 30128 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_312
timestamp 1751532440
transform 1 0 36288 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_314
timestamp 1751532423
transform 1 0 36512 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_317
timestamp 1751532440
transform 1 0 36848 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_319
timestamp 1751532423
transform 1 0 37072 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_353
timestamp 1751532440
transform 1 0 40880 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_357
timestamp 1751532423
transform 1 0 41328 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_375
timestamp 1751532440
transform 1 0 43344 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_384
timestamp 1751532423
transform 1 0 44352 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_387
timestamp 1751532423
transform 1 0 44688 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_392
timestamp 1751532423
transform 1 0 45248 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_414
timestamp 1751532440
transform 1 0 47712 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_416
timestamp 1751532423
transform 1 0 47936 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_419
timestamp 1751532423
transform 1 0 48272 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_5_2
timestamp 1751532312
transform 1 0 1568 0 -1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_10
timestamp 1751532246
transform 1 0 2464 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_14
timestamp 1751532440
transform 1 0 2912 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_16
timestamp 1751532423
transform 1 0 3136 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_44
timestamp 1751532440
transform 1 0 6272 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_64
timestamp 1751532246
transform 1 0 8512 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_68
timestamp 1751532440
transform 1 0 8960 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_90
timestamp 1751532246
transform 1 0 11424 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_94
timestamp 1751532423
transform 1 0 11872 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_135
timestamp 1751532423
transform 1 0 16464 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_142
timestamp 1751532440
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_156
timestamp 1751532423
transform 1 0 18816 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_5_188
timestamp 1751532312
transform 1 0 22400 0 -1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_196
timestamp 1751532440
transform 1 0 23296 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_204
timestamp 1751532246
transform 1 0 24192 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_222
timestamp 1751532246
transform 1 0 26208 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_255
timestamp 1751532440
transform 1 0 29904 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_279
timestamp 1751532423
transform 1 0 32592 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_282
timestamp 1751532440
transform 1 0 32928 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_301
timestamp 1751532440
transform 1 0 35056 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_303
timestamp 1751532423
transform 1 0 35280 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_331
timestamp 1751532440
transform 1 0 38416 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_335
timestamp 1751532423
transform 1 0 38864 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_352
timestamp 1751532423
transform 1 0 40768 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_363
timestamp 1751532423
transform 1 0 42000 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_378
timestamp 1751532423
transform 1 0 43680 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_6_2
timestamp 1751532312
transform 1 0 1568 0 1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_16
timestamp 1751532440
transform 1 0 3136 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_18
timestamp 1751532423
transform 1 0 3360 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_6_55
timestamp 1751532246
transform 1 0 7504 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_59
timestamp 1751532423
transform 1 0 7952 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_94
timestamp 1751532440
transform 1 0 11872 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_114
timestamp 1751532440
transform 1 0 14112 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_123
timestamp 1751532440
transform 1 0 15120 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_125
timestamp 1751532423
transform 1 0 15344 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_128
timestamp 1751532440
transform 1 0 15680 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_157
timestamp 1751532440
transform 1 0 18928 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_161
timestamp 1751532440
transform 1 0 19376 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_165
timestamp 1751532440
transform 1 0 19824 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_173
timestamp 1751532440
transform 1 0 20720 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_234
timestamp 1751532440
transform 1 0 27552 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_236
timestamp 1751532423
transform 1 0 27776 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_247
timestamp 1751532423
transform 1 0 29008 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_254
timestamp 1751532440
transform 1 0 29792 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_258
timestamp 1751532440
transform 1 0 30240 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_289
timestamp 1751532440
transform 1 0 33712 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_300
timestamp 1751532440
transform 1 0 34944 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_317
timestamp 1751532440
transform 1 0 36848 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_331
timestamp 1751532440
transform 1 0 38416 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_333
timestamp 1751532423
transform 1 0 38640 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_351
timestamp 1751532440
transform 1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_353
timestamp 1751532423
transform 1 0 40880 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_364
timestamp 1751532440
transform 1 0 42112 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_368
timestamp 1751532440
transform 1 0 42560 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_370
timestamp 1751532423
transform 1 0 42784 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_29
timestamp 1751532440
transform 1 0 4592 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_51
timestamp 1751532423
transform 1 0 7056 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_78
timestamp 1751532440
transform 1 0 10080 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_80
timestamp 1751532423
transform 1 0 10304 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_117
timestamp 1751532440
transform 1 0 14448 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_131
timestamp 1751532440
transform 1 0 16016 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_135
timestamp 1751532440
transform 1 0 16464 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_139
timestamp 1751532423
transform 1 0 16912 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_142
timestamp 1751532440
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_144
timestamp 1751532423
transform 1 0 17472 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_147
timestamp 1751532440
transform 1 0 17808 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_151
timestamp 1751532440
transform 1 0 18256 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_157
timestamp 1751532423
transform 1 0 18928 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_185
timestamp 1751532440
transform 1 0 22064 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_189
timestamp 1751532423
transform 1 0 22512 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_199
timestamp 1751532423
transform 1 0 23632 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_212
timestamp 1751532440
transform 1 0 25088 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_233
timestamp 1751532440
transform 1 0 27440 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_235
timestamp 1751532423
transform 1 0 27664 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_269
timestamp 1751532423
transform 1 0 31472 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_286
timestamp 1751532440
transform 1 0 33376 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_290
timestamp 1751532440
transform 1 0 33824 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_294
timestamp 1751532440
transform 1 0 34272 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_310
timestamp 1751532440
transform 1 0 36064 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_312
timestamp 1751532423
transform 1 0 36288 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_342
timestamp 1751532423
transform 1 0 39648 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_352
timestamp 1751532423
transform 1 0 40768 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_380
timestamp 1751532246
transform 1 0 43904 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_384
timestamp 1751532423
transform 1 0 44352 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_387
timestamp 1751532440
transform 1 0 44688 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_389
timestamp 1751532423
transform 1 0 44912 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_398
timestamp 1751532423
transform 1 0 45920 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_406
timestamp 1751532440
transform 1 0 46816 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_410
timestamp 1751532440
transform 1 0 47264 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_414
timestamp 1751532246
transform 1 0 47712 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_55
timestamp 1751532246
transform 1 0 7504 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_65
timestamp 1751532423
transform 1 0 8624 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_79
timestamp 1751532440
transform 1 0 10192 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_83
timestamp 1751532246
transform 1 0 10640 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_87
timestamp 1751532440
transform 1 0 11088 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_124
timestamp 1751532440
transform 1 0 15232 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_126
timestamp 1751532423
transform 1 0 15456 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_164
timestamp 1751532423
transform 1 0 19712 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_177
timestamp 1751532440
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_181
timestamp 1751532440
transform 1 0 21616 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_183
timestamp 1751532423
transform 1 0 21840 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_210
timestamp 1751532246
transform 1 0 24864 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_214
timestamp 1751532423
transform 1 0 25312 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_221
timestamp 1751532440
transform 1 0 26096 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_223
timestamp 1751532423
transform 1 0 26320 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_226
timestamp 1751532440
transform 1 0 26656 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_240
timestamp 1751532440
transform 1 0 28224 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_242
timestamp 1751532423
transform 1 0 28448 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_257
timestamp 1751532440
transform 1 0 30128 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_259
timestamp 1751532423
transform 1 0 30352 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_278
timestamp 1751532440
transform 1 0 32480 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_282
timestamp 1751532440
transform 1 0 32928 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_286
timestamp 1751532440
transform 1 0 33376 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_290
timestamp 1751532440
transform 1 0 33824 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_304
timestamp 1751532423
transform 1 0 35392 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_312
timestamp 1751532440
transform 1 0 36288 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_314
timestamp 1751532423
transform 1 0 36512 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_317
timestamp 1751532440
transform 1 0 36848 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_321
timestamp 1751532440
transform 1 0 37296 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_345
timestamp 1751532423
transform 1 0 39984 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_366
timestamp 1751532440
transform 1 0 42336 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_370
timestamp 1751532440
transform 1 0 42784 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_372
timestamp 1751532423
transform 1 0 43008 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_379
timestamp 1751532440
transform 1 0 43792 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_383
timestamp 1751532440
transform 1 0 44240 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_9_2
timestamp 1751532246
transform 1 0 1568 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_9_18
timestamp 1751532246
transform 1 0 3360 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_22
timestamp 1751532423
transform 1 0 3808 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_41
timestamp 1751532440
transform 1 0 5936 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_9_79
timestamp 1751532246
transform 1 0 10192 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_83
timestamp 1751532423
transform 1 0 10640 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_86
timestamp 1751532440
transform 1 0 10976 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_90
timestamp 1751532440
transform 1 0 11424 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_94
timestamp 1751532440
transform 1 0 11872 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_98
timestamp 1751532440
transform 1 0 12320 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_126
timestamp 1751532440
transform 1 0 15456 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_142
timestamp 1751532440
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_153
timestamp 1751532440
transform 1 0 18480 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_155
timestamp 1751532423
transform 1 0 18704 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_160
timestamp 1751532440
transform 1 0 19264 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_162
timestamp 1751532423
transform 1 0 19488 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_190
timestamp 1751532440
transform 1 0 22624 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_9_198
timestamp 1751532246
transform 1 0 23520 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_202
timestamp 1751532440
transform 1 0 23968 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_218
timestamp 1751532440
transform 1 0 25760 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_232
timestamp 1751532440
transform 1 0 27328 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_236
timestamp 1751532440
transform 1 0 27776 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_279
timestamp 1751532423
transform 1 0 32592 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_339
timestamp 1751532440
transform 1 0 39312 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_2
timestamp 1751532440
transform 1 0 1568 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_31
timestamp 1751532440
transform 1 0 4816 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_51
timestamp 1751532246
transform 1 0 7056 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_72
timestamp 1751532440
transform 1 0 9408 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_76
timestamp 1751532440
transform 1 0 9856 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_107
timestamp 1751532440
transform 1 0 13328 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_109
timestamp 1751532423
transform 1 0 13552 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_126
timestamp 1751532440
transform 1 0 15456 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_128
timestamp 1751532423
transform 1 0 15680 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_170
timestamp 1751532423
transform 1 0 20384 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_187
timestamp 1751532423
transform 1 0 22288 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_192
timestamp 1751532440
transform 1 0 22848 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_196
timestamp 1751532246
transform 1 0 23296 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_200
timestamp 1751532440
transform 1 0 23744 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_214
timestamp 1751532440
transform 1 0 25312 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_218
timestamp 1751532423
transform 1 0 25760 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_232
timestamp 1751532440
transform 1 0 27328 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_236
timestamp 1751532246
transform 1 0 27776 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_240
timestamp 1751532440
transform 1 0 28224 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_242
timestamp 1751532423
transform 1 0 28448 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_247
timestamp 1751532246
transform 1 0 29008 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_251
timestamp 1751532423
transform 1 0 29456 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_254
timestamp 1751532440
transform 1 0 29792 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_289
timestamp 1751532440
transform 1 0 33712 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_313
timestamp 1751532440
transform 1 0 36400 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_341
timestamp 1751532246
transform 1 0 39536 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_357
timestamp 1751532440
transform 1 0 41328 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_383
timestamp 1751532440
transform 1 0 44240 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_387
timestamp 1751532440
transform 1 0 44688 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_391
timestamp 1751532423
transform 1 0 45136 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_412
timestamp 1751532440
transform 1 0 47488 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_11_2
timestamp 1751532351
transform 1 0 1568 0 -1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_11_18
timestamp 1751532246
transform 1 0 3360 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_22
timestamp 1751532423
transform 1 0 3808 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_50
timestamp 1751532440
transform 1 0 6944 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_54
timestamp 1751532423
transform 1 0 7392 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_61
timestamp 1751532440
transform 1 0 8176 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_82
timestamp 1751532440
transform 1 0 10528 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_121
timestamp 1751532440
transform 1 0 14896 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_123
timestamp 1751532423
transform 1 0 15120 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_11_133
timestamp 1751532246
transform 1 0 16240 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_137
timestamp 1751532423
transform 1 0 16688 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_11_149
timestamp 1751532246
transform 1 0 18032 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_171
timestamp 1751532440
transform 1 0 20496 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_175
timestamp 1751532440
transform 1 0 20944 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_179
timestamp 1751532423
transform 1 0 21392 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_11_206
timestamp 1751532246
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_11_212
timestamp 1751532246
transform 1 0 25088 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_216
timestamp 1751532423
transform 1 0 25536 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_229
timestamp 1751532440
transform 1 0 26992 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_233
timestamp 1751532440
transform 1 0 27440 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_272
timestamp 1751532440
transform 1 0 31808 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_274
timestamp 1751532423
transform 1 0 32032 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_279
timestamp 1751532423
transform 1 0 32592 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_11_282
timestamp 1751532246
transform 1 0 32928 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_311
timestamp 1751532440
transform 1 0 36176 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_315
timestamp 1751532440
transform 1 0 36624 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_337
timestamp 1751532440
transform 1 0 39088 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_341
timestamp 1751532440
transform 1 0 39536 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_366
timestamp 1751532423
transform 1 0 42336 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_377
timestamp 1751532440
transform 1 0 43568 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_381
timestamp 1751532440
transform 1 0 44016 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_12_2
timestamp 1751532351
transform 1 0 1568 0 1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_12_18
timestamp 1751532312
transform 1 0 3360 0 1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_26
timestamp 1751532440
transform 1 0 4256 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_28
timestamp 1751532423
transform 1 0 4480 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_62
timestamp 1751532423
transform 1 0 8288 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_69
timestamp 1751532423
transform 1 0 9072 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_97
timestamp 1751532440
transform 1 0 12208 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_101
timestamp 1751532440
transform 1 0 12656 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_107
timestamp 1751532423
transform 1 0 13328 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_153
timestamp 1751532440
transform 1 0 18480 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_157
timestamp 1751532246
transform 1 0 18928 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_203
timestamp 1751532440
transform 1 0 24080 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_12_215
timestamp 1751532312
transform 1 0 25424 0 1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_223
timestamp 1751532246
transform 1 0 26320 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_227
timestamp 1751532423
transform 1 0 26768 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_232
timestamp 1751532440
transform 1 0 27328 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_12_236
timestamp 1751532312
transform 1 0 27776 0 1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_244
timestamp 1751532423
transform 1 0 28672 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_257
timestamp 1751532440
transform 1 0 30128 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_259
timestamp 1751532423
transform 1 0 30352 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_290
timestamp 1751532440
transform 1 0 33824 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_294
timestamp 1751532440
transform 1 0 34272 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_303
timestamp 1751532246
transform 1 0 35280 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_317
timestamp 1751532440
transform 1 0 36848 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_370
timestamp 1751532423
transform 1 0 42784 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_13_2
timestamp 1751532312
transform 1 0 1568 0 -1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_10
timestamp 1751532246
transform 1 0 2464 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_13_20
timestamp 1751532312
transform 1 0 3584 0 -1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_28
timestamp 1751532440
transform 1 0 4480 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_30
timestamp 1751532423
transform 1 0 4704 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_50
timestamp 1751532440
transform 1 0 6944 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_88
timestamp 1751532440
transform 1 0 11200 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_90
timestamp 1751532423
transform 1 0 11424 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_118
timestamp 1751532440
transform 1 0 14560 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_142
timestamp 1751532440
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_144
timestamp 1751532423
transform 1 0 17472 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_159
timestamp 1751532423
transform 1 0 19152 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_167
timestamp 1751532440
transform 1 0 20048 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_169
timestamp 1751532423
transform 1 0 20272 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_190
timestamp 1751532440
transform 1 0 22624 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_194
timestamp 1751532246
transform 1 0 23072 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_198
timestamp 1751532423
transform 1 0 23520 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_205
timestamp 1751532246
transform 1 0 24304 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_209
timestamp 1751532423
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_13_235
timestamp 1751532312
transform 1 0 27664 0 -1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_243
timestamp 1751532440
transform 1 0 28560 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_247
timestamp 1751532440
transform 1 0 29008 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_277
timestamp 1751532440
transform 1 0 32368 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_279
timestamp 1751532423
transform 1 0 32592 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_336
timestamp 1751532440
transform 1 0 38976 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_340
timestamp 1751532246
transform 1 0 39424 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_346
timestamp 1751532440
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_352
timestamp 1751532246
transform 1 0 40768 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_356
timestamp 1751532423
transform 1 0 41216 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_382
timestamp 1751532440
transform 1 0 44128 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_415
timestamp 1751532440
transform 1 0 47824 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_419
timestamp 1751532423
transform 1 0 48272 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_2
timestamp 1751532246
transform 1 0 1568 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_33
timestamp 1751532440
transform 1 0 5040 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_37
timestamp 1751532423
transform 1 0 5488 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_52
timestamp 1751532440
transform 1 0 7168 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_54
timestamp 1751532423
transform 1 0 7392 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_107
timestamp 1751532440
transform 1 0 13328 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_109
timestamp 1751532423
transform 1 0 13552 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_158
timestamp 1751532440
transform 1 0 19040 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_174
timestamp 1751532423
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_183
timestamp 1751532440
transform 1 0 21840 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_211
timestamp 1751532246
transform 1 0 24976 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_215
timestamp 1751532440
transform 1 0 25424 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_321
timestamp 1751532440
transform 1 0 37296 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_323
timestamp 1751532423
transform 1 0 37520 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_350
timestamp 1751532440
transform 1 0 40544 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_356
timestamp 1751532440
transform 1 0 41216 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_358
timestamp 1751532423
transform 1 0 41440 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_376
timestamp 1751532440
transform 1 0 43456 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_401
timestamp 1751532440
transform 1 0 46256 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_412
timestamp 1751532440
transform 1 0 47488 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_416
timestamp 1751532440
transform 1 0 47936 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_15_2
timestamp 1751532312
transform 1 0 1568 0 -1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_10
timestamp 1751532246
transform 1 0 2464 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_14
timestamp 1751532440
transform 1 0 2912 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_16
timestamp 1751532423
transform 1 0 3136 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_23
timestamp 1751532423
transform 1 0 3920 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_49
timestamp 1751532423
transform 1 0 6832 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_123
timestamp 1751532246
transform 1 0 15120 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_127
timestamp 1751532423
transform 1 0 15568 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_130
timestamp 1751532440
transform 1 0 15904 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_142
timestamp 1751532440
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_154
timestamp 1751532423
transform 1 0 18592 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_192
timestamp 1751532440
transform 1 0 22848 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_194
timestamp 1751532423
transform 1 0 23072 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_207
timestamp 1751532440
transform 1 0 24528 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_209
timestamp 1751532423
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_212
timestamp 1751532246
transform 1 0 25088 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_216
timestamp 1751532423
transform 1 0 25536 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_219
timestamp 1751532440
transform 1 0 25872 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_223
timestamp 1751532440
transform 1 0 26320 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_227
timestamp 1751532440
transform 1 0 26768 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_229
timestamp 1751532423
transform 1 0 26992 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_240
timestamp 1751532440
transform 1 0 28224 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_244
timestamp 1751532423
transform 1 0 28672 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_319
timestamp 1751532440
transform 1 0 37072 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_352
timestamp 1751532423
transform 1 0 40768 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_390
timestamp 1751532440
transform 1 0 45024 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_392
timestamp 1751532423
transform 1 0 45248 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_2
timestamp 1751532246
transform 1 0 1568 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_6
timestamp 1751532440
transform 1 0 2016 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_37
timestamp 1751532440
transform 1 0 5488 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_39
timestamp 1751532423
transform 1 0 5712 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_58
timestamp 1751532440
transform 1 0 7840 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_60
timestamp 1751532423
transform 1 0 8064 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_68
timestamp 1751532440
transform 1 0 8960 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_70
timestamp 1751532423
transform 1 0 9184 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_117
timestamp 1751532246
transform 1 0 14448 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_173
timestamp 1751532440
transform 1 0 20720 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_181
timestamp 1751532440
transform 1 0 21616 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_183
timestamp 1751532423
transform 1 0 21840 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_202
timestamp 1751532440
transform 1 0 23968 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_204
timestamp 1751532423
transform 1 0 24192 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_217
timestamp 1751532440
transform 1 0 25648 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_219
timestamp 1751532423
transform 1 0 25872 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_240
timestamp 1751532423
transform 1 0 28224 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_247
timestamp 1751532440
transform 1 0 29008 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_249
timestamp 1751532423
transform 1 0 29232 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_260
timestamp 1751532440
transform 1 0 30464 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_307
timestamp 1751532440
transform 1 0 35728 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_311
timestamp 1751532440
transform 1 0 36176 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_321
timestamp 1751532440
transform 1 0 37296 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_323
timestamp 1751532423
transform 1 0 37520 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_351
timestamp 1751532440
transform 1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_353
timestamp 1751532423
transform 1 0 40880 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_387
timestamp 1751532423
transform 1 0 44688 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_406
timestamp 1751532440
transform 1 0 46816 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_415
timestamp 1751532440
transform 1 0 47824 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_419
timestamp 1751532423
transform 1 0 48272 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_17_2
timestamp 1751532351
transform 1 0 1568 0 -1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_17_18
timestamp 1751532246
transform 1 0 3360 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_24
timestamp 1751532440
transform 1 0 4032 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_61
timestamp 1751532423
transform 1 0 8176 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_69
timestamp 1751532423
transform 1 0 9072 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_106
timestamp 1751532423
transform 1 0 13216 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_142
timestamp 1751532440
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_161
timestamp 1751532440
transform 1 0 19376 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_17_192
timestamp 1751532246
transform 1 0 22848 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_208
timestamp 1751532440
transform 1 0 24640 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_222
timestamp 1751532423
transform 1 0 26208 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_235
timestamp 1751532440
transform 1 0 27664 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_237
timestamp 1751532423
transform 1 0 27888 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_248
timestamp 1751532440
transform 1 0 29120 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_252
timestamp 1751532423
transform 1 0 29568 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_344
timestamp 1751532440
transform 1 0 39872 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_348
timestamp 1751532440
transform 1 0 40320 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_419
timestamp 1751532423
transform 1 0 48272 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_18_2
timestamp 1751532351
transform 1 0 1568 0 1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_18
timestamp 1751532246
transform 1 0 3360 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_22
timestamp 1751532440
transform 1 0 3808 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_24
timestamp 1751532423
transform 1 0 4032 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_27
timestamp 1751532440
transform 1 0 4368 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_31
timestamp 1751532440
transform 1 0 4816 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_44
timestamp 1751532423
transform 1 0 6272 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_107
timestamp 1751532440
transform 1 0 13328 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_119
timestamp 1751532440
transform 1 0 14672 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_121
timestamp 1751532423
transform 1 0 14896 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_161
timestamp 1751532440
transform 1 0 19376 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_163
timestamp 1751532423
transform 1 0 19600 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_202
timestamp 1751532440
transform 1 0 23968 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_204
timestamp 1751532423
transform 1 0 24192 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_220
timestamp 1751532440
transform 1 0 25984 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_222
timestamp 1751532423
transform 1 0 26208 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_233
timestamp 1751532440
transform 1 0 27440 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_244
timestamp 1751532423
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_257
timestamp 1751532440
transform 1 0 30128 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_259
timestamp 1751532423
transform 1 0 30352 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_272
timestamp 1751532440
transform 1 0 31808 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_274
timestamp 1751532423
transform 1 0 32032 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_312
timestamp 1751532440
transform 1 0 36288 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_314
timestamp 1751532423
transform 1 0 36512 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_317
timestamp 1751532440
transform 1 0 36848 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_319
timestamp 1751532423
transform 1 0 37072 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_383
timestamp 1751532440
transform 1 0 44240 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_19_2
timestamp 1751532312
transform 1 0 1568 0 -1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_19_10
timestamp 1751532246
transform 1 0 2464 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_14
timestamp 1751532423
transform 1 0 2912 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_52
timestamp 1751532440
transform 1 0 7168 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_56
timestamp 1751532440
transform 1 0 7616 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_67
timestamp 1751532440
transform 1 0 8848 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_69
timestamp 1751532423
transform 1 0 9072 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_72
timestamp 1751532440
transform 1 0 9408 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_74
timestamp 1751532423
transform 1 0 9632 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_110
timestamp 1751532423
transform 1 0 13664 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_173
timestamp 1751532440
transform 1 0 20720 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_209
timestamp 1751532423
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_235
timestamp 1751532440
transform 1 0 27664 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_278
timestamp 1751532440
transform 1 0 32480 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_292
timestamp 1751532440
transform 1 0 34048 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_294
timestamp 1751532423
transform 1 0 34272 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_373
timestamp 1751532440
transform 1 0 43120 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_375
timestamp 1751532423
transform 1 0 43344 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_417
timestamp 1751532440
transform 1 0 48048 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_419
timestamp 1751532423
transform 1 0 48272 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_20_2
timestamp 1751532351
transform 1 0 1568 0 1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_18
timestamp 1751532246
transform 1 0 3360 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_22
timestamp 1751532423
transform 1 0 3808 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_37
timestamp 1751532440
transform 1 0 5488 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_39
timestamp 1751532423
transform 1 0 5712 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_59
timestamp 1751532246
transform 1 0 7952 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_63
timestamp 1751532423
transform 1 0 8400 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_107
timestamp 1751532423
transform 1 0 13328 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_134
timestamp 1751532440
transform 1 0 16352 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_136
timestamp 1751532423
transform 1 0 16576 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_166
timestamp 1751532440
transform 1 0 19936 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_174
timestamp 1751532423
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_181
timestamp 1751532246
transform 1 0 21616 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_185
timestamp 1751532423
transform 1 0 22064 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_188
timestamp 1751532440
transform 1 0 22400 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_192
timestamp 1751532440
transform 1 0 22848 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_216
timestamp 1751532423
transform 1 0 25536 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_234
timestamp 1751532440
transform 1 0 27552 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_238
timestamp 1751532440
transform 1 0 28000 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_242
timestamp 1751532440
transform 1 0 28448 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_244
timestamp 1751532423
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_274
timestamp 1751532423
transform 1 0 32032 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_286
timestamp 1751532440
transform 1 0 33376 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_330
timestamp 1751532440
transform 1 0 38304 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_373
timestamp 1751532440
transform 1 0 43120 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_375
timestamp 1751532423
transform 1 0 43344 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_383
timestamp 1751532440
transform 1 0 44240 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_401
timestamp 1751532440
transform 1 0 46256 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_403
timestamp 1751532423
transform 1 0 46480 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_418
timestamp 1751532440
transform 1 0 48160 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_35
timestamp 1751532440
transform 1 0 5264 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_37
timestamp 1751532423
transform 1 0 5488 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_66
timestamp 1751532440
transform 1 0 8736 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_72
timestamp 1751532440
transform 1 0 9408 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_105
timestamp 1751532423
transform 1 0 13104 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_133
timestamp 1751532423
transform 1 0 16240 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_148
timestamp 1751532440
transform 1 0 17920 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_150
timestamp 1751532423
transform 1 0 18144 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_157
timestamp 1751532423
transform 1 0 18928 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_208
timestamp 1751532440
transform 1 0 24640 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_216
timestamp 1751532423
transform 1 0 25536 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_239
timestamp 1751532440
transform 1 0 28112 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_243
timestamp 1751532440
transform 1 0 28560 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_21_247
timestamp 1751532312
transform 1 0 29008 0 -1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_255
timestamp 1751532440
transform 1 0 29904 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_264
timestamp 1751532440
transform 1 0 30912 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_279
timestamp 1751532423
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_292
timestamp 1751532440
transform 1 0 34048 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_331
timestamp 1751532440
transform 1 0 38416 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_333
timestamp 1751532423
transform 1 0 38640 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_352
timestamp 1751532423
transform 1 0 40768 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_37
timestamp 1751532423
transform 1 0 5488 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_85
timestamp 1751532423
transform 1 0 10864 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_102
timestamp 1751532440
transform 1 0 12768 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_104
timestamp 1751532423
transform 1 0 12992 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_113
timestamp 1751532423
transform 1 0 14000 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_124
timestamp 1751532440
transform 1 0 15232 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_128
timestamp 1751532440
transform 1 0 15680 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_177
timestamp 1751532423
transform 1 0 21168 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_215
timestamp 1751532440
transform 1 0 25424 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_217
timestamp 1751532423
transform 1 0 25648 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_22_253
timestamp 1751532246
transform 1 0 29680 0 1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_257
timestamp 1751532440
transform 1 0 30128 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_290
timestamp 1751532440
transform 1 0 33824 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_313
timestamp 1751532440
transform 1 0 36400 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_356
timestamp 1751532440
transform 1 0 41216 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_2
timestamp 1751532246
transform 1 0 1568 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_12
timestamp 1751532246
transform 1 0 2688 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_16
timestamp 1751532423
transform 1 0 3136 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_59
timestamp 1751532440
transform 1 0 7952 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_67
timestamp 1751532440
transform 1 0 8848 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_69
timestamp 1751532423
transform 1 0 9072 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_72
timestamp 1751532440
transform 1 0 9408 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_107
timestamp 1751532423
transform 1 0 13328 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_128
timestamp 1751532440
transform 1 0 15680 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_132
timestamp 1751532440
transform 1 0 16128 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_136
timestamp 1751532440
transform 1 0 16576 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_142
timestamp 1751532440
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_144
timestamp 1751532423
transform 1 0 17472 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_163
timestamp 1751532246
transform 1 0 19600 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_167
timestamp 1751532423
transform 1 0 20048 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_170
timestamp 1751532440
transform 1 0 20384 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_191
timestamp 1751532440
transform 1 0 22736 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_23_195
timestamp 1751532312
transform 1 0 23184 0 -1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_203
timestamp 1751532423
transform 1 0 24080 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_206
timestamp 1751532440
transform 1 0 24416 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_212
timestamp 1751532440
transform 1 0 25088 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_214
timestamp 1751532423
transform 1 0 25312 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_235
timestamp 1751532440
transform 1 0 27664 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_239
timestamp 1751532440
transform 1 0 28112 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_241
timestamp 1751532423
transform 1 0 28336 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_252
timestamp 1751532423
transform 1 0 29568 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_282
timestamp 1751532440
transform 1 0 32928 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_326
timestamp 1751532440
transform 1 0 37856 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_336
timestamp 1751532440
transform 1 0 38976 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_338
timestamp 1751532423
transform 1 0 39200 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_345
timestamp 1751532440
transform 1 0 39984 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_349
timestamp 1751532423
transform 1 0 40432 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_392
timestamp 1751532440
transform 1 0 45248 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_394
timestamp 1751532423
transform 1 0 45472 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_416
timestamp 1751532440
transform 1 0 47936 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_2
timestamp 1751532440
transform 1 0 1568 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_4
timestamp 1751532423
transform 1 0 1792 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_24_59
timestamp 1751532312
transform 1 0 7952 0 1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_67
timestamp 1751532423
transform 1 0 8848 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_24_75
timestamp 1751532246
transform 1 0 9744 0 1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_79
timestamp 1751532423
transform 1 0 10192 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_102
timestamp 1751532440
transform 1 0 12768 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_104
timestamp 1751532423
transform 1 0 12992 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_137
timestamp 1751532440
transform 1 0 16688 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_141
timestamp 1751532440
transform 1 0 17136 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_143
timestamp 1751532423
transform 1 0 17360 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_24_161
timestamp 1751532246
transform 1 0 19376 0 1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_173
timestamp 1751532440
transform 1 0 20720 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_203
timestamp 1751532440
transform 1 0 24080 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_205
timestamp 1751532423
transform 1 0 24304 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_24_247
timestamp 1751532246
transform 1 0 29008 0 1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_251
timestamp 1751532423
transform 1 0 29456 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_309
timestamp 1751532440
transform 1 0 35952 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_313
timestamp 1751532440
transform 1 0 36400 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_324
timestamp 1751532440
transform 1 0 37632 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_328
timestamp 1751532440
transform 1 0 38080 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_330
timestamp 1751532423
transform 1 0 38304 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_364
timestamp 1751532423
transform 1 0 42112 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_383
timestamp 1751532440
transform 1 0 44240 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_387
timestamp 1751532440
transform 1 0 44688 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_389
timestamp 1751532423
transform 1 0 44912 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_417
timestamp 1751532440
transform 1 0 48048 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_419
timestamp 1751532423
transform 1 0 48272 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_33
timestamp 1751532423
transform 1 0 5040 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_25_66
timestamp 1751532246
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_109
timestamp 1751532440
transform 1 0 13552 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_25_121
timestamp 1751532312
transform 1 0 14896 0 -1 23520
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_139
timestamp 1751532423
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_142
timestamp 1751532440
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_162
timestamp 1751532440
transform 1 0 19488 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_164
timestamp 1751532423
transform 1 0 19712 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_209
timestamp 1751532423
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_25_212
timestamp 1751532246
transform 1 0 25088 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_234
timestamp 1751532440
transform 1 0 27552 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_236
timestamp 1751532423
transform 1 0 27776 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_261
timestamp 1751532440
transform 1 0 30576 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_263
timestamp 1751532423
transform 1 0 30800 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_276
timestamp 1751532440
transform 1 0 32256 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_345
timestamp 1751532440
transform 1 0 39984 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_349
timestamp 1751532423
transform 1 0 40432 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_359
timestamp 1751532440
transform 1 0 41552 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_361
timestamp 1751532423
transform 1 0 41776 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_389
timestamp 1751532440
transform 1 0 44912 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_393
timestamp 1751532423
transform 1 0 45360 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_419
timestamp 1751532423
transform 1 0 48272 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_2
timestamp 1751532440
transform 1 0 1568 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_26_30
timestamp 1751532246
transform 1 0 4704 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_34
timestamp 1751532423
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_26_79
timestamp 1751532312
transform 1 0 10192 0 1 23520
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_26_117
timestamp 1751532246
transform 1 0 14448 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_181
timestamp 1751532440
transform 1 0 21616 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_185
timestamp 1751532440
transform 1 0 22064 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_189
timestamp 1751532440
transform 1 0 22512 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_191
timestamp 1751532423
transform 1 0 22736 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_219
timestamp 1751532423
transform 1 0 25872 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_26_230
timestamp 1751532246
transform 1 0 27104 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_244
timestamp 1751532423
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_257
timestamp 1751532423
transform 1 0 30128 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_295
timestamp 1751532440
transform 1 0 34384 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_297
timestamp 1751532423
transform 1 0 34608 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_324
timestamp 1751532440
transform 1 0 37632 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_341
timestamp 1751532440
transform 1 0 39536 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_361
timestamp 1751532440
transform 1 0 41776 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_365
timestamp 1751532440
transform 1 0 42224 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_369
timestamp 1751532423
transform 1 0 42672 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_383
timestamp 1751532440
transform 1 0 44240 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_404
timestamp 1751532440
transform 1 0 46592 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_417
timestamp 1751532440
transform 1 0 48048 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_419
timestamp 1751532423
transform 1 0 48272 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_2
timestamp 1751532440
transform 1 0 1568 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_4
timestamp 1751532423
transform 1 0 1792 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_55
timestamp 1751532440
transform 1 0 7504 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_67
timestamp 1751532440
transform 1 0 8848 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_69
timestamp 1751532423
transform 1 0 9072 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_79
timestamp 1751532440
transform 1 0 10192 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_81
timestamp 1751532423
transform 1 0 10416 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_27_103
timestamp 1751532246
transform 1 0 12880 0 -1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_107
timestamp 1751532423
transform 1 0 13328 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_27_118
timestamp 1751532246
transform 1 0 14560 0 -1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_122
timestamp 1751532423
transform 1 0 15008 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_129
timestamp 1751532440
transform 1 0 15792 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_137
timestamp 1751532440
transform 1 0 16688 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_139
timestamp 1751532423
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_158
timestamp 1751532440
transform 1 0 19040 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_193
timestamp 1751532423
transform 1 0 22960 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_226
timestamp 1751532440
transform 1 0 26656 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_242
timestamp 1751532440
transform 1 0 28448 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_244
timestamp 1751532423
transform 1 0 28672 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_254
timestamp 1751532440
transform 1 0 29792 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_256
timestamp 1751532423
transform 1 0 30016 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_277
timestamp 1751532440
transform 1 0 32368 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_279
timestamp 1751532423
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_289
timestamp 1751532440
transform 1 0 33712 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_300
timestamp 1751532440
transform 1 0 34944 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_331
timestamp 1751532423
transform 1 0 38416 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_338
timestamp 1751532440
transform 1 0 39200 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_340
timestamp 1751532423
transform 1 0 39424 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_347
timestamp 1751532440
transform 1 0 40208 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_349
timestamp 1751532423
transform 1 0 40432 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_377
timestamp 1751532440
transform 1 0 43568 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_381
timestamp 1751532440
transform 1 0 44016 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_385
timestamp 1751532423
transform 1 0 44464 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_28_2
timestamp 1751532246
transform 1 0 1568 0 1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_6
timestamp 1751532423
transform 1 0 2016 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_34
timestamp 1751532423
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_57
timestamp 1751532440
transform 1 0 7728 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_83
timestamp 1751532440
transform 1 0 10640 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_85
timestamp 1751532423
transform 1 0 10864 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_126
timestamp 1751532440
transform 1 0 15456 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_171
timestamp 1751532440
transform 1 0 20496 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_177
timestamp 1751532440
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_179
timestamp 1751532423
transform 1 0 21392 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_207
timestamp 1751532440
transform 1 0 24528 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_243
timestamp 1751532440
transform 1 0 28560 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_254
timestamp 1751532440
transform 1 0 29792 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_313
timestamp 1751532440
transform 1 0 36400 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_323
timestamp 1751532423
transform 1 0 37520 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_384
timestamp 1751532423
transform 1 0 44352 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_408
timestamp 1751532423
transform 1 0 47040 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_416
timestamp 1751532440
transform 1 0 47936 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_8
timestamp 1751532440
transform 1 0 2240 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_12
timestamp 1751532440
transform 1 0 2688 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_14
timestamp 1751532423
transform 1 0 2912 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_27
timestamp 1751532440
transform 1 0 4368 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_29
timestamp 1751532423
transform 1 0 4592 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_76
timestamp 1751532440
transform 1 0 9856 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_128
timestamp 1751532246
transform 1 0 15680 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_142
timestamp 1751532440
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_166
timestamp 1751532440
transform 1 0 19936 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_168
timestamp 1751532423
transform 1 0 20160 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_187
timestamp 1751532440
transform 1 0 22288 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_191
timestamp 1751532246
transform 1 0 22736 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_195
timestamp 1751532423
transform 1 0 23184 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_236
timestamp 1751532423
transform 1 0 27776 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_268
timestamp 1751532440
transform 1 0 31360 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_272
timestamp 1751532440
transform 1 0 31808 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_276
timestamp 1751532440
transform 1 0 32256 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_294
timestamp 1751532440
transform 1 0 34272 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_298
timestamp 1751532423
transform 1 0 34720 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_326
timestamp 1751532440
transform 1 0 37856 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_343
timestamp 1751532440
transform 1 0 39760 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_347
timestamp 1751532440
transform 1 0 40208 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_349
timestamp 1751532423
transform 1 0 40432 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_365
timestamp 1751532440
transform 1 0 42224 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_418
timestamp 1751532440
transform 1 0 48160 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_30_2
timestamp 1751532312
transform 1 0 1568 0 1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_10
timestamp 1751532423
transform 1 0 2464 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_18
timestamp 1751532440
transform 1 0 3360 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_20
timestamp 1751532423
transform 1 0 3584 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_47
timestamp 1751532440
transform 1 0 6608 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_49
timestamp 1751532423
transform 1 0 6832 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_30_67
timestamp 1751532246
transform 1 0 8848 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_95
timestamp 1751532440
transform 1 0 11984 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_97
timestamp 1751532423
transform 1 0 12208 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_107
timestamp 1751532440
transform 1 0 13328 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_109
timestamp 1751532423
transform 1 0 13552 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_124
timestamp 1751532440
transform 1 0 15232 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_153
timestamp 1751532423
transform 1 0 18480 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_160
timestamp 1751532440
transform 1 0 19264 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_172
timestamp 1751532440
transform 1 0 20608 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_174
timestamp 1751532423
transform 1 0 20832 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_184
timestamp 1751532440
transform 1 0 21952 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_30_199
timestamp 1751532312
transform 1 0 23632 0 1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_230
timestamp 1751532440
transform 1 0 27104 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_265
timestamp 1751532440
transform 1 0 31024 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_314
timestamp 1751532423
transform 1 0 36512 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_30_317
timestamp 1751532246
transform 1 0 36848 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_321
timestamp 1751532423
transform 1 0 37296 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_324
timestamp 1751532440
transform 1 0 37632 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_328
timestamp 1751532440
transform 1 0 38080 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_346
timestamp 1751532423
transform 1 0 40096 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_383
timestamp 1751532440
transform 1 0 44240 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_387
timestamp 1751532440
transform 1 0 44688 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_396
timestamp 1751532423
transform 1 0 45696 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_415
timestamp 1751532440
transform 1 0 47824 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_419
timestamp 1751532423
transform 1 0 48272 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_29
timestamp 1751532423
transform 1 0 4592 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_34
timestamp 1751532423
transform 1 0 5152 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_52
timestamp 1751532440
transform 1 0 7168 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_72
timestamp 1751532423
transform 1 0 9408 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_98
timestamp 1751532440
transform 1 0 12320 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_100
timestamp 1751532423
transform 1 0 12544 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_128
timestamp 1751532246
transform 1 0 15680 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_132
timestamp 1751532440
transform 1 0 16128 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_136
timestamp 1751532440
transform 1 0 16576 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_142
timestamp 1751532423
transform 1 0 17248 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_175
timestamp 1751532440
transform 1 0 20944 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_212
timestamp 1751532440
transform 1 0 25088 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_230
timestamp 1751532440
transform 1 0 27104 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_260
timestamp 1751532440
transform 1 0 30464 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_270
timestamp 1751532246
transform 1 0 31584 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_276
timestamp 1751532440
transform 1 0 32256 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_282
timestamp 1751532440
transform 1 0 32928 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_309
timestamp 1751532246
transform 1 0 35952 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_315
timestamp 1751532440
transform 1 0 36624 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_342
timestamp 1751532423
transform 1 0 39648 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_390
timestamp 1751532440
transform 1 0 45024 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_413
timestamp 1751532423
transform 1 0 47600 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_29
timestamp 1751532440
transform 1 0 4592 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_33
timestamp 1751532440
transform 1 0 5040 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_32_47
timestamp 1751532246
transform 1 0 6608 0 1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_107
timestamp 1751532440
transform 1 0 13328 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_126
timestamp 1751532440
transform 1 0 15456 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_32_134
timestamp 1751532246
transform 1 0 16352 0 1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_138
timestamp 1751532423
transform 1 0 16800 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_141
timestamp 1751532440
transform 1 0 17136 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_166
timestamp 1751532423
transform 1 0 19936 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_174
timestamp 1751532423
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_32_208
timestamp 1751532246
transform 1 0 24640 0 1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_228
timestamp 1751532440
transform 1 0 26880 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_230
timestamp 1751532423
transform 1 0 27104 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_233
timestamp 1751532440
transform 1 0 27440 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_244
timestamp 1751532423
transform 1 0 28672 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_275
timestamp 1751532440
transform 1 0 32144 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_277
timestamp 1751532423
transform 1 0 32368 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_280
timestamp 1751532440
transform 1 0 32704 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_284
timestamp 1751532440
transform 1 0 33152 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_286
timestamp 1751532423
transform 1 0 33376 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_317
timestamp 1751532440
transform 1 0 36848 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_381
timestamp 1751532440
transform 1 0 44016 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_2
timestamp 1751532246
transform 1 0 1568 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_52
timestamp 1751532440
transform 1 0 7168 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_86
timestamp 1751532440
transform 1 0 10976 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_138
timestamp 1751532440
transform 1 0 16800 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_142
timestamp 1751532440
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_177
timestamp 1751532423
transform 1 0 21168 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_198
timestamp 1751532440
transform 1 0 23520 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_202
timestamp 1751532423
transform 1 0 23968 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_222
timestamp 1751532246
transform 1 0 26208 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_228
timestamp 1751532440
transform 1 0 26880 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_257
timestamp 1751532440
transform 1 0 30128 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_259
timestamp 1751532423
transform 1 0 30352 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_276
timestamp 1751532440
transform 1 0 32256 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_282
timestamp 1751532246
transform 1 0 32928 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_302
timestamp 1751532440
transform 1 0 35168 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_306
timestamp 1751532423
transform 1 0 35616 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_339
timestamp 1751532440
transform 1 0 39312 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_362
timestamp 1751532440
transform 1 0 41888 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_366
timestamp 1751532423
transform 1 0 42336 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_394
timestamp 1751532440
transform 1 0 45472 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_411
timestamp 1751532440
transform 1 0 47376 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_413
timestamp 1751532423
transform 1 0 47600 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_34_2
timestamp 1751532312
transform 1 0 1568 0 1 29792
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_10
timestamp 1751532423
transform 1 0 2464 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_32
timestamp 1751532440
transform 1 0 4928 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_34
timestamp 1751532423
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_64
timestamp 1751532423
transform 1 0 8512 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_121
timestamp 1751532423
transform 1 0 14896 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_149
timestamp 1751532440
transform 1 0 18032 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_153
timestamp 1751532423
transform 1 0 18480 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_187
timestamp 1751532440
transform 1 0 22288 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_230
timestamp 1751532440
transform 1 0 27104 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_234
timestamp 1751532423
transform 1 0 27552 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_242
timestamp 1751532440
transform 1 0 28448 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_244
timestamp 1751532423
transform 1 0 28672 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_254
timestamp 1751532440
transform 1 0 29792 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_270
timestamp 1751532440
transform 1 0 31584 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_272
timestamp 1751532423
transform 1 0 31808 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_305
timestamp 1751532440
transform 1 0 35504 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_329
timestamp 1751532440
transform 1 0 38192 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_333
timestamp 1751532423
transform 1 0 38640 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_369
timestamp 1751532440
transform 1 0 42672 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_382
timestamp 1751532440
transform 1 0 44128 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_384
timestamp 1751532423
transform 1 0 44352 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_415
timestamp 1751532440
transform 1 0 47824 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_419
timestamp 1751532423
transform 1 0 48272 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_36
timestamp 1751532440
transform 1 0 5376 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_38
timestamp 1751532423
transform 1 0 5600 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_69
timestamp 1751532423
transform 1 0 9072 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_84
timestamp 1751532440
transform 1 0 10752 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_142
timestamp 1751532440
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_144
timestamp 1751532423
transform 1 0 17472 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_164
timestamp 1751532440
transform 1 0 19712 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_187
timestamp 1751532440
transform 1 0 22288 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_189
timestamp 1751532423
transform 1 0 22512 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_219
timestamp 1751532440
transform 1 0 25872 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_221
timestamp 1751532423
transform 1 0 26096 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_224
timestamp 1751532440
transform 1 0 26432 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_244
timestamp 1751532440
transform 1 0 28672 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_246
timestamp 1751532423
transform 1 0 28896 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_279
timestamp 1751532423
transform 1 0 32592 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_310
timestamp 1751532440
transform 1 0 36064 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_312
timestamp 1751532423
transform 1 0 36288 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_389
timestamp 1751532440
transform 1 0 44912 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_36_2
timestamp 1751532246
transform 1 0 1568 0 1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_12
timestamp 1751532423
transform 1 0 2688 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_34
timestamp 1751532423
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_47
timestamp 1751532440
transform 1 0 6608 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_102
timestamp 1751532440
transform 1 0 12768 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_104
timestamp 1751532423
transform 1 0 12992 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_127
timestamp 1751532440
transform 1 0 15568 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_148
timestamp 1751532440
transform 1 0 17920 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_36_193
timestamp 1751532246
transform 1 0 22960 0 1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_197
timestamp 1751532423
transform 1 0 23408 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_216
timestamp 1751532440
transform 1 0 25536 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_220
timestamp 1751532440
transform 1 0 25984 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_244
timestamp 1751532423
transform 1 0 28672 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_254
timestamp 1751532440
transform 1 0 29792 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_256
timestamp 1751532423
transform 1 0 30016 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_269
timestamp 1751532423
transform 1 0 31472 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_277
timestamp 1751532440
transform 1 0 32368 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_279
timestamp 1751532423
transform 1 0 32592 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_317
timestamp 1751532440
transform 1 0 36848 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_321
timestamp 1751532423
transform 1 0 37296 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_382
timestamp 1751532440
transform 1 0 44128 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_384
timestamp 1751532423
transform 1 0 44352 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_37_2
timestamp 1751532246
transform 1 0 1568 0 -1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_37_12
timestamp 1751532246
transform 1 0 2688 0 -1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_18
timestamp 1751532440
transform 1 0 3360 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_22
timestamp 1751532440
transform 1 0 3808 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_67
timestamp 1751532440
transform 1 0 8848 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_37_69
timestamp 1751532423
transform 1 0 9072 0 -1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_37_78
timestamp 1751532423
transform 1 0 10080 0 -1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_37_158
timestamp 1751532423
transform 1 0 19040 0 -1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_185
timestamp 1751532440
transform 1 0 22064 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_212
timestamp 1751532440
transform 1 0 25088 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_37_269
timestamp 1751532246
transform 1 0 31472 0 -1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_37_273
timestamp 1751532423
transform 1 0 31920 0 -1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_276
timestamp 1751532440
transform 1 0 32256 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_390
timestamp 1751532440
transform 1 0 45024 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_418
timestamp 1751532440
transform 1 0 48160 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_38_29
timestamp 1751532246
transform 1 0 4592 0 1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_37
timestamp 1751532440
transform 1 0 5488 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_97
timestamp 1751532423
transform 1 0 12208 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_131
timestamp 1751532423
transform 1 0 16016 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_156
timestamp 1751532440
transform 1 0 18816 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_38_169
timestamp 1751532246
transform 1 0 20272 0 1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_181
timestamp 1751532423
transform 1 0 21616 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_219
timestamp 1751532440
transform 1 0 25872 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_221
timestamp 1751532423
transform 1 0 26096 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_38_224
timestamp 1751532246
transform 1 0 26432 0 1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_242
timestamp 1751532440
transform 1 0 28448 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_244
timestamp 1751532423
transform 1 0 28672 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_247
timestamp 1751532423
transform 1 0 29008 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_280
timestamp 1751532440
transform 1 0 32704 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_327
timestamp 1751532423
transform 1 0 37968 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_355
timestamp 1751532440
transform 1 0 41104 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_39_2
timestamp 1751532351
transform 1 0 1568 0 -1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_18
timestamp 1751532440
transform 1 0 3360 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_34
timestamp 1751532440
transform 1 0 5152 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_36
timestamp 1751532423
transform 1 0 5376 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_54
timestamp 1751532440
transform 1 0 7392 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_88
timestamp 1751532423
transform 1 0 11200 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_106
timestamp 1751532440
transform 1 0 13216 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_108
timestamp 1751532423
transform 1 0 13440 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_128
timestamp 1751532440
transform 1 0 15680 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_192
timestamp 1751532440
transform 1 0 22848 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_207
timestamp 1751532440
transform 1 0 24528 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_209
timestamp 1751532423
transform 1 0 24752 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_212
timestamp 1751532440
transform 1 0 25088 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_244
timestamp 1751532440
transform 1 0 28672 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_248
timestamp 1751532440
transform 1 0 29120 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_250
timestamp 1751532423
transform 1 0 29344 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_275
timestamp 1751532440
transform 1 0 32144 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_277
timestamp 1751532423
transform 1 0 32368 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_332
timestamp 1751532440
transform 1 0 38528 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_348
timestamp 1751532440
transform 1 0 40320 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_364
timestamp 1751532440
transform 1 0 42112 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_395
timestamp 1751532440
transform 1 0 45584 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_399
timestamp 1751532423
transform 1 0 46032 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_418
timestamp 1751532440
transform 1 0 48160 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_40_2
timestamp 1751532312
transform 1 0 1568 0 1 34496
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_44
timestamp 1751532440
transform 1 0 6272 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_46
timestamp 1751532423
transform 1 0 6496 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_66
timestamp 1751532440
transform 1 0 8736 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_82
timestamp 1751532440
transform 1 0 10528 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_91
timestamp 1751532440
transform 1 0 11536 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_107
timestamp 1751532440
transform 1 0 13328 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_109
timestamp 1751532423
transform 1 0 13552 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_132
timestamp 1751532423
transform 1 0 16128 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_140
timestamp 1751532423
transform 1 0 17024 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_153
timestamp 1751532423
transform 1 0 18480 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_177
timestamp 1751532440
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_179
timestamp 1751532423
transform 1 0 21392 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_199
timestamp 1751532440
transform 1 0 23632 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_201
timestamp 1751532423
transform 1 0 23856 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_230
timestamp 1751532440
transform 1 0 27104 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_232
timestamp 1751532423
transform 1 0 27328 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_40_261
timestamp 1751532246
transform 1 0 30576 0 1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_267
timestamp 1751532440
transform 1 0 31248 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_314
timestamp 1751532423
transform 1 0 36512 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_327
timestamp 1751532440
transform 1 0 37968 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_369
timestamp 1751532440
transform 1 0 42672 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_384
timestamp 1751532423
transform 1 0 44352 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_405
timestamp 1751532423
transform 1 0 46704 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_84
timestamp 1751532423
transform 1 0 10752 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_178
timestamp 1751532440
transform 1 0 21280 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_209
timestamp 1751532423
transform 1 0 24752 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_234
timestamp 1751532440
transform 1 0 27552 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_41_250
timestamp 1751532246
transform 1 0 29344 0 -1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_254
timestamp 1751532423
transform 1 0 29792 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_257
timestamp 1751532440
transform 1 0 30128 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_275
timestamp 1751532440
transform 1 0 32144 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_277
timestamp 1751532423
transform 1 0 32368 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_299
timestamp 1751532440
transform 1 0 34832 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_301
timestamp 1751532423
transform 1 0 35056 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_345
timestamp 1751532440
transform 1 0 39984 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_349
timestamp 1751532423
transform 1 0 40432 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_382
timestamp 1751532423
transform 1 0 44128 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_390
timestamp 1751532423
transform 1 0 45024 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_398
timestamp 1751532423
transform 1 0 45920 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_417
timestamp 1751532440
transform 1 0 48048 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_419
timestamp 1751532423
transform 1 0 48272 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_42_2
timestamp 1751532246
transform 1 0 1568 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_42_12
timestamp 1751532246
transform 1 0 2688 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_16
timestamp 1751532440
transform 1 0 3136 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_37
timestamp 1751532440
transform 1 0 5488 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_41
timestamp 1751532440
transform 1 0 5936 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_58
timestamp 1751532440
transform 1 0 7840 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_87
timestamp 1751532440
transform 1 0 11088 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_103
timestamp 1751532440
transform 1 0 12880 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_114
timestamp 1751532440
transform 1 0 14112 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_118
timestamp 1751532440
transform 1 0 14560 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_120
timestamp 1751532423
transform 1 0 14784 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_191
timestamp 1751532423
transform 1 0 22736 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_247
timestamp 1751532423
transform 1 0 29008 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_262
timestamp 1751532440
transform 1 0 30688 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_264
timestamp 1751532423
transform 1 0 30912 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_296
timestamp 1751532440
transform 1 0 34496 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_298
timestamp 1751532423
transform 1 0 34720 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_311
timestamp 1751532440
transform 1 0 36176 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_344
timestamp 1751532440
transform 1 0 39872 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_368
timestamp 1751532440
transform 1 0 42560 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_383
timestamp 1751532440
transform 1 0 44240 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_62
timestamp 1751532440
transform 1 0 8288 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_66
timestamp 1751532440
transform 1 0 8736 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_72
timestamp 1751532440
transform 1 0 9408 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_86
timestamp 1751532440
transform 1 0 10976 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_90
timestamp 1751532423
transform 1 0 11424 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_115
timestamp 1751532440
transform 1 0 14224 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_121
timestamp 1751532440
transform 1 0 14896 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_43_125
timestamp 1751532246
transform 1 0 15344 0 -1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_129
timestamp 1751532423
transform 1 0 15792 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_138
timestamp 1751532440
transform 1 0 16800 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_43_142
timestamp 1751532246
transform 1 0 17248 0 -1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_165
timestamp 1751532440
transform 1 0 19824 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_195
timestamp 1751532440
transform 1 0 23184 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_205
timestamp 1751532440
transform 1 0 24304 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_207
timestamp 1751532423
transform 1 0 24528 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_212
timestamp 1751532440
transform 1 0 25088 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_214
timestamp 1751532423
transform 1 0 25312 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_227
timestamp 1751532440
transform 1 0 26768 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_229
timestamp 1751532423
transform 1 0 26992 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_244
timestamp 1751532440
transform 1 0 28672 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_43_248
timestamp 1751532246
transform 1 0 29120 0 -1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_252
timestamp 1751532423
transform 1 0 29568 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_255
timestamp 1751532440
transform 1 0 29904 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_259
timestamp 1751532440
transform 1 0 30352 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_263
timestamp 1751532423
transform 1 0 30800 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_278
timestamp 1751532440
transform 1 0 32480 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_309
timestamp 1751532440
transform 1 0 35952 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_352
timestamp 1751532440
transform 1 0 40768 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_372
timestamp 1751532423
transform 1 0 43008 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_379
timestamp 1751532440
transform 1 0 43792 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_388
timestamp 1751532440
transform 1 0 44800 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_390
timestamp 1751532423
transform 1 0 45024 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_419
timestamp 1751532423
transform 1 0 48272 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_44_2
timestamp 1751532246
transform 1 0 1568 0 1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_12
timestamp 1751532440
transform 1 0 2688 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_16
timestamp 1751532440
transform 1 0 3136 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_44_34
timestamp 1751532423
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_37
timestamp 1751532440
transform 1 0 5488 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_44_41
timestamp 1751532246
transform 1 0 5936 0 1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_68
timestamp 1751532440
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_44_107
timestamp 1751532246
transform 1 0 13328 0 1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_140
timestamp 1751532440
transform 1 0 17024 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_144
timestamp 1751532440
transform 1 0 17472 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_148
timestamp 1751532440
transform 1 0 17920 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_44_158
timestamp 1751532246
transform 1 0 19040 0 1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_44_162
timestamp 1751532423
transform 1 0 19488 0 1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_165
timestamp 1751532440
transform 1 0 19824 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_169
timestamp 1751532440
transform 1 0 20272 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_173
timestamp 1751532440
transform 1 0 20720 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_189
timestamp 1751532440
transform 1 0 22512 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_205
timestamp 1751532440
transform 1 0 24304 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_209
timestamp 1751532440
transform 1 0 24752 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_44_211
timestamp 1751532423
transform 1 0 24976 0 1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_214
timestamp 1751532440
transform 1 0 25312 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_44_232
timestamp 1751532423
transform 1 0 27328 0 1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_283
timestamp 1751532440
transform 1 0 33040 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_44_285
timestamp 1751532423
transform 1 0 33264 0 1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_312
timestamp 1751532440
transform 1 0 36288 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_44_314
timestamp 1751532423
transform 1 0 36512 0 1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_348
timestamp 1751532440
transform 1 0 40320 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_44_350
timestamp 1751532423
transform 1 0 40544 0 1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_380
timestamp 1751532440
transform 1 0 43904 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_44_384
timestamp 1751532423
transform 1 0 44352 0 1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_45_2
timestamp 1751532246
transform 1 0 1568 0 -1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_12
timestamp 1751532423
transform 1 0 2688 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_27
timestamp 1751532440
transform 1 0 4368 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_31
timestamp 1751532423
transform 1 0 4816 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_69
timestamp 1751532423
transform 1 0 9072 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_99
timestamp 1751532440
transform 1 0 12432 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_111
timestamp 1751532440
transform 1 0 13776 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_113
timestamp 1751532423
transform 1 0 14000 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_124
timestamp 1751532423
transform 1 0 15232 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_142
timestamp 1751532440
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_171
timestamp 1751532423
transform 1 0 20496 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_190
timestamp 1751532440
transform 1 0 22624 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_194
timestamp 1751532440
transform 1 0 23072 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_196
timestamp 1751532423
transform 1 0 23296 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_233
timestamp 1751532440
transform 1 0 27440 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_251
timestamp 1751532440
transform 1 0 29456 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_253
timestamp 1751532423
transform 1 0 29680 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_264
timestamp 1751532440
transform 1 0 30912 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_278
timestamp 1751532440
transform 1 0 32480 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_296
timestamp 1751532423
transform 1 0 34496 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_321
timestamp 1751532440
transform 1 0 37296 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_347
timestamp 1751532440
transform 1 0 40208 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_349
timestamp 1751532423
transform 1 0 40432 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_369
timestamp 1751532440
transform 1 0 42672 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_417
timestamp 1751532440
transform 1 0 48048 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_419
timestamp 1751532423
transform 1 0 48272 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_46_29
timestamp 1751532246
transform 1 0 4592 0 1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_46_63
timestamp 1751532246
transform 1 0 8400 0 1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_67
timestamp 1751532423
transform 1 0 8848 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_70
timestamp 1751532440
transform 1 0 9184 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_90
timestamp 1751532440
transform 1 0 11424 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_92
timestamp 1751532423
transform 1 0 11648 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_135
timestamp 1751532423
transform 1 0 16464 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_142
timestamp 1751532440
transform 1 0 17248 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_146
timestamp 1751532423
transform 1 0 17696 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_174
timestamp 1751532423
transform 1 0 20832 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_218
timestamp 1751532440
transform 1 0 25760 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_220
timestamp 1751532423
transform 1 0 25984 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_235
timestamp 1751532440
transform 1 0 27664 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_237
timestamp 1751532423
transform 1 0 27888 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_251
timestamp 1751532423
transform 1 0 29456 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_290
timestamp 1751532423
transform 1 0 33824 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_327
timestamp 1751532440
transform 1 0 37968 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_356
timestamp 1751532423
transform 1 0 41216 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_384
timestamp 1751532423
transform 1 0 44352 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_2
timestamp 1751532440
transform 1 0 1568 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_4
timestamp 1751532423
transform 1 0 1792 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_7
timestamp 1751532440
transform 1 0 2128 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_11
timestamp 1751532440
transform 1 0 2576 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_47_38
timestamp 1751532246
transform 1 0 5600 0 -1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_42
timestamp 1751532423
transform 1 0 6048 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_72
timestamp 1751532440
transform 1 0 9408 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_76
timestamp 1751532440
transform 1 0 9856 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_80
timestamp 1751532440
transform 1 0 10304 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_122
timestamp 1751532423
transform 1 0 15008 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_127
timestamp 1751532423
transform 1 0 15568 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_139
timestamp 1751532423
transform 1 0 16912 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_148
timestamp 1751532440
transform 1 0 17920 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_152
timestamp 1751532440
transform 1 0 18368 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_154
timestamp 1751532423
transform 1 0 18592 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_161
timestamp 1751532440
transform 1 0 19376 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_163
timestamp 1751532423
transform 1 0 19600 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_194
timestamp 1751532440
transform 1 0 23072 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_196
timestamp 1751532423
transform 1 0 23296 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_205
timestamp 1751532440
transform 1 0 24304 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_207
timestamp 1751532423
transform 1 0 24528 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_212
timestamp 1751532440
transform 1 0 25088 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_231
timestamp 1751532440
transform 1 0 27216 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_47_249
timestamp 1751532246
transform 1 0 29232 0 -1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_328
timestamp 1751532423
transform 1 0 38080 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_352
timestamp 1751532440
transform 1 0 40768 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_354
timestamp 1751532423
transform 1 0 40992 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_372
timestamp 1751532440
transform 1 0 43008 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_418
timestamp 1751532440
transform 1 0 48160 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_48_2
timestamp 1751532440
transform 1 0 1568 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_48_4
timestamp 1751532423
transform 1 0 1792 0 1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_48_13
timestamp 1751532440
transform 1 0 2800 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_48_15
timestamp 1751532423
transform 1 0 3024 0 1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_48_34
timestamp 1751532423
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_48_78
timestamp 1751532246
transform 1 0 10080 0 1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_48_119
timestamp 1751532423
transform 1 0 14672 0 1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_48_134
timestamp 1751532423
transform 1 0 16352 0 1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_48_221
timestamp 1751532440
transform 1 0 26096 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_48_223
timestamp 1751532423
transform 1 0 26320 0 1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_48_238
timestamp 1751532246
transform 1 0 28000 0 1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_48_242
timestamp 1751532423
transform 1 0 28448 0 1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_48_299
timestamp 1751532440
transform 1 0 34832 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_48_314
timestamp 1751532423
transform 1 0 36512 0 1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_48_327
timestamp 1751532423
transform 1 0 37968 0 1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_48_355
timestamp 1751532423
transform 1 0 41104 0 1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_48_383
timestamp 1751532440
transform 1 0 44240 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_53
timestamp 1751532440
transform 1 0 7280 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_55
timestamp 1751532423
transform 1 0 7504 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_100
timestamp 1751532440
transform 1 0 12544 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_102
timestamp 1751532423
transform 1 0 12768 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_117
timestamp 1751532440
transform 1 0 14448 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_136
timestamp 1751532440
transform 1 0 16576 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_142
timestamp 1751532440
transform 1 0 17248 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_144
timestamp 1751532423
transform 1 0 17472 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_196
timestamp 1751532440
transform 1 0 23296 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_198
timestamp 1751532423
transform 1 0 23520 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_233
timestamp 1751532423
transform 1 0 27440 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_246
timestamp 1751532423
transform 1 0 28896 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_254
timestamp 1751532440
transform 1 0 29792 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_256
timestamp 1751532423
transform 1 0 30016 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_277
timestamp 1751532440
transform 1 0 32368 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_279
timestamp 1751532423
transform 1 0 32592 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_288
timestamp 1751532423
transform 1 0 33600 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_349
timestamp 1751532423
transform 1 0 40432 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_50_8
timestamp 1751532246
transform 1 0 2240 0 1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_50_14
timestamp 1751532440
transform 1 0 2912 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_50_32
timestamp 1751532440
transform 1 0 4928 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_50_34
timestamp 1751532423
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_50_54
timestamp 1751532440
transform 1 0 7392 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_50_63
timestamp 1751532246
transform 1 0 8400 0 1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_50_96
timestamp 1751532440
transform 1 0 12096 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_50_107
timestamp 1751532440
transform 1 0 13328 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_50_109
timestamp 1751532423
transform 1 0 13552 0 1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_50_151
timestamp 1751532440
transform 1 0 18256 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_50_153
timestamp 1751532423
transform 1 0 18480 0 1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_50_160
timestamp 1751532423
transform 1 0 19264 0 1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_50_228
timestamp 1751532440
transform 1 0 26880 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_50_230
timestamp 1751532423
transform 1 0 27104 0 1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_50_247
timestamp 1751532423
transform 1 0 29008 0 1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_50_268
timestamp 1751532423
transform 1 0 31360 0 1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_50_314
timestamp 1751532423
transform 1 0 36512 0 1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_50_324
timestamp 1751532440
transform 1 0 37632 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_50_353
timestamp 1751532423
transform 1 0 40880 0 1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_50_368
timestamp 1751532440
transform 1 0 42560 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_50_382
timestamp 1751532440
transform 1 0 44128 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_50_384
timestamp 1751532423
transform 1 0 44352 0 1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_50_419
timestamp 1751532423
transform 1 0 48272 0 1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_51_2
timestamp 1751532440
transform 1 0 1568 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_51_6
timestamp 1751532440
transform 1 0 2016 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_51_10
timestamp 1751532440
transform 1 0 2464 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_51_14
timestamp 1751532440
transform 1 0 2912 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_51_18
timestamp 1751532440
transform 1 0 3360 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_51_136
timestamp 1751532440
transform 1 0 16576 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_51_142
timestamp 1751532440
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_51_144
timestamp 1751532423
transform 1 0 17472 0 -1 43904
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_51_172
timestamp 1751532423
transform 1 0 20608 0 -1 43904
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_51_216
timestamp 1751532440
transform 1 0 25536 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_51_250
timestamp 1751532423
transform 1 0 29344 0 -1 43904
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_51_366
timestamp 1751532423
transform 1 0 42336 0 -1 43904
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_52_2
timestamp 1751532246
transform 1 0 1568 0 1 43904
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_52_37
timestamp 1751532440
transform 1 0 5488 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_52_39
timestamp 1751532423
transform 1 0 5712 0 1 43904
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_52_89
timestamp 1751532440
transform 1 0 11312 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_52_111
timestamp 1751532423
transform 1 0 13776 0 1 43904
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_52_173
timestamp 1751532440
transform 1 0 20720 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_52_272
timestamp 1751532423
transform 1 0 31808 0 1 43904
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_52_298
timestamp 1751532440
transform 1 0 34720 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_52_300
timestamp 1751532423
transform 1 0 34944 0 1 43904
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_52_342
timestamp 1751532423
transform 1 0 39648 0 1 43904
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_52_384
timestamp 1751532423
transform 1 0 44352 0 1 43904
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_52_419
timestamp 1751532423
transform 1 0 48272 0 1 43904
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_53_2
timestamp 1751532246
transform 1 0 1568 0 -1 45472
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_53_6
timestamp 1751532423
transform 1 0 2016 0 -1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_53_9
timestamp 1751532440
transform 1 0 2352 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_53_13
timestamp 1751532440
transform 1 0 2800 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_53_17
timestamp 1751532440
transform 1 0 3248 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_53_21
timestamp 1751532440
transform 1 0 3696 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_53_25
timestamp 1751532440
transform 1 0 4144 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_53_29
timestamp 1751532440
transform 1 0 4592 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_53_33
timestamp 1751532440
transform 1 0 5040 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_53_41
timestamp 1751532440
transform 1 0 5936 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_53_79
timestamp 1751532423
transform 1 0 10192 0 -1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_53_142
timestamp 1751532440
transform 1 0 17248 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_53_144
timestamp 1751532423
transform 1 0 17472 0 -1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_53_174
timestamp 1751532423
transform 1 0 20832 0 -1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_53_209
timestamp 1751532423
transform 1 0 24752 0 -1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_53_212
timestamp 1751532423
transform 1 0 25088 0 -1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_53_250
timestamp 1751532440
transform 1 0 29344 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_53_252
timestamp 1751532423
transform 1 0 29568 0 -1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_53_282
timestamp 1751532423
transform 1 0 32928 0 -1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_53_310
timestamp 1751532423
transform 1 0 36064 0 -1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_53_364
timestamp 1751532423
transform 1 0 42112 0 -1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_53_392
timestamp 1751532423
transform 1 0 45248 0 -1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_54_2
timestamp 1751532312
transform 1 0 1568 0 1 45472
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_54_10
timestamp 1751532246
transform 1 0 2464 0 1 45472
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_54_14
timestamp 1751532423
transform 1 0 2912 0 1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_54_17
timestamp 1751532440
transform 1 0 3248 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_54_25
timestamp 1751532440
transform 1 0 4144 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_54_27
timestamp 1751532423
transform 1 0 4368 0 1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_54_30
timestamp 1751532440
transform 1 0 4704 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_54_40
timestamp 1751532440
transform 1 0 5824 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_54_42
timestamp 1751532423
transform 1 0 6048 0 1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_54_45
timestamp 1751532440
transform 1 0 6384 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_54_59
timestamp 1751532440
transform 1 0 7952 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_54_67
timestamp 1751532423
transform 1 0 8848 0 1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_54_70
timestamp 1751532246
transform 1 0 9184 0 1 45472
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_54_74
timestamp 1751532423
transform 1 0 9632 0 1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_54_81
timestamp 1751532423
transform 1 0 10416 0 1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_54_104
timestamp 1751532423
transform 1 0 12992 0 1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_54_138
timestamp 1751532423
transform 1 0 16800 0 1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_54_172
timestamp 1751532423
transform 1 0 20608 0 1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_54_212
timestamp 1751532423
transform 1 0 25088 0 1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_54_230
timestamp 1751532440
transform 1 0 27104 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_54_271
timestamp 1751532423
transform 1 0 31696 0 1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input1
timestamp 1751534193
transform 1 0 30128 0 -1 42336
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input2
timestamp 1751534193
transform -1 0 29792 0 1 42336
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input3
timestamp 1751534193
transform -1 0 48384 0 1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input4
timestamp 1751534193
transform -1 0 48384 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input5
timestamp 1751534193
transform -1 0 45360 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input6
timestamp 1751534193
transform -1 0 48384 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input7
timestamp 1751534193
transform -1 0 48384 0 -1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input8
timestamp 1751534193
transform -1 0 48384 0 -1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input9
timestamp 1751534193
transform -1 0 37520 0 1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input10
timestamp 1751534193
transform 1 0 1568 0 1 42336
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input11
timestamp 1751534193
transform 1 0 1568 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output12
timestamp 1751661108
transform -1 0 20384 0 1 45472
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output13
timestamp 1751661108
transform 1 0 21168 0 1 43904
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output14
timestamp 1751661108
transform 1 0 21392 0 1 45472
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output15
timestamp 1751661108
transform 1 0 32032 0 1 45472
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output16
timestamp 1751661108
transform -1 0 34720 0 1 43904
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output17
timestamp 1751661108
transform 1 0 35840 0 1 45472
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output18
timestamp 1751661108
transform 1 0 35056 0 -1 43904
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output19
timestamp 1751661108
transform 1 0 36848 0 1 43904
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output20
timestamp 1751661108
transform 1 0 39648 0 1 45472
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output21
timestamp 1751661108
transform 1 0 39760 0 1 43904
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output22
timestamp 1751661108
transform 1 0 43456 0 1 45472
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output23
timestamp 1751661108
transform -1 0 47488 0 1 43904
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output24
timestamp 1751661108
transform 1 0 44688 0 1 42336
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output25
timestamp 1751661108
transform 1 0 45584 0 -1 42336
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output26
timestamp 1751661108
transform 1 0 13776 0 1 45472
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output27
timestamp 1751661108
transform 1 0 17808 0 -1 43904
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_0_Left_55 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532504
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_0_Right_0
timestamp 1751532504
transform -1 0 48608 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_1_Left_56
timestamp 1751532504
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_1_Right_1
timestamp 1751532504
transform -1 0 48608 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_2_Left_57
timestamp 1751532504
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_2_Right_2
timestamp 1751532504
transform -1 0 48608 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_3_Left_58
timestamp 1751532504
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_3_Right_3
timestamp 1751532504
transform -1 0 48608 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_4_Left_59
timestamp 1751532504
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_4_Right_4
timestamp 1751532504
transform -1 0 48608 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_5_Left_60
timestamp 1751532504
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_5_Right_5
timestamp 1751532504
transform -1 0 48608 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_6_Left_61
timestamp 1751532504
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_6_Right_6
timestamp 1751532504
transform -1 0 48608 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_7_Left_62
timestamp 1751532504
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_7_Right_7
timestamp 1751532504
transform -1 0 48608 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_8_Left_63
timestamp 1751532504
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_8_Right_8
timestamp 1751532504
transform -1 0 48608 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_9_Left_64
timestamp 1751532504
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_9_Right_9
timestamp 1751532504
transform -1 0 48608 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_10_Left_65
timestamp 1751532504
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_10_Right_10
timestamp 1751532504
transform -1 0 48608 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_11_Left_66
timestamp 1751532504
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_11_Right_11
timestamp 1751532504
transform -1 0 48608 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_12_Left_67
timestamp 1751532504
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_12_Right_12
timestamp 1751532504
transform -1 0 48608 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_13_Left_68
timestamp 1751532504
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_13_Right_13
timestamp 1751532504
transform -1 0 48608 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_14_Left_69
timestamp 1751532504
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_14_Right_14
timestamp 1751532504
transform -1 0 48608 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_15_Left_70
timestamp 1751532504
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_15_Right_15
timestamp 1751532504
transform -1 0 48608 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_16_Left_71
timestamp 1751532504
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_16_Right_16
timestamp 1751532504
transform -1 0 48608 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_17_Left_72
timestamp 1751532504
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_17_Right_17
timestamp 1751532504
transform -1 0 48608 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_18_Left_73
timestamp 1751532504
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_18_Right_18
timestamp 1751532504
transform -1 0 48608 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_19_Left_74
timestamp 1751532504
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_19_Right_19
timestamp 1751532504
transform -1 0 48608 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_20_Left_75
timestamp 1751532504
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_20_Right_20
timestamp 1751532504
transform -1 0 48608 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_21_Left_76
timestamp 1751532504
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_21_Right_21
timestamp 1751532504
transform -1 0 48608 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_22_Left_77
timestamp 1751532504
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_22_Right_22
timestamp 1751532504
transform -1 0 48608 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_23_Left_78
timestamp 1751532504
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_23_Right_23
timestamp 1751532504
transform -1 0 48608 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_24_Left_79
timestamp 1751532504
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_24_Right_24
timestamp 1751532504
transform -1 0 48608 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_25_Left_80
timestamp 1751532504
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_25_Right_25
timestamp 1751532504
transform -1 0 48608 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_26_Left_81
timestamp 1751532504
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_26_Right_26
timestamp 1751532504
transform -1 0 48608 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_27_Left_82
timestamp 1751532504
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_27_Right_27
timestamp 1751532504
transform -1 0 48608 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_28_Left_83
timestamp 1751532504
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_28_Right_28
timestamp 1751532504
transform -1 0 48608 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_29_Left_84
timestamp 1751532504
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_29_Right_29
timestamp 1751532504
transform -1 0 48608 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_30_Left_85
timestamp 1751532504
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_30_Right_30
timestamp 1751532504
transform -1 0 48608 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_31_Left_86
timestamp 1751532504
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_31_Right_31
timestamp 1751532504
transform -1 0 48608 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_32_Left_87
timestamp 1751532504
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_32_Right_32
timestamp 1751532504
transform -1 0 48608 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_33_Left_88
timestamp 1751532504
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_33_Right_33
timestamp 1751532504
transform -1 0 48608 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_34_Left_89
timestamp 1751532504
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_34_Right_34
timestamp 1751532504
transform -1 0 48608 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_35_Left_90
timestamp 1751532504
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_35_Right_35
timestamp 1751532504
transform -1 0 48608 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_36_Left_91
timestamp 1751532504
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_36_Right_36
timestamp 1751532504
transform -1 0 48608 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_37_Left_92
timestamp 1751532504
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_37_Right_37
timestamp 1751532504
transform -1 0 48608 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_38_Left_93
timestamp 1751532504
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_38_Right_38
timestamp 1751532504
transform -1 0 48608 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_39_Left_94
timestamp 1751532504
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_39_Right_39
timestamp 1751532504
transform -1 0 48608 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_40_Left_95
timestamp 1751532504
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_40_Right_40
timestamp 1751532504
transform -1 0 48608 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_41_Left_96
timestamp 1751532504
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_41_Right_41
timestamp 1751532504
transform -1 0 48608 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_42_Left_97
timestamp 1751532504
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_42_Right_42
timestamp 1751532504
transform -1 0 48608 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_43_Left_98
timestamp 1751532504
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_43_Right_43
timestamp 1751532504
transform -1 0 48608 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_44_Left_99
timestamp 1751532504
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_44_Right_44
timestamp 1751532504
transform -1 0 48608 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_45_Left_100
timestamp 1751532504
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_45_Right_45
timestamp 1751532504
transform -1 0 48608 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_46_Left_101
timestamp 1751532504
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_46_Right_46
timestamp 1751532504
transform -1 0 48608 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_47_Left_102
timestamp 1751532504
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_47_Right_47
timestamp 1751532504
transform -1 0 48608 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_48_Left_103
timestamp 1751532504
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_48_Right_48
timestamp 1751532504
transform -1 0 48608 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_49_Left_104
timestamp 1751532504
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_49_Right_49
timestamp 1751532504
transform -1 0 48608 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_50_Left_105
timestamp 1751532504
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_50_Right_50
timestamp 1751532504
transform -1 0 48608 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_51_Left_106
timestamp 1751532504
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_51_Right_51
timestamp 1751532504
transform -1 0 48608 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_52_Left_107
timestamp 1751532504
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_52_Right_52
timestamp 1751532504
transform -1 0 48608 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_53_Left_108
timestamp 1751532504
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_53_Right_53
timestamp 1751532504
transform -1 0 48608 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_54_Left_109
timestamp 1751532504
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_54_Right_54
timestamp 1751532504
transform -1 0 48608 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_110
timestamp 1751532504
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_111
timestamp 1751532504
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_112
timestamp 1751532504
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_113
timestamp 1751532504
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_114
timestamp 1751532504
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_115
timestamp 1751532504
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_116
timestamp 1751532504
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_117
timestamp 1751532504
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_118
timestamp 1751532504
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_119
timestamp 1751532504
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_120
timestamp 1751532504
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_121
timestamp 1751532504
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_122
timestamp 1751532504
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_123
timestamp 1751532504
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_124
timestamp 1751532504
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_125
timestamp 1751532504
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_126
timestamp 1751532504
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_127
timestamp 1751532504
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_128
timestamp 1751532504
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_129
timestamp 1751532504
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_130
timestamp 1751532504
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_131
timestamp 1751532504
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_132
timestamp 1751532504
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_133
timestamp 1751532504
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_134
timestamp 1751532504
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_135
timestamp 1751532504
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_136
timestamp 1751532504
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_137
timestamp 1751532504
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_138
timestamp 1751532504
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_139
timestamp 1751532504
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_140
timestamp 1751532504
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_141
timestamp 1751532504
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_142
timestamp 1751532504
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_143
timestamp 1751532504
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_144
timestamp 1751532504
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_145
timestamp 1751532504
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_146
timestamp 1751532504
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_147
timestamp 1751532504
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_148
timestamp 1751532504
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_149
timestamp 1751532504
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_150
timestamp 1751532504
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_151
timestamp 1751532504
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_152
timestamp 1751532504
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_153
timestamp 1751532504
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_154
timestamp 1751532504
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_155
timestamp 1751532504
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_156
timestamp 1751532504
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_157
timestamp 1751532504
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_158
timestamp 1751532504
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_159
timestamp 1751532504
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_160
timestamp 1751532504
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_161
timestamp 1751532504
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_162
timestamp 1751532504
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_163
timestamp 1751532504
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_164
timestamp 1751532504
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_165
timestamp 1751532504
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_166
timestamp 1751532504
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_167
timestamp 1751532504
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_168
timestamp 1751532504
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_169
timestamp 1751532504
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_170
timestamp 1751532504
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_171
timestamp 1751532504
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_172
timestamp 1751532504
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_173
timestamp 1751532504
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_174
timestamp 1751532504
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_175
timestamp 1751532504
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_176
timestamp 1751532504
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_177
timestamp 1751532504
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_178
timestamp 1751532504
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_179
timestamp 1751532504
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_180
timestamp 1751532504
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_181
timestamp 1751532504
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_182
timestamp 1751532504
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_183
timestamp 1751532504
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_184
timestamp 1751532504
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_185
timestamp 1751532504
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_186
timestamp 1751532504
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_187
timestamp 1751532504
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_188
timestamp 1751532504
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_189
timestamp 1751532504
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_190
timestamp 1751532504
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_191
timestamp 1751532504
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_192
timestamp 1751532504
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_193
timestamp 1751532504
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_194
timestamp 1751532504
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_195
timestamp 1751532504
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_196
timestamp 1751532504
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_197
timestamp 1751532504
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_198
timestamp 1751532504
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_199
timestamp 1751532504
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_200
timestamp 1751532504
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_201
timestamp 1751532504
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_202
timestamp 1751532504
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_203
timestamp 1751532504
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_204
timestamp 1751532504
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_205
timestamp 1751532504
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_206
timestamp 1751532504
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_207
timestamp 1751532504
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_208
timestamp 1751532504
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_209
timestamp 1751532504
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_210
timestamp 1751532504
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_211
timestamp 1751532504
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_212
timestamp 1751532504
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_213
timestamp 1751532504
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_214
timestamp 1751532504
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_215
timestamp 1751532504
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_216
timestamp 1751532504
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_217
timestamp 1751532504
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_218
timestamp 1751532504
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_219
timestamp 1751532504
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_220
timestamp 1751532504
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_221
timestamp 1751532504
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_222
timestamp 1751532504
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_223
timestamp 1751532504
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_224
timestamp 1751532504
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_225
timestamp 1751532504
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_226
timestamp 1751532504
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_227
timestamp 1751532504
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_228
timestamp 1751532504
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_229
timestamp 1751532504
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_230
timestamp 1751532504
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_231
timestamp 1751532504
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_232
timestamp 1751532504
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_233
timestamp 1751532504
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_234
timestamp 1751532504
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_235
timestamp 1751532504
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_236
timestamp 1751532504
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_237
timestamp 1751532504
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_238
timestamp 1751532504
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_239
timestamp 1751532504
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_240
timestamp 1751532504
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_241
timestamp 1751532504
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_242
timestamp 1751532504
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_243
timestamp 1751532504
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_244
timestamp 1751532504
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_245
timestamp 1751532504
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_246
timestamp 1751532504
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_247
timestamp 1751532504
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_248
timestamp 1751532504
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_249
timestamp 1751532504
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_250
timestamp 1751532504
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_251
timestamp 1751532504
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_252
timestamp 1751532504
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_253
timestamp 1751532504
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_25_254
timestamp 1751532504
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_25_255
timestamp 1751532504
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_25_256
timestamp 1751532504
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_25_257
timestamp 1751532504
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_25_258
timestamp 1751532504
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_259
timestamp 1751532504
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_260
timestamp 1751532504
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_261
timestamp 1751532504
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_262
timestamp 1751532504
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_263
timestamp 1751532504
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_264
timestamp 1751532504
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_27_265
timestamp 1751532504
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_27_266
timestamp 1751532504
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_27_267
timestamp 1751532504
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_27_268
timestamp 1751532504
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_27_269
timestamp 1751532504
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_270
timestamp 1751532504
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_271
timestamp 1751532504
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_272
timestamp 1751532504
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_273
timestamp 1751532504
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_274
timestamp 1751532504
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_275
timestamp 1751532504
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_29_276
timestamp 1751532504
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_29_277
timestamp 1751532504
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_29_278
timestamp 1751532504
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_29_279
timestamp 1751532504
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_29_280
timestamp 1751532504
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_281
timestamp 1751532504
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_282
timestamp 1751532504
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_283
timestamp 1751532504
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_284
timestamp 1751532504
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_285
timestamp 1751532504
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_286
timestamp 1751532504
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_31_287
timestamp 1751532504
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_31_288
timestamp 1751532504
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_31_289
timestamp 1751532504
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_31_290
timestamp 1751532504
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_31_291
timestamp 1751532504
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_292
timestamp 1751532504
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_293
timestamp 1751532504
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_294
timestamp 1751532504
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_295
timestamp 1751532504
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_296
timestamp 1751532504
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_297
timestamp 1751532504
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_33_298
timestamp 1751532504
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_33_299
timestamp 1751532504
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_33_300
timestamp 1751532504
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_33_301
timestamp 1751532504
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_33_302
timestamp 1751532504
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_303
timestamp 1751532504
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_304
timestamp 1751532504
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_305
timestamp 1751532504
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_306
timestamp 1751532504
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_307
timestamp 1751532504
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_308
timestamp 1751532504
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_35_309
timestamp 1751532504
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_35_310
timestamp 1751532504
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_35_311
timestamp 1751532504
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_35_312
timestamp 1751532504
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_35_313
timestamp 1751532504
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_314
timestamp 1751532504
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_315
timestamp 1751532504
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_316
timestamp 1751532504
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_317
timestamp 1751532504
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_318
timestamp 1751532504
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_319
timestamp 1751532504
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_37_320
timestamp 1751532504
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_37_321
timestamp 1751532504
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_37_322
timestamp 1751532504
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_37_323
timestamp 1751532504
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_37_324
timestamp 1751532504
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_38_325
timestamp 1751532504
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_38_326
timestamp 1751532504
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_38_327
timestamp 1751532504
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_38_328
timestamp 1751532504
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_38_329
timestamp 1751532504
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_38_330
timestamp 1751532504
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_39_331
timestamp 1751532504
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_39_332
timestamp 1751532504
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_39_333
timestamp 1751532504
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_39_334
timestamp 1751532504
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_39_335
timestamp 1751532504
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_40_336
timestamp 1751532504
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_40_337
timestamp 1751532504
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_40_338
timestamp 1751532504
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_40_339
timestamp 1751532504
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_40_340
timestamp 1751532504
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_40_341
timestamp 1751532504
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_41_342
timestamp 1751532504
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_41_343
timestamp 1751532504
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_41_344
timestamp 1751532504
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_41_345
timestamp 1751532504
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_41_346
timestamp 1751532504
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_347
timestamp 1751532504
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_348
timestamp 1751532504
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_349
timestamp 1751532504
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_350
timestamp 1751532504
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_351
timestamp 1751532504
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_352
timestamp 1751532504
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_43_353
timestamp 1751532504
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_43_354
timestamp 1751532504
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_43_355
timestamp 1751532504
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_43_356
timestamp 1751532504
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_43_357
timestamp 1751532504
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_44_358
timestamp 1751532504
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_44_359
timestamp 1751532504
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_44_360
timestamp 1751532504
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_44_361
timestamp 1751532504
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_44_362
timestamp 1751532504
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_44_363
timestamp 1751532504
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_45_364
timestamp 1751532504
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_45_365
timestamp 1751532504
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_45_366
timestamp 1751532504
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_45_367
timestamp 1751532504
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_45_368
timestamp 1751532504
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_46_369
timestamp 1751532504
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_46_370
timestamp 1751532504
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_46_371
timestamp 1751532504
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_46_372
timestamp 1751532504
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_46_373
timestamp 1751532504
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_46_374
timestamp 1751532504
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_47_375
timestamp 1751532504
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_47_376
timestamp 1751532504
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_47_377
timestamp 1751532504
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_47_378
timestamp 1751532504
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_47_379
timestamp 1751532504
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_48_380
timestamp 1751532504
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_48_381
timestamp 1751532504
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_48_382
timestamp 1751532504
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_48_383
timestamp 1751532504
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_48_384
timestamp 1751532504
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_48_385
timestamp 1751532504
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_386
timestamp 1751532504
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_387
timestamp 1751532504
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_388
timestamp 1751532504
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_389
timestamp 1751532504
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_390
timestamp 1751532504
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_50_391
timestamp 1751532504
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_50_392
timestamp 1751532504
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_50_393
timestamp 1751532504
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_50_394
timestamp 1751532504
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_50_395
timestamp 1751532504
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_50_396
timestamp 1751532504
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_51_397
timestamp 1751532504
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_51_398
timestamp 1751532504
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_51_399
timestamp 1751532504
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_51_400
timestamp 1751532504
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_51_401
timestamp 1751532504
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_52_402
timestamp 1751532504
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_52_403
timestamp 1751532504
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_52_404
timestamp 1751532504
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_52_405
timestamp 1751532504
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_52_406
timestamp 1751532504
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_52_407
timestamp 1751532504
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_53_408
timestamp 1751532504
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_53_409
timestamp 1751532504
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_53_410
timestamp 1751532504
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_53_411
timestamp 1751532504
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_53_412
timestamp 1751532504
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_54_413
timestamp 1751532504
transform 1 0 5152 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_54_414
timestamp 1751532504
transform 1 0 8960 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_54_415
timestamp 1751532504
transform 1 0 12768 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_54_416
timestamp 1751532504
transform 1 0 16576 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_54_417
timestamp 1751532504
transform 1 0 20384 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_54_418
timestamp 1751532504
transform 1 0 24192 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_54_419
timestamp 1751532504
transform 1 0 28000 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_54_420
timestamp 1751532504
transform 1 0 31808 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_54_421
timestamp 1751532504
transform 1 0 35616 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_54_422
timestamp 1751532504
transform 1 0 39424 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_54_423
timestamp 1751532504
transform 1 0 43232 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_54_424
timestamp 1751532504
transform 1 0 47040 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_sn76489_28 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532612
transform 1 0 3696 0 1 45472
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_sn76489_29
timestamp 1751532612
transform 1 0 5376 0 1 45472
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_sn76489_30
timestamp 1751532612
transform 1 0 6832 0 1 45472
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_sn76489_31
timestamp 1751532612
transform 1 0 8400 0 1 45472
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_sn76489_32
timestamp 1751532612
transform 1 0 9968 0 1 45472
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_sn76489_33
timestamp 1751532612
transform -1 0 11648 0 1 45472
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_sn76489_34
timestamp 1751532612
transform 1 0 13328 0 1 43904
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_sn76489_35
timestamp 1751532612
transform -1 0 12096 0 1 45472
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_sn76489_36
timestamp 1751532612
transform 1 0 24080 0 1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_sn76489_37
timestamp 1751532612
transform -1 0 25648 0 1 45472
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_sn76489_38
timestamp 1751532612
transform 1 0 31248 0 1 45472
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_sn76489_39
timestamp 1751532612
transform 1 0 29792 0 1 43904
box -86 -86 534 870
<< labels >>
flabel metal3 s 49200 42112 50000 42224 0 FreeSans 448 0 0 0 custom_settings[0]
port 0 nsew signal input
flabel metal3 s 49200 47040 50000 47152 0 FreeSans 448 0 0 0 custom_settings[1]
port 1 nsew signal input
flabel metal3 s 49200 2688 50000 2800 0 FreeSans 448 0 0 0 io_in_1[0]
port 2 nsew signal input
flabel metal3 s 49200 7616 50000 7728 0 FreeSans 448 0 0 0 io_in_1[1]
port 3 nsew signal input
flabel metal3 s 49200 12544 50000 12656 0 FreeSans 448 0 0 0 io_in_1[2]
port 4 nsew signal input
flabel metal3 s 49200 17472 50000 17584 0 FreeSans 448 0 0 0 io_in_1[3]
port 5 nsew signal input
flabel metal3 s 49200 22400 50000 22512 0 FreeSans 448 0 0 0 io_in_1[4]
port 6 nsew signal input
flabel metal3 s 49200 27328 50000 27440 0 FreeSans 448 0 0 0 io_in_1[5]
port 7 nsew signal input
flabel metal3 s 49200 32256 50000 32368 0 FreeSans 448 0 0 0 io_in_1[6]
port 8 nsew signal input
flabel metal3 s 49200 37184 50000 37296 0 FreeSans 448 0 0 0 io_in_1[7]
port 9 nsew signal input
flabel metal3 s 0 41440 800 41552 0 FreeSans 448 0 0 0 io_in_2
port 10 nsew signal input
flabel metal2 s 3584 49200 3696 50000 0 FreeSans 448 90 0 0 io_out[0]
port 11 nsew signal output
flabel metal2 s 19264 49200 19376 50000 0 FreeSans 448 90 0 0 io_out[10]
port 12 nsew signal output
flabel metal2 s 20832 49200 20944 50000 0 FreeSans 448 90 0 0 io_out[11]
port 13 nsew signal output
flabel metal2 s 22400 49200 22512 50000 0 FreeSans 448 90 0 0 io_out[12]
port 14 nsew signal output
flabel metal2 s 23968 49200 24080 50000 0 FreeSans 448 90 0 0 io_out[13]
port 15 nsew signal output
flabel metal2 s 25536 49200 25648 50000 0 FreeSans 448 90 0 0 io_out[14]
port 16 nsew signal output
flabel metal2 s 27104 49200 27216 50000 0 FreeSans 448 90 0 0 io_out[15]
port 17 nsew signal output
flabel metal2 s 28672 49200 28784 50000 0 FreeSans 448 90 0 0 io_out[16]
port 18 nsew signal output
flabel metal2 s 30240 49200 30352 50000 0 FreeSans 448 90 0 0 io_out[17]
port 19 nsew signal output
flabel metal2 s 31808 49200 31920 50000 0 FreeSans 448 90 0 0 io_out[18]
port 20 nsew signal output
flabel metal2 s 33376 49200 33488 50000 0 FreeSans 448 90 0 0 io_out[19]
port 21 nsew signal output
flabel metal2 s 5152 49200 5264 50000 0 FreeSans 448 90 0 0 io_out[1]
port 22 nsew signal output
flabel metal2 s 34944 49200 35056 50000 0 FreeSans 448 90 0 0 io_out[20]
port 23 nsew signal output
flabel metal2 s 36512 49200 36624 50000 0 FreeSans 448 90 0 0 io_out[21]
port 24 nsew signal output
flabel metal2 s 38080 49200 38192 50000 0 FreeSans 448 90 0 0 io_out[22]
port 25 nsew signal output
flabel metal2 s 39648 49200 39760 50000 0 FreeSans 448 90 0 0 io_out[23]
port 26 nsew signal output
flabel metal2 s 41216 49200 41328 50000 0 FreeSans 448 90 0 0 io_out[24]
port 27 nsew signal output
flabel metal2 s 42784 49200 42896 50000 0 FreeSans 448 90 0 0 io_out[25]
port 28 nsew signal output
flabel metal2 s 44352 49200 44464 50000 0 FreeSans 448 90 0 0 io_out[26]
port 29 nsew signal output
flabel metal2 s 45920 49200 46032 50000 0 FreeSans 448 90 0 0 io_out[27]
port 30 nsew signal output
flabel metal2 s 6720 49200 6832 50000 0 FreeSans 448 90 0 0 io_out[2]
port 31 nsew signal output
flabel metal2 s 8288 49200 8400 50000 0 FreeSans 448 90 0 0 io_out[3]
port 32 nsew signal output
flabel metal2 s 9856 49200 9968 50000 0 FreeSans 448 90 0 0 io_out[4]
port 33 nsew signal output
flabel metal2 s 11424 49200 11536 50000 0 FreeSans 448 90 0 0 io_out[5]
port 34 nsew signal output
flabel metal2 s 12992 49200 13104 50000 0 FreeSans 448 90 0 0 io_out[6]
port 35 nsew signal output
flabel metal2 s 14560 49200 14672 50000 0 FreeSans 448 90 0 0 io_out[7]
port 36 nsew signal output
flabel metal2 s 16128 49200 16240 50000 0 FreeSans 448 90 0 0 io_out[8]
port 37 nsew signal output
flabel metal2 s 17696 49200 17808 50000 0 FreeSans 448 90 0 0 io_out[9]
port 38 nsew signal output
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 rst_n
port 39 nsew signal input
flabel metal4 s 4448 3076 4768 46316 0 FreeSans 1280 90 0 0 vdd
port 40 nsew power bidirectional
flabel metal4 s 35168 3076 35488 46316 0 FreeSans 1280 90 0 0 vdd
port 40 nsew power bidirectional
flabel metal4 s 19808 3076 20128 46316 0 FreeSans 1280 90 0 0 vss
port 41 nsew ground bidirectional
flabel metal3 s 0 8288 800 8400 0 FreeSans 448 0 0 0 wb_clk_i
port 42 nsew signal input
rlabel metal1 24976 46256 24976 46256 0 vdd
rlabel metal1 24976 45472 24976 45472 0 vss
rlabel metal2 43400 34384 43400 34384 0 _0000_
rlabel metal2 46200 36792 46200 36792 0 _0001_
rlabel metal3 43848 39368 43848 39368 0 _0002_
rlabel metal2 46200 30576 46200 30576 0 _0003_
rlabel metal2 47656 30688 47656 30688 0 _0004_
rlabel metal3 23464 7672 23464 7672 0 _0005_
rlabel metal3 23240 5880 23240 5880 0 _0006_
rlabel metal3 21560 5880 21560 5880 0 _0007_
rlabel metal2 21112 7616 21112 7616 0 _0008_
rlabel metal2 28504 8624 28504 8624 0 _0009_
rlabel metal2 27384 7056 27384 7056 0 _0010_
rlabel metal2 27048 5488 27048 5488 0 _0011_
rlabel metal2 27160 3920 27160 3920 0 _0012_
rlabel metal3 35504 18312 35504 18312 0 _0013_
rlabel metal2 36232 15736 36232 15736 0 _0014_
rlabel metal2 33208 17304 33208 17304 0 _0015_
rlabel metal2 33768 16464 33768 16464 0 _0016_
rlabel metal2 30576 20552 30576 20552 0 _0017_
rlabel metal2 33544 23688 33544 23688 0 _0018_
rlabel metal2 37576 24976 37576 24976 0 _0019_
rlabel metal3 36120 26320 36120 26320 0 _0020_
rlabel metal2 26712 32088 26712 32088 0 _0021_
rlabel metal3 26264 34832 26264 34832 0 _0022_
rlabel metal2 23688 36848 23688 36848 0 _0023_
rlabel metal2 23632 39704 23632 39704 0 _0024_
rlabel metal2 23576 43120 23576 43120 0 _0025_
rlabel metal2 26040 45360 26040 45360 0 _0026_
rlabel metal3 23800 44520 23800 44520 0 _0027_
rlabel metal2 2408 27440 2408 27440 0 _0028_
rlabel metal3 5040 28728 5040 28728 0 _0029_
rlabel metal2 2352 30968 2352 30968 0 _0030_
rlabel metal2 2352 32760 2352 32760 0 _0031_
rlabel metal2 7000 35952 7000 35952 0 _0032_
rlabel metal2 10192 37352 10192 37352 0 _0033_
rlabel metal2 2352 39032 2352 39032 0 _0034_
rlabel metal2 2408 41608 2408 41608 0 _0035_
rlabel metal2 3080 43960 3080 43960 0 _0036_
rlabel metal2 7112 45080 7112 45080 0 _0037_
rlabel metal2 11144 45360 11144 45360 0 _0038_
rlabel metal2 7224 33040 7224 33040 0 _0039_
rlabel metal3 7560 30296 7560 30296 0 _0040_
rlabel metal3 9576 33432 9576 33432 0 _0041_
rlabel metal2 2352 35672 2352 35672 0 _0042_
rlabel metal2 2352 37240 2352 37240 0 _0043_
rlabel metal3 7952 38808 7952 38808 0 _0044_
rlabel metal2 6608 40600 6608 40600 0 _0045_
rlabel metal2 9688 42448 9688 42448 0 _0046_
rlabel metal3 18144 40600 18144 40600 0 _0047_
rlabel metal2 16856 40712 16856 40712 0 _0048_
rlabel metal2 12376 45360 12376 45360 0 _0049_
rlabel metal2 14112 16744 14112 16744 0 _0050_
rlabel metal3 9968 15176 9968 15176 0 _0051_
rlabel metal2 9688 15736 9688 15736 0 _0052_
rlabel metal3 5376 16744 5376 16744 0 _0053_
rlabel metal2 3080 15792 3080 15792 0 _0054_
rlabel metal2 3136 13944 3136 13944 0 _0055_
rlabel metal2 4816 12152 4816 12152 0 _0056_
rlabel metal2 2912 10808 2912 10808 0 _0057_
rlabel metal2 2408 10136 2408 10136 0 _0058_
rlabel metal2 2688 8456 2688 8456 0 _0059_
rlabel metal2 4144 6888 4144 6888 0 _0060_
rlabel metal2 5656 6160 5656 6160 0 _0061_
rlabel metal3 8792 6104 8792 6104 0 _0062_
rlabel metal3 10416 8344 10416 8344 0 _0063_
rlabel metal2 8232 10248 8232 10248 0 _0064_
rlabel metal2 11368 13272 11368 13272 0 _0065_
rlabel metal2 41664 21560 41664 21560 0 _0066_
rlabel metal2 44016 23128 44016 23128 0 _0067_
rlabel metal2 41496 26040 41496 26040 0 _0068_
rlabel metal2 39256 23464 39256 23464 0 _0069_
rlabel metal2 35784 23240 35784 23240 0 _0070_
rlabel metal2 34496 21000 34496 21000 0 _0071_
rlabel metal2 35784 19936 35784 19936 0 _0072_
rlabel metal2 38472 25816 38472 25816 0 _0073_
rlabel metal2 23240 30296 23240 30296 0 _0074_
rlabel metal2 22568 33656 22568 33656 0 _0075_
rlabel metal2 15848 30520 15848 30520 0 _0076_
rlabel metal2 14840 35952 14840 35952 0 _0077_
rlabel metal2 16464 36568 16464 36568 0 _0078_
rlabel metal3 18480 38248 18480 38248 0 _0079_
rlabel metal2 18648 39928 18648 39928 0 _0080_
rlabel metal2 18424 42224 18424 42224 0 _0081_
rlabel metal2 18536 45024 18536 45024 0 _0082_
rlabel metal3 19712 41384 19712 41384 0 _0083_
rlabel metal2 37240 18368 37240 18368 0 _0084_
rlabel metal2 43008 19880 43008 19880 0 _0085_
rlabel metal3 45304 18312 45304 18312 0 _0086_
rlabel metal2 46536 17136 46536 17136 0 _0087_
rlabel metal2 46424 12040 46424 12040 0 _0088_
rlabel metal3 44688 10584 44688 10584 0 _0089_
rlabel metal2 47544 15456 47544 15456 0 _0090_
rlabel metal2 46256 9912 46256 9912 0 _0091_
rlabel metal3 41328 10584 41328 10584 0 _0092_
rlabel metal3 38192 13048 38192 13048 0 _0093_
rlabel metal2 39032 20608 39032 20608 0 _0094_
rlabel metal2 38696 6832 38696 6832 0 _0095_
rlabel metal3 44912 8232 44912 8232 0 _0096_
rlabel metal3 46312 7336 46312 7336 0 _0097_
rlabel metal3 46760 5208 46760 5208 0 _0098_
rlabel metal3 42448 4200 42448 4200 0 _0099_
rlabel metal2 41832 8624 41832 8624 0 _0100_
rlabel metal2 37688 3640 37688 3640 0 _0101_
rlabel metal2 34552 3640 34552 3640 0 _0102_
rlabel metal2 38136 8400 38136 8400 0 _0103_
rlabel metal2 33768 11312 33768 11312 0 _0104_
rlabel metal3 5096 18312 5096 18312 0 _0105_
rlabel metal2 35504 6776 35504 6776 0 _0106_
rlabel metal2 24248 4760 24248 4760 0 _0107_
rlabel metal2 20440 3808 20440 3808 0 _0108_
rlabel metal2 16296 4200 16296 4200 0 _0109_
rlabel metal2 10920 6384 10920 6384 0 _0110_
rlabel metal2 16408 10024 16408 10024 0 _0111_
rlabel metal2 12712 4648 12712 4648 0 _0112_
rlabel metal3 11592 9016 11592 9016 0 _0113_
rlabel metal2 10920 11312 10920 11312 0 _0114_
rlabel metal2 16296 13496 16296 13496 0 _0115_
rlabel metal2 10248 18592 10248 18592 0 _0116_
rlabel metal2 42504 28784 42504 28784 0 _0117_
rlabel metal2 39424 28056 39424 28056 0 _0118_
rlabel metal2 35112 32816 35112 32816 0 _0119_
rlabel metal3 35448 34328 35448 34328 0 _0120_
rlabel metal2 33768 40656 33768 40656 0 _0121_
rlabel metal2 33768 41944 33768 41944 0 _0122_
rlabel metal2 33096 42280 33096 42280 0 _0123_
rlabel metal2 38696 42308 38696 42308 0 _0124_
rlabel metal2 43064 44408 43064 44408 0 _0125_
rlabel metal2 41608 41720 41608 41720 0 _0126_
rlabel metal2 46032 39928 46032 39928 0 _0127_
rlabel metal2 46312 42000 46312 42000 0 _0128_
rlabel metal2 46200 45136 46200 45136 0 _0129_
rlabel metal2 30520 44744 30520 44744 0 _0130_
rlabel metal2 44632 29624 44632 29624 0 _0131_
rlabel metal2 42952 31248 42952 31248 0 _0132_
rlabel metal2 36232 30520 36232 30520 0 _0133_
rlabel metal2 38920 33544 38920 33544 0 _0134_
rlabel metal2 39256 35224 39256 35224 0 _0135_
rlabel metal2 41832 35952 41832 35952 0 _0136_
rlabel metal2 38416 37240 38416 37240 0 _0137_
rlabel metal3 39480 39032 39480 39032 0 _0138_
rlabel metal2 39312 39368 39312 39368 0 _0139_
rlabel metal2 42168 39536 42168 39536 0 _0140_
rlabel metal3 45976 39592 45976 39592 0 _0141_
rlabel metal2 46200 37800 46200 37800 0 _0142_
rlabel metal2 44184 32816 44184 32816 0 _0143_
rlabel metal2 41944 41608 41944 41608 0 _0144_
rlabel metal2 7224 17864 7224 17864 0 _0145_
rlabel metal2 39256 14728 39256 14728 0 _0146_
rlabel metal3 38304 16072 38304 16072 0 _0147_
rlabel metal3 34328 15288 34328 15288 0 _0148_
rlabel metal2 36232 13888 36232 13888 0 _0149_
rlabel metal2 31472 11480 31472 11480 0 _0150_
rlabel metal2 31864 13300 31864 13300 0 _0151_
rlabel metal2 31528 9016 31528 9016 0 _0152_
rlabel metal2 31080 7056 31080 7056 0 _0153_
rlabel metal2 30408 5096 30408 5096 0 _0154_
rlabel metal2 29624 4704 29624 4704 0 _0155_
rlabel metal3 29344 9912 29344 9912 0 _0156_
rlabel metal3 29176 12152 29176 12152 0 _0157_
rlabel metal2 21224 9184 21224 9184 0 _0158_
rlabel metal2 19544 11760 19544 11760 0 _0159_
rlabel metal2 18088 8400 18088 8400 0 _0160_
rlabel metal2 21784 10696 21784 10696 0 _0161_
rlabel metal3 13104 12040 13104 12040 0 _0162_
rlabel metal2 12376 14056 12376 14056 0 _0163_
rlabel metal2 20104 24808 20104 24808 0 _0164_
rlabel metal3 17024 24920 17024 24920 0 _0165_
rlabel metal2 16576 26488 16576 26488 0 _0166_
rlabel metal2 17976 23464 17976 23464 0 _0167_
rlabel metal2 26600 22680 26600 22680 0 _0168_
rlabel metal2 24472 23408 24472 23408 0 _0169_
rlabel metal2 26600 20440 26600 20440 0 _0170_
rlabel metal3 22512 24920 22512 24920 0 _0171_
rlabel metal2 1848 20496 1848 20496 0 _0172_
rlabel metal2 2352 21784 2352 21784 0 _0173_
rlabel metal2 8904 21112 8904 21112 0 _0174_
rlabel metal3 5152 19880 5152 19880 0 _0175_
rlabel metal2 10528 21560 10528 21560 0 _0176_
rlabel metal3 10024 23128 10024 23128 0 _0177_
rlabel metal3 9744 19432 9744 19432 0 _0178_
rlabel metal2 17080 24248 17080 24248 0 _0179_
rlabel metal3 44688 20888 44688 20888 0 _0180_
rlabel metal3 46872 20552 46872 20552 0 _0181_
rlabel metal2 45864 22792 45864 22792 0 _0182_
rlabel metal2 46200 25312 46200 25312 0 _0183_
rlabel metal2 43288 25928 43288 25928 0 _0184_
rlabel metal2 42840 28448 42840 28448 0 _0185_
rlabel metal2 47544 28952 47544 28952 0 _0186_
rlabel metal2 16072 17976 16072 17976 0 _0187_
rlabel metal2 19544 15904 19544 15904 0 _0188_
rlabel metal3 17248 14616 17248 14616 0 _0189_
rlabel metal2 28168 18816 28168 18816 0 _0190_
rlabel metal2 29288 18032 29288 18032 0 _0191_
rlabel metal3 12488 15512 12488 15512 0 _0192_
rlabel metal2 2968 34552 2968 34552 0 _0193_
rlabel metal2 2688 35224 2688 35224 0 _0194_
rlabel metal3 17024 20552 17024 20552 0 _0195_
rlabel metal2 3248 42336 3248 42336 0 _0196_
rlabel metal3 4536 35784 4536 35784 0 _0197_
rlabel metal3 3276 36456 3276 36456 0 _0198_
rlabel metal2 4928 37352 4928 37352 0 _0199_
rlabel metal2 4088 34356 4088 34356 0 _0200_
rlabel metal2 4984 35644 4984 35644 0 _0201_
rlabel metal2 4452 38024 4452 38024 0 _0202_
rlabel metal2 4424 36624 4424 36624 0 _0203_
rlabel metal3 3220 38024 3220 38024 0 _0204_
rlabel metal2 7756 39536 7756 39536 0 _0205_
rlabel metal2 6860 39368 6860 39368 0 _0206_
rlabel metal2 8232 38743 8232 38743 0 _0207_
rlabel metal3 8260 37352 8260 37352 0 _0208_
rlabel metal2 8960 38696 8960 38696 0 _0209_
rlabel metal3 9912 41272 9912 41272 0 _0210_
rlabel metal3 8288 41048 8288 41048 0 _0211_
rlabel metal2 8344 41202 8344 41202 0 _0212_
rlabel metal2 7280 40712 7280 40712 0 _0213_
rlabel metal2 7896 42392 7896 42392 0 _0214_
rlabel metal2 7000 40656 7000 40656 0 _0215_
rlabel metal2 12040 41664 12040 41664 0 _0216_
rlabel metal2 12600 40802 12600 40802 0 _0217_
rlabel metal2 10696 41627 10696 41627 0 _0218_
rlabel metal2 11536 41664 11536 41664 0 _0219_
rlabel metal2 10024 42056 10024 42056 0 _0220_
rlabel metal2 42392 22792 42392 22792 0 _0221_
rlabel metal2 15344 40656 15344 40656 0 _0222_
rlabel metal2 16072 41440 16072 41440 0 _0223_
rlabel metal2 11816 40656 11816 40656 0 _0224_
rlabel metal2 15848 39984 15848 39984 0 _0225_
rlabel metal2 16296 40059 16296 40059 0 _0226_
rlabel metal2 15922 41850 15922 41850 0 _0227_
rlabel metal2 16520 40460 16520 40460 0 _0228_
rlabel metal2 15960 43596 15960 43596 0 _0229_
rlabel metal2 14308 42952 14308 42952 0 _0230_
rlabel metal2 16184 42784 16184 42784 0 _0231_
rlabel metal2 15960 42644 15960 42644 0 _0232_
rlabel metal3 17724 42728 17724 42728 0 _0233_
rlabel metal3 16800 42728 16800 42728 0 _0234_
rlabel metal2 17192 40824 17192 40824 0 _0235_
rlabel metal2 15288 43176 15288 43176 0 _0236_
rlabel metal2 15624 44268 15624 44268 0 _0237_
rlabel metal2 14392 17024 14392 17024 0 _0238_
rlabel metal3 11480 15064 11480 15064 0 _0239_
rlabel metal2 32424 19572 32424 19572 0 _0240_
rlabel metal3 30548 18200 30548 18200 0 _0241_
rlabel metal2 33040 18284 33040 18284 0 _0242_
rlabel metal2 33208 18648 33208 18648 0 _0243_
rlabel metal2 32872 19754 32872 19754 0 _0244_
rlabel metal2 32648 19082 32648 19082 0 _0245_
rlabel metal2 8344 18151 8344 18151 0 _0246_
rlabel metal3 7448 15400 7448 15400 0 _0247_
rlabel metal3 7112 13496 7112 13496 0 _0248_
rlabel metal2 12544 18200 12544 18200 0 _0249_
rlabel metal2 8596 16632 8596 16632 0 _0250_
rlabel metal2 8568 7986 8568 7986 0 _0251_
rlabel metal2 15428 15960 15428 15960 0 _0252_
rlabel metal2 7560 11256 7560 11256 0 _0253_
rlabel metal2 9744 13608 9744 13608 0 _0254_
rlabel metal3 9240 13608 9240 13608 0 _0255_
rlabel metal2 8232 15456 8232 15456 0 _0256_
rlabel metal3 8064 15288 8064 15288 0 _0257_
rlabel metal3 9212 15288 9212 15288 0 _0258_
rlabel metal2 4984 15344 4984 15344 0 _0259_
rlabel metal2 7336 15938 7336 15938 0 _0260_
rlabel metal2 6440 16108 6440 16108 0 _0261_
rlabel metal2 6664 15624 6664 15624 0 _0262_
rlabel metal2 5096 16576 5096 16576 0 _0263_
rlabel metal2 5320 15245 5320 15245 0 _0264_
rlabel metal2 5656 15204 5656 15204 0 _0265_
rlabel metal3 4480 15288 4480 15288 0 _0266_
rlabel metal2 9016 9722 9016 9722 0 _0267_
rlabel metal2 6328 13571 6328 13571 0 _0268_
rlabel metal2 6664 14028 6664 14028 0 _0269_
rlabel metal3 4760 13720 4760 13720 0 _0270_
rlabel metal2 5992 11290 5992 11290 0 _0271_
rlabel metal2 6104 12180 6104 12180 0 _0272_
rlabel metal3 7224 13048 7224 13048 0 _0273_
rlabel metal2 5208 12824 5208 12824 0 _0274_
rlabel metal3 5488 9016 5488 9016 0 _0275_
rlabel metal2 5208 10541 5208 10541 0 _0276_
rlabel metal3 6216 11480 6216 11480 0 _0277_
rlabel metal2 3304 10696 3304 10696 0 _0278_
rlabel metal2 5992 9716 5992 9716 0 _0279_
rlabel metal2 9856 9576 9856 9576 0 _0280_
rlabel metal3 6832 9912 6832 9912 0 _0281_
rlabel metal2 2632 10304 2632 10304 0 _0282_
rlabel metal2 5488 9044 5488 9044 0 _0283_
rlabel metal3 6384 8904 6384 8904 0 _0284_
rlabel metal2 3080 8344 3080 8344 0 _0285_
rlabel metal2 6104 8268 6104 8268 0 _0286_
rlabel metal2 6328 7504 6328 7504 0 _0287_
rlabel metal2 4536 6776 4536 6776 0 _0288_
rlabel metal3 8512 11368 8512 11368 0 _0289_
rlabel metal2 8008 6621 8008 6621 0 _0290_
rlabel metal2 7000 7532 7000 7532 0 _0291_
rlabel metal2 5208 7168 5208 7168 0 _0292_
rlabel metal2 8680 8120 8680 8120 0 _0293_
rlabel metal2 10248 7392 10248 7392 0 _0294_
rlabel metal2 10024 6328 10024 6328 0 _0295_
rlabel metal3 7896 8904 7896 8904 0 _0296_
rlabel metal2 8848 9912 8848 9912 0 _0297_
rlabel metal2 8904 9100 8904 9100 0 _0298_
rlabel metal2 9688 10836 9688 10836 0 _0299_
rlabel metal2 8568 11704 8568 11704 0 _0300_
rlabel metal2 8568 10500 8568 10500 0 _0301_
rlabel metal3 12124 16632 12124 16632 0 _0302_
rlabel metal2 10808 14616 10808 14616 0 _0303_
rlabel metal2 9874 12451 9874 12451 0 _0304_
rlabel metal2 10248 12656 10248 12656 0 _0305_
rlabel metal3 46620 21672 46620 21672 0 _0306_
rlabel metal2 47376 25480 47376 25480 0 _0307_
rlabel metal2 46648 26964 46648 26964 0 _0308_
rlabel metal2 47824 26348 47824 26348 0 _0309_
rlabel metal2 47684 25704 47684 25704 0 _0310_
rlabel via2 47432 26278 47432 26278 0 _0311_
rlabel metal2 44632 24024 44632 24024 0 _0312_
rlabel metal2 37184 15624 37184 15624 0 _0313_
rlabel metal2 16296 10248 16296 10248 0 _0314_
rlabel metal2 44072 20895 44072 20895 0 _0315_
rlabel metal2 43960 21224 43960 21224 0 _0316_
rlabel metal2 43960 22400 43960 22400 0 _0317_
rlabel metal2 42056 22064 42056 22064 0 _0318_
rlabel metal2 42896 24024 42896 24024 0 _0319_
rlabel metal2 43288 24808 43288 24808 0 _0320_
rlabel metal2 42952 22764 42952 22764 0 _0321_
rlabel metal2 40712 23856 40712 23856 0 _0322_
rlabel metal2 41384 24659 41384 24659 0 _0323_
rlabel metal2 41608 24584 41608 24584 0 _0324_
rlabel metal2 41608 25564 41608 25564 0 _0325_
rlabel metal2 40544 23884 40544 23884 0 _0326_
rlabel metal2 40964 23240 40964 23240 0 _0327_
rlabel metal2 40208 24696 40208 24696 0 _0328_
rlabel metal2 36120 23954 36120 23954 0 _0329_
rlabel metal2 37072 22176 37072 22176 0 _0330_
rlabel metal2 35336 23856 35336 23856 0 _0331_
rlabel metal2 35672 20888 35672 20888 0 _0332_
rlabel metal3 35308 22344 35308 22344 0 _0333_
rlabel metal2 35448 20888 35448 20888 0 _0334_
rlabel metal2 35028 20776 35028 20776 0 _0335_
rlabel metal3 35952 19992 35952 19992 0 _0336_
rlabel metal2 36092 20104 36092 20104 0 _0337_
rlabel metal2 39368 27160 39368 27160 0 _0338_
rlabel metal2 45528 26208 45528 26208 0 _0339_
rlabel metal2 41272 26208 41272 26208 0 _0340_
rlabel metal2 40992 26600 40992 26600 0 _0341_
rlabel metal2 38920 26320 38920 26320 0 _0342_
rlabel metal2 25760 29428 25760 29428 0 _0343_
rlabel metal2 24696 31024 24696 31024 0 _0344_
rlabel metal2 24864 33068 24864 33068 0 _0345_
rlabel metal3 24976 29512 24976 29512 0 _0346_
rlabel metal3 23772 30968 23772 30968 0 _0347_
rlabel metal3 24416 32648 24416 32648 0 _0348_
rlabel metal2 23912 30744 23912 30744 0 _0349_
rlabel metal2 24584 31844 24584 31844 0 _0350_
rlabel metal2 22596 32648 22596 32648 0 _0351_
rlabel metal2 25032 33768 25032 33768 0 _0352_
rlabel metal2 23688 33992 23688 33992 0 _0353_
rlabel metal3 17836 32536 17836 32536 0 _0354_
rlabel metal2 17416 31808 17416 31808 0 _0355_
rlabel metal2 18088 32051 18088 32051 0 _0356_
rlabel metal2 16744 29680 16744 29680 0 _0357_
rlabel metal2 16520 29680 16520 29680 0 _0358_
rlabel metal2 16156 29512 16156 29512 0 _0359_
rlabel metal2 17332 33320 17332 33320 0 _0360_
rlabel metal2 16296 34132 16296 34132 0 _0361_
rlabel metal2 16520 33236 16520 33236 0 _0362_
rlabel metal3 17388 34776 17388 34776 0 _0363_
rlabel metal2 16968 33656 16968 33656 0 _0364_
rlabel metal2 18480 35840 18480 35840 0 _0365_
rlabel metal2 19208 35243 19208 35243 0 _0366_
rlabel metal2 21056 36064 21056 36064 0 _0367_
rlabel metal3 18816 37240 18816 37240 0 _0368_
rlabel metal2 20440 36512 20440 36512 0 _0369_
rlabel metal2 18928 37156 18928 37156 0 _0370_
rlabel metal2 20664 37352 20664 37352 0 _0371_
rlabel metal3 22232 37240 22232 37240 0 _0372_
rlabel metal2 21672 36232 21672 36232 0 _0373_
rlabel metal3 21700 36456 21700 36456 0 _0374_
rlabel metal2 23184 41804 23184 41804 0 _0375_
rlabel metal2 22232 36792 22232 36792 0 _0376_
rlabel metal3 20860 36680 20860 36680 0 _0377_
rlabel metal3 20748 39592 20748 39592 0 _0378_
rlabel metal2 22456 39144 22456 39144 0 _0379_
rlabel metal2 21112 38886 21112 38886 0 _0380_
rlabel metal2 22008 38771 22008 38771 0 _0381_
rlabel metal3 22232 40376 22232 40376 0 _0382_
rlabel metal2 19320 40264 19320 40264 0 _0383_
rlabel metal3 23072 41944 23072 41944 0 _0384_
rlabel metal2 21840 41076 21840 41076 0 _0385_
rlabel metal3 23548 41160 23548 41160 0 _0386_
rlabel metal2 23016 41496 23016 41496 0 _0387_
rlabel metal2 22736 41440 22736 41440 0 _0388_
rlabel metal2 21784 42672 21784 42672 0 _0389_
rlabel metal2 22904 43400 22904 43400 0 _0390_
rlabel metal2 22680 43302 22680 43302 0 _0391_
rlabel metal2 23996 43624 23996 43624 0 _0392_
rlabel metal2 23128 43960 23128 43960 0 _0393_
rlabel metal2 24444 44184 24444 44184 0 _0394_
rlabel metal2 21000 44520 21000 44520 0 _0395_
rlabel metal3 21784 42840 21784 42840 0 _0396_
rlabel metal2 20104 41664 20104 41664 0 _0397_
rlabel metal2 38024 10192 38024 10192 0 _0398_
rlabel metal2 39032 11256 39032 11256 0 _0399_
rlabel metal2 40824 17808 40824 17808 0 _0400_
rlabel metal2 43288 16184 43288 16184 0 _0401_
rlabel metal2 43736 16800 43736 16800 0 _0402_
rlabel metal2 42448 14056 42448 14056 0 _0403_
rlabel metal3 42728 13608 42728 13608 0 _0404_
rlabel metal2 42504 14168 42504 14168 0 _0405_
rlabel metal2 40936 15960 40936 15960 0 _0406_
rlabel metal3 39704 18312 39704 18312 0 _0407_
rlabel metal2 34664 23408 34664 23408 0 _0408_
rlabel metal3 39816 18424 39816 18424 0 _0409_
rlabel metal2 41328 18480 41328 18480 0 _0410_
rlabel metal2 24248 10948 24248 10948 0 _0411_
rlabel metal2 43736 18564 43736 18564 0 _0412_
rlabel metal2 42392 15624 42392 15624 0 _0413_
rlabel metal2 42056 18144 42056 18144 0 _0414_
rlabel metal2 42168 18704 42168 18704 0 _0415_
rlabel metal2 43736 17584 43736 17584 0 _0416_
rlabel metal2 44520 19936 44520 19936 0 _0417_
rlabel metal3 44352 19208 44352 19208 0 _0418_
rlabel metal2 44100 19432 44100 19432 0 _0419_
rlabel metal2 44072 19740 44072 19740 0 _0420_
rlabel metal3 44296 17640 44296 17640 0 _0421_
rlabel metal2 43960 18132 43960 18132 0 _0422_
rlabel metal2 44884 16856 44884 16856 0 _0423_
rlabel metal2 45976 19488 45976 19488 0 _0424_
rlabel metal3 45500 19208 45500 19208 0 _0425_
rlabel metal2 44718 18668 44718 18668 0 _0426_
rlabel metal2 43400 6104 43400 6104 0 _0427_
rlabel metal2 45416 16452 45416 16452 0 _0428_
rlabel metal2 44744 15702 44744 15702 0 _0429_
rlabel metal2 44296 15624 44296 15624 0 _0430_
rlabel metal2 44856 14280 44856 14280 0 _0431_
rlabel metal2 44912 16072 44912 16072 0 _0432_
rlabel metal3 45556 16296 45556 16296 0 _0433_
rlabel metal3 18368 3528 18368 3528 0 _0434_
rlabel metal3 47656 16072 47656 16072 0 _0435_
rlabel metal3 47348 16856 47348 16856 0 _0436_
rlabel via1 46398 16872 46398 16872 0 _0437_
rlabel metal2 43400 15344 43400 15344 0 _0438_
rlabel metal2 45752 13776 45752 13776 0 _0439_
rlabel metal2 45864 12852 45864 12852 0 _0440_
rlabel metal2 45752 13132 45752 13132 0 _0441_
rlabel metal2 48160 12376 48160 12376 0 _0442_
rlabel metal2 46510 12396 46510 12396 0 _0443_
rlabel metal2 40824 11088 40824 11088 0 _0444_
rlabel metal2 43960 15624 43960 15624 0 _0445_
rlabel metal2 44156 15848 44156 15848 0 _0446_
rlabel metal2 43848 11522 43848 11522 0 _0447_
rlabel metal2 40264 10976 40264 10976 0 _0448_
rlabel metal2 42840 11256 42840 11256 0 _0449_
rlabel metal2 42952 11508 42952 11508 0 _0450_
rlabel metal3 43176 13720 43176 13720 0 _0451_
rlabel metal3 45528 15176 45528 15176 0 _0452_
rlabel metal2 45192 12096 45192 12096 0 _0453_
rlabel metal2 47376 15176 47376 15176 0 _0454_
rlabel metal2 46468 15772 46468 15772 0 _0455_
rlabel metal2 41160 12712 41160 12712 0 _0456_
rlabel metal3 46032 12152 46032 12152 0 _0457_
rlabel metal2 45864 11573 45864 11573 0 _0458_
rlabel metal3 45444 11928 45444 11928 0 _0459_
rlabel metal2 47544 6272 47544 6272 0 _0460_
rlabel metal3 47628 10584 47628 10584 0 _0461_
rlabel metal2 46510 11292 46510 11292 0 _0462_
rlabel metal2 41272 12342 41272 12342 0 _0463_
rlabel metal3 41020 12152 41020 12152 0 _0464_
rlabel metal2 41832 12103 41832 12103 0 _0465_
rlabel metal2 40600 11284 40600 11284 0 _0466_
rlabel metal3 39704 19992 39704 19992 0 _0467_
rlabel metal3 40516 9800 40516 9800 0 _0468_
rlabel metal2 40936 10724 40936 10724 0 _0469_
rlabel metal3 16184 11368 16184 11368 0 _0470_
rlabel metal3 37128 12152 37128 12152 0 _0471_
rlabel metal2 37772 12152 37772 12152 0 _0472_
rlabel metal2 37352 13048 37352 13048 0 _0473_
rlabel metal3 21224 15960 21224 15960 0 _0474_
rlabel metal2 37884 11928 37884 11928 0 _0475_
rlabel metal2 38696 17304 38696 17304 0 _0476_
rlabel metal2 40040 19712 40040 19712 0 _0477_
rlabel metal2 39928 19852 39928 19852 0 _0478_
rlabel metal2 37940 5880 37940 5880 0 _0479_
rlabel metal3 40992 7448 40992 7448 0 _0480_
rlabel metal2 40040 7924 40040 7924 0 _0481_
rlabel metal2 39704 7784 39704 7784 0 _0482_
rlabel metal2 41384 6216 41384 6216 0 _0483_
rlabel metal2 39816 7000 39816 7000 0 _0484_
rlabel metal2 39256 6804 39256 6804 0 _0485_
rlabel metal2 39592 8120 39592 8120 0 _0486_
rlabel metal2 37520 5880 37520 5880 0 _0487_
rlabel metal2 37296 6048 37296 6048 0 _0488_
rlabel metal2 43120 5656 43120 5656 0 _0489_
rlabel metal3 42504 5880 42504 5880 0 _0490_
rlabel metal2 42616 7392 42616 7392 0 _0491_
rlabel metal2 42728 7476 42728 7476 0 _0492_
rlabel metal2 43456 7784 43456 7784 0 _0493_
rlabel metal2 46368 4312 46368 4312 0 _0494_
rlabel metal2 46704 6888 46704 6888 0 _0495_
rlabel metal2 44158 8383 44158 8383 0 _0496_
rlabel metal3 43568 6664 43568 6664 0 _0497_
rlabel metal2 44072 7140 44072 7140 0 _0498_
rlabel metal2 44016 6048 44016 6048 0 _0499_
rlabel metal2 46956 5992 46956 5992 0 _0500_
rlabel metal2 45012 7524 45012 7524 0 _0501_
rlabel via2 43960 5088 43960 5088 0 _0502_
rlabel metal2 44856 4788 44856 4788 0 _0503_
rlabel metal3 42336 5208 42336 5208 0 _0504_
rlabel metal2 45136 5320 45136 5320 0 _0505_
rlabel metal2 45528 6188 45528 6188 0 _0506_
rlabel metal2 47432 6048 47432 6048 0 _0507_
rlabel via2 45838 5896 45838 5896 0 _0508_
rlabel metal3 40488 5880 40488 5880 0 _0509_
rlabel metal2 40376 5012 40376 5012 0 _0510_
rlabel metal2 42224 4060 42224 4060 0 _0511_
rlabel metal2 41720 4732 41720 4732 0 _0512_
rlabel metal3 24500 3640 24500 3640 0 _0513_
rlabel metal3 44996 3528 44996 3528 0 _0514_
rlabel metal2 41440 4396 41440 4396 0 _0515_
rlabel metal2 40040 5824 40040 5824 0 _0516_
rlabel via1 41515 5080 41515 5080 0 _0517_
rlabel metal2 41272 5432 41272 5432 0 _0518_
rlabel metal2 40320 9184 40320 9184 0 _0519_
rlabel metal2 42000 8484 42000 8484 0 _0520_
rlabel metal2 46172 3304 46172 3304 0 _0521_
rlabel metal3 40432 5096 40432 5096 0 _0522_
rlabel via2 37128 3509 37128 3509 0 _0523_
rlabel metal3 40264 5488 40264 5488 0 _0524_
rlabel metal2 25480 3696 25480 3696 0 _0525_
rlabel metal2 38808 4088 38808 4088 0 _0526_
rlabel metal2 39816 3780 39816 3780 0 _0527_
rlabel metal3 34832 5768 34832 5768 0 _0528_
rlabel metal2 34888 5264 34888 5264 0 _0529_
rlabel metal2 33992 4013 33992 4013 0 _0530_
rlabel metal2 34244 5656 34244 5656 0 _0531_
rlabel metal2 35672 5376 35672 5376 0 _0532_
rlabel metal2 34638 3452 34638 3452 0 _0533_
rlabel metal2 35000 9486 35000 9486 0 _0534_
rlabel metal2 35672 8512 35672 8512 0 _0535_
rlabel metal3 35224 11256 35224 11256 0 _0536_
rlabel metal3 36456 8344 36456 8344 0 _0537_
rlabel metal2 38696 9912 38696 9912 0 _0538_
rlabel metal2 38584 9324 38584 9324 0 _0539_
rlabel metal2 35168 11508 35168 11508 0 _0540_
rlabel metal3 34608 11368 34608 11368 0 _0541_
rlabel metal3 34692 11592 34692 11592 0 _0542_
rlabel metal2 6888 17995 6888 17995 0 _0543_
rlabel metal3 46872 19152 46872 19152 0 _0544_
rlabel metal2 6020 17864 6020 17864 0 _0545_
rlabel metal2 6160 18676 6160 18676 0 _0546_
rlabel metal2 33740 7560 33740 7560 0 _0547_
rlabel metal2 18424 4816 18424 4816 0 _0548_
rlabel metal2 18536 6524 18536 6524 0 _0549_
rlabel metal3 17472 11480 17472 11480 0 _0550_
rlabel metal2 17864 6552 17864 6552 0 _0551_
rlabel metal2 18312 6328 18312 6328 0 _0552_
rlabel metal2 19656 6608 19656 6608 0 _0553_
rlabel metal2 24808 4592 24808 4592 0 _0554_
rlabel metal2 34776 7672 34776 7672 0 _0555_
rlabel metal3 35364 8232 35364 8232 0 _0556_
rlabel metal2 24528 4312 24528 4312 0 _0557_
rlabel metal2 23240 5124 23240 5124 0 _0558_
rlabel metal2 24332 4200 24332 4200 0 _0559_
rlabel metal3 25620 3528 25620 3528 0 _0560_
rlabel metal2 25436 4216 25436 4216 0 _0561_
rlabel metal3 19656 5096 19656 5096 0 _0562_
rlabel metal2 19320 4200 19320 4200 0 _0563_
rlabel metal2 19208 3836 19208 3836 0 _0564_
rlabel metal3 19740 3304 19740 3304 0 _0565_
rlabel metal2 22456 3864 22456 3864 0 _0566_
rlabel metal3 22596 4424 22596 4424 0 _0567_
rlabel metal2 20956 3623 20956 3623 0 _0568_
rlabel metal2 15400 4676 15400 4676 0 _0569_
rlabel via2 16520 5887 16520 5887 0 _0570_
rlabel metal2 15624 5040 15624 5040 0 _0571_
rlabel metal2 15512 5096 15512 5096 0 _0572_
rlabel metal2 15148 5880 15148 5880 0 _0573_
rlabel metal2 16072 4396 16072 4396 0 _0574_
rlabel metal2 17864 3584 17864 3584 0 _0575_
rlabel metal3 16940 3528 16940 3528 0 _0576_
rlabel metal2 16382 4388 16382 4388 0 _0577_
rlabel metal2 15960 8736 15960 8736 0 _0578_
rlabel metal3 13384 7336 13384 7336 0 _0579_
rlabel metal2 13160 6300 13160 6300 0 _0580_
rlabel metal2 13944 6860 13944 6860 0 _0581_
rlabel metal2 12880 5096 12880 5096 0 _0582_
rlabel via1 12535 5896 12535 5896 0 _0583_
rlabel metal3 17472 7448 17472 7448 0 _0584_
rlabel metal2 15940 7224 15940 7224 0 _0585_
rlabel metal2 16128 7560 16128 7560 0 _0586_
rlabel metal2 17892 10696 17892 10696 0 _0587_
rlabel metal2 16912 10780 16912 10780 0 _0588_
rlabel metal2 15288 6216 15288 6216 0 _0589_
rlabel metal2 14448 5068 14448 5068 0 _0590_
rlabel metal2 15176 6832 15176 6832 0 _0591_
rlabel metal2 13972 3528 13972 3528 0 _0592_
rlabel metal2 13676 4796 13676 4796 0 _0593_
rlabel metal2 13832 9912 13832 9912 0 _0594_
rlabel metal2 12600 9268 12600 9268 0 _0595_
rlabel metal3 14140 10024 14140 10024 0 _0596_
rlabel metal3 13076 8232 13076 8232 0 _0597_
rlabel metal2 11872 9604 11872 9604 0 _0598_
rlabel metal2 15624 9408 15624 9408 0 _0599_
rlabel metal2 14392 10528 14392 10528 0 _0600_
rlabel metal2 13384 10668 13384 10668 0 _0601_
rlabel metal2 15232 10864 15232 10864 0 _0602_
rlabel metal2 16016 11648 16016 11648 0 _0603_
rlabel via2 15150 11351 15150 11351 0 _0604_
rlabel metal2 14952 13272 14952 13272 0 _0605_
rlabel metal2 15176 13328 15176 13328 0 _0606_
rlabel metal3 18396 13720 18396 13720 0 _0607_
rlabel metal2 16912 13636 16912 13636 0 _0608_
rlabel metal3 13272 16072 13272 16072 0 _0609_
rlabel metal3 13412 15288 13412 15288 0 _0610_
rlabel metal2 45640 23296 45640 23296 0 _0611_
rlabel metal3 35438 28616 35438 28616 0 _0612_
rlabel metal3 40488 30184 40488 30184 0 _0613_
rlabel metal2 41384 29876 41384 29876 0 _0614_
rlabel metal2 41160 27776 41160 27776 0 _0615_
rlabel metal2 41160 28476 41160 28476 0 _0616_
rlabel metal2 36344 29512 36344 29512 0 _0617_
rlabel metal2 37220 29484 37220 29484 0 _0618_
rlabel metal2 37464 29008 37464 29008 0 _0619_
rlabel metal2 38304 27832 38304 27832 0 _0620_
rlabel metal3 37912 27832 37912 27832 0 _0621_
rlabel metal2 38892 27832 38892 27832 0 _0622_
rlabel metal3 34076 31752 34076 31752 0 _0623_
rlabel metal2 34552 30968 34552 30968 0 _0624_
rlabel metal2 33972 31108 33972 31108 0 _0625_
rlabel metal3 34878 30968 34878 30968 0 _0626_
rlabel metal2 39032 32480 39032 32480 0 _0627_
rlabel metal2 36344 31136 36344 31136 0 _0628_
rlabel metal2 38808 29736 38808 29736 0 _0629_
rlabel metal2 33768 30800 33768 30800 0 _0630_
rlabel metal2 35448 40544 35448 40544 0 _0631_
rlabel metal2 33656 32088 33656 32088 0 _0632_
rlabel metal2 33404 31864 33404 31864 0 _0633_
rlabel metal2 36568 34384 36568 34384 0 _0634_
rlabel metal2 33972 33600 33972 33600 0 _0635_
rlabel metal2 35691 34048 35691 34048 0 _0636_
rlabel metal2 35504 33880 35504 33880 0 _0637_
rlabel metal3 35672 33320 35672 33320 0 _0638_
rlabel metal2 34720 33824 34720 33824 0 _0639_
rlabel metal3 37240 35000 37240 35000 0 _0640_
rlabel metal2 37296 34104 37296 34104 0 _0641_
rlabel metal2 34552 39480 34552 39480 0 _0642_
rlabel metal2 35336 39088 35336 39088 0 _0643_
rlabel metal2 35112 38920 35112 38920 0 _0644_
rlabel metal3 35700 38808 35700 38808 0 _0645_
rlabel metal2 36232 38668 36232 38668 0 _0646_
rlabel metal3 35504 38920 35504 38920 0 _0647_
rlabel metal2 34944 41944 34944 41944 0 _0648_
rlabel metal3 37184 41832 37184 41832 0 _0649_
rlabel metal2 37016 41847 37016 41847 0 _0650_
rlabel metal3 36372 41384 36372 41384 0 _0651_
rlabel metal3 37576 42056 37576 42056 0 _0652_
rlabel metal2 34328 42056 34328 42056 0 _0653_
rlabel metal2 38080 43652 38080 43652 0 _0654_
rlabel metal3 36400 44184 36400 44184 0 _0655_
rlabel metal2 36680 45388 36680 45388 0 _0656_
rlabel metal3 36876 45864 36876 45864 0 _0657_
rlabel metal2 42448 42980 42448 42980 0 _0658_
rlabel metal2 38920 45640 38920 45640 0 _0659_
rlabel metal2 33656 45360 33656 45360 0 _0660_
rlabel metal2 40180 42168 40180 42168 0 _0661_
rlabel metal2 42504 44688 42504 44688 0 _0662_
rlabel metal3 39032 44800 39032 44800 0 _0663_
rlabel metal2 40488 43064 40488 43064 0 _0664_
rlabel metal2 40264 40936 40264 40936 0 _0665_
rlabel metal2 40124 40152 40124 40152 0 _0666_
rlabel metal2 42168 43792 42168 43792 0 _0667_
rlabel metal2 41104 43624 41104 43624 0 _0668_
rlabel metal2 43288 44337 43288 44337 0 _0669_
rlabel metal2 47544 44856 47544 44856 0 _0670_
rlabel metal2 42280 42952 42280 42952 0 _0671_
rlabel metal2 48048 43960 48048 43960 0 _0672_
rlabel metal2 42616 40880 42616 40880 0 _0673_
rlabel metal2 43960 41365 43960 41365 0 _0674_
rlabel metal2 43456 42700 43456 42700 0 _0675_
rlabel metal2 41832 41104 41832 41104 0 _0676_
rlabel via2 41496 41152 41496 41152 0 _0677_
rlabel metal4 46424 40656 46424 40656 0 _0678_
rlabel metal3 46088 40376 46088 40376 0 _0679_
rlabel metal3 46872 37240 46872 37240 0 _0680_
rlabel metal2 25088 22092 25088 22092 0 _0681_
rlabel metal2 46256 39368 46256 39368 0 _0682_
rlabel metal2 44016 42336 44016 42336 0 _0683_
rlabel metal3 46648 43624 46648 43624 0 _0684_
rlabel metal2 43064 43247 43064 43247 0 _0685_
rlabel metal3 45920 43512 45920 43512 0 _0686_
rlabel metal2 47404 37240 47404 37240 0 _0687_
rlabel metal2 47600 45752 47600 45752 0 _0688_
rlabel metal2 48048 36792 48048 36792 0 _0689_
rlabel metal2 45416 35756 45416 35756 0 _0690_
rlabel metal2 17696 44856 17696 44856 0 _0691_
rlabel metal2 44632 40656 44632 40656 0 _0692_
rlabel metal2 41272 38024 41272 38024 0 _0693_
rlabel metal2 43512 30332 43512 30332 0 _0694_
rlabel metal2 43736 30072 43736 30072 0 _0695_
rlabel metal2 43624 30604 43624 30604 0 _0696_
rlabel metal2 43008 37240 43008 37240 0 _0697_
rlabel metal2 41496 33992 41496 33992 0 _0698_
rlabel metal2 42308 33544 42308 33544 0 _0699_
rlabel metal2 39704 31024 39704 31024 0 _0700_
rlabel metal2 38976 30352 38976 30352 0 _0701_
rlabel metal2 39704 34216 39704 34216 0 _0702_
rlabel metal2 41720 35154 41720 35154 0 _0703_
rlabel via2 41944 34874 41944 34874 0 _0704_
rlabel metal2 40432 31360 40432 31360 0 _0705_
rlabel metal2 39144 33544 39144 33544 0 _0706_
rlabel metal2 38808 33152 38808 33152 0 _0707_
rlabel metal3 40488 32536 40488 32536 0 _0708_
rlabel metal2 39592 32760 39592 32760 0 _0709_
rlabel metal3 40460 34104 40460 34104 0 _0710_
rlabel metal3 37688 35672 37688 35672 0 _0711_
rlabel metal2 42448 35168 42448 35168 0 _0712_
rlabel metal2 38136 35616 38136 35616 0 _0713_
rlabel metal2 40824 35728 40824 35728 0 _0714_
rlabel metal2 43512 40152 43512 40152 0 _0715_
rlabel metal2 35224 36568 35224 36568 0 _0716_
rlabel metal2 39480 35784 39480 35784 0 _0717_
rlabel metal3 40628 35672 40628 35672 0 _0718_
rlabel metal2 39704 40432 39704 40432 0 _0719_
rlabel metal2 40348 36680 40348 36680 0 _0720_
rlabel metal3 37352 37128 37352 37128 0 _0721_
rlabel metal2 38360 37884 38360 37884 0 _0722_
rlabel metal2 41720 39116 41720 39116 0 _0723_
rlabel metal2 44408 38766 44408 38766 0 _0724_
rlabel metal2 42112 38304 42112 38304 0 _0725_
rlabel metal2 38584 39536 38584 39536 0 _0726_
rlabel metal2 39592 38976 39592 38976 0 _0727_
rlabel metal2 37128 39144 37128 39144 0 _0728_
rlabel metal2 39480 40432 39480 40432 0 _0729_
rlabel metal2 39172 40152 39172 40152 0 _0730_
rlabel metal2 42420 38920 42420 38920 0 _0731_
rlabel metal3 42224 40376 42224 40376 0 _0732_
rlabel metal2 42784 40600 42784 40600 0 _0733_
rlabel metal2 45948 38920 45948 38920 0 _0734_
rlabel metal2 44408 39816 44408 39816 0 _0735_
rlabel metal3 45472 35560 45472 35560 0 _0736_
rlabel metal3 45247 38808 45247 38808 0 _0737_
rlabel metal3 47376 38808 47376 38808 0 _0738_
rlabel metal2 47488 38976 47488 38976 0 _0739_
rlabel metal2 43400 31962 43400 31962 0 _0740_
rlabel metal3 44324 31976 44324 31976 0 _0741_
rlabel metal3 39900 14504 39900 14504 0 _0742_
rlabel metal2 19208 16800 19208 16800 0 _0743_
rlabel metal2 22008 18368 22008 18368 0 _0744_
rlabel metal2 25928 14784 25928 14784 0 _0745_
rlabel metal2 19656 19432 19656 19432 0 _0746_
rlabel metal2 19320 19244 19320 19244 0 _0747_
rlabel metal2 19432 17276 19432 17276 0 _0748_
rlabel metal2 26712 13776 26712 13776 0 _0749_
rlabel metal2 26824 13580 26824 13580 0 _0750_
rlabel metal2 39704 14364 39704 14364 0 _0751_
rlabel metal2 23408 12236 23408 12236 0 _0752_
rlabel metal2 29512 14280 29512 14280 0 _0753_
rlabel metal2 29624 14280 29624 14280 0 _0754_
rlabel metal2 38920 13972 38920 13972 0 _0755_
rlabel metal2 40992 14364 40992 14364 0 _0756_
rlabel metal3 25704 14504 25704 14504 0 _0757_
rlabel metal2 37968 14420 37968 14420 0 _0758_
rlabel metal2 34720 16716 34720 16716 0 _0759_
rlabel metal3 31472 16296 31472 16296 0 _0760_
rlabel metal2 36904 14028 36904 14028 0 _0761_
rlabel metal2 36064 13804 36064 13804 0 _0762_
rlabel metal2 32368 12488 32368 12488 0 _0763_
rlabel metal2 22400 15624 22400 15624 0 _0764_
rlabel metal2 22904 12992 22904 12992 0 _0765_
rlabel metal2 25984 13272 25984 13272 0 _0766_
rlabel metal3 32844 12936 32844 12936 0 _0767_
rlabel metal2 24976 20692 24976 20692 0 _0768_
rlabel metal2 20608 16296 20608 16296 0 _0769_
rlabel metal2 23576 12096 23576 12096 0 _0770_
rlabel metal3 28448 12936 28448 12936 0 _0771_
rlabel metal2 21392 15736 21392 15736 0 _0772_
rlabel metal2 22568 20132 22568 20132 0 _0773_
rlabel metal2 22120 17556 22120 17556 0 _0774_
rlabel metal2 16968 17136 16968 17136 0 _0775_
rlabel metal2 20104 17696 20104 17696 0 _0776_
rlabel metal2 22456 17080 22456 17080 0 _0777_
rlabel metal2 22568 16884 22568 16884 0 _0778_
rlabel metal2 30800 7532 30800 7532 0 _0779_
rlabel metal2 32844 9016 32844 9016 0 _0780_
rlabel metal2 20440 18984 20440 18984 0 _0781_
rlabel metal2 22008 17080 22008 17080 0 _0782_
rlabel metal2 33208 5488 33208 5488 0 _0783_
rlabel metal2 31864 9016 31864 9016 0 _0784_
rlabel metal2 32396 6104 32396 6104 0 _0785_
rlabel metal2 31360 7392 31360 7392 0 _0786_
rlabel metal2 32704 5600 32704 5600 0 _0787_
rlabel metal3 30659 12152 30659 12152 0 _0788_
rlabel metal3 32284 5880 32284 5880 0 _0789_
rlabel metal2 32060 4312 32060 4312 0 _0790_
rlabel metal2 31192 4536 31192 4536 0 _0791_
rlabel metal2 32172 10584 32172 10584 0 _0792_
rlabel metal2 30016 10108 30016 10108 0 _0793_
rlabel metal2 30492 11592 30492 11592 0 _0794_
rlabel metal2 31528 12208 31528 12208 0 _0795_
rlabel metal2 20496 8568 20496 8568 0 _0796_
rlabel metal2 19544 14000 19544 14000 0 _0797_
rlabel metal2 19432 13804 19432 13804 0 _0798_
rlabel via2 20104 9781 20104 9781 0 _0799_
rlabel metal3 21224 12936 21224 12936 0 _0800_
rlabel metal2 20832 9996 20832 9996 0 _0801_
rlabel metal2 19180 10808 19180 10808 0 _0802_
rlabel metal2 19712 12292 19712 12292 0 _0803_
rlabel metal2 18732 9240 18732 9240 0 _0804_
rlabel metal2 21672 12544 21672 12544 0 _0805_
rlabel metal2 19600 10164 19600 10164 0 _0806_
rlabel metal2 21336 11480 21336 11480 0 _0807_
rlabel metal2 22456 14224 22456 14224 0 _0808_
rlabel metal2 22176 11676 22176 11676 0 _0809_
rlabel metal2 13944 12236 13944 12236 0 _0810_
rlabel metal2 21728 13328 21728 13328 0 _0811_
rlabel metal2 14280 14364 14280 14364 0 _0812_
rlabel metal2 20524 13496 20524 13496 0 _0813_
rlabel metal2 19096 20552 19096 20552 0 _0814_
rlabel metal2 18312 21784 18312 21784 0 _0815_
rlabel metal2 18872 19488 18872 19488 0 _0816_
rlabel metal2 18088 20496 18088 20496 0 _0817_
rlabel metal3 18760 25480 18760 25480 0 _0818_
rlabel metal3 18200 20776 18200 20776 0 _0819_
rlabel metal2 18676 21672 18676 21672 0 _0820_
rlabel metal2 19880 25536 19880 25536 0 _0821_
rlabel metal2 17808 22428 17808 22428 0 _0822_
rlabel metal2 18396 22568 18396 22568 0 _0823_
rlabel metal2 17864 24640 17864 24640 0 _0824_
rlabel metal2 17808 20468 17808 20468 0 _0825_
rlabel metal2 18368 21168 18368 21168 0 _0826_
rlabel metal3 17472 26264 17472 26264 0 _0827_
rlabel metal2 22792 22960 22792 22960 0 _0828_
rlabel metal2 19460 21000 19460 21000 0 _0829_
rlabel metal3 18480 23128 18480 23128 0 _0830_
rlabel metal2 23128 20832 23128 20832 0 _0831_
rlabel metal2 22120 20300 22120 20300 0 _0832_
rlabel metal3 21728 21560 21728 21560 0 _0833_
rlabel metal2 22680 18275 22680 18275 0 _0834_
rlabel metal2 25704 21056 25704 21056 0 _0835_
rlabel metal2 24920 22232 24920 22232 0 _0836_
rlabel metal2 25850 21803 25850 21803 0 _0837_
rlabel metal2 26264 22064 26264 22064 0 _0838_
rlabel metal2 23406 22624 23406 22624 0 _0839_
rlabel metal2 24136 22848 24136 22848 0 _0840_
rlabel metal2 26114 20291 26114 20291 0 _0841_
rlabel metal2 26824 19936 26824 19936 0 _0842_
rlabel metal2 22541 22344 22541 22344 0 _0843_
rlabel via1 22494 23146 22494 23146 0 _0844_
rlabel metal2 22120 23856 22120 23856 0 _0845_
rlabel metal2 15904 19096 15904 19096 0 _0846_
rlabel metal2 14728 19376 14728 19376 0 _0847_
rlabel metal2 15736 19152 15736 19152 0 _0848_
rlabel metal2 15736 20048 15736 20048 0 _0849_
rlabel metal2 15624 19404 15624 19404 0 _0850_
rlabel metal2 15288 19712 15288 19712 0 _0851_
rlabel via1 6518 20010 6518 20010 0 _0852_
rlabel metal2 2184 19880 2184 19880 0 _0853_
rlabel metal3 13020 19096 13020 19096 0 _0854_
rlabel metal2 5880 21280 5880 21280 0 _0855_
rlabel metal3 11788 20104 11788 20104 0 _0856_
rlabel metal3 8792 21448 8792 21448 0 _0857_
rlabel metal2 15456 19544 15456 19544 0 _0858_
rlabel metal3 8008 19992 8008 19992 0 _0859_
rlabel metal2 21672 19936 21672 19936 0 _0860_
rlabel metal2 20664 19404 20664 19404 0 _0861_
rlabel metal2 21896 20384 21896 20384 0 _0862_
rlabel metal2 15848 22288 15848 22288 0 _0863_
rlabel metal2 15214 21635 15214 21635 0 _0864_
rlabel metal2 14840 21616 14840 21616 0 _0865_
rlabel metal3 14644 22344 14644 22344 0 _0866_
rlabel metal2 10136 23240 10136 23240 0 _0867_
rlabel metal3 14532 20776 14532 20776 0 _0868_
rlabel metal2 9352 20048 9352 20048 0 _0869_
rlabel via1 16465 23128 16465 23128 0 _0870_
rlabel metal2 16016 23016 16016 23016 0 _0871_
rlabel metal3 47936 21560 47936 21560 0 _0872_
rlabel metal2 47292 21672 47292 21672 0 _0873_
rlabel metal2 46536 21784 46536 21784 0 _0874_
rlabel metal2 46312 23184 46312 23184 0 _0875_
rlabel metal2 45304 23632 45304 23632 0 _0876_
rlabel metal2 45864 24234 45864 24234 0 _0877_
rlabel metal2 46200 23744 46200 23744 0 _0878_
rlabel metal2 46312 25004 46312 25004 0 _0879_
rlabel metal2 45640 25928 45640 25928 0 _0880_
rlabel metal2 46816 26040 46816 26040 0 _0881_
rlabel metal2 43736 25704 43736 25704 0 _0882_
rlabel metal2 46292 27608 46292 27608 0 _0883_
rlabel metal3 45500 25704 45500 25704 0 _0884_
rlabel metal2 46032 26488 46032 26488 0 _0885_
rlabel metal2 45164 27272 45164 27272 0 _0886_
rlabel metal2 46536 28168 46536 28168 0 _0887_
rlabel metal2 46620 29400 46620 29400 0 _0888_
rlabel metal2 23408 18172 23408 18172 0 _0889_
rlabel metal2 22568 15288 22568 15288 0 _0890_
rlabel metal2 18536 15560 18536 15560 0 _0891_
rlabel metal2 28028 15400 28028 15400 0 _0892_
rlabel metal2 28924 16968 28924 16968 0 _0893_
rlabel metal2 26096 18032 26096 18032 0 _0894_
rlabel metal2 13944 16520 13944 16520 0 _0895_
rlabel metal3 24864 23240 24864 23240 0 _0896_
rlabel metal2 26824 22960 26824 22960 0 _0897_
rlabel metal2 25816 24836 25816 24836 0 _0898_
rlabel metal3 26852 23912 26852 23912 0 _0899_
rlabel metal3 25648 24696 25648 24696 0 _0900_
rlabel metal2 26376 25368 26376 25368 0 _0901_
rlabel metal2 28504 28504 28504 28504 0 _0902_
rlabel metal3 26320 24808 26320 24808 0 _0903_
rlabel metal2 32312 19936 32312 19936 0 _0904_
rlabel metal2 30520 25396 30520 25396 0 _0905_
rlabel metal3 27496 26264 27496 26264 0 _0906_
rlabel metal2 29512 23604 29512 23604 0 _0907_
rlabel metal2 29344 23128 29344 23128 0 _0908_
rlabel metal2 29792 25256 29792 25256 0 _0909_
rlabel via2 29288 27034 29288 27034 0 _0910_
rlabel metal2 30240 25368 30240 25368 0 _0911_
rlabel metal2 29176 26516 29176 26516 0 _0912_
rlabel metal2 23352 24416 23352 24416 0 _0913_
rlabel metal2 29288 32928 29288 32928 0 _0914_
rlabel metal2 16744 25424 16744 25424 0 _0915_
rlabel metal2 21224 26264 21224 26264 0 _0916_
rlabel metal2 21224 26488 21224 26488 0 _0917_
rlabel via1 20496 35686 20496 35686 0 _0918_
rlabel metal3 18928 25816 18928 25816 0 _0919_
rlabel metal2 18312 28644 18312 28644 0 _0920_
rlabel metal2 18312 31102 18312 31102 0 _0921_
rlabel metal2 20776 34524 20776 34524 0 _0922_
rlabel metal3 20636 28616 20636 28616 0 _0923_
rlabel metal2 19880 29512 19880 29512 0 _0924_
rlabel metal3 20048 32536 20048 32536 0 _0925_
rlabel metal2 18872 28840 18872 28840 0 _0926_
rlabel metal2 20440 31024 20440 31024 0 _0927_
rlabel metal2 21448 28672 21448 28672 0 _0928_
rlabel metal2 19404 29512 19404 29512 0 _0929_
rlabel metal2 19432 32844 19432 32844 0 _0930_
rlabel metal2 21224 32704 21224 32704 0 _0931_
rlabel metal3 31360 32648 31360 32648 0 _0932_
rlabel metal3 30744 34048 30744 34048 0 _0933_
rlabel metal2 13608 21280 13608 21280 0 _0934_
rlabel metal2 13328 20776 13328 20776 0 _0935_
rlabel metal2 13440 15932 13440 15932 0 _0936_
rlabel metal2 13272 27440 13272 27440 0 _0937_
rlabel metal2 15624 28448 15624 28448 0 _0938_
rlabel metal2 11816 24808 11816 24808 0 _0939_
rlabel metal2 12600 22596 12600 22596 0 _0940_
rlabel metal2 15176 25648 15176 25648 0 _0941_
rlabel metal2 12600 24808 12600 24808 0 _0942_
rlabel metal2 12544 25424 12544 25424 0 _0943_
rlabel metal2 10808 24920 10808 24920 0 _0944_
rlabel metal2 11144 23632 11144 23632 0 _0945_
rlabel metal3 12712 25368 12712 25368 0 _0946_
rlabel metal2 13590 25760 13590 25760 0 _0947_
rlabel metal3 13048 31976 13048 31976 0 _0948_
rlabel metal2 2856 22400 2856 22400 0 _0949_
rlabel metal2 2408 24696 2408 24696 0 _0950_
rlabel metal2 3192 25396 3192 25396 0 _0951_
rlabel metal2 3192 24752 3192 24752 0 _0952_
rlabel metal2 2408 25312 2408 25312 0 _0953_
rlabel metal2 5992 25991 5992 25991 0 _0954_
rlabel metal2 6552 23184 6552 23184 0 _0955_
rlabel metal3 6608 25480 6608 25480 0 _0956_
rlabel metal2 5880 26264 5880 26264 0 _0957_
rlabel metal2 6664 23324 6664 23324 0 _0958_
rlabel metal2 4536 22260 4536 22260 0 _0959_
rlabel metal2 9464 24640 9464 24640 0 _0960_
rlabel metal2 7560 25592 7560 25592 0 _0961_
rlabel metal2 6888 26236 6888 26236 0 _0962_
rlabel metal2 14392 32620 14392 32620 0 _0963_
rlabel metal2 11480 25844 11480 25844 0 _0964_
rlabel metal2 10584 27737 10584 27737 0 _0965_
rlabel metal2 14314 26058 14314 26058 0 _0966_
rlabel metal2 11256 27916 11256 27916 0 _0967_
rlabel metal2 11368 28714 11368 28714 0 _0968_
rlabel metal2 10276 26488 10276 26488 0 _0969_
rlabel metal2 9016 28448 9016 28448 0 _0970_
rlabel metal2 8848 30016 8848 30016 0 _0971_
rlabel metal3 4088 22904 4088 22904 0 _0972_
rlabel metal2 4312 19712 4312 19712 0 _0973_
rlabel metal2 4872 23940 4872 23940 0 _0974_
rlabel metal2 4592 23828 4592 23828 0 _0975_
rlabel metal3 5040 24024 5040 24024 0 _0976_
rlabel metal3 8792 26264 8792 26264 0 _0977_
rlabel metal2 7000 24724 7000 24724 0 _0978_
rlabel metal2 5544 29120 5544 29120 0 _0979_
rlabel metal2 4760 22176 4760 22176 0 _0980_
rlabel metal2 7224 22848 7224 22848 0 _0981_
rlabel metal2 6832 24920 6832 24920 0 _0982_
rlabel metal2 4872 25956 4872 25956 0 _0983_
rlabel metal2 5768 27664 5768 27664 0 _0984_
rlabel metal2 12488 27132 12488 27132 0 _0985_
rlabel metal2 14168 26488 14168 26488 0 _0986_
rlabel metal3 10752 27160 10752 27160 0 _0987_
rlabel metal2 9352 27496 9352 27496 0 _0988_
rlabel metal2 9464 29400 9464 29400 0 _0989_
rlabel metal3 12152 30968 12152 30968 0 _0990_
rlabel metal2 15176 33152 15176 33152 0 _0991_
rlabel metal2 2072 23576 2072 23576 0 _0992_
rlabel metal2 3752 26320 3752 26320 0 _0993_
rlabel metal2 6104 23240 6104 23240 0 _0994_
rlabel metal2 4984 24192 4984 24192 0 _0995_
rlabel via1 4097 26376 4097 26376 0 _0996_
rlabel metal2 6160 31752 6160 31752 0 _0997_
rlabel metal2 15008 27328 15008 27328 0 _0998_
rlabel metal2 15568 24920 15568 24920 0 _0999_
rlabel metal3 14784 29400 14784 29400 0 _1000_
rlabel metal2 15512 28672 15512 28672 0 _1001_
rlabel metal2 14840 27608 14840 27608 0 _1002_
rlabel via1 14778 29412 14778 29412 0 _1003_
rlabel metal2 15176 30968 15176 30968 0 _1004_
rlabel metal2 15060 33469 15060 33469 0 _1005_
rlabel via2 13832 33301 13832 33301 0 _1006_
rlabel metal2 15848 33516 15848 33516 0 _1007_
rlabel metal2 31192 33600 31192 33600 0 _1008_
rlabel metal3 32480 34104 32480 34104 0 _1009_
rlabel metal2 21336 31696 21336 31696 0 _1010_
rlabel metal3 19852 30856 19852 30856 0 _1011_
rlabel metal2 21560 33600 21560 33600 0 _1012_
rlabel metal2 18648 26572 18648 26572 0 _1013_
rlabel metal2 20384 26264 20384 26264 0 _1014_
rlabel metal2 21896 30100 21896 30100 0 _1015_
rlabel metal2 20664 40768 20664 40768 0 _1016_
rlabel metal2 21614 31388 21614 31388 0 _1017_
rlabel metal2 25144 31528 25144 31528 0 _1018_
rlabel metal2 24808 31612 24808 31612 0 _1019_
rlabel metal2 25312 24556 25312 24556 0 _1020_
rlabel metal2 28504 24388 28504 24388 0 _1021_
rlabel metal2 29288 25004 29288 25004 0 _1022_
rlabel metal2 26600 26572 26600 26572 0 _1023_
rlabel metal2 24808 23296 24808 23296 0 _1024_
rlabel metal2 28056 25676 28056 25676 0 _1025_
rlabel via1 30912 24713 30912 24713 0 _1026_
rlabel metal2 31136 24780 31136 24780 0 _1027_
rlabel metal2 30856 25704 30856 25704 0 _1028_
rlabel metal2 10920 30548 10920 30548 0 _1029_
rlabel metal2 10808 31332 10808 31332 0 _1030_
rlabel metal2 14616 30464 14616 30464 0 _1031_
rlabel metal2 15288 30576 15288 30576 0 _1032_
rlabel metal2 31976 34356 31976 34356 0 _1033_
rlabel metal3 30072 30968 30072 30968 0 _1034_
rlabel metal2 32068 30912 32068 30912 0 _1035_
rlabel metal3 32704 30968 32704 30968 0 _1036_
rlabel metal3 20440 26936 20440 26936 0 _1037_
rlabel metal3 23268 28616 23268 28616 0 _1038_
rlabel metal2 23688 28308 23688 28308 0 _1039_
rlabel metal2 23128 27090 23128 27090 0 _1040_
rlabel metal2 23016 28672 23016 28672 0 _1041_
rlabel via2 26040 27839 26040 27839 0 _1042_
rlabel metal2 28112 25480 28112 25480 0 _1043_
rlabel metal2 25368 26460 25368 26460 0 _1044_
rlabel metal2 27552 27552 27552 27552 0 _1045_
rlabel metal2 30968 27776 30968 27776 0 _1046_
rlabel metal3 32480 24696 32480 24696 0 _1047_
rlabel metal2 30184 29624 30184 29624 0 _1048_
rlabel metal2 10294 28840 10294 28840 0 _1049_
rlabel metal3 21000 29624 21000 29624 0 _1050_
rlabel metal2 23436 27272 23436 27272 0 _1051_
rlabel metal2 31732 29596 31732 29596 0 _1052_
rlabel metal2 30968 31052 30968 31052 0 _1053_
rlabel metal2 30632 30268 30632 30268 0 _1054_
rlabel metal2 22456 28728 22456 28728 0 _1055_
rlabel metal2 22680 29344 22680 29344 0 _1056_
rlabel metal2 21224 34188 21224 34188 0 _1057_
rlabel metal3 22036 29400 22036 29400 0 _1058_
rlabel metal2 23240 29120 23240 29120 0 _1059_
rlabel metal2 29624 28392 29624 28392 0 _1060_
rlabel metal2 25480 28448 25480 28448 0 _1061_
rlabel metal2 28840 27888 28840 27888 0 _1062_
rlabel metal2 29288 28168 29288 28168 0 _1063_
rlabel metal2 33264 22344 33264 22344 0 _1064_
rlabel metal2 5880 29478 5880 29478 0 _1065_
rlabel metal3 9482 28616 9482 28616 0 _1066_
rlabel metal3 21224 26488 21224 26488 0 _1067_
rlabel metal2 34644 29176 34644 29176 0 _1068_
rlabel metal3 32872 29400 32872 29400 0 _1069_
rlabel metal2 32424 30220 32424 30220 0 _1070_
rlabel metal2 33096 32928 33096 32928 0 _1071_
rlabel metal3 33432 35672 33432 35672 0 _1072_
rlabel metal2 21840 27720 21840 27720 0 _1073_
rlabel metal2 23800 33320 23800 33320 0 _1074_
rlabel metal2 29596 25704 29596 25704 0 _1075_
rlabel via3 28158 31752 28158 31752 0 _1076_
rlabel metal3 28784 34216 28784 34216 0 _1077_
rlabel metal2 7952 22932 7952 22932 0 _1078_
rlabel metal2 5992 23212 5992 23212 0 _1079_
rlabel metal2 8540 23240 8540 23240 0 _1080_
rlabel metal2 10920 27916 10920 27916 0 _1081_
rlabel metal2 15176 28112 15176 28112 0 _1082_
rlabel metal2 12040 34804 12040 34804 0 _1083_
rlabel metal2 5936 36120 5936 36120 0 _1084_
rlabel metal3 11704 36456 11704 36456 0 _1085_
rlabel metal2 14112 33796 14112 33796 0 _1086_
rlabel metal2 14672 34272 14672 34272 0 _1087_
rlabel metal3 18088 35112 18088 35112 0 _1088_
rlabel metal2 30744 35728 30744 35728 0 _1089_
rlabel metal2 29960 33880 29960 33880 0 _1090_
rlabel metal2 32004 33208 32004 33208 0 _1091_
rlabel metal2 29680 33824 29680 33824 0 _1092_
rlabel metal2 31620 35504 31620 35504 0 _1093_
rlabel metal3 32648 36456 32648 36456 0 _1094_
rlabel metal2 34328 36596 34328 36596 0 _1095_
rlabel metal2 35560 36288 35560 36288 0 _1096_
rlabel metal2 35028 37352 35028 37352 0 _1097_
rlabel metal2 33432 35924 33432 35924 0 _1098_
rlabel metal3 32452 36568 32452 36568 0 _1099_
rlabel metal2 26516 27272 26516 27272 0 _1100_
rlabel metal2 26264 35616 26264 35616 0 _1101_
rlabel metal2 20440 40768 20440 40768 0 _1102_
rlabel metal2 19777 34832 19777 34832 0 _1103_
rlabel metal2 19656 35280 19656 35280 0 _1104_
rlabel metal2 29064 36120 29064 36120 0 _1105_
rlabel metal2 9240 24780 9240 24780 0 _1106_
rlabel metal2 9968 25116 9968 25116 0 _1107_
rlabel metal2 10360 25872 10360 25872 0 _1108_
rlabel metal2 11760 26432 11760 26432 0 _1109_
rlabel metal3 14448 26824 14448 26824 0 _1110_
rlabel metal2 11908 35392 11908 35392 0 _1111_
rlabel metal3 12376 35672 12376 35672 0 _1112_
rlabel metal2 12544 35140 12544 35140 0 _1113_
rlabel metal2 12376 34300 12376 34300 0 _1114_
rlabel metal2 12824 35168 12824 35168 0 _1115_
rlabel metal3 21112 35672 21112 35672 0 _1116_
rlabel metal2 31528 36553 31528 36553 0 _1117_
rlabel metal2 28168 33068 28168 33068 0 _1118_
rlabel metal2 31752 35924 31752 35924 0 _1119_
rlabel metal3 33086 37240 33086 37240 0 _1120_
rlabel metal3 34776 37240 34776 37240 0 _1121_
rlabel metal2 32368 38752 32368 38752 0 _1122_
rlabel metal3 32928 38808 32928 38808 0 _1123_
rlabel metal2 21392 33460 21392 33460 0 _1124_
rlabel metal2 21896 34160 21896 34160 0 _1125_
rlabel metal2 21540 37380 21540 37380 0 _1126_
rlabel metal2 28504 26488 28504 26488 0 _1127_
rlabel metal2 26824 35672 26824 35672 0 _1128_
rlabel metal3 28784 37352 28784 37352 0 _1129_
rlabel metal2 8288 25172 8288 25172 0 _1130_
rlabel metal3 8876 24696 8876 24696 0 _1131_
rlabel metal3 8344 24808 8344 24808 0 _1132_
rlabel metal2 8820 25704 8820 25704 0 _1133_
rlabel metal2 15400 28336 15400 28336 0 _1134_
rlabel metal2 14616 27384 14616 27384 0 _1135_
rlabel metal2 11900 39368 11900 39368 0 _1136_
rlabel metal2 14280 37632 14280 37632 0 _1137_
rlabel metal3 12936 39592 12936 39592 0 _1138_
rlabel metal2 14616 38108 14616 38108 0 _1139_
rlabel metal2 13608 36932 13608 36932 0 _1140_
rlabel metal2 11312 39144 11312 39144 0 _1141_
rlabel metal2 12040 37023 12040 37023 0 _1142_
rlabel metal3 13216 37240 13216 37240 0 _1143_
rlabel metal2 12376 37184 12376 37184 0 _1144_
rlabel metal2 15828 38304 15828 38304 0 _1145_
rlabel via2 28056 38009 28056 38009 0 _1146_
rlabel metal3 31472 38024 31472 38024 0 _1147_
rlabel metal2 31780 38808 31780 38808 0 _1148_
rlabel metal2 31920 38696 31920 38696 0 _1149_
rlabel metal2 34216 38416 34216 38416 0 _1150_
rlabel via2 21000 34118 21000 34118 0 _1151_
rlabel metal2 22212 39284 22212 39284 0 _1152_
rlabel via2 25256 26281 25256 26281 0 _1153_
rlabel metal2 25592 26348 25592 26348 0 _1154_
rlabel metal2 25592 27888 25592 27888 0 _1155_
rlabel metal3 28224 39592 28224 39592 0 _1156_
rlabel metal2 28168 39536 28168 39536 0 _1157_
rlabel metal2 7560 26404 7560 26404 0 _1158_
rlabel metal2 8344 26544 8344 26544 0 _1159_
rlabel metal2 13160 40544 13160 40544 0 _1160_
rlabel metal2 12152 39928 12152 39928 0 _1161_
rlabel metal2 13272 39508 13272 39508 0 _1162_
rlabel metal3 13944 38808 13944 38808 0 _1163_
rlabel metal2 15120 38696 15120 38696 0 _1164_
rlabel metal2 15156 39340 15156 39340 0 _1165_
rlabel metal2 15400 39424 15400 39424 0 _1166_
rlabel metal3 29848 38808 29848 38808 0 _1167_
rlabel metal2 26488 37199 26488 37199 0 _1168_
rlabel metal2 29960 38752 29960 38752 0 _1169_
rlabel metal3 31248 39592 31248 39592 0 _1170_
rlabel metal2 32284 38248 32284 38248 0 _1171_
rlabel metal2 31808 39508 31808 39508 0 _1172_
rlabel metal2 37184 39676 37184 39676 0 _1173_
rlabel metal3 35476 39592 35476 39592 0 _1174_
rlabel metal2 36568 39984 36568 39984 0 _1175_
rlabel metal2 30744 39004 30744 39004 0 _1176_
rlabel metal2 31416 40096 31416 40096 0 _1177_
rlabel via1 21662 41944 21662 41944 0 _1178_
rlabel metal2 26132 41888 26132 41888 0 _1179_
rlabel metal2 27776 40376 27776 40376 0 _1180_
rlabel metal2 12852 37352 12852 37352 0 _1181_
rlabel metal2 12600 38892 12600 38892 0 _1182_
rlabel metal2 13608 40432 13608 40432 0 _1183_
rlabel metal2 3052 44968 3052 44968 0 _1184_
rlabel metal2 15828 40964 15828 40964 0 _1185_
rlabel metal2 14484 40572 14484 40572 0 _1186_
rlabel metal3 18088 40880 18088 40880 0 _1187_
rlabel metal2 30184 40460 30184 40460 0 _1188_
rlabel metal2 26068 26376 26068 26376 0 _1189_
rlabel metal2 29176 40992 29176 40992 0 _1190_
rlabel metal3 29176 41944 29176 41944 0 _1191_
rlabel metal2 29624 41468 29624 41468 0 _1192_
rlabel metal3 31630 41160 31630 41160 0 _1193_
rlabel metal4 36904 39312 36904 39312 0 _1194_
rlabel via2 30520 40391 30520 40391 0 _1195_
rlabel metal2 30912 40488 30912 40488 0 _1196_
rlabel metal2 22344 42840 22344 42840 0 _1197_
rlabel metal3 22764 42504 22764 42504 0 _1198_
rlabel metal2 26824 42784 26824 42784 0 _1199_
rlabel metal2 27272 42728 27272 42728 0 _1200_
rlabel metal3 9912 25536 9912 25536 0 _1201_
rlabel via1 11918 43512 11918 43512 0 _1202_
rlabel metal2 12376 43512 12376 43512 0 _1203_
rlabel metal2 14504 42467 14504 42467 0 _1204_
rlabel metal2 13720 43232 13720 43232 0 _1205_
rlabel metal3 29960 42952 29960 42952 0 _1206_
rlabel metal2 21560 41364 21560 41364 0 _1207_
rlabel metal2 30836 42476 30836 42476 0 _1208_
rlabel metal2 31844 42140 31844 42140 0 _1209_
rlabel metal2 43736 42644 43736 42644 0 _1210_
rlabel metal3 31668 42952 31668 42952 0 _1211_
rlabel metal3 30744 43512 30744 43512 0 _1212_
rlabel via2 28280 43527 28280 43527 0 _1213_
rlabel metal2 31752 43064 31752 43064 0 _1214_
rlabel metal2 10584 43176 10584 43176 0 _1215_
rlabel via2 12600 42720 12600 42720 0 _1216_
rlabel metal3 21112 43456 21112 43456 0 _1217_
rlabel metal2 29960 43568 29960 43568 0 _1218_
rlabel metal2 32010 43418 32010 43418 0 _1219_
rlabel metal3 31724 43400 31724 43400 0 _1220_
rlabel metal2 34440 43400 34440 43400 0 _1221_
rlabel metal2 45248 22904 45248 22904 0 _1222_
rlabel metal2 39704 23576 39704 23576 0 _1223_
rlabel metal2 39032 24024 39032 24024 0 _1224_
rlabel metal3 44912 39928 44912 39928 0 _1225_
rlabel metal2 43792 37240 43792 37240 0 _1226_
rlabel metal2 42280 36554 42280 36554 0 _1227_
rlabel metal2 44744 30912 44744 30912 0 _1228_
rlabel metal3 43596 34888 43596 34888 0 _1229_
rlabel metal2 38360 22176 38360 22176 0 _1230_
rlabel metal2 38864 26824 38864 26824 0 _1231_
rlabel metal3 44464 33320 44464 33320 0 _1232_
rlabel metal2 47040 30184 47040 30184 0 _1233_
rlabel metal3 47264 35560 47264 35560 0 _1234_
rlabel metal2 47320 35280 47320 35280 0 _1235_
rlabel metal2 45304 37464 45304 37464 0 _1236_
rlabel metal2 46872 34061 46872 34061 0 _1237_
rlabel metal2 46536 34440 46536 34440 0 _1238_
rlabel metal3 45976 39144 45976 39144 0 _1239_
rlabel metal2 46536 30400 46536 30400 0 _1240_
rlabel metal2 47544 30736 47544 30736 0 _1241_
rlabel metal2 24752 19292 24752 19292 0 _1242_
rlabel metal2 20048 18424 20048 18424 0 _1243_
rlabel metal2 18536 19152 18536 19152 0 _1244_
rlabel metal2 24612 18200 24612 18200 0 _1245_
rlabel metal2 26040 9296 26040 9296 0 _1246_
rlabel metal2 25592 18816 25592 18816 0 _1247_
rlabel metal2 23800 19040 23800 19040 0 _1248_
rlabel metal2 26824 17864 26824 17864 0 _1249_
rlabel metal2 26600 15736 26600 15736 0 _1250_
rlabel metal2 25368 7616 25368 7616 0 _1251_
rlabel metal2 25536 21560 25536 21560 0 _1252_
rlabel metal2 26712 11032 26712 11032 0 _1253_
rlabel metal2 17864 19880 17864 19880 0 _1254_
rlabel metal2 20440 22848 20440 22848 0 _1255_
rlabel metal3 16520 22344 16520 22344 0 _1256_
rlabel metal2 25514 7747 25514 7747 0 _1257_
rlabel metal3 25032 7448 25032 7448 0 _1258_
rlabel metal2 24304 6580 24304 6580 0 _1259_
rlabel metal2 23744 17192 23744 17192 0 _1260_
rlabel metal2 24024 12432 24024 12432 0 _1261_
rlabel metal2 22568 9856 22568 9856 0 _1262_
rlabel metal2 26040 12488 26040 12488 0 _1263_
rlabel metal2 16632 15792 16632 15792 0 _1264_
rlabel metal2 22680 14224 22680 14224 0 _1265_
rlabel metal2 22624 15988 22624 15988 0 _1266_
rlabel metal2 23968 6972 23968 6972 0 _1267_
rlabel metal2 21476 5320 21476 5320 0 _1268_
rlabel metal2 23464 13048 23464 13048 0 _1269_
rlabel metal2 22736 9884 22736 9884 0 _1270_
rlabel metal2 22400 6972 22400 6972 0 _1271_
rlabel metal2 22148 7672 22148 7672 0 _1272_
rlabel metal2 21532 13608 21532 13608 0 _1273_
rlabel metal2 25424 16296 25424 16296 0 _1274_
rlabel metal2 24696 9296 24696 9296 0 _1275_
rlabel metal2 21280 8540 21280 8540 0 _1276_
rlabel metal2 26320 19208 26320 19208 0 _1277_
rlabel metal2 26488 18312 26488 18312 0 _1278_
rlabel metal2 26600 17080 26600 17080 0 _1279_
rlabel metal3 27160 9800 27160 9800 0 _1280_
rlabel via1 27551 9744 27551 9744 0 _1281_
rlabel metal2 28168 9072 28168 9072 0 _1282_
rlabel metal3 28420 6664 28420 6664 0 _1283_
rlabel metal2 27048 9016 27048 9016 0 _1284_
rlabel metal2 27216 6972 27216 6972 0 _1285_
rlabel metal2 27720 5348 27720 5348 0 _1286_
rlabel metal2 26880 5460 26880 5460 0 _1287_
rlabel metal2 27832 3416 27832 3416 0 _1288_
rlabel metal2 26712 5544 26712 5544 0 _1289_
rlabel metal2 24360 17136 24360 17136 0 _1290_
rlabel metal2 25760 17360 25760 17360 0 _1291_
rlabel metal2 28168 17696 28168 17696 0 _1292_
rlabel metal2 33656 17052 33656 17052 0 _1293_
rlabel metal3 25844 15176 25844 15176 0 _1294_
rlabel metal3 31528 17640 31528 17640 0 _1295_
rlabel metal2 35168 18424 35168 18424 0 _1296_
rlabel metal2 36904 15596 36904 15596 0 _1297_
rlabel metal3 30632 15288 30632 15288 0 _1298_
rlabel metal2 29680 15848 29680 15848 0 _1299_
rlabel metal3 34132 15176 34132 15176 0 _1300_
rlabel metal2 33880 16940 33880 16940 0 _1301_
rlabel via3 29708 15176 29708 15176 0 _1302_
rlabel metal2 28560 15932 28560 15932 0 _1303_
rlabel metal3 31920 16072 31920 16072 0 _1304_
rlabel metal2 48272 21336 48272 21336 0 _1305_
rlabel metal2 43960 20642 43960 20642 0 _1306_
rlabel metal2 31752 20818 31752 20818 0 _1307_
rlabel metal2 31472 22708 31472 22708 0 _1308_
rlabel metal3 31136 20776 31136 20776 0 _1309_
rlabel metal2 31640 23296 31640 23296 0 _1310_
rlabel metal2 31752 23688 31752 23688 0 _1311_
rlabel metal3 31696 23800 31696 23800 0 _1312_
rlabel metal2 23744 15288 23744 15288 0 _1313_
rlabel metal2 23408 15176 23408 15176 0 _1314_
rlabel metal2 32564 22314 32564 22314 0 _1315_
rlabel metal2 31360 25032 31360 25032 0 _1316_
rlabel metal2 34440 25704 34440 25704 0 _1317_
rlabel metal2 34776 25685 34776 25685 0 _1318_
rlabel metal2 34804 24808 34804 24808 0 _1319_
rlabel metal2 16408 19432 16408 19432 0 _1320_
rlabel metal2 16744 20216 16744 20216 0 _1321_
rlabel metal2 44380 24920 44380 24920 0 _1322_
rlabel metal2 35896 25368 35896 25368 0 _1323_
rlabel metal2 36540 25480 36540 25480 0 _1324_
rlabel metal2 31808 27048 31808 27048 0 _1325_
rlabel metal2 35224 26992 35224 26992 0 _1326_
rlabel metal2 33992 26628 33992 26628 0 _1327_
rlabel metal3 35420 27048 35420 27048 0 _1328_
rlabel metal2 36008 27160 36008 27160 0 _1329_
rlabel metal2 36288 27552 36288 27552 0 _1330_
rlabel metal3 28728 31752 28728 31752 0 _1331_
rlabel metal2 29288 31696 29288 31696 0 _1332_
rlabel metal3 29316 31976 29316 31976 0 _1333_
rlabel metal2 27832 31248 27832 31248 0 _1334_
rlabel metal2 27048 31808 27048 31808 0 _1335_
rlabel metal2 25704 35463 25704 35463 0 _1336_
rlabel metal2 24584 34776 24584 34776 0 _1337_
rlabel metal2 26824 34748 26824 34748 0 _1338_
rlabel metal2 19488 3332 19488 3332 0 _1339_
rlabel metal3 22624 16296 22624 16296 0 _1340_
rlabel metal2 26292 34104 26292 34104 0 _1341_
rlabel metal2 25928 34384 25928 34384 0 _1342_
rlabel metal2 26376 37464 26376 37464 0 _1343_
rlabel metal2 26152 37087 26152 37087 0 _1344_
rlabel metal2 26600 37856 26600 37856 0 _1345_
rlabel metal3 25284 40600 25284 40600 0 _1346_
rlabel metal2 26712 36904 26712 36904 0 _1347_
rlabel metal2 24248 37576 24248 37576 0 _1348_
rlabel metal2 39592 41888 39592 41888 0 _1349_
rlabel metal3 16464 38808 16464 38808 0 _1350_
rlabel metal2 2968 31808 2968 31808 0 _1351_
rlabel metal2 26488 40320 26488 40320 0 _1352_
rlabel metal2 26712 40264 26712 40264 0 _1353_
rlabel metal3 24752 41272 24752 41272 0 _1354_
rlabel via1 25738 40394 25738 40394 0 _1355_
rlabel metal2 24248 40152 24248 40152 0 _1356_
rlabel metal2 25256 42616 25256 42616 0 _1357_
rlabel metal2 26376 41440 26376 41440 0 _1358_
rlabel metal2 26152 40936 26152 40936 0 _1359_
rlabel metal2 24248 41627 24248 41627 0 _1360_
rlabel metal2 26206 42700 26206 42700 0 _1361_
rlabel metal2 24472 43512 24472 43512 0 _1362_
rlabel metal2 29680 45864 29680 45864 0 _1363_
rlabel metal2 28840 46004 28840 46004 0 _1364_
rlabel metal2 25928 44352 25928 44352 0 _1365_
rlabel metal2 26264 44044 26264 44044 0 _1366_
rlabel metal2 26768 44632 26768 44632 0 _1367_
rlabel metal2 25704 45136 25704 45136 0 _1368_
rlabel metal2 26488 45976 26488 45976 0 _1369_
rlabel metal2 28616 44576 28616 44576 0 _1370_
rlabel metal2 28448 44296 28448 44296 0 _1371_
rlabel metal3 26796 44296 26796 44296 0 _1372_
rlabel metal2 6832 27916 6832 27916 0 _1373_
rlabel metal2 3080 29540 3080 29540 0 _1374_
rlabel metal2 2856 27152 2856 27152 0 _1375_
rlabel metal2 4872 29008 4872 29008 0 _1376_
rlabel metal2 5068 27272 5068 27272 0 _1377_
rlabel metal2 6496 28812 6496 28812 0 _1378_
rlabel metal2 2856 30128 2856 30128 0 _1379_
rlabel metal2 3304 29484 3304 29484 0 _1380_
rlabel metal2 3080 30400 3080 30400 0 _1381_
rlabel metal2 3304 31444 3304 31444 0 _1382_
rlabel metal2 4480 31668 4480 31668 0 _1383_
rlabel metal3 2856 31752 2856 31752 0 _1384_
rlabel metal2 5992 34048 5992 34048 0 _1385_
rlabel metal2 4312 31976 4312 31976 0 _1386_
rlabel metal2 6104 32256 6104 32256 0 _1387_
rlabel metal2 7168 34272 7168 34272 0 _1388_
rlabel metal2 5824 34216 5824 34216 0 _1389_
rlabel metal2 2632 33488 2632 33488 0 _1390_
rlabel metal2 10472 34888 10472 34888 0 _1391_
rlabel metal3 8960 34888 8960 34888 0 _1392_
rlabel via1 6271 32536 6271 32536 0 _1393_
rlabel metal2 7560 34356 7560 34356 0 _1394_
rlabel metal2 8148 35112 8148 35112 0 _1395_
rlabel metal2 7112 35448 7112 35448 0 _1396_
rlabel metal2 7140 36456 7140 36456 0 _1397_
rlabel metal3 10584 39032 10584 39032 0 _1398_
rlabel metal2 9884 39368 9884 39368 0 _1399_
rlabel metal2 10696 37324 10696 37324 0 _1400_
rlabel metal2 38864 24136 38864 24136 0 _1401_
rlabel metal3 10052 36680 10052 36680 0 _1402_
rlabel metal2 9800 37940 9800 37940 0 _1403_
rlabel metal2 2968 39088 2968 39088 0 _1404_
rlabel metal3 5096 39592 5096 39592 0 _1405_
rlabel metal2 5880 39690 5880 39690 0 _1406_
rlabel metal2 4872 40712 4872 40712 0 _1407_
rlabel metal2 2912 40656 2912 40656 0 _1408_
rlabel metal3 5712 39704 5712 39704 0 _1409_
rlabel metal2 2576 38808 2576 38808 0 _1410_
rlabel metal2 4312 42560 4312 42560 0 _1411_
rlabel via1 3640 42720 3640 42720 0 _1412_
rlabel metal2 3640 41846 3640 41846 0 _1413_
rlabel metal2 4704 42560 4704 42560 0 _1414_
rlabel metal2 3416 41076 3416 41076 0 _1415_
rlabel metal2 16632 37744 16632 37744 0 _1416_
rlabel metal2 5488 43512 5488 43512 0 _1417_
rlabel metal2 5992 44408 5992 44408 0 _1418_
rlabel metal2 7112 41804 7112 41804 0 _1419_
rlabel metal2 5712 43008 5712 43008 0 _1420_
rlabel via2 7448 43531 7448 43531 0 _1421_
rlabel metal2 7224 43456 7224 43456 0 _1422_
rlabel metal2 4424 43568 4424 43568 0 _1423_
rlabel metal2 10024 44618 10024 44618 0 _1424_
rlabel metal2 9940 43400 9940 43400 0 _1425_
rlabel metal2 8568 43624 8568 43624 0 _1426_
rlabel metal2 7896 43736 7896 43736 0 _1427_
rlabel metal2 7476 44296 7476 44296 0 _1428_
rlabel metal2 8176 43624 8176 43624 0 _1429_
rlabel metal2 6860 44520 6860 44520 0 _1430_
rlabel metal3 9072 44296 9072 44296 0 _1431_
rlabel metal2 9800 44772 9800 44772 0 _1432_
rlabel metal2 8120 32213 8120 32213 0 _1433_
rlabel metal3 9072 30968 9072 30968 0 _1434_
rlabel metal2 7560 32648 7560 32648 0 _1435_
rlabel metal2 8064 30968 8064 30968 0 _1436_
rlabel metal2 6440 31024 6440 31024 0 _1437_
rlabel metal3 6496 30968 6496 30968 0 _1438_
rlabel metal2 8456 30912 8456 30912 0 _1439_
rlabel metal2 9800 31696 9800 31696 0 _1440_
rlabel metal2 10388 31696 10388 31696 0 _1441_
rlabel metal2 9324 31864 9324 31864 0 _1442_
rlabel metal2 10920 34552 10920 34552 0 _1443_
rlabel metal2 9128 34440 9128 34440 0 _1444_
rlabel metal2 5152 35672 5152 35672 0 _1445_
rlabel via2 40936 16869 40936 16869 0 clknet_0_wb_clk_i
rlabel metal2 3304 7896 3304 7896 0 clknet_4_0_0_wb_clk_i
rlabel metal3 46928 15288 46928 15288 0 clknet_4_10_0_wb_clk_i
rlabel metal2 44744 21560 44744 21560 0 clknet_4_11_0_wb_clk_i
rlabel metal2 25256 44576 25256 44576 0 clknet_4_12_0_wb_clk_i
rlabel metal2 45416 44380 45416 44380 0 clknet_4_13_0_wb_clk_i
rlabel metal2 48244 25592 48244 25592 0 clknet_4_14_0_wb_clk_i
rlabel metal2 23688 39368 23688 39368 0 clknet_4_15_0_wb_clk_i
rlabel metal2 1624 21952 1624 21952 0 clknet_4_1_0_wb_clk_i
rlabel metal2 17696 15288 17696 15288 0 clknet_4_2_0_wb_clk_i
rlabel metal3 22428 23912 22428 23912 0 clknet_4_3_0_wb_clk_i
rlabel metal2 2128 29680 2128 29680 0 clknet_4_4_0_wb_clk_i
rlabel metal2 2100 44072 2100 44072 0 clknet_4_5_0_wb_clk_i
rlabel metal3 20076 25368 20076 25368 0 clknet_4_6_0_wb_clk_i
rlabel metal2 22848 42728 22848 42728 0 clknet_4_7_0_wb_clk_i
rlabel metal2 26656 4312 26656 4312 0 clknet_4_8_0_wb_clk_i
rlabel metal2 25928 22344 25928 22344 0 clknet_4_9_0_wb_clk_i
rlabel metal2 30184 42056 30184 42056 0 custom_settings[0]
rlabel metal2 29736 42952 29736 42952 0 custom_settings[1]
rlabel metal3 39130 2744 39130 2744 0 io_in_1[0]
rlabel metal2 48328 8176 48328 8176 0 io_in_1[1]
rlabel metal2 48328 11256 48328 11256 0 io_in_1[2]
rlabel metal3 48986 17528 48986 17528 0 io_in_1[3]
rlabel metal3 49042 22456 49042 22456 0 io_in_1[4]
rlabel metal3 46648 16184 46648 16184 0 io_in_1[5]
rlabel metal3 46704 29400 46704 29400 0 io_in_1[6]
rlabel metal3 49336 37968 49336 37968 0 io_in_1[7]
rlabel metal2 1988 44968 1988 44968 0 io_in_2
rlabel metal2 19320 47698 19320 47698 0 io_out[10]
rlabel metal2 20888 46914 20888 46914 0 io_out[11]
rlabel metal2 22456 47698 22456 47698 0 io_out[12]
rlabel metal2 30296 47698 30296 47698 0 io_out[17]
rlabel metal2 32312 44800 32312 44800 0 io_out[18]
rlabel metal2 33432 47698 33432 47698 0 io_out[19]
rlabel metal2 35000 47810 35000 47810 0 io_out[20]
rlabel metal2 38024 44912 38024 44912 0 io_out[21]
rlabel metal2 38136 47698 38136 47698 0 io_out[22]
rlabel metal2 39704 46914 39704 46914 0 io_out[23]
rlabel metal2 41272 47306 41272 47306 0 io_out[24]
rlabel metal3 44240 44520 44240 44520 0 io_out[25]
rlabel metal2 44408 47194 44408 47194 0 io_out[26]
rlabel metal2 45976 47418 45976 47418 0 io_out[27]
rlabel metal2 16184 47586 16184 47586 0 io_out[8]
rlabel metal2 17752 47810 17752 47810 0 io_out[9]
rlabel metal2 47208 25424 47208 25424 0 net1
rlabel metal3 1736 42504 1736 42504 0 net10
rlabel metal2 19964 22456 19964 22456 0 net11
rlabel via2 20104 45850 20104 45850 0 net12
rlabel metal2 21336 44562 21336 44562 0 net13
rlabel metal2 21336 45752 21336 45752 0 net14
rlabel metal3 31584 45864 31584 45864 0 net15
rlabel metal2 33320 42504 33320 42504 0 net16
rlabel metal2 34328 40936 34328 40936 0 net17
rlabel metal2 36232 40572 36232 40572 0 net18
rlabel metal2 36680 42028 36680 42028 0 net19
rlabel metal2 40936 42616 40936 42616 0 net2
rlabel metal2 36456 45332 36456 45332 0 net20
rlabel via1 38817 43512 38817 43512 0 net21
rlabel metal2 43512 44444 43512 44444 0 net22
rlabel metal2 23408 40936 23408 40936 0 net23
rlabel metal2 42728 43471 42728 43471 0 net24
rlabel metal2 2800 43176 2800 43176 0 net25
rlabel metal2 12712 44968 12712 44968 0 net26
rlabel metal3 16520 44688 16520 44688 0 net27
rlabel metal2 3920 46004 3920 46004 0 net28
rlabel metal2 5600 45948 5600 45948 0 net29
rlabel metal2 23912 16520 23912 16520 0 net3
rlabel metal2 7056 46004 7056 46004 0 net30
rlabel metal2 8624 45780 8624 45780 0 net31
rlabel metal2 10192 45780 10192 45780 0 net32
rlabel metal2 11424 46004 11424 46004 0 net33
rlabel metal2 13468 44072 13468 44072 0 net34
rlabel metal2 11872 45724 11872 45724 0 net35
rlabel metal2 24304 41076 24304 41076 0 net36
rlabel metal2 25424 46004 25424 46004 0 net37
rlabel metal2 31472 45724 31472 45724 0 net38
rlabel metal2 30016 44436 30016 44436 0 net39
rlabel metal3 27048 11536 27048 11536 0 net4
rlabel metal2 44968 17248 44968 17248 0 net5
rlabel metal3 46760 20328 46760 20328 0 net6
rlabel metal2 47992 27552 47992 27552 0 net7
rlabel metal2 46648 25368 46648 25368 0 net8
rlabel metal2 20300 21784 20300 21784 0 net9
rlabel metal2 1680 26264 1680 26264 0 rst_n
rlabel metal2 34608 41160 34608 41160 0 tt_um_rejunity_sn76489.DAC_clk
rlabel metal4 30408 40992 30408 40992 0 tt_um_rejunity_sn76489.DAC_dat
rlabel metal2 32984 43624 32984 43624 0 tt_um_rejunity_sn76489.DAC_le
rlabel metal2 12488 23128 12488 23128 0 tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[0\]
rlabel metal2 11812 22437 11812 22437 0 tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[1\]
rlabel metal2 12040 20440 12040 20440 0 tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[2\]
rlabel metal2 15176 24360 15176 24360 0 tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[3\]
rlabel metal2 12544 19208 12544 19208 0 tt_um_rejunity_sn76489.chan\[0\].attenuation.in
rlabel metal2 2184 22064 2184 22064 0 tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[0\]
rlabel via1 2628 23893 2628 23893 0 tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[1\]
rlabel metal3 9688 22344 9688 22344 0 tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[2\]
rlabel metal2 6664 19488 6664 19488 0 tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[3\]
rlabel metal2 7784 19208 7784 19208 0 tt_um_rejunity_sn76489.chan\[1\].attenuation.in
rlabel metal2 30028 23781 30028 23781 0 tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[0\]
rlabel metal3 25872 23128 25872 23128 0 tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[1\]
rlabel metal2 28616 20888 28616 20888 0 tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[2\]
rlabel metal2 26148 24005 26148 24005 0 tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[3\]
rlabel metal2 34216 22344 34216 22344 0 tt_um_rejunity_sn76489.chan\[2\].attenuation.in
rlabel metal2 21784 26264 21784 26264 0 tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[0\]
rlabel metal2 18704 26040 18704 26040 0 tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[1\]
rlabel metal2 17976 27496 17976 27496 0 tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[2\]
rlabel metal2 19320 23352 19320 23352 0 tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[3\]
rlabel metal2 18984 26432 18984 26432 0 tt_um_rejunity_sn76489.chan\[3\].attenuation.in
rlabel metal2 45640 21448 45640 21448 0 tt_um_rejunity_sn76489.clk_counter\[0\]
rlabel metal3 45752 21112 45752 21112 0 tt_um_rejunity_sn76489.clk_counter\[1\]
rlabel metal3 47376 22232 47376 22232 0 tt_um_rejunity_sn76489.clk_counter\[2\]
rlabel metal3 46480 24808 46480 24808 0 tt_um_rejunity_sn76489.clk_counter\[3\]
rlabel metal3 46256 25480 46256 25480 0 tt_um_rejunity_sn76489.clk_counter\[4\]
rlabel metal2 46872 27440 46872 27440 0 tt_um_rejunity_sn76489.clk_counter\[5\]
rlabel metal3 45752 27832 45752 27832 0 tt_um_rejunity_sn76489.clk_counter\[6\]
rlabel metal2 32088 20048 32088 20048 0 tt_um_rejunity_sn76489.control_noise\[0\]\[0\]
rlabel metal2 31808 19992 31808 19992 0 tt_um_rejunity_sn76489.control_noise\[0\]\[1\]
rlabel metal3 13664 17640 13664 17640 0 tt_um_rejunity_sn76489.control_noise\[0\]\[2\]
rlabel metal2 25256 7280 25256 7280 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[0\]
rlabel metal2 24528 5992 24528 5992 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[1\]
rlabel metal2 20328 5208 20328 5208 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[2\]
rlabel metal3 20608 7448 20608 7448 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[3\]
rlabel metal2 19320 8848 19320 8848 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[4\]
rlabel metal2 18928 10584 18928 10584 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[5\]
rlabel metal2 16184 8064 16184 8064 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[6\]
rlabel metal2 20552 10920 20552 10920 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[7\]
rlabel metal2 13496 11312 13496 11312 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[8\]
rlabel metal3 14280 14504 14280 14504 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[9\]
rlabel metal2 38920 8344 38920 8344 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[0\]
rlabel metal2 41048 7336 41048 7336 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[1\]
rlabel metal2 42392 6440 42392 6440 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[2\]
rlabel metal2 40712 4872 40712 4872 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[3\]
rlabel metal2 38920 6440 38920 6440 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[4\]
rlabel metal2 39032 5936 39032 5936 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[5\]
rlabel metal2 32536 5152 32536 5152 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[6\]
rlabel metal2 32424 4536 32424 4536 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[7\]
rlabel metal2 32536 10416 32536 10416 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[8\]
rlabel metal3 32564 12040 32564 12040 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[9\]
rlabel metal2 39592 18256 39592 18256 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[0\]
rlabel metal2 41384 17472 41384 17472 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[1\]
rlabel metal2 42504 17528 42504 17528 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[2\]
rlabel metal2 42280 15904 42280 15904 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[3\]
rlabel metal2 40264 15148 40264 15148 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[4\]
rlabel metal3 40768 15960 40768 15960 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[5\]
rlabel metal2 41608 15960 41608 15960 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[6\]
rlabel metal2 42728 13720 42728 13720 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[7\]
rlabel metal2 41048 12656 41048 12656 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[8\]
rlabel metal2 35672 13160 35672 13160 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[9\]
rlabel metal2 8344 32480 8344 32480 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[0\]
rlabel metal3 13328 44296 13328 44296 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[10\]
rlabel metal3 8792 30184 8792 30184 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[1\]
rlabel metal2 11116 31696 11116 31696 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[2\]
rlabel metal2 3416 34720 3416 34720 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[3\]
rlabel metal3 5152 37240 5152 37240 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[4\]
rlabel metal2 7000 39256 7000 39256 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[5\]
rlabel metal2 8232 40992 8232 40992 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[6\]
rlabel metal3 11256 41160 11256 41160 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[7\]
rlabel via2 15624 41160 15624 41160 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[8\]
rlabel metal2 15064 42896 15064 42896 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[9\]
rlabel metal2 4536 27832 4536 27832 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[0\]
rlabel metal2 13104 45192 13104 45192 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[10\]
rlabel metal2 2800 29316 2800 29316 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[1\]
rlabel metal2 4256 30968 4256 30968 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[2\]
rlabel metal2 4312 32536 4312 32536 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[3\]
rlabel metal2 9520 35756 9520 35756 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[4\]
rlabel metal2 11312 39508 11312 39508 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[5\]
rlabel metal2 4312 39760 4312 39760 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[6\]
rlabel metal3 5152 41944 5152 41944 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[7\]
rlabel metal2 4984 43960 4984 43960 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[8\]
rlabel metal2 9520 45080 9520 45080 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[9\]
rlabel metal2 32704 21672 32704 21672 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[0\]
rlabel metal2 24472 45528 24472 45528 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[10\]
rlabel metal3 33236 23576 33236 23576 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[1\]
rlabel metal2 35672 24920 35672 24920 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[2\]
rlabel metal2 35112 26544 35112 26544 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[3\]
rlabel metal2 28000 32424 28000 32424 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[4\]
rlabel metal3 25172 35560 25172 35560 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[5\]
rlabel metal2 25928 36456 25928 36456 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[6\]
rlabel metal2 25480 40040 25480 40040 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[7\]
rlabel metal2 25480 43176 25480 43176 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[8\]
rlabel metal2 29176 44688 29176 44688 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[9\]
rlabel metal3 39760 26264 39760 26264 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[0\]
rlabel metal2 16968 45024 16968 45024 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[10\]
rlabel metal3 24976 30072 24976 30072 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[1\]
rlabel metal2 24696 32872 24696 32872 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[2\]
rlabel metal2 17808 32228 17808 32228 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[3\]
rlabel metal2 17248 34916 17248 34916 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[4\]
rlabel metal2 18816 35756 18816 35756 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[5\]
rlabel metal2 20440 37184 20440 37184 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[6\]
rlabel metal3 20832 40376 20832 40376 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[7\]
rlabel metal2 20664 41944 20664 41944 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[8\]
rlabel metal2 19992 43232 19992 43232 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[9\]
rlabel metal3 18424 17640 18424 17640 0 tt_um_rejunity_sn76489.latch_control_reg\[0\]
rlabel metal2 21280 16072 21280 16072 0 tt_um_rejunity_sn76489.latch_control_reg\[1\]
rlabel metal2 17304 16016 17304 16016 0 tt_um_rejunity_sn76489.latch_control_reg\[2\]
rlabel metal2 43512 21168 43512 21168 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[0\]
rlabel metal2 42168 22736 42168 22736 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[1\]
rlabel metal2 43400 25032 43400 25032 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[2\]
rlabel metal2 41496 23520 41496 23520 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[3\]
rlabel metal2 37464 22008 37464 22008 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[4\]
rlabel metal2 34440 22064 34440 22064 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[5\]
rlabel metal2 33880 19656 33880 19656 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[6\]
rlabel metal2 7168 7448 7168 7448 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[10\]
rlabel metal2 9744 6552 9744 6552 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[11\]
rlabel metal3 8008 8232 8008 8232 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[12\]
rlabel metal2 9240 10584 9240 10584 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[13\]
rlabel metal2 9520 12152 9520 12152 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[14\]
rlabel metal2 12880 16856 12880 16856 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[1\]
rlabel metal2 7672 16408 7672 16408 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[2\]
rlabel metal3 5600 15960 5600 15960 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[3\]
rlabel metal3 5432 14504 5432 14504 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[4\]
rlabel metal2 7224 12600 7224 12600 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[5\]
rlabel metal3 5096 11368 5096 11368 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[6\]
rlabel metal3 5600 9800 5600 9800 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[7\]
rlabel metal3 4256 8232 4256 8232 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[8\]
rlabel metal2 5992 8288 5992 8288 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[9\]
rlabel metal2 15624 16408 15624 16408 0 tt_um_rejunity_sn76489.noise\[0\].gen.restart_noise
rlabel metal2 9072 16856 9072 16856 0 tt_um_rejunity_sn76489.noise\[0\].gen.signal_edge.previous_signal_state_0
rlabel metal2 40600 29064 40600 29064 0 tt_um_rejunity_sn76489.pwm.accumulator\[0\]
rlabel metal2 44520 40880 44520 40880 0 tt_um_rejunity_sn76489.pwm.accumulator\[10\]
rlabel metal2 44184 42392 44184 42392 0 tt_um_rejunity_sn76489.pwm.accumulator\[11\]
rlabel metal2 20720 45864 20720 45864 0 tt_um_rejunity_sn76489.pwm.accumulator\[12\]
rlabel metal2 37464 28616 37464 28616 0 tt_um_rejunity_sn76489.pwm.accumulator\[1\]
rlabel metal2 33208 32760 33208 32760 0 tt_um_rejunity_sn76489.pwm.accumulator\[2\]
rlabel metal2 36176 34888 36176 34888 0 tt_um_rejunity_sn76489.pwm.accumulator\[3\]
rlabel metal3 35280 40376 35280 40376 0 tt_um_rejunity_sn76489.pwm.accumulator\[4\]
rlabel metal2 34776 41832 34776 41832 0 tt_um_rejunity_sn76489.pwm.accumulator\[5\]
rlabel metal2 36288 44940 36288 44940 0 tt_um_rejunity_sn76489.pwm.accumulator\[6\]
rlabel metal2 40320 44968 40320 44968 0 tt_um_rejunity_sn76489.pwm.accumulator\[7\]
rlabel metal3 44044 44296 44044 44296 0 tt_um_rejunity_sn76489.pwm.accumulator\[8\]
rlabel metal2 43512 41216 43512 41216 0 tt_um_rejunity_sn76489.pwm.accumulator\[9\]
rlabel metal2 44856 36456 44856 36456 0 tt_um_rejunity_sn76489.spi_dac_i_2.counter\[0\]
rlabel metal2 47768 36030 47768 36030 0 tt_um_rejunity_sn76489.spi_dac_i_2.counter\[1\]
rlabel metal2 47880 34216 47880 34216 0 tt_um_rejunity_sn76489.spi_dac_i_2.counter\[2\]
rlabel metal2 45640 32760 45640 32760 0 tt_um_rejunity_sn76489.spi_dac_i_2.counter\[3\]
rlabel metal2 48048 32676 48048 32676 0 tt_um_rejunity_sn76489.spi_dac_i_2.counter\[4\]
rlabel metal2 41272 31846 41272 31846 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[0\]
rlabel metal3 46144 38248 46144 38248 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[10\]
rlabel via2 43064 31734 43064 31734 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[11\]
rlabel metal2 40712 31668 40712 31668 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[1\]
rlabel metal2 40880 33432 40880 33432 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[2\]
rlabel metal2 42168 35098 42168 35098 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[3\]
rlabel via2 41160 36438 41160 36438 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[4\]
rlabel metal2 40264 37408 40264 37408 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[5\]
rlabel metal2 41720 38118 41720 38118 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[6\]
rlabel metal3 40936 38696 40936 38696 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[7\]
rlabel metal2 44072 39368 44072 39368 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[8\]
rlabel metal2 45640 39172 45640 39172 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[9\]
rlabel metal2 26040 6586 26040 6586 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[0\]
rlabel metal2 26040 3304 26040 3304 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[1\]
rlabel metal2 20048 5012 20048 5012 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[2\]
rlabel metal3 18452 5096 18452 5096 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[3\]
rlabel metal2 13888 7588 13888 7588 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[4\]
rlabel metal2 18350 7410 18350 7410 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[5\]
rlabel metal2 15792 6468 15792 6468 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[6\]
rlabel metal2 14504 8792 14504 8792 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[7\]
rlabel metal2 16408 11032 16408 11032 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[8\]
rlabel metal3 16716 13720 16716 13720 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[9\]
rlabel metal2 39198 8092 39198 8092 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[0\]
rlabel metal2 46312 6832 46312 6832 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[1\]
rlabel metal2 45696 7336 45696 7336 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[2\]
rlabel metal2 42979 5096 42979 5096 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[3\]
rlabel metal2 41272 5775 41272 5775 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[4\]
rlabel metal2 39928 9072 39928 9072 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[5\]
rlabel metal2 39424 4424 39424 4424 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[6\]
rlabel metal2 40936 5768 40936 5768 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[7\]
rlabel metal2 39312 9128 39312 9128 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[8\]
rlabel metal2 35672 11424 35672 11424 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[9\]
rlabel metal2 43848 17326 43848 17326 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[0\]
rlabel metal2 44072 17360 44072 17360 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[1\]
rlabel metal2 44856 18816 44856 18816 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[2\]
rlabel metal2 48104 17192 48104 17192 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[3\]
rlabel metal2 43624 13798 43624 13798 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[4\]
rlabel metal2 43546 15250 43546 15250 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[5\]
rlabel metal2 45640 15736 45640 15736 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[6\]
rlabel metal2 47768 10472 47768 10472 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[7\]
rlabel metal2 40376 11144 40376 11144 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[8\]
rlabel metal2 40600 12712 40600 12712 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[9\]
rlabel metal3 504 8120 504 8120 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
