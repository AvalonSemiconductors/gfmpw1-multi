* NGSPICE file created from diceroll.ext - technology: gf180mcuD

.subckt diceroll io_in io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] rst_n vdd vss wb_clk_i
.ends

