VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_ay8913
  CLASS BLOCK ;
  FOREIGN wrapped_ay8913 ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN custom_settings[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 250.880 300.000 251.440 ;
    END
  END custom_settings[0]
  PIN custom_settings[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 280.000 300.000 280.560 ;
    END
  END custom_settings[1]
  PIN io_in_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 17.920 300.000 18.480 ;
    END
  END io_in_1[0]
  PIN io_in_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 47.040 300.000 47.600 ;
    END
  END io_in_1[1]
  PIN io_in_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 76.160 300.000 76.720 ;
    END
  END io_in_1[2]
  PIN io_in_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 105.280 300.000 105.840 ;
    END
  END io_in_1[3]
  PIN io_in_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 134.400 300.000 134.960 ;
    END
  END io_in_1[4]
  PIN io_in_1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 163.520 300.000 164.080 ;
    END
  END io_in_1[5]
  PIN io_in_1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 192.640 300.000 193.200 ;
    END
  END io_in_1[6]
  PIN io_in_1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 221.760 300.000 222.320 ;
    END
  END io_in_1[7]
  PIN io_in_2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 187.040 296.000 187.600 300.000 ;
    END
  END io_in_2[0]
  PIN io_in_2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 296.000 262.640 300.000 ;
    END
  END io_in_2[1]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 0.000 14.000 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 0.000 114.800 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 0.000 124.880 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 0.000 134.960 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 0.000 145.040 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 0.000 155.120 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 0.000 165.200 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 174.720 0.000 175.280 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 0.000 185.360 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 0.000 195.440 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 0.000 205.520 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 0.000 24.080 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 215.040 0.000 215.600 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 0.000 225.680 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 235.200 0.000 235.760 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 245.280 0.000 245.840 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 255.360 0.000 255.920 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.440 0.000 266.000 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 0.000 276.080 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 285.600 0.000 286.160 4.000 ;
    END
  END io_out[27]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 0.000 34.160 4.000 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 0.000 44.240 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 0.000 54.320 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 0.000 64.400 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 0.000 74.480 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 0.000 84.560 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 0.000 94.640 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 0.000 104.720 4.000 ;
    END
  END io_out[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 112.000 296.000 112.560 300.000 ;
    END
  END rst_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 282.540 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 282.540 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 296.000 37.520 300.000 ;
    END
  END wb_clk_i
  OBS
      LAYER Pwell ;
        RECT 6.290 280.480 293.310 282.670 ;
      LAYER Nwell ;
        RECT 6.290 276.285 293.310 280.480 ;
        RECT 6.290 276.160 91.665 276.285 ;
      LAYER Pwell ;
        RECT 6.290 272.640 293.310 276.160 ;
      LAYER Nwell ;
        RECT 6.290 272.515 91.105 272.640 ;
        RECT 6.290 268.445 293.310 272.515 ;
        RECT 6.290 268.320 165.800 268.445 ;
      LAYER Pwell ;
        RECT 6.290 264.800 293.310 268.320 ;
      LAYER Nwell ;
        RECT 6.290 260.605 293.310 264.800 ;
        RECT 6.290 260.480 79.905 260.605 ;
      LAYER Pwell ;
        RECT 6.290 256.960 293.310 260.480 ;
      LAYER Nwell ;
        RECT 6.290 256.835 175.105 256.960 ;
        RECT 6.290 252.765 293.310 256.835 ;
        RECT 6.290 252.640 117.425 252.765 ;
      LAYER Pwell ;
        RECT 6.290 249.120 293.310 252.640 ;
      LAYER Nwell ;
        RECT 6.290 248.995 66.120 249.120 ;
        RECT 6.290 244.925 293.310 248.995 ;
        RECT 6.290 244.800 81.025 244.925 ;
      LAYER Pwell ;
        RECT 6.290 241.280 293.310 244.800 ;
      LAYER Nwell ;
        RECT 6.290 241.155 34.545 241.280 ;
        RECT 6.290 237.085 293.310 241.155 ;
        RECT 6.290 236.960 132.695 237.085 ;
      LAYER Pwell ;
        RECT 6.290 233.440 293.310 236.960 ;
      LAYER Nwell ;
        RECT 6.290 233.315 30.280 233.440 ;
        RECT 6.290 229.245 293.310 233.315 ;
        RECT 6.290 229.120 240.065 229.245 ;
      LAYER Pwell ;
        RECT 6.290 225.600 293.310 229.120 ;
      LAYER Nwell ;
        RECT 6.290 225.475 80.505 225.600 ;
        RECT 6.290 221.405 293.310 225.475 ;
        RECT 6.290 221.280 91.105 221.405 ;
      LAYER Pwell ;
        RECT 6.290 217.760 293.310 221.280 ;
      LAYER Nwell ;
        RECT 6.290 217.635 33.080 217.760 ;
        RECT 6.290 213.565 293.310 217.635 ;
        RECT 6.290 213.440 125.825 213.565 ;
      LAYER Pwell ;
        RECT 6.290 209.920 293.310 213.440 ;
      LAYER Nwell ;
        RECT 6.290 209.795 63.665 209.920 ;
        RECT 6.290 205.725 293.310 209.795 ;
        RECT 6.290 205.600 46.305 205.725 ;
      LAYER Pwell ;
        RECT 6.290 202.080 293.310 205.600 ;
      LAYER Nwell ;
        RECT 6.290 201.955 60.865 202.080 ;
        RECT 6.290 197.885 293.310 201.955 ;
        RECT 6.290 197.760 12.705 197.885 ;
      LAYER Pwell ;
        RECT 6.290 194.240 293.310 197.760 ;
      LAYER Nwell ;
        RECT 6.290 194.115 12.705 194.240 ;
        RECT 6.290 190.045 293.310 194.115 ;
        RECT 6.290 189.920 85.505 190.045 ;
      LAYER Pwell ;
        RECT 6.290 186.400 293.310 189.920 ;
      LAYER Nwell ;
        RECT 6.290 186.275 66.465 186.400 ;
        RECT 6.290 182.205 293.310 186.275 ;
        RECT 6.290 182.080 12.705 182.205 ;
      LAYER Pwell ;
        RECT 6.290 178.560 293.310 182.080 ;
      LAYER Nwell ;
        RECT 6.290 178.435 103.425 178.560 ;
        RECT 6.290 174.365 293.310 178.435 ;
        RECT 6.290 174.240 51.560 174.365 ;
      LAYER Pwell ;
        RECT 6.290 170.720 293.310 174.240 ;
      LAYER Nwell ;
        RECT 6.290 170.595 62.545 170.720 ;
        RECT 6.290 166.525 293.310 170.595 ;
        RECT 6.290 166.400 12.705 166.525 ;
      LAYER Pwell ;
        RECT 6.290 162.880 293.310 166.400 ;
      LAYER Nwell ;
        RECT 6.290 162.755 12.705 162.880 ;
        RECT 6.290 158.685 293.310 162.755 ;
        RECT 6.290 158.560 59.400 158.685 ;
      LAYER Pwell ;
        RECT 6.290 155.040 293.310 158.560 ;
      LAYER Nwell ;
        RECT 6.290 154.915 69.265 155.040 ;
        RECT 6.290 150.845 293.310 154.915 ;
        RECT 6.290 150.720 12.705 150.845 ;
      LAYER Pwell ;
        RECT 6.290 147.200 293.310 150.720 ;
      LAYER Nwell ;
        RECT 6.290 147.075 110.705 147.200 ;
        RECT 6.290 143.005 293.310 147.075 ;
        RECT 6.290 142.880 92.225 143.005 ;
      LAYER Pwell ;
        RECT 6.290 139.360 293.310 142.880 ;
      LAYER Nwell ;
        RECT 6.290 139.235 12.705 139.360 ;
        RECT 6.290 135.040 293.310 139.235 ;
      LAYER Pwell ;
        RECT 6.290 131.520 293.310 135.040 ;
      LAYER Nwell ;
        RECT 6.290 131.395 63.880 131.520 ;
        RECT 6.290 127.325 293.310 131.395 ;
        RECT 6.290 127.200 44.065 127.325 ;
      LAYER Pwell ;
        RECT 6.290 123.680 293.310 127.200 ;
      LAYER Nwell ;
        RECT 6.290 123.555 12.705 123.680 ;
        RECT 6.290 119.485 293.310 123.555 ;
        RECT 6.290 119.360 93.345 119.485 ;
      LAYER Pwell ;
        RECT 6.290 115.840 293.310 119.360 ;
      LAYER Nwell ;
        RECT 6.290 115.715 12.705 115.840 ;
        RECT 6.290 111.645 293.310 115.715 ;
        RECT 6.290 111.520 37.345 111.645 ;
      LAYER Pwell ;
        RECT 6.290 108.000 293.310 111.520 ;
      LAYER Nwell ;
        RECT 6.290 107.875 169.505 108.000 ;
        RECT 6.290 103.805 293.310 107.875 ;
        RECT 6.290 103.680 12.705 103.805 ;
      LAYER Pwell ;
        RECT 6.290 100.160 293.310 103.680 ;
      LAYER Nwell ;
        RECT 6.290 100.035 51.905 100.160 ;
        RECT 6.290 95.965 293.310 100.035 ;
        RECT 6.290 95.840 84.040 95.965 ;
      LAYER Pwell ;
        RECT 6.290 92.320 293.310 95.840 ;
      LAYER Nwell ;
        RECT 6.290 92.195 31.960 92.320 ;
        RECT 6.290 88.125 293.310 92.195 ;
        RECT 6.290 88.000 12.705 88.125 ;
      LAYER Pwell ;
        RECT 6.290 84.480 293.310 88.000 ;
      LAYER Nwell ;
        RECT 6.290 84.355 106.440 84.480 ;
        RECT 6.290 80.285 293.310 84.355 ;
        RECT 6.290 80.160 53.800 80.285 ;
      LAYER Pwell ;
        RECT 6.290 76.640 293.310 80.160 ;
      LAYER Nwell ;
        RECT 6.290 76.515 27.825 76.640 ;
        RECT 6.290 72.445 293.310 76.515 ;
        RECT 6.290 72.320 12.705 72.445 ;
      LAYER Pwell ;
        RECT 6.290 68.800 293.310 72.320 ;
      LAYER Nwell ;
        RECT 6.290 68.675 55.825 68.800 ;
        RECT 6.290 64.605 293.310 68.675 ;
        RECT 6.290 64.480 35.665 64.605 ;
      LAYER Pwell ;
        RECT 6.290 60.960 293.310 64.480 ;
      LAYER Nwell ;
        RECT 6.290 60.835 100.065 60.960 ;
        RECT 6.290 56.765 293.310 60.835 ;
        RECT 6.290 56.640 12.705 56.765 ;
      LAYER Pwell ;
        RECT 6.290 53.120 293.310 56.640 ;
      LAYER Nwell ;
        RECT 6.290 52.995 98.385 53.120 ;
        RECT 6.290 48.925 293.310 52.995 ;
        RECT 6.290 48.800 14.945 48.925 ;
      LAYER Pwell ;
        RECT 6.290 45.280 293.310 48.800 ;
      LAYER Nwell ;
        RECT 6.290 45.155 91.105 45.280 ;
        RECT 6.290 41.085 293.310 45.155 ;
        RECT 6.290 40.960 95.800 41.085 ;
      LAYER Pwell ;
        RECT 6.290 37.440 293.310 40.960 ;
      LAYER Nwell ;
        RECT 6.290 37.315 60.305 37.440 ;
        RECT 6.290 33.245 293.310 37.315 ;
        RECT 6.290 33.120 39.240 33.245 ;
      LAYER Pwell ;
        RECT 6.290 29.600 293.310 33.120 ;
      LAYER Nwell ;
        RECT 6.290 29.475 191.345 29.600 ;
        RECT 6.290 25.405 293.310 29.475 ;
        RECT 6.290 25.280 53.585 25.405 ;
      LAYER Pwell ;
        RECT 6.290 21.760 293.310 25.280 ;
      LAYER Nwell ;
        RECT 6.290 21.635 54.705 21.760 ;
        RECT 6.290 17.565 293.310 21.635 ;
        RECT 6.290 17.440 222.145 17.565 ;
      LAYER Pwell ;
        RECT 6.290 15.250 293.310 17.440 ;
      LAYER Metal1 ;
        RECT 6.720 8.550 292.880 282.540 ;
      LAYER Metal2 ;
        RECT 9.100 295.700 36.660 296.000 ;
        RECT 37.820 295.700 111.700 296.000 ;
        RECT 112.860 295.700 186.740 296.000 ;
        RECT 187.900 295.700 261.780 296.000 ;
        RECT 262.940 295.700 291.620 296.000 ;
        RECT 9.100 4.300 291.620 295.700 ;
        RECT 9.100 3.500 13.140 4.300 ;
        RECT 14.300 3.500 23.220 4.300 ;
        RECT 24.380 3.500 33.300 4.300 ;
        RECT 34.460 3.500 43.380 4.300 ;
        RECT 44.540 3.500 53.460 4.300 ;
        RECT 54.620 3.500 63.540 4.300 ;
        RECT 64.700 3.500 73.620 4.300 ;
        RECT 74.780 3.500 83.700 4.300 ;
        RECT 84.860 3.500 93.780 4.300 ;
        RECT 94.940 3.500 103.860 4.300 ;
        RECT 105.020 3.500 113.940 4.300 ;
        RECT 115.100 3.500 124.020 4.300 ;
        RECT 125.180 3.500 134.100 4.300 ;
        RECT 135.260 3.500 144.180 4.300 ;
        RECT 145.340 3.500 154.260 4.300 ;
        RECT 155.420 3.500 164.340 4.300 ;
        RECT 165.500 3.500 174.420 4.300 ;
        RECT 175.580 3.500 184.500 4.300 ;
        RECT 185.660 3.500 194.580 4.300 ;
        RECT 195.740 3.500 204.660 4.300 ;
        RECT 205.820 3.500 214.740 4.300 ;
        RECT 215.900 3.500 224.820 4.300 ;
        RECT 225.980 3.500 234.900 4.300 ;
        RECT 236.060 3.500 244.980 4.300 ;
        RECT 246.140 3.500 255.060 4.300 ;
        RECT 256.220 3.500 265.140 4.300 ;
        RECT 266.300 3.500 275.220 4.300 ;
        RECT 276.380 3.500 285.300 4.300 ;
        RECT 286.460 3.500 291.620 4.300 ;
      LAYER Metal3 ;
        RECT 9.050 280.860 296.000 282.380 ;
        RECT 9.050 279.700 295.700 280.860 ;
        RECT 9.050 251.740 296.000 279.700 ;
        RECT 9.050 250.580 295.700 251.740 ;
        RECT 9.050 222.620 296.000 250.580 ;
        RECT 9.050 221.460 295.700 222.620 ;
        RECT 9.050 193.500 296.000 221.460 ;
        RECT 9.050 192.340 295.700 193.500 ;
        RECT 9.050 164.380 296.000 192.340 ;
        RECT 9.050 163.220 295.700 164.380 ;
        RECT 9.050 135.260 296.000 163.220 ;
        RECT 9.050 134.100 295.700 135.260 ;
        RECT 9.050 106.140 296.000 134.100 ;
        RECT 9.050 104.980 295.700 106.140 ;
        RECT 9.050 77.020 296.000 104.980 ;
        RECT 9.050 75.860 295.700 77.020 ;
        RECT 9.050 47.900 296.000 75.860 ;
        RECT 9.050 46.740 295.700 47.900 ;
        RECT 9.050 18.780 296.000 46.740 ;
        RECT 9.050 17.620 295.700 18.780 ;
        RECT 9.050 15.540 296.000 17.620 ;
      LAYER Metal4 ;
        RECT 43.260 35.930 98.740 279.910 ;
        RECT 100.940 35.930 175.540 279.910 ;
        RECT 177.740 35.930 252.340 279.910 ;
        RECT 254.540 35.930 272.580 279.910 ;
  END
END wrapped_ay8913
END LIBRARY

