magic
tech gf180mcuD
magscale 1 5
timestamp 1702046838
<< obsm1 >>
rect 672 1538 69328 63142
<< metal2 >>
rect 224 64600 280 65000
rect 672 64600 728 65000
rect 1120 64600 1176 65000
rect 1568 64600 1624 65000
rect 2016 64600 2072 65000
rect 2464 64600 2520 65000
rect 2912 64600 2968 65000
rect 3360 64600 3416 65000
rect 3808 64600 3864 65000
rect 4256 64600 4312 65000
rect 4704 64600 4760 65000
rect 5152 64600 5208 65000
rect 5600 64600 5656 65000
rect 6048 64600 6104 65000
rect 6496 64600 6552 65000
rect 6944 64600 7000 65000
rect 7392 64600 7448 65000
rect 7840 64600 7896 65000
rect 8288 64600 8344 65000
rect 8736 64600 8792 65000
rect 9184 64600 9240 65000
rect 9632 64600 9688 65000
rect 10080 64600 10136 65000
rect 10528 64600 10584 65000
rect 10976 64600 11032 65000
rect 11424 64600 11480 65000
rect 11872 64600 11928 65000
rect 12320 64600 12376 65000
rect 12768 64600 12824 65000
rect 13216 64600 13272 65000
rect 13664 64600 13720 65000
rect 14112 64600 14168 65000
rect 14560 64600 14616 65000
rect 15008 64600 15064 65000
rect 15456 64600 15512 65000
rect 15904 64600 15960 65000
rect 16352 64600 16408 65000
rect 16800 64600 16856 65000
rect 17248 64600 17304 65000
rect 17696 64600 17752 65000
rect 18144 64600 18200 65000
rect 18592 64600 18648 65000
rect 19040 64600 19096 65000
rect 19488 64600 19544 65000
rect 19936 64600 19992 65000
rect 20384 64600 20440 65000
rect 20832 64600 20888 65000
rect 21280 64600 21336 65000
rect 21728 64600 21784 65000
rect 22176 64600 22232 65000
rect 22624 64600 22680 65000
rect 23072 64600 23128 65000
rect 23520 64600 23576 65000
rect 23968 64600 24024 65000
rect 24416 64600 24472 65000
rect 24864 64600 24920 65000
rect 25312 64600 25368 65000
rect 25760 64600 25816 65000
rect 26208 64600 26264 65000
rect 26656 64600 26712 65000
rect 27104 64600 27160 65000
rect 27552 64600 27608 65000
rect 28000 64600 28056 65000
rect 28448 64600 28504 65000
rect 28896 64600 28952 65000
rect 29344 64600 29400 65000
rect 29792 64600 29848 65000
rect 30240 64600 30296 65000
rect 30688 64600 30744 65000
rect 31136 64600 31192 65000
rect 31584 64600 31640 65000
rect 32032 64600 32088 65000
rect 32480 64600 32536 65000
rect 32928 64600 32984 65000
rect 33376 64600 33432 65000
rect 33824 64600 33880 65000
rect 34272 64600 34328 65000
rect 34720 64600 34776 65000
rect 35168 64600 35224 65000
rect 35616 64600 35672 65000
rect 36064 64600 36120 65000
rect 36512 64600 36568 65000
rect 36960 64600 37016 65000
rect 37408 64600 37464 65000
rect 37856 64600 37912 65000
rect 38304 64600 38360 65000
rect 38752 64600 38808 65000
rect 39200 64600 39256 65000
rect 39648 64600 39704 65000
rect 40096 64600 40152 65000
rect 40544 64600 40600 65000
rect 40992 64600 41048 65000
rect 41440 64600 41496 65000
rect 41888 64600 41944 65000
rect 42336 64600 42392 65000
rect 42784 64600 42840 65000
rect 43232 64600 43288 65000
rect 43680 64600 43736 65000
rect 44128 64600 44184 65000
rect 44576 64600 44632 65000
rect 45024 64600 45080 65000
rect 45472 64600 45528 65000
rect 45920 64600 45976 65000
rect 46368 64600 46424 65000
rect 46816 64600 46872 65000
rect 47264 64600 47320 65000
rect 47712 64600 47768 65000
rect 48160 64600 48216 65000
rect 48608 64600 48664 65000
rect 49056 64600 49112 65000
rect 49504 64600 49560 65000
rect 49952 64600 50008 65000
rect 50400 64600 50456 65000
rect 50848 64600 50904 65000
rect 51296 64600 51352 65000
rect 51744 64600 51800 65000
rect 52192 64600 52248 65000
rect 52640 64600 52696 65000
rect 53088 64600 53144 65000
rect 53536 64600 53592 65000
rect 53984 64600 54040 65000
rect 54432 64600 54488 65000
rect 54880 64600 54936 65000
rect 55328 64600 55384 65000
rect 55776 64600 55832 65000
rect 56224 64600 56280 65000
rect 56672 64600 56728 65000
rect 57120 64600 57176 65000
rect 57568 64600 57624 65000
rect 58016 64600 58072 65000
rect 58464 64600 58520 65000
rect 58912 64600 58968 65000
rect 59360 64600 59416 65000
rect 59808 64600 59864 65000
rect 60256 64600 60312 65000
rect 60704 64600 60760 65000
rect 61152 64600 61208 65000
rect 61600 64600 61656 65000
rect 62048 64600 62104 65000
rect 62496 64600 62552 65000
rect 62944 64600 63000 65000
rect 63392 64600 63448 65000
rect 63840 64600 63896 65000
rect 64288 64600 64344 65000
rect 64736 64600 64792 65000
rect 65184 64600 65240 65000
rect 65632 64600 65688 65000
rect 66080 64600 66136 65000
rect 66528 64600 66584 65000
rect 66976 64600 67032 65000
rect 67424 64600 67480 65000
rect 67872 64600 67928 65000
rect 68320 64600 68376 65000
rect 68768 64600 68824 65000
rect 69216 64600 69272 65000
rect 69664 64600 69720 65000
rect 3360 0 3416 400
rect 3808 0 3864 400
rect 4256 0 4312 400
rect 4704 0 4760 400
rect 5152 0 5208 400
rect 5600 0 5656 400
rect 6048 0 6104 400
rect 6496 0 6552 400
rect 6944 0 7000 400
rect 7392 0 7448 400
rect 7840 0 7896 400
rect 8288 0 8344 400
rect 8736 0 8792 400
rect 9184 0 9240 400
rect 9632 0 9688 400
rect 10080 0 10136 400
rect 10528 0 10584 400
rect 10976 0 11032 400
rect 11424 0 11480 400
rect 11872 0 11928 400
rect 12320 0 12376 400
rect 12768 0 12824 400
rect 13216 0 13272 400
rect 13664 0 13720 400
rect 14112 0 14168 400
rect 14560 0 14616 400
rect 15008 0 15064 400
rect 15456 0 15512 400
rect 15904 0 15960 400
rect 16352 0 16408 400
rect 16800 0 16856 400
rect 17248 0 17304 400
rect 17696 0 17752 400
rect 18144 0 18200 400
rect 18592 0 18648 400
rect 19040 0 19096 400
rect 19488 0 19544 400
rect 19936 0 19992 400
rect 20384 0 20440 400
rect 20832 0 20888 400
rect 21280 0 21336 400
rect 21728 0 21784 400
rect 22176 0 22232 400
rect 22624 0 22680 400
rect 23072 0 23128 400
rect 23520 0 23576 400
rect 23968 0 24024 400
rect 24416 0 24472 400
rect 24864 0 24920 400
rect 25312 0 25368 400
rect 25760 0 25816 400
rect 26208 0 26264 400
rect 26656 0 26712 400
rect 27104 0 27160 400
rect 27552 0 27608 400
rect 28000 0 28056 400
rect 28448 0 28504 400
rect 28896 0 28952 400
rect 29344 0 29400 400
rect 29792 0 29848 400
rect 30240 0 30296 400
rect 30688 0 30744 400
rect 31136 0 31192 400
rect 31584 0 31640 400
rect 32032 0 32088 400
rect 32480 0 32536 400
rect 32928 0 32984 400
rect 33376 0 33432 400
rect 33824 0 33880 400
rect 34272 0 34328 400
rect 34720 0 34776 400
rect 35168 0 35224 400
rect 35616 0 35672 400
rect 36064 0 36120 400
rect 36512 0 36568 400
rect 36960 0 37016 400
rect 37408 0 37464 400
rect 37856 0 37912 400
rect 38304 0 38360 400
rect 38752 0 38808 400
rect 39200 0 39256 400
rect 39648 0 39704 400
rect 40096 0 40152 400
rect 40544 0 40600 400
rect 40992 0 41048 400
rect 41440 0 41496 400
rect 41888 0 41944 400
rect 42336 0 42392 400
rect 42784 0 42840 400
rect 43232 0 43288 400
rect 43680 0 43736 400
rect 44128 0 44184 400
rect 44576 0 44632 400
rect 45024 0 45080 400
rect 45472 0 45528 400
rect 45920 0 45976 400
rect 46368 0 46424 400
rect 46816 0 46872 400
rect 47264 0 47320 400
rect 47712 0 47768 400
rect 48160 0 48216 400
rect 48608 0 48664 400
rect 49056 0 49112 400
rect 49504 0 49560 400
rect 49952 0 50008 400
rect 50400 0 50456 400
rect 50848 0 50904 400
rect 51296 0 51352 400
rect 51744 0 51800 400
rect 52192 0 52248 400
rect 52640 0 52696 400
rect 53088 0 53144 400
rect 53536 0 53592 400
rect 53984 0 54040 400
rect 54432 0 54488 400
rect 54880 0 54936 400
rect 55328 0 55384 400
rect 55776 0 55832 400
rect 56224 0 56280 400
rect 56672 0 56728 400
rect 57120 0 57176 400
rect 57568 0 57624 400
rect 58016 0 58072 400
rect 58464 0 58520 400
rect 58912 0 58968 400
rect 59360 0 59416 400
rect 59808 0 59864 400
rect 60256 0 60312 400
rect 60704 0 60760 400
rect 61152 0 61208 400
rect 61600 0 61656 400
rect 62048 0 62104 400
rect 62496 0 62552 400
rect 62944 0 63000 400
rect 63392 0 63448 400
rect 63840 0 63896 400
rect 64288 0 64344 400
rect 64736 0 64792 400
rect 65184 0 65240 400
rect 65632 0 65688 400
rect 66080 0 66136 400
rect 66528 0 66584 400
<< obsm2 >>
rect 310 64570 642 64666
rect 758 64570 1090 64666
rect 1206 64570 1538 64666
rect 1654 64570 1986 64666
rect 2102 64570 2434 64666
rect 2550 64570 2882 64666
rect 2998 64570 3330 64666
rect 3446 64570 3778 64666
rect 3894 64570 4226 64666
rect 4342 64570 4674 64666
rect 4790 64570 5122 64666
rect 5238 64570 5570 64666
rect 5686 64570 6018 64666
rect 6134 64570 6466 64666
rect 6582 64570 6914 64666
rect 7030 64570 7362 64666
rect 7478 64570 7810 64666
rect 7926 64570 8258 64666
rect 8374 64570 8706 64666
rect 8822 64570 9154 64666
rect 9270 64570 9602 64666
rect 9718 64570 10050 64666
rect 10166 64570 10498 64666
rect 10614 64570 10946 64666
rect 11062 64570 11394 64666
rect 11510 64570 11842 64666
rect 11958 64570 12290 64666
rect 12406 64570 12738 64666
rect 12854 64570 13186 64666
rect 13302 64570 13634 64666
rect 13750 64570 14082 64666
rect 14198 64570 14530 64666
rect 14646 64570 14978 64666
rect 15094 64570 15426 64666
rect 15542 64570 15874 64666
rect 15990 64570 16322 64666
rect 16438 64570 16770 64666
rect 16886 64570 17218 64666
rect 17334 64570 17666 64666
rect 17782 64570 18114 64666
rect 18230 64570 18562 64666
rect 18678 64570 19010 64666
rect 19126 64570 19458 64666
rect 19574 64570 19906 64666
rect 20022 64570 20354 64666
rect 20470 64570 20802 64666
rect 20918 64570 21250 64666
rect 21366 64570 21698 64666
rect 21814 64570 22146 64666
rect 22262 64570 22594 64666
rect 22710 64570 23042 64666
rect 23158 64570 23490 64666
rect 23606 64570 23938 64666
rect 24054 64570 24386 64666
rect 24502 64570 24834 64666
rect 24950 64570 25282 64666
rect 25398 64570 25730 64666
rect 25846 64570 26178 64666
rect 26294 64570 26626 64666
rect 26742 64570 27074 64666
rect 27190 64570 27522 64666
rect 27638 64570 27970 64666
rect 28086 64570 28418 64666
rect 28534 64570 28866 64666
rect 28982 64570 29314 64666
rect 29430 64570 29762 64666
rect 29878 64570 30210 64666
rect 30326 64570 30658 64666
rect 30774 64570 31106 64666
rect 31222 64570 31554 64666
rect 31670 64570 32002 64666
rect 32118 64570 32450 64666
rect 32566 64570 32898 64666
rect 33014 64570 33346 64666
rect 33462 64570 33794 64666
rect 33910 64570 34242 64666
rect 34358 64570 34690 64666
rect 34806 64570 35138 64666
rect 35254 64570 35586 64666
rect 35702 64570 36034 64666
rect 36150 64570 36482 64666
rect 36598 64570 36930 64666
rect 37046 64570 37378 64666
rect 37494 64570 37826 64666
rect 37942 64570 38274 64666
rect 38390 64570 38722 64666
rect 38838 64570 39170 64666
rect 39286 64570 39618 64666
rect 39734 64570 40066 64666
rect 40182 64570 40514 64666
rect 40630 64570 40962 64666
rect 41078 64570 41410 64666
rect 41526 64570 41858 64666
rect 41974 64570 42306 64666
rect 42422 64570 42754 64666
rect 42870 64570 43202 64666
rect 43318 64570 43650 64666
rect 43766 64570 44098 64666
rect 44214 64570 44546 64666
rect 44662 64570 44994 64666
rect 45110 64570 45442 64666
rect 45558 64570 45890 64666
rect 46006 64570 46338 64666
rect 46454 64570 46786 64666
rect 46902 64570 47234 64666
rect 47350 64570 47682 64666
rect 47798 64570 48130 64666
rect 48246 64570 48578 64666
rect 48694 64570 49026 64666
rect 49142 64570 49474 64666
rect 49590 64570 49922 64666
rect 50038 64570 50370 64666
rect 50486 64570 50818 64666
rect 50934 64570 51266 64666
rect 51382 64570 51714 64666
rect 51830 64570 52162 64666
rect 52278 64570 52610 64666
rect 52726 64570 53058 64666
rect 53174 64570 53506 64666
rect 53622 64570 53954 64666
rect 54070 64570 54402 64666
rect 54518 64570 54850 64666
rect 54966 64570 55298 64666
rect 55414 64570 55746 64666
rect 55862 64570 56194 64666
rect 56310 64570 56642 64666
rect 56758 64570 57090 64666
rect 57206 64570 57538 64666
rect 57654 64570 57986 64666
rect 58102 64570 58434 64666
rect 58550 64570 58882 64666
rect 58998 64570 59330 64666
rect 59446 64570 59778 64666
rect 59894 64570 60226 64666
rect 60342 64570 60674 64666
rect 60790 64570 61122 64666
rect 61238 64570 61570 64666
rect 61686 64570 62018 64666
rect 62134 64570 62466 64666
rect 62582 64570 62914 64666
rect 63030 64570 63362 64666
rect 63478 64570 63810 64666
rect 63926 64570 64258 64666
rect 64374 64570 64706 64666
rect 64822 64570 65154 64666
rect 65270 64570 65602 64666
rect 65718 64570 66050 64666
rect 66166 64570 66498 64666
rect 66614 64570 66946 64666
rect 67062 64570 67394 64666
rect 67510 64570 67842 64666
rect 67958 64570 68290 64666
rect 68406 64570 68738 64666
rect 68854 64570 69186 64666
rect 69302 64570 69634 64666
rect 238 430 69706 64570
rect 238 350 3330 430
rect 3446 350 3778 430
rect 3894 350 4226 430
rect 4342 350 4674 430
rect 4790 350 5122 430
rect 5238 350 5570 430
rect 5686 350 6018 430
rect 6134 350 6466 430
rect 6582 350 6914 430
rect 7030 350 7362 430
rect 7478 350 7810 430
rect 7926 350 8258 430
rect 8374 350 8706 430
rect 8822 350 9154 430
rect 9270 350 9602 430
rect 9718 350 10050 430
rect 10166 350 10498 430
rect 10614 350 10946 430
rect 11062 350 11394 430
rect 11510 350 11842 430
rect 11958 350 12290 430
rect 12406 350 12738 430
rect 12854 350 13186 430
rect 13302 350 13634 430
rect 13750 350 14082 430
rect 14198 350 14530 430
rect 14646 350 14978 430
rect 15094 350 15426 430
rect 15542 350 15874 430
rect 15990 350 16322 430
rect 16438 350 16770 430
rect 16886 350 17218 430
rect 17334 350 17666 430
rect 17782 350 18114 430
rect 18230 350 18562 430
rect 18678 350 19010 430
rect 19126 350 19458 430
rect 19574 350 19906 430
rect 20022 350 20354 430
rect 20470 350 20802 430
rect 20918 350 21250 430
rect 21366 350 21698 430
rect 21814 350 22146 430
rect 22262 350 22594 430
rect 22710 350 23042 430
rect 23158 350 23490 430
rect 23606 350 23938 430
rect 24054 350 24386 430
rect 24502 350 24834 430
rect 24950 350 25282 430
rect 25398 350 25730 430
rect 25846 350 26178 430
rect 26294 350 26626 430
rect 26742 350 27074 430
rect 27190 350 27522 430
rect 27638 350 27970 430
rect 28086 350 28418 430
rect 28534 350 28866 430
rect 28982 350 29314 430
rect 29430 350 29762 430
rect 29878 350 30210 430
rect 30326 350 30658 430
rect 30774 350 31106 430
rect 31222 350 31554 430
rect 31670 350 32002 430
rect 32118 350 32450 430
rect 32566 350 32898 430
rect 33014 350 33346 430
rect 33462 350 33794 430
rect 33910 350 34242 430
rect 34358 350 34690 430
rect 34806 350 35138 430
rect 35254 350 35586 430
rect 35702 350 36034 430
rect 36150 350 36482 430
rect 36598 350 36930 430
rect 37046 350 37378 430
rect 37494 350 37826 430
rect 37942 350 38274 430
rect 38390 350 38722 430
rect 38838 350 39170 430
rect 39286 350 39618 430
rect 39734 350 40066 430
rect 40182 350 40514 430
rect 40630 350 40962 430
rect 41078 350 41410 430
rect 41526 350 41858 430
rect 41974 350 42306 430
rect 42422 350 42754 430
rect 42870 350 43202 430
rect 43318 350 43650 430
rect 43766 350 44098 430
rect 44214 350 44546 430
rect 44662 350 44994 430
rect 45110 350 45442 430
rect 45558 350 45890 430
rect 46006 350 46338 430
rect 46454 350 46786 430
rect 46902 350 47234 430
rect 47350 350 47682 430
rect 47798 350 48130 430
rect 48246 350 48578 430
rect 48694 350 49026 430
rect 49142 350 49474 430
rect 49590 350 49922 430
rect 50038 350 50370 430
rect 50486 350 50818 430
rect 50934 350 51266 430
rect 51382 350 51714 430
rect 51830 350 52162 430
rect 52278 350 52610 430
rect 52726 350 53058 430
rect 53174 350 53506 430
rect 53622 350 53954 430
rect 54070 350 54402 430
rect 54518 350 54850 430
rect 54966 350 55298 430
rect 55414 350 55746 430
rect 55862 350 56194 430
rect 56310 350 56642 430
rect 56758 350 57090 430
rect 57206 350 57538 430
rect 57654 350 57986 430
rect 58102 350 58434 430
rect 58550 350 58882 430
rect 58998 350 59330 430
rect 59446 350 59778 430
rect 59894 350 60226 430
rect 60342 350 60674 430
rect 60790 350 61122 430
rect 61238 350 61570 430
rect 61686 350 62018 430
rect 62134 350 62466 430
rect 62582 350 62914 430
rect 63030 350 63362 430
rect 63478 350 63810 430
rect 63926 350 64258 430
rect 64374 350 64706 430
rect 64822 350 65154 430
rect 65270 350 65602 430
rect 65718 350 66050 430
rect 66166 350 66498 430
rect 66614 350 69706 430
<< metal3 >>
rect 69600 63168 70000 63224
rect 69600 62608 70000 62664
rect 69600 62048 70000 62104
rect 69600 61488 70000 61544
rect 69600 60928 70000 60984
rect 0 60704 400 60760
rect 69600 60368 70000 60424
rect 0 60144 400 60200
rect 69600 59808 70000 59864
rect 0 59584 400 59640
rect 69600 59248 70000 59304
rect 0 59024 400 59080
rect 69600 58688 70000 58744
rect 0 58464 400 58520
rect 69600 58128 70000 58184
rect 0 57904 400 57960
rect 69600 57568 70000 57624
rect 0 57344 400 57400
rect 69600 57008 70000 57064
rect 0 56784 400 56840
rect 69600 56448 70000 56504
rect 0 56224 400 56280
rect 69600 55888 70000 55944
rect 0 55664 400 55720
rect 69600 55328 70000 55384
rect 0 55104 400 55160
rect 69600 54768 70000 54824
rect 0 54544 400 54600
rect 69600 54208 70000 54264
rect 0 53984 400 54040
rect 69600 53648 70000 53704
rect 0 53424 400 53480
rect 69600 53088 70000 53144
rect 0 52864 400 52920
rect 69600 52528 70000 52584
rect 0 52304 400 52360
rect 69600 51968 70000 52024
rect 0 51744 400 51800
rect 69600 51408 70000 51464
rect 0 51184 400 51240
rect 69600 50848 70000 50904
rect 0 50624 400 50680
rect 69600 50288 70000 50344
rect 0 50064 400 50120
rect 69600 49728 70000 49784
rect 0 49504 400 49560
rect 69600 49168 70000 49224
rect 0 48944 400 49000
rect 69600 48608 70000 48664
rect 0 48384 400 48440
rect 69600 48048 70000 48104
rect 0 47824 400 47880
rect 69600 47488 70000 47544
rect 0 47264 400 47320
rect 69600 46928 70000 46984
rect 0 46704 400 46760
rect 69600 46368 70000 46424
rect 0 46144 400 46200
rect 69600 45808 70000 45864
rect 0 45584 400 45640
rect 69600 45248 70000 45304
rect 0 45024 400 45080
rect 69600 44688 70000 44744
rect 0 44464 400 44520
rect 69600 44128 70000 44184
rect 0 43904 400 43960
rect 69600 43568 70000 43624
rect 0 43344 400 43400
rect 69600 43008 70000 43064
rect 0 42784 400 42840
rect 69600 42448 70000 42504
rect 0 42224 400 42280
rect 69600 41888 70000 41944
rect 0 41664 400 41720
rect 69600 41328 70000 41384
rect 0 41104 400 41160
rect 69600 40768 70000 40824
rect 0 40544 400 40600
rect 69600 40208 70000 40264
rect 0 39984 400 40040
rect 69600 39648 70000 39704
rect 0 39424 400 39480
rect 69600 39088 70000 39144
rect 0 38864 400 38920
rect 69600 38528 70000 38584
rect 0 38304 400 38360
rect 69600 37968 70000 38024
rect 0 37744 400 37800
rect 69600 37408 70000 37464
rect 0 37184 400 37240
rect 69600 36848 70000 36904
rect 0 36624 400 36680
rect 69600 36288 70000 36344
rect 0 36064 400 36120
rect 69600 35728 70000 35784
rect 0 35504 400 35560
rect 69600 35168 70000 35224
rect 0 34944 400 35000
rect 69600 34608 70000 34664
rect 0 34384 400 34440
rect 69600 34048 70000 34104
rect 0 33824 400 33880
rect 69600 33488 70000 33544
rect 0 33264 400 33320
rect 69600 32928 70000 32984
rect 0 32704 400 32760
rect 69600 32368 70000 32424
rect 0 32144 400 32200
rect 69600 31808 70000 31864
rect 0 31584 400 31640
rect 69600 31248 70000 31304
rect 0 31024 400 31080
rect 69600 30688 70000 30744
rect 0 30464 400 30520
rect 69600 30128 70000 30184
rect 0 29904 400 29960
rect 69600 29568 70000 29624
rect 0 29344 400 29400
rect 69600 29008 70000 29064
rect 0 28784 400 28840
rect 69600 28448 70000 28504
rect 0 28224 400 28280
rect 69600 27888 70000 27944
rect 0 27664 400 27720
rect 69600 27328 70000 27384
rect 0 27104 400 27160
rect 69600 26768 70000 26824
rect 0 26544 400 26600
rect 69600 26208 70000 26264
rect 0 25984 400 26040
rect 69600 25648 70000 25704
rect 0 25424 400 25480
rect 69600 25088 70000 25144
rect 0 24864 400 24920
rect 69600 24528 70000 24584
rect 0 24304 400 24360
rect 69600 23968 70000 24024
rect 0 23744 400 23800
rect 69600 23408 70000 23464
rect 0 23184 400 23240
rect 69600 22848 70000 22904
rect 0 22624 400 22680
rect 69600 22288 70000 22344
rect 0 22064 400 22120
rect 69600 21728 70000 21784
rect 0 21504 400 21560
rect 69600 21168 70000 21224
rect 0 20944 400 21000
rect 69600 20608 70000 20664
rect 0 20384 400 20440
rect 69600 20048 70000 20104
rect 0 19824 400 19880
rect 69600 19488 70000 19544
rect 0 19264 400 19320
rect 69600 18928 70000 18984
rect 0 18704 400 18760
rect 69600 18368 70000 18424
rect 0 18144 400 18200
rect 69600 17808 70000 17864
rect 0 17584 400 17640
rect 69600 17248 70000 17304
rect 0 17024 400 17080
rect 69600 16688 70000 16744
rect 0 16464 400 16520
rect 69600 16128 70000 16184
rect 0 15904 400 15960
rect 69600 15568 70000 15624
rect 0 15344 400 15400
rect 69600 15008 70000 15064
rect 0 14784 400 14840
rect 69600 14448 70000 14504
rect 0 14224 400 14280
rect 69600 13888 70000 13944
rect 0 13664 400 13720
rect 69600 13328 70000 13384
rect 0 13104 400 13160
rect 69600 12768 70000 12824
rect 0 12544 400 12600
rect 69600 12208 70000 12264
rect 0 11984 400 12040
rect 69600 11648 70000 11704
rect 0 11424 400 11480
rect 69600 11088 70000 11144
rect 0 10864 400 10920
rect 69600 10528 70000 10584
rect 0 10304 400 10360
rect 69600 9968 70000 10024
rect 0 9744 400 9800
rect 69600 9408 70000 9464
rect 0 9184 400 9240
rect 69600 8848 70000 8904
rect 0 8624 400 8680
rect 69600 8288 70000 8344
rect 0 8064 400 8120
rect 69600 7728 70000 7784
rect 0 7504 400 7560
rect 69600 7168 70000 7224
rect 0 6944 400 7000
rect 69600 6608 70000 6664
rect 0 6384 400 6440
rect 69600 6048 70000 6104
rect 0 5824 400 5880
rect 69600 5488 70000 5544
rect 0 5264 400 5320
rect 69600 4928 70000 4984
rect 0 4704 400 4760
rect 69600 4368 70000 4424
rect 0 4144 400 4200
rect 69600 3808 70000 3864
rect 69600 3248 70000 3304
rect 69600 2688 70000 2744
rect 69600 2128 70000 2184
rect 69600 1568 70000 1624
<< obsm3 >>
rect 233 63254 69650 63434
rect 233 63138 69570 63254
rect 233 62694 69650 63138
rect 233 62578 69570 62694
rect 233 62134 69650 62578
rect 233 62018 69570 62134
rect 233 61574 69650 62018
rect 233 61458 69570 61574
rect 233 61014 69650 61458
rect 233 60898 69570 61014
rect 233 60790 69650 60898
rect 430 60674 69650 60790
rect 233 60454 69650 60674
rect 233 60338 69570 60454
rect 233 60230 69650 60338
rect 430 60114 69650 60230
rect 233 59894 69650 60114
rect 233 59778 69570 59894
rect 233 59670 69650 59778
rect 430 59554 69650 59670
rect 233 59334 69650 59554
rect 233 59218 69570 59334
rect 233 59110 69650 59218
rect 430 58994 69650 59110
rect 233 58774 69650 58994
rect 233 58658 69570 58774
rect 233 58550 69650 58658
rect 430 58434 69650 58550
rect 233 58214 69650 58434
rect 233 58098 69570 58214
rect 233 57990 69650 58098
rect 430 57874 69650 57990
rect 233 57654 69650 57874
rect 233 57538 69570 57654
rect 233 57430 69650 57538
rect 430 57314 69650 57430
rect 233 57094 69650 57314
rect 233 56978 69570 57094
rect 233 56870 69650 56978
rect 430 56754 69650 56870
rect 233 56534 69650 56754
rect 233 56418 69570 56534
rect 233 56310 69650 56418
rect 430 56194 69650 56310
rect 233 55974 69650 56194
rect 233 55858 69570 55974
rect 233 55750 69650 55858
rect 430 55634 69650 55750
rect 233 55414 69650 55634
rect 233 55298 69570 55414
rect 233 55190 69650 55298
rect 430 55074 69650 55190
rect 233 54854 69650 55074
rect 233 54738 69570 54854
rect 233 54630 69650 54738
rect 430 54514 69650 54630
rect 233 54294 69650 54514
rect 233 54178 69570 54294
rect 233 54070 69650 54178
rect 430 53954 69650 54070
rect 233 53734 69650 53954
rect 233 53618 69570 53734
rect 233 53510 69650 53618
rect 430 53394 69650 53510
rect 233 53174 69650 53394
rect 233 53058 69570 53174
rect 233 52950 69650 53058
rect 430 52834 69650 52950
rect 233 52614 69650 52834
rect 233 52498 69570 52614
rect 233 52390 69650 52498
rect 430 52274 69650 52390
rect 233 52054 69650 52274
rect 233 51938 69570 52054
rect 233 51830 69650 51938
rect 430 51714 69650 51830
rect 233 51494 69650 51714
rect 233 51378 69570 51494
rect 233 51270 69650 51378
rect 430 51154 69650 51270
rect 233 50934 69650 51154
rect 233 50818 69570 50934
rect 233 50710 69650 50818
rect 430 50594 69650 50710
rect 233 50374 69650 50594
rect 233 50258 69570 50374
rect 233 50150 69650 50258
rect 430 50034 69650 50150
rect 233 49814 69650 50034
rect 233 49698 69570 49814
rect 233 49590 69650 49698
rect 430 49474 69650 49590
rect 233 49254 69650 49474
rect 233 49138 69570 49254
rect 233 49030 69650 49138
rect 430 48914 69650 49030
rect 233 48694 69650 48914
rect 233 48578 69570 48694
rect 233 48470 69650 48578
rect 430 48354 69650 48470
rect 233 48134 69650 48354
rect 233 48018 69570 48134
rect 233 47910 69650 48018
rect 430 47794 69650 47910
rect 233 47574 69650 47794
rect 233 47458 69570 47574
rect 233 47350 69650 47458
rect 430 47234 69650 47350
rect 233 47014 69650 47234
rect 233 46898 69570 47014
rect 233 46790 69650 46898
rect 430 46674 69650 46790
rect 233 46454 69650 46674
rect 233 46338 69570 46454
rect 233 46230 69650 46338
rect 430 46114 69650 46230
rect 233 45894 69650 46114
rect 233 45778 69570 45894
rect 233 45670 69650 45778
rect 430 45554 69650 45670
rect 233 45334 69650 45554
rect 233 45218 69570 45334
rect 233 45110 69650 45218
rect 430 44994 69650 45110
rect 233 44774 69650 44994
rect 233 44658 69570 44774
rect 233 44550 69650 44658
rect 430 44434 69650 44550
rect 233 44214 69650 44434
rect 233 44098 69570 44214
rect 233 43990 69650 44098
rect 430 43874 69650 43990
rect 233 43654 69650 43874
rect 233 43538 69570 43654
rect 233 43430 69650 43538
rect 430 43314 69650 43430
rect 233 43094 69650 43314
rect 233 42978 69570 43094
rect 233 42870 69650 42978
rect 430 42754 69650 42870
rect 233 42534 69650 42754
rect 233 42418 69570 42534
rect 233 42310 69650 42418
rect 430 42194 69650 42310
rect 233 41974 69650 42194
rect 233 41858 69570 41974
rect 233 41750 69650 41858
rect 430 41634 69650 41750
rect 233 41414 69650 41634
rect 233 41298 69570 41414
rect 233 41190 69650 41298
rect 430 41074 69650 41190
rect 233 40854 69650 41074
rect 233 40738 69570 40854
rect 233 40630 69650 40738
rect 430 40514 69650 40630
rect 233 40294 69650 40514
rect 233 40178 69570 40294
rect 233 40070 69650 40178
rect 430 39954 69650 40070
rect 233 39734 69650 39954
rect 233 39618 69570 39734
rect 233 39510 69650 39618
rect 430 39394 69650 39510
rect 233 39174 69650 39394
rect 233 39058 69570 39174
rect 233 38950 69650 39058
rect 430 38834 69650 38950
rect 233 38614 69650 38834
rect 233 38498 69570 38614
rect 233 38390 69650 38498
rect 430 38274 69650 38390
rect 233 38054 69650 38274
rect 233 37938 69570 38054
rect 233 37830 69650 37938
rect 430 37714 69650 37830
rect 233 37494 69650 37714
rect 233 37378 69570 37494
rect 233 37270 69650 37378
rect 430 37154 69650 37270
rect 233 36934 69650 37154
rect 233 36818 69570 36934
rect 233 36710 69650 36818
rect 430 36594 69650 36710
rect 233 36374 69650 36594
rect 233 36258 69570 36374
rect 233 36150 69650 36258
rect 430 36034 69650 36150
rect 233 35814 69650 36034
rect 233 35698 69570 35814
rect 233 35590 69650 35698
rect 430 35474 69650 35590
rect 233 35254 69650 35474
rect 233 35138 69570 35254
rect 233 35030 69650 35138
rect 430 34914 69650 35030
rect 233 34694 69650 34914
rect 233 34578 69570 34694
rect 233 34470 69650 34578
rect 430 34354 69650 34470
rect 233 34134 69650 34354
rect 233 34018 69570 34134
rect 233 33910 69650 34018
rect 430 33794 69650 33910
rect 233 33574 69650 33794
rect 233 33458 69570 33574
rect 233 33350 69650 33458
rect 430 33234 69650 33350
rect 233 33014 69650 33234
rect 233 32898 69570 33014
rect 233 32790 69650 32898
rect 430 32674 69650 32790
rect 233 32454 69650 32674
rect 233 32338 69570 32454
rect 233 32230 69650 32338
rect 430 32114 69650 32230
rect 233 31894 69650 32114
rect 233 31778 69570 31894
rect 233 31670 69650 31778
rect 430 31554 69650 31670
rect 233 31334 69650 31554
rect 233 31218 69570 31334
rect 233 31110 69650 31218
rect 430 30994 69650 31110
rect 233 30774 69650 30994
rect 233 30658 69570 30774
rect 233 30550 69650 30658
rect 430 30434 69650 30550
rect 233 30214 69650 30434
rect 233 30098 69570 30214
rect 233 29990 69650 30098
rect 430 29874 69650 29990
rect 233 29654 69650 29874
rect 233 29538 69570 29654
rect 233 29430 69650 29538
rect 430 29314 69650 29430
rect 233 29094 69650 29314
rect 233 28978 69570 29094
rect 233 28870 69650 28978
rect 430 28754 69650 28870
rect 233 28534 69650 28754
rect 233 28418 69570 28534
rect 233 28310 69650 28418
rect 430 28194 69650 28310
rect 233 27974 69650 28194
rect 233 27858 69570 27974
rect 233 27750 69650 27858
rect 430 27634 69650 27750
rect 233 27414 69650 27634
rect 233 27298 69570 27414
rect 233 27190 69650 27298
rect 430 27074 69650 27190
rect 233 26854 69650 27074
rect 233 26738 69570 26854
rect 233 26630 69650 26738
rect 430 26514 69650 26630
rect 233 26294 69650 26514
rect 233 26178 69570 26294
rect 233 26070 69650 26178
rect 430 25954 69650 26070
rect 233 25734 69650 25954
rect 233 25618 69570 25734
rect 233 25510 69650 25618
rect 430 25394 69650 25510
rect 233 25174 69650 25394
rect 233 25058 69570 25174
rect 233 24950 69650 25058
rect 430 24834 69650 24950
rect 233 24614 69650 24834
rect 233 24498 69570 24614
rect 233 24390 69650 24498
rect 430 24274 69650 24390
rect 233 24054 69650 24274
rect 233 23938 69570 24054
rect 233 23830 69650 23938
rect 430 23714 69650 23830
rect 233 23494 69650 23714
rect 233 23378 69570 23494
rect 233 23270 69650 23378
rect 430 23154 69650 23270
rect 233 22934 69650 23154
rect 233 22818 69570 22934
rect 233 22710 69650 22818
rect 430 22594 69650 22710
rect 233 22374 69650 22594
rect 233 22258 69570 22374
rect 233 22150 69650 22258
rect 430 22034 69650 22150
rect 233 21814 69650 22034
rect 233 21698 69570 21814
rect 233 21590 69650 21698
rect 430 21474 69650 21590
rect 233 21254 69650 21474
rect 233 21138 69570 21254
rect 233 21030 69650 21138
rect 430 20914 69650 21030
rect 233 20694 69650 20914
rect 233 20578 69570 20694
rect 233 20470 69650 20578
rect 430 20354 69650 20470
rect 233 20134 69650 20354
rect 233 20018 69570 20134
rect 233 19910 69650 20018
rect 430 19794 69650 19910
rect 233 19574 69650 19794
rect 233 19458 69570 19574
rect 233 19350 69650 19458
rect 430 19234 69650 19350
rect 233 19014 69650 19234
rect 233 18898 69570 19014
rect 233 18790 69650 18898
rect 430 18674 69650 18790
rect 233 18454 69650 18674
rect 233 18338 69570 18454
rect 233 18230 69650 18338
rect 430 18114 69650 18230
rect 233 17894 69650 18114
rect 233 17778 69570 17894
rect 233 17670 69650 17778
rect 430 17554 69650 17670
rect 233 17334 69650 17554
rect 233 17218 69570 17334
rect 233 17110 69650 17218
rect 430 16994 69650 17110
rect 233 16774 69650 16994
rect 233 16658 69570 16774
rect 233 16550 69650 16658
rect 430 16434 69650 16550
rect 233 16214 69650 16434
rect 233 16098 69570 16214
rect 233 15990 69650 16098
rect 430 15874 69650 15990
rect 233 15654 69650 15874
rect 233 15538 69570 15654
rect 233 15430 69650 15538
rect 430 15314 69650 15430
rect 233 15094 69650 15314
rect 233 14978 69570 15094
rect 233 14870 69650 14978
rect 430 14754 69650 14870
rect 233 14534 69650 14754
rect 233 14418 69570 14534
rect 233 14310 69650 14418
rect 430 14194 69650 14310
rect 233 13974 69650 14194
rect 233 13858 69570 13974
rect 233 13750 69650 13858
rect 430 13634 69650 13750
rect 233 13414 69650 13634
rect 233 13298 69570 13414
rect 233 13190 69650 13298
rect 430 13074 69650 13190
rect 233 12854 69650 13074
rect 233 12738 69570 12854
rect 233 12630 69650 12738
rect 430 12514 69650 12630
rect 233 12294 69650 12514
rect 233 12178 69570 12294
rect 233 12070 69650 12178
rect 430 11954 69650 12070
rect 233 11734 69650 11954
rect 233 11618 69570 11734
rect 233 11510 69650 11618
rect 430 11394 69650 11510
rect 233 11174 69650 11394
rect 233 11058 69570 11174
rect 233 10950 69650 11058
rect 430 10834 69650 10950
rect 233 10614 69650 10834
rect 233 10498 69570 10614
rect 233 10390 69650 10498
rect 430 10274 69650 10390
rect 233 10054 69650 10274
rect 233 9938 69570 10054
rect 233 9830 69650 9938
rect 430 9714 69650 9830
rect 233 9494 69650 9714
rect 233 9378 69570 9494
rect 233 9270 69650 9378
rect 430 9154 69650 9270
rect 233 8934 69650 9154
rect 233 8818 69570 8934
rect 233 8710 69650 8818
rect 430 8594 69650 8710
rect 233 8374 69650 8594
rect 233 8258 69570 8374
rect 233 8150 69650 8258
rect 430 8034 69650 8150
rect 233 7814 69650 8034
rect 233 7698 69570 7814
rect 233 7590 69650 7698
rect 430 7474 69650 7590
rect 233 7254 69650 7474
rect 233 7138 69570 7254
rect 233 7030 69650 7138
rect 430 6914 69650 7030
rect 233 6694 69650 6914
rect 233 6578 69570 6694
rect 233 6470 69650 6578
rect 430 6354 69650 6470
rect 233 6134 69650 6354
rect 233 6018 69570 6134
rect 233 5910 69650 6018
rect 430 5794 69650 5910
rect 233 5574 69650 5794
rect 233 5458 69570 5574
rect 233 5350 69650 5458
rect 430 5234 69650 5350
rect 233 5014 69650 5234
rect 233 4898 69570 5014
rect 233 4790 69650 4898
rect 430 4674 69650 4790
rect 233 4454 69650 4674
rect 233 4338 69570 4454
rect 233 4230 69650 4338
rect 430 4114 69650 4230
rect 233 3894 69650 4114
rect 233 3778 69570 3894
rect 233 3334 69650 3778
rect 233 3218 69570 3334
rect 233 2774 69650 3218
rect 233 2658 69570 2774
rect 233 2214 69650 2658
rect 233 2098 69570 2214
rect 233 1654 69650 2098
rect 233 1538 69570 1654
rect 233 798 69650 1538
<< metal4 >>
rect 2224 1538 2384 63142
rect 9904 1538 10064 63142
rect 17584 1538 17744 63142
rect 25264 1538 25424 63142
rect 32944 1538 33104 63142
rect 40624 1538 40784 63142
rect 48304 1538 48464 63142
rect 55984 1538 56144 63142
rect 63664 1538 63824 63142
<< obsm4 >>
rect 1022 1801 2194 62879
rect 2414 1801 9874 62879
rect 10094 1801 17554 62879
rect 17774 1801 25234 62879
rect 25454 1801 32914 62879
rect 33134 1801 40594 62879
rect 40814 1801 48274 62879
rect 48494 1801 55954 62879
rect 56174 1801 63634 62879
rect 63854 1801 68082 62879
<< labels >>
rlabel metal2 s 28000 64600 28056 65000 6 ay8913_do[0]
port 1 nsew signal input
rlabel metal2 s 32480 64600 32536 65000 6 ay8913_do[10]
port 2 nsew signal input
rlabel metal2 s 32928 64600 32984 65000 6 ay8913_do[11]
port 3 nsew signal input
rlabel metal2 s 33376 64600 33432 65000 6 ay8913_do[12]
port 4 nsew signal input
rlabel metal2 s 33824 64600 33880 65000 6 ay8913_do[13]
port 5 nsew signal input
rlabel metal2 s 34272 64600 34328 65000 6 ay8913_do[14]
port 6 nsew signal input
rlabel metal2 s 34720 64600 34776 65000 6 ay8913_do[15]
port 7 nsew signal input
rlabel metal2 s 35168 64600 35224 65000 6 ay8913_do[16]
port 8 nsew signal input
rlabel metal2 s 35616 64600 35672 65000 6 ay8913_do[17]
port 9 nsew signal input
rlabel metal2 s 36064 64600 36120 65000 6 ay8913_do[18]
port 10 nsew signal input
rlabel metal2 s 36512 64600 36568 65000 6 ay8913_do[19]
port 11 nsew signal input
rlabel metal2 s 28448 64600 28504 65000 6 ay8913_do[1]
port 12 nsew signal input
rlabel metal2 s 36960 64600 37016 65000 6 ay8913_do[20]
port 13 nsew signal input
rlabel metal2 s 37408 64600 37464 65000 6 ay8913_do[21]
port 14 nsew signal input
rlabel metal2 s 37856 64600 37912 65000 6 ay8913_do[22]
port 15 nsew signal input
rlabel metal2 s 38304 64600 38360 65000 6 ay8913_do[23]
port 16 nsew signal input
rlabel metal2 s 38752 64600 38808 65000 6 ay8913_do[24]
port 17 nsew signal input
rlabel metal2 s 39200 64600 39256 65000 6 ay8913_do[25]
port 18 nsew signal input
rlabel metal2 s 39648 64600 39704 65000 6 ay8913_do[26]
port 19 nsew signal input
rlabel metal2 s 40096 64600 40152 65000 6 ay8913_do[27]
port 20 nsew signal input
rlabel metal2 s 28896 64600 28952 65000 6 ay8913_do[2]
port 21 nsew signal input
rlabel metal2 s 29344 64600 29400 65000 6 ay8913_do[3]
port 22 nsew signal input
rlabel metal2 s 29792 64600 29848 65000 6 ay8913_do[4]
port 23 nsew signal input
rlabel metal2 s 30240 64600 30296 65000 6 ay8913_do[5]
port 24 nsew signal input
rlabel metal2 s 30688 64600 30744 65000 6 ay8913_do[6]
port 25 nsew signal input
rlabel metal2 s 31136 64600 31192 65000 6 ay8913_do[7]
port 26 nsew signal input
rlabel metal2 s 31584 64600 31640 65000 6 ay8913_do[8]
port 27 nsew signal input
rlabel metal2 s 32032 64600 32088 65000 6 ay8913_do[9]
port 28 nsew signal input
rlabel metal2 s 19488 64600 19544 65000 6 blinker_do[0]
port 29 nsew signal input
rlabel metal2 s 19936 64600 19992 65000 6 blinker_do[1]
port 30 nsew signal input
rlabel metal2 s 20384 64600 20440 65000 6 blinker_do[2]
port 31 nsew signal input
rlabel metal3 s 69600 21728 70000 21784 6 custom_settings[0]
port 32 nsew signal output
rlabel metal3 s 69600 27328 70000 27384 6 custom_settings[10]
port 33 nsew signal output
rlabel metal3 s 69600 27888 70000 27944 6 custom_settings[11]
port 34 nsew signal output
rlabel metal3 s 69600 28448 70000 28504 6 custom_settings[12]
port 35 nsew signal output
rlabel metal3 s 69600 29008 70000 29064 6 custom_settings[13]
port 36 nsew signal output
rlabel metal3 s 69600 29568 70000 29624 6 custom_settings[14]
port 37 nsew signal output
rlabel metal3 s 69600 30128 70000 30184 6 custom_settings[15]
port 38 nsew signal output
rlabel metal3 s 69600 30688 70000 30744 6 custom_settings[16]
port 39 nsew signal output
rlabel metal3 s 69600 31248 70000 31304 6 custom_settings[17]
port 40 nsew signal output
rlabel metal3 s 69600 31808 70000 31864 6 custom_settings[18]
port 41 nsew signal output
rlabel metal3 s 69600 32368 70000 32424 6 custom_settings[19]
port 42 nsew signal output
rlabel metal3 s 69600 22288 70000 22344 6 custom_settings[1]
port 43 nsew signal output
rlabel metal3 s 69600 32928 70000 32984 6 custom_settings[20]
port 44 nsew signal output
rlabel metal3 s 69600 33488 70000 33544 6 custom_settings[21]
port 45 nsew signal output
rlabel metal3 s 69600 34048 70000 34104 6 custom_settings[22]
port 46 nsew signal output
rlabel metal3 s 69600 34608 70000 34664 6 custom_settings[23]
port 47 nsew signal output
rlabel metal3 s 69600 35168 70000 35224 6 custom_settings[24]
port 48 nsew signal output
rlabel metal3 s 69600 35728 70000 35784 6 custom_settings[25]
port 49 nsew signal output
rlabel metal3 s 69600 36288 70000 36344 6 custom_settings[26]
port 50 nsew signal output
rlabel metal3 s 69600 36848 70000 36904 6 custom_settings[27]
port 51 nsew signal output
rlabel metal3 s 69600 37408 70000 37464 6 custom_settings[28]
port 52 nsew signal output
rlabel metal3 s 69600 37968 70000 38024 6 custom_settings[29]
port 53 nsew signal output
rlabel metal3 s 69600 22848 70000 22904 6 custom_settings[2]
port 54 nsew signal output
rlabel metal3 s 69600 38528 70000 38584 6 custom_settings[30]
port 55 nsew signal output
rlabel metal3 s 69600 39088 70000 39144 6 custom_settings[31]
port 56 nsew signal output
rlabel metal3 s 69600 23408 70000 23464 6 custom_settings[3]
port 57 nsew signal output
rlabel metal3 s 69600 23968 70000 24024 6 custom_settings[4]
port 58 nsew signal output
rlabel metal3 s 69600 24528 70000 24584 6 custom_settings[5]
port 59 nsew signal output
rlabel metal3 s 69600 25088 70000 25144 6 custom_settings[6]
port 60 nsew signal output
rlabel metal3 s 69600 25648 70000 25704 6 custom_settings[7]
port 61 nsew signal output
rlabel metal3 s 69600 26208 70000 26264 6 custom_settings[8]
port 62 nsew signal output
rlabel metal3 s 69600 26768 70000 26824 6 custom_settings[9]
port 63 nsew signal output
rlabel metal3 s 0 57344 400 57400 6 hellorld_do
port 64 nsew signal input
rlabel metal2 s 224 64600 280 65000 6 io_in_0
port 65 nsew signal input
rlabel metal3 s 0 4144 400 4200 6 io_oeb[0]
port 66 nsew signal output
rlabel metal3 s 0 9744 400 9800 6 io_oeb[10]
port 67 nsew signal output
rlabel metal3 s 0 10304 400 10360 6 io_oeb[11]
port 68 nsew signal output
rlabel metal3 s 0 10864 400 10920 6 io_oeb[12]
port 69 nsew signal output
rlabel metal3 s 0 11424 400 11480 6 io_oeb[13]
port 70 nsew signal output
rlabel metal3 s 0 11984 400 12040 6 io_oeb[14]
port 71 nsew signal output
rlabel metal3 s 0 12544 400 12600 6 io_oeb[15]
port 72 nsew signal output
rlabel metal3 s 0 13104 400 13160 6 io_oeb[16]
port 73 nsew signal output
rlabel metal3 s 0 13664 400 13720 6 io_oeb[17]
port 74 nsew signal output
rlabel metal3 s 0 14224 400 14280 6 io_oeb[18]
port 75 nsew signal output
rlabel metal3 s 0 14784 400 14840 6 io_oeb[19]
port 76 nsew signal output
rlabel metal3 s 0 4704 400 4760 6 io_oeb[1]
port 77 nsew signal output
rlabel metal3 s 0 15344 400 15400 6 io_oeb[20]
port 78 nsew signal output
rlabel metal3 s 0 15904 400 15960 6 io_oeb[21]
port 79 nsew signal output
rlabel metal3 s 0 16464 400 16520 6 io_oeb[22]
port 80 nsew signal output
rlabel metal3 s 0 17024 400 17080 6 io_oeb[23]
port 81 nsew signal output
rlabel metal3 s 0 17584 400 17640 6 io_oeb[24]
port 82 nsew signal output
rlabel metal3 s 0 18144 400 18200 6 io_oeb[25]
port 83 nsew signal output
rlabel metal3 s 0 18704 400 18760 6 io_oeb[26]
port 84 nsew signal output
rlabel metal3 s 0 19264 400 19320 6 io_oeb[27]
port 85 nsew signal output
rlabel metal3 s 0 19824 400 19880 6 io_oeb[28]
port 86 nsew signal output
rlabel metal3 s 0 20384 400 20440 6 io_oeb[29]
port 87 nsew signal output
rlabel metal3 s 0 5264 400 5320 6 io_oeb[2]
port 88 nsew signal output
rlabel metal3 s 0 20944 400 21000 6 io_oeb[30]
port 89 nsew signal output
rlabel metal3 s 0 21504 400 21560 6 io_oeb[31]
port 90 nsew signal output
rlabel metal3 s 0 22064 400 22120 6 io_oeb[32]
port 91 nsew signal output
rlabel metal3 s 0 22624 400 22680 6 io_oeb[33]
port 92 nsew signal output
rlabel metal3 s 0 23184 400 23240 6 io_oeb[34]
port 93 nsew signal output
rlabel metal3 s 0 23744 400 23800 6 io_oeb[35]
port 94 nsew signal output
rlabel metal3 s 0 24304 400 24360 6 io_oeb[36]
port 95 nsew signal output
rlabel metal3 s 0 24864 400 24920 6 io_oeb[37]
port 96 nsew signal output
rlabel metal3 s 0 5824 400 5880 6 io_oeb[3]
port 97 nsew signal output
rlabel metal3 s 0 6384 400 6440 6 io_oeb[4]
port 98 nsew signal output
rlabel metal3 s 0 6944 400 7000 6 io_oeb[5]
port 99 nsew signal output
rlabel metal3 s 0 7504 400 7560 6 io_oeb[6]
port 100 nsew signal output
rlabel metal3 s 0 8064 400 8120 6 io_oeb[7]
port 101 nsew signal output
rlabel metal3 s 0 8624 400 8680 6 io_oeb[8]
port 102 nsew signal output
rlabel metal3 s 0 9184 400 9240 6 io_oeb[9]
port 103 nsew signal output
rlabel metal2 s 672 64600 728 65000 6 io_out[0]
port 104 nsew signal output
rlabel metal2 s 5152 64600 5208 65000 6 io_out[10]
port 105 nsew signal output
rlabel metal2 s 5600 64600 5656 65000 6 io_out[11]
port 106 nsew signal output
rlabel metal2 s 6048 64600 6104 65000 6 io_out[12]
port 107 nsew signal output
rlabel metal2 s 6496 64600 6552 65000 6 io_out[13]
port 108 nsew signal output
rlabel metal2 s 6944 64600 7000 65000 6 io_out[14]
port 109 nsew signal output
rlabel metal2 s 7392 64600 7448 65000 6 io_out[15]
port 110 nsew signal output
rlabel metal2 s 7840 64600 7896 65000 6 io_out[16]
port 111 nsew signal output
rlabel metal2 s 8288 64600 8344 65000 6 io_out[17]
port 112 nsew signal output
rlabel metal2 s 8736 64600 8792 65000 6 io_out[18]
port 113 nsew signal output
rlabel metal2 s 9184 64600 9240 65000 6 io_out[19]
port 114 nsew signal output
rlabel metal2 s 1120 64600 1176 65000 6 io_out[1]
port 115 nsew signal output
rlabel metal2 s 9632 64600 9688 65000 6 io_out[20]
port 116 nsew signal output
rlabel metal2 s 10080 64600 10136 65000 6 io_out[21]
port 117 nsew signal output
rlabel metal2 s 10528 64600 10584 65000 6 io_out[22]
port 118 nsew signal output
rlabel metal2 s 10976 64600 11032 65000 6 io_out[23]
port 119 nsew signal output
rlabel metal2 s 11424 64600 11480 65000 6 io_out[24]
port 120 nsew signal output
rlabel metal2 s 11872 64600 11928 65000 6 io_out[25]
port 121 nsew signal output
rlabel metal2 s 12320 64600 12376 65000 6 io_out[26]
port 122 nsew signal output
rlabel metal2 s 12768 64600 12824 65000 6 io_out[27]
port 123 nsew signal output
rlabel metal2 s 13216 64600 13272 65000 6 io_out[28]
port 124 nsew signal output
rlabel metal2 s 13664 64600 13720 65000 6 io_out[29]
port 125 nsew signal output
rlabel metal2 s 1568 64600 1624 65000 6 io_out[2]
port 126 nsew signal output
rlabel metal2 s 14112 64600 14168 65000 6 io_out[30]
port 127 nsew signal output
rlabel metal2 s 14560 64600 14616 65000 6 io_out[31]
port 128 nsew signal output
rlabel metal2 s 15008 64600 15064 65000 6 io_out[32]
port 129 nsew signal output
rlabel metal2 s 15456 64600 15512 65000 6 io_out[33]
port 130 nsew signal output
rlabel metal2 s 15904 64600 15960 65000 6 io_out[34]
port 131 nsew signal output
rlabel metal2 s 16352 64600 16408 65000 6 io_out[35]
port 132 nsew signal output
rlabel metal2 s 16800 64600 16856 65000 6 io_out[36]
port 133 nsew signal output
rlabel metal2 s 17248 64600 17304 65000 6 io_out[37]
port 134 nsew signal output
rlabel metal2 s 2016 64600 2072 65000 6 io_out[3]
port 135 nsew signal output
rlabel metal2 s 2464 64600 2520 65000 6 io_out[4]
port 136 nsew signal output
rlabel metal2 s 2912 64600 2968 65000 6 io_out[5]
port 137 nsew signal output
rlabel metal2 s 3360 64600 3416 65000 6 io_out[6]
port 138 nsew signal output
rlabel metal2 s 3808 64600 3864 65000 6 io_out[7]
port 139 nsew signal output
rlabel metal2 s 4256 64600 4312 65000 6 io_out[8]
port 140 nsew signal output
rlabel metal2 s 4704 64600 4760 65000 6 io_out[9]
port 141 nsew signal output
rlabel metal2 s 17696 64600 17752 65000 6 irq[0]
port 142 nsew signal output
rlabel metal2 s 18144 64600 18200 65000 6 irq[1]
port 143 nsew signal output
rlabel metal2 s 18592 64600 18648 65000 6 irq[2]
port 144 nsew signal output
rlabel metal3 s 0 39424 400 39480 6 mc14500_do[0]
port 145 nsew signal input
rlabel metal3 s 0 45024 400 45080 6 mc14500_do[10]
port 146 nsew signal input
rlabel metal3 s 0 45584 400 45640 6 mc14500_do[11]
port 147 nsew signal input
rlabel metal3 s 0 46144 400 46200 6 mc14500_do[12]
port 148 nsew signal input
rlabel metal3 s 0 46704 400 46760 6 mc14500_do[13]
port 149 nsew signal input
rlabel metal3 s 0 47264 400 47320 6 mc14500_do[14]
port 150 nsew signal input
rlabel metal3 s 0 47824 400 47880 6 mc14500_do[15]
port 151 nsew signal input
rlabel metal3 s 0 48384 400 48440 6 mc14500_do[16]
port 152 nsew signal input
rlabel metal3 s 0 48944 400 49000 6 mc14500_do[17]
port 153 nsew signal input
rlabel metal3 s 0 49504 400 49560 6 mc14500_do[18]
port 154 nsew signal input
rlabel metal3 s 0 50064 400 50120 6 mc14500_do[19]
port 155 nsew signal input
rlabel metal3 s 0 39984 400 40040 6 mc14500_do[1]
port 156 nsew signal input
rlabel metal3 s 0 50624 400 50680 6 mc14500_do[20]
port 157 nsew signal input
rlabel metal3 s 0 51184 400 51240 6 mc14500_do[21]
port 158 nsew signal input
rlabel metal3 s 0 51744 400 51800 6 mc14500_do[22]
port 159 nsew signal input
rlabel metal3 s 0 52304 400 52360 6 mc14500_do[23]
port 160 nsew signal input
rlabel metal3 s 0 52864 400 52920 6 mc14500_do[24]
port 161 nsew signal input
rlabel metal3 s 0 53424 400 53480 6 mc14500_do[25]
port 162 nsew signal input
rlabel metal3 s 0 53984 400 54040 6 mc14500_do[26]
port 163 nsew signal input
rlabel metal3 s 0 54544 400 54600 6 mc14500_do[27]
port 164 nsew signal input
rlabel metal3 s 0 55104 400 55160 6 mc14500_do[28]
port 165 nsew signal input
rlabel metal3 s 0 55664 400 55720 6 mc14500_do[29]
port 166 nsew signal input
rlabel metal3 s 0 40544 400 40600 6 mc14500_do[2]
port 167 nsew signal input
rlabel metal3 s 0 56224 400 56280 6 mc14500_do[30]
port 168 nsew signal input
rlabel metal3 s 0 41104 400 41160 6 mc14500_do[3]
port 169 nsew signal input
rlabel metal3 s 0 41664 400 41720 6 mc14500_do[4]
port 170 nsew signal input
rlabel metal3 s 0 42224 400 42280 6 mc14500_do[5]
port 171 nsew signal input
rlabel metal3 s 0 42784 400 42840 6 mc14500_do[6]
port 172 nsew signal input
rlabel metal3 s 0 43344 400 43400 6 mc14500_do[7]
port 173 nsew signal input
rlabel metal3 s 0 43904 400 43960 6 mc14500_do[8]
port 174 nsew signal input
rlabel metal3 s 0 44464 400 44520 6 mc14500_do[9]
port 175 nsew signal input
rlabel metal2 s 21280 64600 21336 65000 6 mc14500_sram_addr[0]
port 176 nsew signal input
rlabel metal2 s 21728 64600 21784 65000 6 mc14500_sram_addr[1]
port 177 nsew signal input
rlabel metal2 s 22176 64600 22232 65000 6 mc14500_sram_addr[2]
port 178 nsew signal input
rlabel metal2 s 22624 64600 22680 65000 6 mc14500_sram_addr[3]
port 179 nsew signal input
rlabel metal2 s 23072 64600 23128 65000 6 mc14500_sram_addr[4]
port 180 nsew signal input
rlabel metal2 s 23520 64600 23576 65000 6 mc14500_sram_addr[5]
port 181 nsew signal input
rlabel metal2 s 27552 64600 27608 65000 6 mc14500_sram_gwe
port 182 nsew signal input
rlabel metal2 s 23968 64600 24024 65000 6 mc14500_sram_in[0]
port 183 nsew signal input
rlabel metal2 s 24416 64600 24472 65000 6 mc14500_sram_in[1]
port 184 nsew signal input
rlabel metal2 s 24864 64600 24920 65000 6 mc14500_sram_in[2]
port 185 nsew signal input
rlabel metal2 s 25312 64600 25368 65000 6 mc14500_sram_in[3]
port 186 nsew signal input
rlabel metal2 s 25760 64600 25816 65000 6 mc14500_sram_in[4]
port 187 nsew signal input
rlabel metal2 s 26208 64600 26264 65000 6 mc14500_sram_in[5]
port 188 nsew signal input
rlabel metal2 s 26656 64600 26712 65000 6 mc14500_sram_in[6]
port 189 nsew signal input
rlabel metal2 s 27104 64600 27160 65000 6 mc14500_sram_in[7]
port 190 nsew signal input
rlabel metal2 s 40544 64600 40600 65000 6 pdp11_do[0]
port 191 nsew signal input
rlabel metal2 s 49504 64600 49560 65000 6 pdp11_do[10]
port 192 nsew signal input
rlabel metal2 s 50400 64600 50456 65000 6 pdp11_do[11]
port 193 nsew signal input
rlabel metal2 s 51296 64600 51352 65000 6 pdp11_do[12]
port 194 nsew signal input
rlabel metal2 s 52192 64600 52248 65000 6 pdp11_do[13]
port 195 nsew signal input
rlabel metal2 s 53088 64600 53144 65000 6 pdp11_do[14]
port 196 nsew signal input
rlabel metal2 s 53984 64600 54040 65000 6 pdp11_do[15]
port 197 nsew signal input
rlabel metal2 s 54880 64600 54936 65000 6 pdp11_do[16]
port 198 nsew signal input
rlabel metal2 s 55776 64600 55832 65000 6 pdp11_do[17]
port 199 nsew signal input
rlabel metal2 s 56672 64600 56728 65000 6 pdp11_do[18]
port 200 nsew signal input
rlabel metal2 s 57568 64600 57624 65000 6 pdp11_do[19]
port 201 nsew signal input
rlabel metal2 s 41440 64600 41496 65000 6 pdp11_do[1]
port 202 nsew signal input
rlabel metal2 s 58464 64600 58520 65000 6 pdp11_do[20]
port 203 nsew signal input
rlabel metal2 s 59360 64600 59416 65000 6 pdp11_do[21]
port 204 nsew signal input
rlabel metal2 s 60256 64600 60312 65000 6 pdp11_do[22]
port 205 nsew signal input
rlabel metal2 s 61152 64600 61208 65000 6 pdp11_do[23]
port 206 nsew signal input
rlabel metal2 s 62048 64600 62104 65000 6 pdp11_do[24]
port 207 nsew signal input
rlabel metal2 s 62944 64600 63000 65000 6 pdp11_do[25]
port 208 nsew signal input
rlabel metal2 s 63840 64600 63896 65000 6 pdp11_do[26]
port 209 nsew signal input
rlabel metal2 s 64736 64600 64792 65000 6 pdp11_do[27]
port 210 nsew signal input
rlabel metal2 s 65632 64600 65688 65000 6 pdp11_do[28]
port 211 nsew signal input
rlabel metal2 s 66528 64600 66584 65000 6 pdp11_do[29]
port 212 nsew signal input
rlabel metal2 s 42336 64600 42392 65000 6 pdp11_do[2]
port 213 nsew signal input
rlabel metal2 s 67424 64600 67480 65000 6 pdp11_do[30]
port 214 nsew signal input
rlabel metal2 s 68320 64600 68376 65000 6 pdp11_do[31]
port 215 nsew signal input
rlabel metal2 s 69216 64600 69272 65000 6 pdp11_do[32]
port 216 nsew signal input
rlabel metal2 s 43232 64600 43288 65000 6 pdp11_do[3]
port 217 nsew signal input
rlabel metal2 s 44128 64600 44184 65000 6 pdp11_do[4]
port 218 nsew signal input
rlabel metal2 s 45024 64600 45080 65000 6 pdp11_do[5]
port 219 nsew signal input
rlabel metal2 s 45920 64600 45976 65000 6 pdp11_do[6]
port 220 nsew signal input
rlabel metal2 s 46816 64600 46872 65000 6 pdp11_do[7]
port 221 nsew signal input
rlabel metal2 s 47712 64600 47768 65000 6 pdp11_do[8]
port 222 nsew signal input
rlabel metal2 s 48608 64600 48664 65000 6 pdp11_do[9]
port 223 nsew signal input
rlabel metal2 s 40992 64600 41048 65000 6 pdp11_oeb[0]
port 224 nsew signal input
rlabel metal2 s 49952 64600 50008 65000 6 pdp11_oeb[10]
port 225 nsew signal input
rlabel metal2 s 50848 64600 50904 65000 6 pdp11_oeb[11]
port 226 nsew signal input
rlabel metal2 s 51744 64600 51800 65000 6 pdp11_oeb[12]
port 227 nsew signal input
rlabel metal2 s 52640 64600 52696 65000 6 pdp11_oeb[13]
port 228 nsew signal input
rlabel metal2 s 53536 64600 53592 65000 6 pdp11_oeb[14]
port 229 nsew signal input
rlabel metal2 s 54432 64600 54488 65000 6 pdp11_oeb[15]
port 230 nsew signal input
rlabel metal2 s 55328 64600 55384 65000 6 pdp11_oeb[16]
port 231 nsew signal input
rlabel metal2 s 56224 64600 56280 65000 6 pdp11_oeb[17]
port 232 nsew signal input
rlabel metal2 s 57120 64600 57176 65000 6 pdp11_oeb[18]
port 233 nsew signal input
rlabel metal2 s 58016 64600 58072 65000 6 pdp11_oeb[19]
port 234 nsew signal input
rlabel metal2 s 41888 64600 41944 65000 6 pdp11_oeb[1]
port 235 nsew signal input
rlabel metal2 s 58912 64600 58968 65000 6 pdp11_oeb[20]
port 236 nsew signal input
rlabel metal2 s 59808 64600 59864 65000 6 pdp11_oeb[21]
port 237 nsew signal input
rlabel metal2 s 60704 64600 60760 65000 6 pdp11_oeb[22]
port 238 nsew signal input
rlabel metal2 s 61600 64600 61656 65000 6 pdp11_oeb[23]
port 239 nsew signal input
rlabel metal2 s 62496 64600 62552 65000 6 pdp11_oeb[24]
port 240 nsew signal input
rlabel metal2 s 63392 64600 63448 65000 6 pdp11_oeb[25]
port 241 nsew signal input
rlabel metal2 s 64288 64600 64344 65000 6 pdp11_oeb[26]
port 242 nsew signal input
rlabel metal2 s 65184 64600 65240 65000 6 pdp11_oeb[27]
port 243 nsew signal input
rlabel metal2 s 66080 64600 66136 65000 6 pdp11_oeb[28]
port 244 nsew signal input
rlabel metal2 s 66976 64600 67032 65000 6 pdp11_oeb[29]
port 245 nsew signal input
rlabel metal2 s 42784 64600 42840 65000 6 pdp11_oeb[2]
port 246 nsew signal input
rlabel metal2 s 67872 64600 67928 65000 6 pdp11_oeb[30]
port 247 nsew signal input
rlabel metal2 s 68768 64600 68824 65000 6 pdp11_oeb[31]
port 248 nsew signal input
rlabel metal2 s 69664 64600 69720 65000 6 pdp11_oeb[32]
port 249 nsew signal input
rlabel metal2 s 43680 64600 43736 65000 6 pdp11_oeb[3]
port 250 nsew signal input
rlabel metal2 s 44576 64600 44632 65000 6 pdp11_oeb[4]
port 251 nsew signal input
rlabel metal2 s 45472 64600 45528 65000 6 pdp11_oeb[5]
port 252 nsew signal input
rlabel metal2 s 46368 64600 46424 65000 6 pdp11_oeb[6]
port 253 nsew signal input
rlabel metal2 s 47264 64600 47320 65000 6 pdp11_oeb[7]
port 254 nsew signal input
rlabel metal2 s 48160 64600 48216 65000 6 pdp11_oeb[8]
port 255 nsew signal input
rlabel metal2 s 49056 64600 49112 65000 6 pdp11_oeb[9]
port 256 nsew signal input
rlabel metal2 s 45472 0 45528 400 6 qcpu_do[0]
port 257 nsew signal input
rlabel metal2 s 49952 0 50008 400 6 qcpu_do[10]
port 258 nsew signal input
rlabel metal2 s 50400 0 50456 400 6 qcpu_do[11]
port 259 nsew signal input
rlabel metal2 s 50848 0 50904 400 6 qcpu_do[12]
port 260 nsew signal input
rlabel metal2 s 51296 0 51352 400 6 qcpu_do[13]
port 261 nsew signal input
rlabel metal2 s 51744 0 51800 400 6 qcpu_do[14]
port 262 nsew signal input
rlabel metal2 s 52192 0 52248 400 6 qcpu_do[15]
port 263 nsew signal input
rlabel metal2 s 52640 0 52696 400 6 qcpu_do[16]
port 264 nsew signal input
rlabel metal2 s 53088 0 53144 400 6 qcpu_do[17]
port 265 nsew signal input
rlabel metal2 s 53536 0 53592 400 6 qcpu_do[18]
port 266 nsew signal input
rlabel metal2 s 53984 0 54040 400 6 qcpu_do[19]
port 267 nsew signal input
rlabel metal2 s 45920 0 45976 400 6 qcpu_do[1]
port 268 nsew signal input
rlabel metal2 s 54432 0 54488 400 6 qcpu_do[20]
port 269 nsew signal input
rlabel metal2 s 54880 0 54936 400 6 qcpu_do[21]
port 270 nsew signal input
rlabel metal2 s 55328 0 55384 400 6 qcpu_do[22]
port 271 nsew signal input
rlabel metal2 s 55776 0 55832 400 6 qcpu_do[23]
port 272 nsew signal input
rlabel metal2 s 56224 0 56280 400 6 qcpu_do[24]
port 273 nsew signal input
rlabel metal2 s 56672 0 56728 400 6 qcpu_do[25]
port 274 nsew signal input
rlabel metal2 s 57120 0 57176 400 6 qcpu_do[26]
port 275 nsew signal input
rlabel metal2 s 57568 0 57624 400 6 qcpu_do[27]
port 276 nsew signal input
rlabel metal2 s 58016 0 58072 400 6 qcpu_do[28]
port 277 nsew signal input
rlabel metal2 s 58464 0 58520 400 6 qcpu_do[29]
port 278 nsew signal input
rlabel metal2 s 46368 0 46424 400 6 qcpu_do[2]
port 279 nsew signal input
rlabel metal2 s 58912 0 58968 400 6 qcpu_do[30]
port 280 nsew signal input
rlabel metal2 s 59360 0 59416 400 6 qcpu_do[31]
port 281 nsew signal input
rlabel metal2 s 59808 0 59864 400 6 qcpu_do[32]
port 282 nsew signal input
rlabel metal2 s 46816 0 46872 400 6 qcpu_do[3]
port 283 nsew signal input
rlabel metal2 s 47264 0 47320 400 6 qcpu_do[4]
port 284 nsew signal input
rlabel metal2 s 47712 0 47768 400 6 qcpu_do[5]
port 285 nsew signal input
rlabel metal2 s 48160 0 48216 400 6 qcpu_do[6]
port 286 nsew signal input
rlabel metal2 s 48608 0 48664 400 6 qcpu_do[7]
port 287 nsew signal input
rlabel metal2 s 49056 0 49112 400 6 qcpu_do[8]
port 288 nsew signal input
rlabel metal2 s 49504 0 49560 400 6 qcpu_do[9]
port 289 nsew signal input
rlabel metal3 s 69600 39648 70000 39704 6 qcpu_oeb[0]
port 290 nsew signal input
rlabel metal3 s 69600 45248 70000 45304 6 qcpu_oeb[10]
port 291 nsew signal input
rlabel metal3 s 69600 45808 70000 45864 6 qcpu_oeb[11]
port 292 nsew signal input
rlabel metal3 s 69600 46368 70000 46424 6 qcpu_oeb[12]
port 293 nsew signal input
rlabel metal3 s 69600 46928 70000 46984 6 qcpu_oeb[13]
port 294 nsew signal input
rlabel metal3 s 69600 47488 70000 47544 6 qcpu_oeb[14]
port 295 nsew signal input
rlabel metal3 s 69600 48048 70000 48104 6 qcpu_oeb[15]
port 296 nsew signal input
rlabel metal3 s 69600 48608 70000 48664 6 qcpu_oeb[16]
port 297 nsew signal input
rlabel metal3 s 69600 49168 70000 49224 6 qcpu_oeb[17]
port 298 nsew signal input
rlabel metal3 s 69600 49728 70000 49784 6 qcpu_oeb[18]
port 299 nsew signal input
rlabel metal3 s 69600 50288 70000 50344 6 qcpu_oeb[19]
port 300 nsew signal input
rlabel metal3 s 69600 40208 70000 40264 6 qcpu_oeb[1]
port 301 nsew signal input
rlabel metal3 s 69600 50848 70000 50904 6 qcpu_oeb[20]
port 302 nsew signal input
rlabel metal3 s 69600 51408 70000 51464 6 qcpu_oeb[21]
port 303 nsew signal input
rlabel metal3 s 69600 51968 70000 52024 6 qcpu_oeb[22]
port 304 nsew signal input
rlabel metal3 s 69600 52528 70000 52584 6 qcpu_oeb[23]
port 305 nsew signal input
rlabel metal3 s 69600 53088 70000 53144 6 qcpu_oeb[24]
port 306 nsew signal input
rlabel metal3 s 69600 53648 70000 53704 6 qcpu_oeb[25]
port 307 nsew signal input
rlabel metal3 s 69600 54208 70000 54264 6 qcpu_oeb[26]
port 308 nsew signal input
rlabel metal3 s 69600 54768 70000 54824 6 qcpu_oeb[27]
port 309 nsew signal input
rlabel metal3 s 69600 55328 70000 55384 6 qcpu_oeb[28]
port 310 nsew signal input
rlabel metal3 s 69600 55888 70000 55944 6 qcpu_oeb[29]
port 311 nsew signal input
rlabel metal3 s 69600 40768 70000 40824 6 qcpu_oeb[2]
port 312 nsew signal input
rlabel metal3 s 69600 56448 70000 56504 6 qcpu_oeb[30]
port 313 nsew signal input
rlabel metal3 s 69600 57008 70000 57064 6 qcpu_oeb[31]
port 314 nsew signal input
rlabel metal3 s 69600 57568 70000 57624 6 qcpu_oeb[32]
port 315 nsew signal input
rlabel metal3 s 69600 41328 70000 41384 6 qcpu_oeb[3]
port 316 nsew signal input
rlabel metal3 s 69600 41888 70000 41944 6 qcpu_oeb[4]
port 317 nsew signal input
rlabel metal3 s 69600 42448 70000 42504 6 qcpu_oeb[5]
port 318 nsew signal input
rlabel metal3 s 69600 43008 70000 43064 6 qcpu_oeb[6]
port 319 nsew signal input
rlabel metal3 s 69600 43568 70000 43624 6 qcpu_oeb[7]
port 320 nsew signal input
rlabel metal3 s 69600 44128 70000 44184 6 qcpu_oeb[8]
port 321 nsew signal input
rlabel metal3 s 69600 44688 70000 44744 6 qcpu_oeb[9]
port 322 nsew signal input
rlabel metal2 s 60256 0 60312 400 6 qcpu_sram_addr[0]
port 323 nsew signal input
rlabel metal2 s 60704 0 60760 400 6 qcpu_sram_addr[1]
port 324 nsew signal input
rlabel metal2 s 61152 0 61208 400 6 qcpu_sram_addr[2]
port 325 nsew signal input
rlabel metal2 s 61600 0 61656 400 6 qcpu_sram_addr[3]
port 326 nsew signal input
rlabel metal2 s 62048 0 62104 400 6 qcpu_sram_addr[4]
port 327 nsew signal input
rlabel metal2 s 62496 0 62552 400 6 qcpu_sram_addr[5]
port 328 nsew signal input
rlabel metal2 s 62944 0 63000 400 6 qcpu_sram_gwe
port 329 nsew signal input
rlabel metal2 s 63392 0 63448 400 6 qcpu_sram_in[0]
port 330 nsew signal input
rlabel metal2 s 63840 0 63896 400 6 qcpu_sram_in[1]
port 331 nsew signal input
rlabel metal2 s 64288 0 64344 400 6 qcpu_sram_in[2]
port 332 nsew signal input
rlabel metal2 s 64736 0 64792 400 6 qcpu_sram_in[3]
port 333 nsew signal input
rlabel metal2 s 65184 0 65240 400 6 qcpu_sram_in[4]
port 334 nsew signal input
rlabel metal2 s 65632 0 65688 400 6 qcpu_sram_in[5]
port 335 nsew signal input
rlabel metal2 s 66080 0 66136 400 6 qcpu_sram_in[6]
port 336 nsew signal input
rlabel metal2 s 66528 0 66584 400 6 qcpu_sram_in[7]
port 337 nsew signal input
rlabel metal3 s 69600 58128 70000 58184 6 qcpu_sram_out[0]
port 338 nsew signal output
rlabel metal3 s 69600 58688 70000 58744 6 qcpu_sram_out[1]
port 339 nsew signal output
rlabel metal3 s 69600 59248 70000 59304 6 qcpu_sram_out[2]
port 340 nsew signal output
rlabel metal3 s 69600 59808 70000 59864 6 qcpu_sram_out[3]
port 341 nsew signal output
rlabel metal3 s 69600 60368 70000 60424 6 qcpu_sram_out[4]
port 342 nsew signal output
rlabel metal3 s 69600 60928 70000 60984 6 qcpu_sram_out[5]
port 343 nsew signal output
rlabel metal3 s 69600 61488 70000 61544 6 qcpu_sram_out[6]
port 344 nsew signal output
rlabel metal3 s 69600 62048 70000 62104 6 qcpu_sram_out[7]
port 345 nsew signal output
rlabel metal3 s 69600 62608 70000 62664 6 rst_ay8913
port 346 nsew signal output
rlabel metal2 s 19040 64600 19096 65000 6 rst_blinker
port 347 nsew signal output
rlabel metal3 s 0 56784 400 56840 6 rst_hellorld
port 348 nsew signal output
rlabel metal3 s 0 38864 400 38920 6 rst_mc14500
port 349 nsew signal output
rlabel metal3 s 69600 63168 70000 63224 6 rst_pdp11
port 350 nsew signal output
rlabel metal3 s 0 38304 400 38360 6 rst_qcpu
port 351 nsew signal output
rlabel metal3 s 0 25424 400 25480 6 rst_sid
port 352 nsew signal output
rlabel metal2 s 20832 64600 20888 65000 6 rst_sn76489
port 353 nsew signal output
rlabel metal3 s 0 57904 400 57960 6 rst_tbb1143
port 354 nsew signal output
rlabel metal3 s 0 25984 400 26040 6 sid_do[0]
port 355 nsew signal input
rlabel metal3 s 0 31584 400 31640 6 sid_do[10]
port 356 nsew signal input
rlabel metal3 s 0 32144 400 32200 6 sid_do[11]
port 357 nsew signal input
rlabel metal3 s 0 32704 400 32760 6 sid_do[12]
port 358 nsew signal input
rlabel metal3 s 0 33264 400 33320 6 sid_do[13]
port 359 nsew signal input
rlabel metal3 s 0 33824 400 33880 6 sid_do[14]
port 360 nsew signal input
rlabel metal3 s 0 34384 400 34440 6 sid_do[15]
port 361 nsew signal input
rlabel metal3 s 0 34944 400 35000 6 sid_do[16]
port 362 nsew signal input
rlabel metal3 s 0 35504 400 35560 6 sid_do[17]
port 363 nsew signal input
rlabel metal3 s 0 36064 400 36120 6 sid_do[18]
port 364 nsew signal input
rlabel metal3 s 0 36624 400 36680 6 sid_do[19]
port 365 nsew signal input
rlabel metal3 s 0 26544 400 26600 6 sid_do[1]
port 366 nsew signal input
rlabel metal3 s 0 37184 400 37240 6 sid_do[20]
port 367 nsew signal input
rlabel metal3 s 0 27104 400 27160 6 sid_do[2]
port 368 nsew signal input
rlabel metal3 s 0 27664 400 27720 6 sid_do[3]
port 369 nsew signal input
rlabel metal3 s 0 28224 400 28280 6 sid_do[4]
port 370 nsew signal input
rlabel metal3 s 0 28784 400 28840 6 sid_do[5]
port 371 nsew signal input
rlabel metal3 s 0 29344 400 29400 6 sid_do[6]
port 372 nsew signal input
rlabel metal3 s 0 29904 400 29960 6 sid_do[7]
port 373 nsew signal input
rlabel metal3 s 0 30464 400 30520 6 sid_do[8]
port 374 nsew signal input
rlabel metal3 s 0 31024 400 31080 6 sid_do[9]
port 375 nsew signal input
rlabel metal3 s 0 37744 400 37800 6 sid_oeb
port 376 nsew signal input
rlabel metal2 s 32928 0 32984 400 6 sn76489_do[0]
port 377 nsew signal input
rlabel metal2 s 37408 0 37464 400 6 sn76489_do[10]
port 378 nsew signal input
rlabel metal2 s 37856 0 37912 400 6 sn76489_do[11]
port 379 nsew signal input
rlabel metal2 s 38304 0 38360 400 6 sn76489_do[12]
port 380 nsew signal input
rlabel metal2 s 38752 0 38808 400 6 sn76489_do[13]
port 381 nsew signal input
rlabel metal2 s 39200 0 39256 400 6 sn76489_do[14]
port 382 nsew signal input
rlabel metal2 s 39648 0 39704 400 6 sn76489_do[15]
port 383 nsew signal input
rlabel metal2 s 40096 0 40152 400 6 sn76489_do[16]
port 384 nsew signal input
rlabel metal2 s 40544 0 40600 400 6 sn76489_do[17]
port 385 nsew signal input
rlabel metal2 s 40992 0 41048 400 6 sn76489_do[18]
port 386 nsew signal input
rlabel metal2 s 41440 0 41496 400 6 sn76489_do[19]
port 387 nsew signal input
rlabel metal2 s 33376 0 33432 400 6 sn76489_do[1]
port 388 nsew signal input
rlabel metal2 s 41888 0 41944 400 6 sn76489_do[20]
port 389 nsew signal input
rlabel metal2 s 42336 0 42392 400 6 sn76489_do[21]
port 390 nsew signal input
rlabel metal2 s 42784 0 42840 400 6 sn76489_do[22]
port 391 nsew signal input
rlabel metal2 s 43232 0 43288 400 6 sn76489_do[23]
port 392 nsew signal input
rlabel metal2 s 43680 0 43736 400 6 sn76489_do[24]
port 393 nsew signal input
rlabel metal2 s 44128 0 44184 400 6 sn76489_do[25]
port 394 nsew signal input
rlabel metal2 s 44576 0 44632 400 6 sn76489_do[26]
port 395 nsew signal input
rlabel metal2 s 45024 0 45080 400 6 sn76489_do[27]
port 396 nsew signal input
rlabel metal2 s 33824 0 33880 400 6 sn76489_do[2]
port 397 nsew signal input
rlabel metal2 s 34272 0 34328 400 6 sn76489_do[3]
port 398 nsew signal input
rlabel metal2 s 34720 0 34776 400 6 sn76489_do[4]
port 399 nsew signal input
rlabel metal2 s 35168 0 35224 400 6 sn76489_do[5]
port 400 nsew signal input
rlabel metal2 s 35616 0 35672 400 6 sn76489_do[6]
port 401 nsew signal input
rlabel metal2 s 36064 0 36120 400 6 sn76489_do[7]
port 402 nsew signal input
rlabel metal2 s 36512 0 36568 400 6 sn76489_do[8]
port 403 nsew signal input
rlabel metal2 s 36960 0 37016 400 6 sn76489_do[9]
port 404 nsew signal input
rlabel metal3 s 0 58464 400 58520 6 tbb1143_do[0]
port 405 nsew signal input
rlabel metal3 s 0 59024 400 59080 6 tbb1143_do[1]
port 406 nsew signal input
rlabel metal3 s 0 59584 400 59640 6 tbb1143_do[2]
port 407 nsew signal input
rlabel metal3 s 0 60144 400 60200 6 tbb1143_do[3]
port 408 nsew signal input
rlabel metal3 s 0 60704 400 60760 6 tbb1143_do[4]
port 409 nsew signal input
rlabel metal4 s 2224 1538 2384 63142 6 vdd
port 410 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 63142 6 vdd
port 410 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 63142 6 vdd
port 410 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 63142 6 vdd
port 410 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 63142 6 vdd
port 410 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 63142 6 vss
port 411 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 63142 6 vss
port 411 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 63142 6 vss
port 411 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 63142 6 vss
port 411 nsew ground bidirectional
rlabel metal2 s 3360 0 3416 400 6 wb_clk_i
port 412 nsew signal input
rlabel metal2 s 3808 0 3864 400 6 wb_rst_i
port 413 nsew signal input
rlabel metal3 s 69600 21168 70000 21224 6 wbs_ack_o
port 414 nsew signal output
rlabel metal2 s 4256 0 4312 400 6 wbs_adr_i[0]
port 415 nsew signal input
rlabel metal2 s 8736 0 8792 400 6 wbs_adr_i[10]
port 416 nsew signal input
rlabel metal2 s 9184 0 9240 400 6 wbs_adr_i[11]
port 417 nsew signal input
rlabel metal2 s 9632 0 9688 400 6 wbs_adr_i[12]
port 418 nsew signal input
rlabel metal2 s 10080 0 10136 400 6 wbs_adr_i[13]
port 419 nsew signal input
rlabel metal2 s 10528 0 10584 400 6 wbs_adr_i[14]
port 420 nsew signal input
rlabel metal2 s 10976 0 11032 400 6 wbs_adr_i[15]
port 421 nsew signal input
rlabel metal2 s 11424 0 11480 400 6 wbs_adr_i[16]
port 422 nsew signal input
rlabel metal2 s 11872 0 11928 400 6 wbs_adr_i[17]
port 423 nsew signal input
rlabel metal2 s 12320 0 12376 400 6 wbs_adr_i[18]
port 424 nsew signal input
rlabel metal2 s 12768 0 12824 400 6 wbs_adr_i[19]
port 425 nsew signal input
rlabel metal2 s 4704 0 4760 400 6 wbs_adr_i[1]
port 426 nsew signal input
rlabel metal2 s 13216 0 13272 400 6 wbs_adr_i[20]
port 427 nsew signal input
rlabel metal2 s 13664 0 13720 400 6 wbs_adr_i[21]
port 428 nsew signal input
rlabel metal2 s 14112 0 14168 400 6 wbs_adr_i[22]
port 429 nsew signal input
rlabel metal2 s 14560 0 14616 400 6 wbs_adr_i[23]
port 430 nsew signal input
rlabel metal2 s 15008 0 15064 400 6 wbs_adr_i[24]
port 431 nsew signal input
rlabel metal2 s 15456 0 15512 400 6 wbs_adr_i[25]
port 432 nsew signal input
rlabel metal2 s 15904 0 15960 400 6 wbs_adr_i[26]
port 433 nsew signal input
rlabel metal2 s 16352 0 16408 400 6 wbs_adr_i[27]
port 434 nsew signal input
rlabel metal2 s 16800 0 16856 400 6 wbs_adr_i[28]
port 435 nsew signal input
rlabel metal2 s 17248 0 17304 400 6 wbs_adr_i[29]
port 436 nsew signal input
rlabel metal2 s 5152 0 5208 400 6 wbs_adr_i[2]
port 437 nsew signal input
rlabel metal2 s 17696 0 17752 400 6 wbs_adr_i[30]
port 438 nsew signal input
rlabel metal2 s 18144 0 18200 400 6 wbs_adr_i[31]
port 439 nsew signal input
rlabel metal2 s 5600 0 5656 400 6 wbs_adr_i[3]
port 440 nsew signal input
rlabel metal2 s 6048 0 6104 400 6 wbs_adr_i[4]
port 441 nsew signal input
rlabel metal2 s 6496 0 6552 400 6 wbs_adr_i[5]
port 442 nsew signal input
rlabel metal2 s 6944 0 7000 400 6 wbs_adr_i[6]
port 443 nsew signal input
rlabel metal2 s 7392 0 7448 400 6 wbs_adr_i[7]
port 444 nsew signal input
rlabel metal2 s 7840 0 7896 400 6 wbs_adr_i[8]
port 445 nsew signal input
rlabel metal2 s 8288 0 8344 400 6 wbs_adr_i[9]
port 446 nsew signal input
rlabel metal3 s 69600 20048 70000 20104 6 wbs_cyc_i
port 447 nsew signal input
rlabel metal2 s 18592 0 18648 400 6 wbs_dat_i[0]
port 448 nsew signal input
rlabel metal2 s 23072 0 23128 400 6 wbs_dat_i[10]
port 449 nsew signal input
rlabel metal2 s 23520 0 23576 400 6 wbs_dat_i[11]
port 450 nsew signal input
rlabel metal2 s 23968 0 24024 400 6 wbs_dat_i[12]
port 451 nsew signal input
rlabel metal2 s 24416 0 24472 400 6 wbs_dat_i[13]
port 452 nsew signal input
rlabel metal2 s 24864 0 24920 400 6 wbs_dat_i[14]
port 453 nsew signal input
rlabel metal2 s 25312 0 25368 400 6 wbs_dat_i[15]
port 454 nsew signal input
rlabel metal2 s 25760 0 25816 400 6 wbs_dat_i[16]
port 455 nsew signal input
rlabel metal2 s 26208 0 26264 400 6 wbs_dat_i[17]
port 456 nsew signal input
rlabel metal2 s 26656 0 26712 400 6 wbs_dat_i[18]
port 457 nsew signal input
rlabel metal2 s 27104 0 27160 400 6 wbs_dat_i[19]
port 458 nsew signal input
rlabel metal2 s 19040 0 19096 400 6 wbs_dat_i[1]
port 459 nsew signal input
rlabel metal2 s 27552 0 27608 400 6 wbs_dat_i[20]
port 460 nsew signal input
rlabel metal2 s 28000 0 28056 400 6 wbs_dat_i[21]
port 461 nsew signal input
rlabel metal2 s 28448 0 28504 400 6 wbs_dat_i[22]
port 462 nsew signal input
rlabel metal2 s 28896 0 28952 400 6 wbs_dat_i[23]
port 463 nsew signal input
rlabel metal2 s 29344 0 29400 400 6 wbs_dat_i[24]
port 464 nsew signal input
rlabel metal2 s 29792 0 29848 400 6 wbs_dat_i[25]
port 465 nsew signal input
rlabel metal2 s 30240 0 30296 400 6 wbs_dat_i[26]
port 466 nsew signal input
rlabel metal2 s 30688 0 30744 400 6 wbs_dat_i[27]
port 467 nsew signal input
rlabel metal2 s 31136 0 31192 400 6 wbs_dat_i[28]
port 468 nsew signal input
rlabel metal2 s 31584 0 31640 400 6 wbs_dat_i[29]
port 469 nsew signal input
rlabel metal2 s 19488 0 19544 400 6 wbs_dat_i[2]
port 470 nsew signal input
rlabel metal2 s 32032 0 32088 400 6 wbs_dat_i[30]
port 471 nsew signal input
rlabel metal2 s 32480 0 32536 400 6 wbs_dat_i[31]
port 472 nsew signal input
rlabel metal2 s 19936 0 19992 400 6 wbs_dat_i[3]
port 473 nsew signal input
rlabel metal2 s 20384 0 20440 400 6 wbs_dat_i[4]
port 474 nsew signal input
rlabel metal2 s 20832 0 20888 400 6 wbs_dat_i[5]
port 475 nsew signal input
rlabel metal2 s 21280 0 21336 400 6 wbs_dat_i[6]
port 476 nsew signal input
rlabel metal2 s 21728 0 21784 400 6 wbs_dat_i[7]
port 477 nsew signal input
rlabel metal2 s 22176 0 22232 400 6 wbs_dat_i[8]
port 478 nsew signal input
rlabel metal2 s 22624 0 22680 400 6 wbs_dat_i[9]
port 479 nsew signal input
rlabel metal3 s 69600 1568 70000 1624 6 wbs_dat_o[0]
port 480 nsew signal output
rlabel metal3 s 69600 7168 70000 7224 6 wbs_dat_o[10]
port 481 nsew signal output
rlabel metal3 s 69600 7728 70000 7784 6 wbs_dat_o[11]
port 482 nsew signal output
rlabel metal3 s 69600 8288 70000 8344 6 wbs_dat_o[12]
port 483 nsew signal output
rlabel metal3 s 69600 8848 70000 8904 6 wbs_dat_o[13]
port 484 nsew signal output
rlabel metal3 s 69600 9408 70000 9464 6 wbs_dat_o[14]
port 485 nsew signal output
rlabel metal3 s 69600 9968 70000 10024 6 wbs_dat_o[15]
port 486 nsew signal output
rlabel metal3 s 69600 10528 70000 10584 6 wbs_dat_o[16]
port 487 nsew signal output
rlabel metal3 s 69600 11088 70000 11144 6 wbs_dat_o[17]
port 488 nsew signal output
rlabel metal3 s 69600 11648 70000 11704 6 wbs_dat_o[18]
port 489 nsew signal output
rlabel metal3 s 69600 12208 70000 12264 6 wbs_dat_o[19]
port 490 nsew signal output
rlabel metal3 s 69600 2128 70000 2184 6 wbs_dat_o[1]
port 491 nsew signal output
rlabel metal3 s 69600 12768 70000 12824 6 wbs_dat_o[20]
port 492 nsew signal output
rlabel metal3 s 69600 13328 70000 13384 6 wbs_dat_o[21]
port 493 nsew signal output
rlabel metal3 s 69600 13888 70000 13944 6 wbs_dat_o[22]
port 494 nsew signal output
rlabel metal3 s 69600 14448 70000 14504 6 wbs_dat_o[23]
port 495 nsew signal output
rlabel metal3 s 69600 15008 70000 15064 6 wbs_dat_o[24]
port 496 nsew signal output
rlabel metal3 s 69600 15568 70000 15624 6 wbs_dat_o[25]
port 497 nsew signal output
rlabel metal3 s 69600 16128 70000 16184 6 wbs_dat_o[26]
port 498 nsew signal output
rlabel metal3 s 69600 16688 70000 16744 6 wbs_dat_o[27]
port 499 nsew signal output
rlabel metal3 s 69600 17248 70000 17304 6 wbs_dat_o[28]
port 500 nsew signal output
rlabel metal3 s 69600 17808 70000 17864 6 wbs_dat_o[29]
port 501 nsew signal output
rlabel metal3 s 69600 2688 70000 2744 6 wbs_dat_o[2]
port 502 nsew signal output
rlabel metal3 s 69600 18368 70000 18424 6 wbs_dat_o[30]
port 503 nsew signal output
rlabel metal3 s 69600 18928 70000 18984 6 wbs_dat_o[31]
port 504 nsew signal output
rlabel metal3 s 69600 3248 70000 3304 6 wbs_dat_o[3]
port 505 nsew signal output
rlabel metal3 s 69600 3808 70000 3864 6 wbs_dat_o[4]
port 506 nsew signal output
rlabel metal3 s 69600 4368 70000 4424 6 wbs_dat_o[5]
port 507 nsew signal output
rlabel metal3 s 69600 4928 70000 4984 6 wbs_dat_o[6]
port 508 nsew signal output
rlabel metal3 s 69600 5488 70000 5544 6 wbs_dat_o[7]
port 509 nsew signal output
rlabel metal3 s 69600 6048 70000 6104 6 wbs_dat_o[8]
port 510 nsew signal output
rlabel metal3 s 69600 6608 70000 6664 6 wbs_dat_o[9]
port 511 nsew signal output
rlabel metal3 s 69600 20608 70000 20664 6 wbs_stb_i
port 512 nsew signal input
rlabel metal3 s 69600 19488 70000 19544 6 wbs_we_i
port 513 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 70000 65000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9076072
string GDS_FILE /run/media/tholin/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/gfmpw1-multi/openlane/Multiplexer/runs/23_12_08_15_40/results/signoff/multiplexer.magic.gds
string GDS_START 398754
<< end >>

