VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO multiplexer
  CLASS BLOCK ;
  FOREIGN multiplexer ;
  ORIGIN 0.000 0.000 ;
  SIZE 650.000 BY 600.000 ;
  PIN ay8913_do[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 484.960 596.000 485.520 600.000 ;
    END
  END ay8913_do[0]
  PIN ay8913_do[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 529.760 596.000 530.320 600.000 ;
    END
  END ay8913_do[10]
  PIN ay8913_do[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 534.240 596.000 534.800 600.000 ;
    END
  END ay8913_do[11]
  PIN ay8913_do[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 538.720 596.000 539.280 600.000 ;
    END
  END ay8913_do[12]
  PIN ay8913_do[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 543.200 596.000 543.760 600.000 ;
    END
  END ay8913_do[13]
  PIN ay8913_do[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 547.680 596.000 548.240 600.000 ;
    END
  END ay8913_do[14]
  PIN ay8913_do[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 552.160 596.000 552.720 600.000 ;
    END
  END ay8913_do[15]
  PIN ay8913_do[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 556.640 596.000 557.200 600.000 ;
    END
  END ay8913_do[16]
  PIN ay8913_do[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 561.120 596.000 561.680 600.000 ;
    END
  END ay8913_do[17]
  PIN ay8913_do[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 565.600 596.000 566.160 600.000 ;
    END
  END ay8913_do[18]
  PIN ay8913_do[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 570.080 596.000 570.640 600.000 ;
    END
  END ay8913_do[19]
  PIN ay8913_do[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 489.440 596.000 490.000 600.000 ;
    END
  END ay8913_do[1]
  PIN ay8913_do[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 574.560 596.000 575.120 600.000 ;
    END
  END ay8913_do[20]
  PIN ay8913_do[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 579.040 596.000 579.600 600.000 ;
    END
  END ay8913_do[21]
  PIN ay8913_do[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 583.520 596.000 584.080 600.000 ;
    END
  END ay8913_do[22]
  PIN ay8913_do[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 588.000 596.000 588.560 600.000 ;
    END
  END ay8913_do[23]
  PIN ay8913_do[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 592.480 596.000 593.040 600.000 ;
    END
  END ay8913_do[24]
  PIN ay8913_do[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 596.960 596.000 597.520 600.000 ;
    END
  END ay8913_do[25]
  PIN ay8913_do[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 601.440 596.000 602.000 600.000 ;
    END
  END ay8913_do[26]
  PIN ay8913_do[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 605.920 596.000 606.480 600.000 ;
    END
  END ay8913_do[27]
  PIN ay8913_do[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 493.920 596.000 494.480 600.000 ;
    END
  END ay8913_do[2]
  PIN ay8913_do[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 498.400 596.000 498.960 600.000 ;
    END
  END ay8913_do[3]
  PIN ay8913_do[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 502.880 596.000 503.440 600.000 ;
    END
  END ay8913_do[4]
  PIN ay8913_do[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 507.360 596.000 507.920 600.000 ;
    END
  END ay8913_do[5]
  PIN ay8913_do[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 511.840 596.000 512.400 600.000 ;
    END
  END ay8913_do[6]
  PIN ay8913_do[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 516.320 596.000 516.880 600.000 ;
    END
  END ay8913_do[7]
  PIN ay8913_do[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 520.800 596.000 521.360 600.000 ;
    END
  END ay8913_do[8]
  PIN ay8913_do[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 525.280 596.000 525.840 600.000 ;
    END
  END ay8913_do[9]
  PIN blinker_do[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 399.840 596.000 400.400 600.000 ;
    END
  END blinker_do[0]
  PIN blinker_do[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 404.320 596.000 404.880 600.000 ;
    END
  END blinker_do[1]
  PIN blinker_do[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 408.800 596.000 409.360 600.000 ;
    END
  END blinker_do[2]
  PIN custom_settings[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 198.240 650.000 198.800 ;
    END
  END custom_settings[0]
  PIN custom_settings[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 243.040 650.000 243.600 ;
    END
  END custom_settings[10]
  PIN custom_settings[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 247.520 650.000 248.080 ;
    END
  END custom_settings[11]
  PIN custom_settings[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 252.000 650.000 252.560 ;
    END
  END custom_settings[12]
  PIN custom_settings[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 256.480 650.000 257.040 ;
    END
  END custom_settings[13]
  PIN custom_settings[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 260.960 650.000 261.520 ;
    END
  END custom_settings[14]
  PIN custom_settings[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 265.440 650.000 266.000 ;
    END
  END custom_settings[15]
  PIN custom_settings[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 269.920 650.000 270.480 ;
    END
  END custom_settings[16]
  PIN custom_settings[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 274.400 650.000 274.960 ;
    END
  END custom_settings[17]
  PIN custom_settings[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 278.880 650.000 279.440 ;
    END
  END custom_settings[18]
  PIN custom_settings[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 283.360 650.000 283.920 ;
    END
  END custom_settings[19]
  PIN custom_settings[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 202.720 650.000 203.280 ;
    END
  END custom_settings[1]
  PIN custom_settings[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 287.840 650.000 288.400 ;
    END
  END custom_settings[20]
  PIN custom_settings[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 292.320 650.000 292.880 ;
    END
  END custom_settings[21]
  PIN custom_settings[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 296.800 650.000 297.360 ;
    END
  END custom_settings[22]
  PIN custom_settings[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 301.280 650.000 301.840 ;
    END
  END custom_settings[23]
  PIN custom_settings[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 305.760 650.000 306.320 ;
    END
  END custom_settings[24]
  PIN custom_settings[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 310.240 650.000 310.800 ;
    END
  END custom_settings[25]
  PIN custom_settings[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 314.720 650.000 315.280 ;
    END
  END custom_settings[26]
  PIN custom_settings[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 319.200 650.000 319.760 ;
    END
  END custom_settings[27]
  PIN custom_settings[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 323.680 650.000 324.240 ;
    END
  END custom_settings[28]
  PIN custom_settings[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 328.160 650.000 328.720 ;
    END
  END custom_settings[29]
  PIN custom_settings[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 207.200 650.000 207.760 ;
    END
  END custom_settings[2]
  PIN custom_settings[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 332.640 650.000 333.200 ;
    END
  END custom_settings[30]
  PIN custom_settings[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 337.120 650.000 337.680 ;
    END
  END custom_settings[31]
  PIN custom_settings[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 211.680 650.000 212.240 ;
    END
  END custom_settings[3]
  PIN custom_settings[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 216.160 650.000 216.720 ;
    END
  END custom_settings[4]
  PIN custom_settings[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 220.640 650.000 221.200 ;
    END
  END custom_settings[5]
  PIN custom_settings[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 225.120 650.000 225.680 ;
    END
  END custom_settings[6]
  PIN custom_settings[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 229.600 650.000 230.160 ;
    END
  END custom_settings[7]
  PIN custom_settings[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 234.080 650.000 234.640 ;
    END
  END custom_settings[8]
  PIN custom_settings[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 238.560 650.000 239.120 ;
    END
  END custom_settings[9]
  PIN hellorld_do
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 565.600 4.000 566.160 ;
    END
  END hellorld_do
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 41.440 596.000 42.000 600.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 86.240 596.000 86.800 600.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 596.000 91.280 600.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 596.000 95.760 600.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 99.680 596.000 100.240 600.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 596.000 104.720 600.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 108.640 596.000 109.200 600.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 113.120 596.000 113.680 600.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 596.000 118.160 600.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 122.080 596.000 122.640 600.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 126.560 596.000 127.120 600.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 45.920 596.000 46.480 600.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 596.000 131.600 600.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 135.520 596.000 136.080 600.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 140.000 596.000 140.560 600.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 596.000 145.040 600.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 148.960 596.000 149.520 600.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 153.440 596.000 154.000 600.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 596.000 158.480 600.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 162.400 596.000 162.960 600.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 166.880 596.000 167.440 600.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 596.000 171.920 600.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 596.000 50.960 600.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 175.840 596.000 176.400 600.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 180.320 596.000 180.880 600.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 596.000 185.360 600.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 189.280 596.000 189.840 600.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 193.760 596.000 194.320 600.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 198.240 596.000 198.800 600.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 202.720 596.000 203.280 600.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 207.200 596.000 207.760 600.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 54.880 596.000 55.440 600.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 59.360 596.000 59.920 600.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 596.000 64.400 600.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 68.320 596.000 68.880 600.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 72.800 596.000 73.360 600.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 596.000 77.840 600.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 81.760 596.000 82.320 600.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 33.600 4.000 34.160 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 89.600 4.000 90.160 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 95.200 4.000 95.760 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 100.800 4.000 101.360 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 106.400 4.000 106.960 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 112.000 4.000 112.560 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 117.600 4.000 118.160 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 123.200 4.000 123.760 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 128.800 4.000 129.360 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 134.400 4.000 134.960 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 140.000 4.000 140.560 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 39.200 4.000 39.760 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 145.600 4.000 146.160 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 151.200 4.000 151.760 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 156.800 4.000 157.360 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 162.400 4.000 162.960 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 168.000 4.000 168.560 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 173.600 4.000 174.160 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 179.200 4.000 179.760 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 184.800 4.000 185.360 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 190.400 4.000 190.960 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 196.000 4.000 196.560 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 44.800 4.000 45.360 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 201.600 4.000 202.160 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 207.200 4.000 207.760 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 212.800 4.000 213.360 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 218.400 4.000 218.960 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 224.000 4.000 224.560 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 229.600 4.000 230.160 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 235.200 4.000 235.760 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 240.800 4.000 241.360 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 50.400 4.000 50.960 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 56.000 4.000 56.560 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 61.600 4.000 62.160 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 67.200 4.000 67.760 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 72.800 4.000 73.360 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 78.400 4.000 78.960 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 84.000 4.000 84.560 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 596.000 212.240 600.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 256.480 596.000 257.040 600.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 260.960 596.000 261.520 600.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 265.440 596.000 266.000 600.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 269.920 596.000 270.480 600.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 274.400 596.000 274.960 600.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 278.880 596.000 279.440 600.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 283.360 596.000 283.920 600.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 287.840 596.000 288.400 600.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 292.320 596.000 292.880 600.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 296.800 596.000 297.360 600.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 216.160 596.000 216.720 600.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 301.280 596.000 301.840 600.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 305.760 596.000 306.320 600.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 310.240 596.000 310.800 600.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 314.720 596.000 315.280 600.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 319.200 596.000 319.760 600.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 323.680 596.000 324.240 600.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 328.160 596.000 328.720 600.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 332.640 596.000 333.200 600.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 337.120 596.000 337.680 600.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 341.600 596.000 342.160 600.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 220.640 596.000 221.200 600.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 346.080 596.000 346.640 600.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 350.560 596.000 351.120 600.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 355.040 596.000 355.600 600.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 359.520 596.000 360.080 600.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 364.000 596.000 364.560 600.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 368.480 596.000 369.040 600.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 372.960 596.000 373.520 600.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 377.440 596.000 378.000 600.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 596.000 225.680 600.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 229.600 596.000 230.160 600.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 234.080 596.000 234.640 600.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 238.560 596.000 239.120 600.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 243.040 596.000 243.600 600.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 247.520 596.000 248.080 600.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 596.000 252.560 600.000 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 381.920 596.000 382.480 600.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 386.400 596.000 386.960 600.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 390.880 596.000 391.440 600.000 ;
    END
  END irq[2]
  PIN mc14500_do[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 386.400 4.000 386.960 ;
    END
  END mc14500_do[0]
  PIN mc14500_do[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 442.400 4.000 442.960 ;
    END
  END mc14500_do[10]
  PIN mc14500_do[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 448.000 4.000 448.560 ;
    END
  END mc14500_do[11]
  PIN mc14500_do[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 453.600 4.000 454.160 ;
    END
  END mc14500_do[12]
  PIN mc14500_do[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 459.200 4.000 459.760 ;
    END
  END mc14500_do[13]
  PIN mc14500_do[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 464.800 4.000 465.360 ;
    END
  END mc14500_do[14]
  PIN mc14500_do[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 470.400 4.000 470.960 ;
    END
  END mc14500_do[15]
  PIN mc14500_do[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 476.000 4.000 476.560 ;
    END
  END mc14500_do[16]
  PIN mc14500_do[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 481.600 4.000 482.160 ;
    END
  END mc14500_do[17]
  PIN mc14500_do[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 487.200 4.000 487.760 ;
    END
  END mc14500_do[18]
  PIN mc14500_do[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 492.800 4.000 493.360 ;
    END
  END mc14500_do[19]
  PIN mc14500_do[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 392.000 4.000 392.560 ;
    END
  END mc14500_do[1]
  PIN mc14500_do[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 498.400 4.000 498.960 ;
    END
  END mc14500_do[20]
  PIN mc14500_do[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 504.000 4.000 504.560 ;
    END
  END mc14500_do[21]
  PIN mc14500_do[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 509.600 4.000 510.160 ;
    END
  END mc14500_do[22]
  PIN mc14500_do[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 515.200 4.000 515.760 ;
    END
  END mc14500_do[23]
  PIN mc14500_do[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 520.800 4.000 521.360 ;
    END
  END mc14500_do[24]
  PIN mc14500_do[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 526.400 4.000 526.960 ;
    END
  END mc14500_do[25]
  PIN mc14500_do[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 532.000 4.000 532.560 ;
    END
  END mc14500_do[26]
  PIN mc14500_do[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 537.600 4.000 538.160 ;
    END
  END mc14500_do[27]
  PIN mc14500_do[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 543.200 4.000 543.760 ;
    END
  END mc14500_do[28]
  PIN mc14500_do[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 548.800 4.000 549.360 ;
    END
  END mc14500_do[29]
  PIN mc14500_do[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 397.600 4.000 398.160 ;
    END
  END mc14500_do[2]
  PIN mc14500_do[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 554.400 4.000 554.960 ;
    END
  END mc14500_do[30]
  PIN mc14500_do[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 403.200 4.000 403.760 ;
    END
  END mc14500_do[3]
  PIN mc14500_do[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 408.800 4.000 409.360 ;
    END
  END mc14500_do[4]
  PIN mc14500_do[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 414.400 4.000 414.960 ;
    END
  END mc14500_do[5]
  PIN mc14500_do[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 420.000 4.000 420.560 ;
    END
  END mc14500_do[6]
  PIN mc14500_do[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 425.600 4.000 426.160 ;
    END
  END mc14500_do[7]
  PIN mc14500_do[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 431.200 4.000 431.760 ;
    END
  END mc14500_do[8]
  PIN mc14500_do[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 436.800 4.000 437.360 ;
    END
  END mc14500_do[9]
  PIN mc14500_sram_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 417.760 596.000 418.320 600.000 ;
    END
  END mc14500_sram_addr[0]
  PIN mc14500_sram_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 422.240 596.000 422.800 600.000 ;
    END
  END mc14500_sram_addr[1]
  PIN mc14500_sram_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 426.720 596.000 427.280 600.000 ;
    END
  END mc14500_sram_addr[2]
  PIN mc14500_sram_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 431.200 596.000 431.760 600.000 ;
    END
  END mc14500_sram_addr[3]
  PIN mc14500_sram_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 435.680 596.000 436.240 600.000 ;
    END
  END mc14500_sram_addr[4]
  PIN mc14500_sram_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 440.160 596.000 440.720 600.000 ;
    END
  END mc14500_sram_addr[5]
  PIN mc14500_sram_gwe
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 480.480 596.000 481.040 600.000 ;
    END
  END mc14500_sram_gwe
  PIN mc14500_sram_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 444.640 596.000 445.200 600.000 ;
    END
  END mc14500_sram_in[0]
  PIN mc14500_sram_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 449.120 596.000 449.680 600.000 ;
    END
  END mc14500_sram_in[1]
  PIN mc14500_sram_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 453.600 596.000 454.160 600.000 ;
    END
  END mc14500_sram_in[2]
  PIN mc14500_sram_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 458.080 596.000 458.640 600.000 ;
    END
  END mc14500_sram_in[3]
  PIN mc14500_sram_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 462.560 596.000 463.120 600.000 ;
    END
  END mc14500_sram_in[4]
  PIN mc14500_sram_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 467.040 596.000 467.600 600.000 ;
    END
  END mc14500_sram_in[5]
  PIN mc14500_sram_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 471.520 596.000 472.080 600.000 ;
    END
  END mc14500_sram_in[6]
  PIN mc14500_sram_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 476.000 596.000 476.560 600.000 ;
    END
  END mc14500_sram_in[7]
  PIN qcpu_do[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 446.880 0.000 447.440 4.000 ;
    END
  END qcpu_do[0]
  PIN qcpu_do[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 491.680 0.000 492.240 4.000 ;
    END
  END qcpu_do[10]
  PIN qcpu_do[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 496.160 0.000 496.720 4.000 ;
    END
  END qcpu_do[11]
  PIN qcpu_do[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 500.640 0.000 501.200 4.000 ;
    END
  END qcpu_do[12]
  PIN qcpu_do[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 505.120 0.000 505.680 4.000 ;
    END
  END qcpu_do[13]
  PIN qcpu_do[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 509.600 0.000 510.160 4.000 ;
    END
  END qcpu_do[14]
  PIN qcpu_do[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 514.080 0.000 514.640 4.000 ;
    END
  END qcpu_do[15]
  PIN qcpu_do[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 518.560 0.000 519.120 4.000 ;
    END
  END qcpu_do[16]
  PIN qcpu_do[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 523.040 0.000 523.600 4.000 ;
    END
  END qcpu_do[17]
  PIN qcpu_do[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 527.520 0.000 528.080 4.000 ;
    END
  END qcpu_do[18]
  PIN qcpu_do[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 532.000 0.000 532.560 4.000 ;
    END
  END qcpu_do[19]
  PIN qcpu_do[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 451.360 0.000 451.920 4.000 ;
    END
  END qcpu_do[1]
  PIN qcpu_do[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 536.480 0.000 537.040 4.000 ;
    END
  END qcpu_do[20]
  PIN qcpu_do[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 540.960 0.000 541.520 4.000 ;
    END
  END qcpu_do[21]
  PIN qcpu_do[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 545.440 0.000 546.000 4.000 ;
    END
  END qcpu_do[22]
  PIN qcpu_do[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 549.920 0.000 550.480 4.000 ;
    END
  END qcpu_do[23]
  PIN qcpu_do[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 554.400 0.000 554.960 4.000 ;
    END
  END qcpu_do[24]
  PIN qcpu_do[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 558.880 0.000 559.440 4.000 ;
    END
  END qcpu_do[25]
  PIN qcpu_do[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 563.360 0.000 563.920 4.000 ;
    END
  END qcpu_do[26]
  PIN qcpu_do[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 567.840 0.000 568.400 4.000 ;
    END
  END qcpu_do[27]
  PIN qcpu_do[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 572.320 0.000 572.880 4.000 ;
    END
  END qcpu_do[28]
  PIN qcpu_do[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 576.800 0.000 577.360 4.000 ;
    END
  END qcpu_do[29]
  PIN qcpu_do[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 455.840 0.000 456.400 4.000 ;
    END
  END qcpu_do[2]
  PIN qcpu_do[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 581.280 0.000 581.840 4.000 ;
    END
  END qcpu_do[30]
  PIN qcpu_do[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 585.760 0.000 586.320 4.000 ;
    END
  END qcpu_do[31]
  PIN qcpu_do[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 590.240 0.000 590.800 4.000 ;
    END
  END qcpu_do[32]
  PIN qcpu_do[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 460.320 0.000 460.880 4.000 ;
    END
  END qcpu_do[3]
  PIN qcpu_do[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 464.800 0.000 465.360 4.000 ;
    END
  END qcpu_do[4]
  PIN qcpu_do[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 469.280 0.000 469.840 4.000 ;
    END
  END qcpu_do[5]
  PIN qcpu_do[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 473.760 0.000 474.320 4.000 ;
    END
  END qcpu_do[6]
  PIN qcpu_do[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 478.240 0.000 478.800 4.000 ;
    END
  END qcpu_do[7]
  PIN qcpu_do[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 482.720 0.000 483.280 4.000 ;
    END
  END qcpu_do[8]
  PIN qcpu_do[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 487.200 0.000 487.760 4.000 ;
    END
  END qcpu_do[9]
  PIN qcpu_oeb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 341.600 650.000 342.160 ;
    END
  END qcpu_oeb[0]
  PIN qcpu_oeb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 386.400 650.000 386.960 ;
    END
  END qcpu_oeb[10]
  PIN qcpu_oeb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 390.880 650.000 391.440 ;
    END
  END qcpu_oeb[11]
  PIN qcpu_oeb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 395.360 650.000 395.920 ;
    END
  END qcpu_oeb[12]
  PIN qcpu_oeb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 399.840 650.000 400.400 ;
    END
  END qcpu_oeb[13]
  PIN qcpu_oeb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 404.320 650.000 404.880 ;
    END
  END qcpu_oeb[14]
  PIN qcpu_oeb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 408.800 650.000 409.360 ;
    END
  END qcpu_oeb[15]
  PIN qcpu_oeb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 413.280 650.000 413.840 ;
    END
  END qcpu_oeb[16]
  PIN qcpu_oeb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 417.760 650.000 418.320 ;
    END
  END qcpu_oeb[17]
  PIN qcpu_oeb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 422.240 650.000 422.800 ;
    END
  END qcpu_oeb[18]
  PIN qcpu_oeb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 426.720 650.000 427.280 ;
    END
  END qcpu_oeb[19]
  PIN qcpu_oeb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 346.080 650.000 346.640 ;
    END
  END qcpu_oeb[1]
  PIN qcpu_oeb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 431.200 650.000 431.760 ;
    END
  END qcpu_oeb[20]
  PIN qcpu_oeb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 435.680 650.000 436.240 ;
    END
  END qcpu_oeb[21]
  PIN qcpu_oeb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 440.160 650.000 440.720 ;
    END
  END qcpu_oeb[22]
  PIN qcpu_oeb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 444.640 650.000 445.200 ;
    END
  END qcpu_oeb[23]
  PIN qcpu_oeb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 449.120 650.000 449.680 ;
    END
  END qcpu_oeb[24]
  PIN qcpu_oeb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 453.600 650.000 454.160 ;
    END
  END qcpu_oeb[25]
  PIN qcpu_oeb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 458.080 650.000 458.640 ;
    END
  END qcpu_oeb[26]
  PIN qcpu_oeb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 462.560 650.000 463.120 ;
    END
  END qcpu_oeb[27]
  PIN qcpu_oeb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 467.040 650.000 467.600 ;
    END
  END qcpu_oeb[28]
  PIN qcpu_oeb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 471.520 650.000 472.080 ;
    END
  END qcpu_oeb[29]
  PIN qcpu_oeb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 350.560 650.000 351.120 ;
    END
  END qcpu_oeb[2]
  PIN qcpu_oeb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 476.000 650.000 476.560 ;
    END
  END qcpu_oeb[30]
  PIN qcpu_oeb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 480.480 650.000 481.040 ;
    END
  END qcpu_oeb[31]
  PIN qcpu_oeb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 484.960 650.000 485.520 ;
    END
  END qcpu_oeb[32]
  PIN qcpu_oeb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 355.040 650.000 355.600 ;
    END
  END qcpu_oeb[3]
  PIN qcpu_oeb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 359.520 650.000 360.080 ;
    END
  END qcpu_oeb[4]
  PIN qcpu_oeb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 364.000 650.000 364.560 ;
    END
  END qcpu_oeb[5]
  PIN qcpu_oeb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 368.480 650.000 369.040 ;
    END
  END qcpu_oeb[6]
  PIN qcpu_oeb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 372.960 650.000 373.520 ;
    END
  END qcpu_oeb[7]
  PIN qcpu_oeb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 377.440 650.000 378.000 ;
    END
  END qcpu_oeb[8]
  PIN qcpu_oeb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 381.920 650.000 382.480 ;
    END
  END qcpu_oeb[9]
  PIN qcpu_sram_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 594.720 0.000 595.280 4.000 ;
    END
  END qcpu_sram_addr[0]
  PIN qcpu_sram_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 599.200 0.000 599.760 4.000 ;
    END
  END qcpu_sram_addr[1]
  PIN qcpu_sram_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 603.680 0.000 604.240 4.000 ;
    END
  END qcpu_sram_addr[2]
  PIN qcpu_sram_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 608.160 0.000 608.720 4.000 ;
    END
  END qcpu_sram_addr[3]
  PIN qcpu_sram_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 612.640 0.000 613.200 4.000 ;
    END
  END qcpu_sram_addr[4]
  PIN qcpu_sram_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 617.120 0.000 617.680 4.000 ;
    END
  END qcpu_sram_addr[5]
  PIN qcpu_sram_gwe
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 621.600 0.000 622.160 4.000 ;
    END
  END qcpu_sram_gwe
  PIN qcpu_sram_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 489.440 650.000 490.000 ;
    END
  END qcpu_sram_in[0]
  PIN qcpu_sram_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 493.920 650.000 494.480 ;
    END
  END qcpu_sram_in[1]
  PIN qcpu_sram_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 498.400 650.000 498.960 ;
    END
  END qcpu_sram_in[2]
  PIN qcpu_sram_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 502.880 650.000 503.440 ;
    END
  END qcpu_sram_in[3]
  PIN qcpu_sram_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 507.360 650.000 507.920 ;
    END
  END qcpu_sram_in[4]
  PIN qcpu_sram_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 511.840 650.000 512.400 ;
    END
  END qcpu_sram_in[5]
  PIN qcpu_sram_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 516.320 650.000 516.880 ;
    END
  END qcpu_sram_in[6]
  PIN qcpu_sram_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 520.800 650.000 521.360 ;
    END
  END qcpu_sram_in[7]
  PIN qcpu_sram_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 525.280 650.000 525.840 ;
    END
  END qcpu_sram_out[0]
  PIN qcpu_sram_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 529.760 650.000 530.320 ;
    END
  END qcpu_sram_out[1]
  PIN qcpu_sram_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 534.240 650.000 534.800 ;
    END
  END qcpu_sram_out[2]
  PIN qcpu_sram_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 538.720 650.000 539.280 ;
    END
  END qcpu_sram_out[3]
  PIN qcpu_sram_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 543.200 650.000 543.760 ;
    END
  END qcpu_sram_out[4]
  PIN qcpu_sram_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 547.680 650.000 548.240 ;
    END
  END qcpu_sram_out[5]
  PIN qcpu_sram_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 552.160 650.000 552.720 ;
    END
  END qcpu_sram_out[6]
  PIN qcpu_sram_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 556.640 650.000 557.200 ;
    END
  END qcpu_sram_out[7]
  PIN rst_ay8913
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 561.120 650.000 561.680 ;
    END
  END rst_ay8913
  PIN rst_blinker
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 395.360 596.000 395.920 600.000 ;
    END
  END rst_blinker
  PIN rst_hellorld
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 560.000 4.000 560.560 ;
    END
  END rst_hellorld
  PIN rst_mc14500
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 380.800 4.000 381.360 ;
    END
  END rst_mc14500
  PIN rst_qcpu
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 375.200 4.000 375.760 ;
    END
  END rst_qcpu
  PIN rst_sid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 246.400 4.000 246.960 ;
    END
  END rst_sid
  PIN rst_sn76489
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 413.280 596.000 413.840 600.000 ;
    END
  END rst_sn76489
  PIN sid_do[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 252.000 4.000 252.560 ;
    END
  END sid_do[0]
  PIN sid_do[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 308.000 4.000 308.560 ;
    END
  END sid_do[10]
  PIN sid_do[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 313.600 4.000 314.160 ;
    END
  END sid_do[11]
  PIN sid_do[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 319.200 4.000 319.760 ;
    END
  END sid_do[12]
  PIN sid_do[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 324.800 4.000 325.360 ;
    END
  END sid_do[13]
  PIN sid_do[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 330.400 4.000 330.960 ;
    END
  END sid_do[14]
  PIN sid_do[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 336.000 4.000 336.560 ;
    END
  END sid_do[15]
  PIN sid_do[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 341.600 4.000 342.160 ;
    END
  END sid_do[16]
  PIN sid_do[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 347.200 4.000 347.760 ;
    END
  END sid_do[17]
  PIN sid_do[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 352.800 4.000 353.360 ;
    END
  END sid_do[18]
  PIN sid_do[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 358.400 4.000 358.960 ;
    END
  END sid_do[19]
  PIN sid_do[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 257.600 4.000 258.160 ;
    END
  END sid_do[1]
  PIN sid_do[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 364.000 4.000 364.560 ;
    END
  END sid_do[20]
  PIN sid_do[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 263.200 4.000 263.760 ;
    END
  END sid_do[2]
  PIN sid_do[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 268.800 4.000 269.360 ;
    END
  END sid_do[3]
  PIN sid_do[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 274.400 4.000 274.960 ;
    END
  END sid_do[4]
  PIN sid_do[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 280.000 4.000 280.560 ;
    END
  END sid_do[5]
  PIN sid_do[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 285.600 4.000 286.160 ;
    END
  END sid_do[6]
  PIN sid_do[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 291.200 4.000 291.760 ;
    END
  END sid_do[7]
  PIN sid_do[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 296.800 4.000 297.360 ;
    END
  END sid_do[8]
  PIN sid_do[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 302.400 4.000 302.960 ;
    END
  END sid_do[9]
  PIN sid_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 369.600 4.000 370.160 ;
    END
  END sid_oeb
  PIN sn76489_do[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 321.440 0.000 322.000 4.000 ;
    END
  END sn76489_do[0]
  PIN sn76489_do[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 366.240 0.000 366.800 4.000 ;
    END
  END sn76489_do[10]
  PIN sn76489_do[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 370.720 0.000 371.280 4.000 ;
    END
  END sn76489_do[11]
  PIN sn76489_do[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 375.200 0.000 375.760 4.000 ;
    END
  END sn76489_do[12]
  PIN sn76489_do[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 379.680 0.000 380.240 4.000 ;
    END
  END sn76489_do[13]
  PIN sn76489_do[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 384.160 0.000 384.720 4.000 ;
    END
  END sn76489_do[14]
  PIN sn76489_do[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 388.640 0.000 389.200 4.000 ;
    END
  END sn76489_do[15]
  PIN sn76489_do[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 393.120 0.000 393.680 4.000 ;
    END
  END sn76489_do[16]
  PIN sn76489_do[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 397.600 0.000 398.160 4.000 ;
    END
  END sn76489_do[17]
  PIN sn76489_do[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 402.080 0.000 402.640 4.000 ;
    END
  END sn76489_do[18]
  PIN sn76489_do[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 406.560 0.000 407.120 4.000 ;
    END
  END sn76489_do[19]
  PIN sn76489_do[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 325.920 0.000 326.480 4.000 ;
    END
  END sn76489_do[1]
  PIN sn76489_do[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 411.040 0.000 411.600 4.000 ;
    END
  END sn76489_do[20]
  PIN sn76489_do[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 415.520 0.000 416.080 4.000 ;
    END
  END sn76489_do[21]
  PIN sn76489_do[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 420.000 0.000 420.560 4.000 ;
    END
  END sn76489_do[22]
  PIN sn76489_do[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 424.480 0.000 425.040 4.000 ;
    END
  END sn76489_do[23]
  PIN sn76489_do[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 428.960 0.000 429.520 4.000 ;
    END
  END sn76489_do[24]
  PIN sn76489_do[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 433.440 0.000 434.000 4.000 ;
    END
  END sn76489_do[25]
  PIN sn76489_do[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 437.920 0.000 438.480 4.000 ;
    END
  END sn76489_do[26]
  PIN sn76489_do[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 442.400 0.000 442.960 4.000 ;
    END
  END sn76489_do[27]
  PIN sn76489_do[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 330.400 0.000 330.960 4.000 ;
    END
  END sn76489_do[2]
  PIN sn76489_do[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 334.880 0.000 335.440 4.000 ;
    END
  END sn76489_do[3]
  PIN sn76489_do[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 339.360 0.000 339.920 4.000 ;
    END
  END sn76489_do[4]
  PIN sn76489_do[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 343.840 0.000 344.400 4.000 ;
    END
  END sn76489_do[5]
  PIN sn76489_do[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 348.320 0.000 348.880 4.000 ;
    END
  END sn76489_do[6]
  PIN sn76489_do[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 352.800 0.000 353.360 4.000 ;
    END
  END sn76489_do[7]
  PIN sn76489_do[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 357.280 0.000 357.840 4.000 ;
    END
  END sn76489_do[8]
  PIN sn76489_do[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 361.760 0.000 362.320 4.000 ;
    END
  END sn76489_do[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 584.380 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 584.380 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 25.760 0.000 26.320 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 0.000 30.800 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 193.760 650.000 194.320 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 34.720 0.000 35.280 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 79.520 0.000 80.080 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 0.000 84.560 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 88.480 0.000 89.040 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 92.960 0.000 93.520 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 0.000 98.000 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 101.920 0.000 102.480 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 106.400 0.000 106.960 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 0.000 111.440 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 115.360 0.000 115.920 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 119.840 0.000 120.400 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 39.200 0.000 39.760 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 0.000 124.880 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 128.800 0.000 129.360 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 133.280 0.000 133.840 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 0.000 138.320 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 142.240 0.000 142.800 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 146.720 0.000 147.280 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 0.000 151.760 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 155.680 0.000 156.240 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 160.160 0.000 160.720 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 0.000 165.200 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 0.000 44.240 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 169.120 0.000 169.680 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 173.600 0.000 174.160 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 48.160 0.000 48.720 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 52.640 0.000 53.200 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 0.000 57.680 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 61.600 0.000 62.160 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 66.080 0.000 66.640 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 0.000 71.120 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 75.040 0.000 75.600 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 184.800 650.000 185.360 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 0.000 178.640 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 222.880 0.000 223.440 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 227.360 0.000 227.920 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 231.840 0.000 232.400 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 236.320 0.000 236.880 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 240.800 0.000 241.360 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 245.280 0.000 245.840 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 249.760 0.000 250.320 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 254.240 0.000 254.800 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 0.000 259.280 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 263.200 0.000 263.760 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 182.560 0.000 183.120 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 267.680 0.000 268.240 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 272.160 0.000 272.720 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 276.640 0.000 277.200 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 281.120 0.000 281.680 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 285.600 0.000 286.160 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 290.080 0.000 290.640 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 294.560 0.000 295.120 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 299.040 0.000 299.600 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 303.520 0.000 304.080 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 308.000 0.000 308.560 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 187.040 0.000 187.600 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 312.480 0.000 313.040 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 316.960 0.000 317.520 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 0.000 192.080 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 196.000 0.000 196.560 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 200.480 0.000 201.040 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 0.000 205.520 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 209.440 0.000 210.000 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 213.920 0.000 214.480 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 0.000 218.960 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 36.960 650.000 37.520 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 81.760 650.000 82.320 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 86.240 650.000 86.800 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 90.720 650.000 91.280 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 95.200 650.000 95.760 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 99.680 650.000 100.240 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 104.160 650.000 104.720 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 108.640 650.000 109.200 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 113.120 650.000 113.680 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 117.600 650.000 118.160 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 122.080 650.000 122.640 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 41.440 650.000 42.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 126.560 650.000 127.120 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 131.040 650.000 131.600 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 135.520 650.000 136.080 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 140.000 650.000 140.560 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 144.480 650.000 145.040 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 148.960 650.000 149.520 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 153.440 650.000 154.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 157.920 650.000 158.480 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 162.400 650.000 162.960 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 166.880 650.000 167.440 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 45.920 650.000 46.480 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 171.360 650.000 171.920 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 175.840 650.000 176.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 50.400 650.000 50.960 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 54.880 650.000 55.440 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 59.360 650.000 59.920 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 63.840 650.000 64.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 68.320 650.000 68.880 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 72.800 650.000 73.360 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 77.280 650.000 77.840 ;
    END
  END wbs_dat_o[9]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 189.280 650.000 189.840 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 646.000 180.320 650.000 180.880 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 14.150 642.880 586.730 ;
      LAYER Metal2 ;
        RECT 5.740 595.700 41.140 596.820 ;
        RECT 42.300 595.700 45.620 596.820 ;
        RECT 46.780 595.700 50.100 596.820 ;
        RECT 51.260 595.700 54.580 596.820 ;
        RECT 55.740 595.700 59.060 596.820 ;
        RECT 60.220 595.700 63.540 596.820 ;
        RECT 64.700 595.700 68.020 596.820 ;
        RECT 69.180 595.700 72.500 596.820 ;
        RECT 73.660 595.700 76.980 596.820 ;
        RECT 78.140 595.700 81.460 596.820 ;
        RECT 82.620 595.700 85.940 596.820 ;
        RECT 87.100 595.700 90.420 596.820 ;
        RECT 91.580 595.700 94.900 596.820 ;
        RECT 96.060 595.700 99.380 596.820 ;
        RECT 100.540 595.700 103.860 596.820 ;
        RECT 105.020 595.700 108.340 596.820 ;
        RECT 109.500 595.700 112.820 596.820 ;
        RECT 113.980 595.700 117.300 596.820 ;
        RECT 118.460 595.700 121.780 596.820 ;
        RECT 122.940 595.700 126.260 596.820 ;
        RECT 127.420 595.700 130.740 596.820 ;
        RECT 131.900 595.700 135.220 596.820 ;
        RECT 136.380 595.700 139.700 596.820 ;
        RECT 140.860 595.700 144.180 596.820 ;
        RECT 145.340 595.700 148.660 596.820 ;
        RECT 149.820 595.700 153.140 596.820 ;
        RECT 154.300 595.700 157.620 596.820 ;
        RECT 158.780 595.700 162.100 596.820 ;
        RECT 163.260 595.700 166.580 596.820 ;
        RECT 167.740 595.700 171.060 596.820 ;
        RECT 172.220 595.700 175.540 596.820 ;
        RECT 176.700 595.700 180.020 596.820 ;
        RECT 181.180 595.700 184.500 596.820 ;
        RECT 185.660 595.700 188.980 596.820 ;
        RECT 190.140 595.700 193.460 596.820 ;
        RECT 194.620 595.700 197.940 596.820 ;
        RECT 199.100 595.700 202.420 596.820 ;
        RECT 203.580 595.700 206.900 596.820 ;
        RECT 208.060 595.700 211.380 596.820 ;
        RECT 212.540 595.700 215.860 596.820 ;
        RECT 217.020 595.700 220.340 596.820 ;
        RECT 221.500 595.700 224.820 596.820 ;
        RECT 225.980 595.700 229.300 596.820 ;
        RECT 230.460 595.700 233.780 596.820 ;
        RECT 234.940 595.700 238.260 596.820 ;
        RECT 239.420 595.700 242.740 596.820 ;
        RECT 243.900 595.700 247.220 596.820 ;
        RECT 248.380 595.700 251.700 596.820 ;
        RECT 252.860 595.700 256.180 596.820 ;
        RECT 257.340 595.700 260.660 596.820 ;
        RECT 261.820 595.700 265.140 596.820 ;
        RECT 266.300 595.700 269.620 596.820 ;
        RECT 270.780 595.700 274.100 596.820 ;
        RECT 275.260 595.700 278.580 596.820 ;
        RECT 279.740 595.700 283.060 596.820 ;
        RECT 284.220 595.700 287.540 596.820 ;
        RECT 288.700 595.700 292.020 596.820 ;
        RECT 293.180 595.700 296.500 596.820 ;
        RECT 297.660 595.700 300.980 596.820 ;
        RECT 302.140 595.700 305.460 596.820 ;
        RECT 306.620 595.700 309.940 596.820 ;
        RECT 311.100 595.700 314.420 596.820 ;
        RECT 315.580 595.700 318.900 596.820 ;
        RECT 320.060 595.700 323.380 596.820 ;
        RECT 324.540 595.700 327.860 596.820 ;
        RECT 329.020 595.700 332.340 596.820 ;
        RECT 333.500 595.700 336.820 596.820 ;
        RECT 337.980 595.700 341.300 596.820 ;
        RECT 342.460 595.700 345.780 596.820 ;
        RECT 346.940 595.700 350.260 596.820 ;
        RECT 351.420 595.700 354.740 596.820 ;
        RECT 355.900 595.700 359.220 596.820 ;
        RECT 360.380 595.700 363.700 596.820 ;
        RECT 364.860 595.700 368.180 596.820 ;
        RECT 369.340 595.700 372.660 596.820 ;
        RECT 373.820 595.700 377.140 596.820 ;
        RECT 378.300 595.700 381.620 596.820 ;
        RECT 382.780 595.700 386.100 596.820 ;
        RECT 387.260 595.700 390.580 596.820 ;
        RECT 391.740 595.700 395.060 596.820 ;
        RECT 396.220 595.700 399.540 596.820 ;
        RECT 400.700 595.700 404.020 596.820 ;
        RECT 405.180 595.700 408.500 596.820 ;
        RECT 409.660 595.700 412.980 596.820 ;
        RECT 414.140 595.700 417.460 596.820 ;
        RECT 418.620 595.700 421.940 596.820 ;
        RECT 423.100 595.700 426.420 596.820 ;
        RECT 427.580 595.700 430.900 596.820 ;
        RECT 432.060 595.700 435.380 596.820 ;
        RECT 436.540 595.700 439.860 596.820 ;
        RECT 441.020 595.700 444.340 596.820 ;
        RECT 445.500 595.700 448.820 596.820 ;
        RECT 449.980 595.700 453.300 596.820 ;
        RECT 454.460 595.700 457.780 596.820 ;
        RECT 458.940 595.700 462.260 596.820 ;
        RECT 463.420 595.700 466.740 596.820 ;
        RECT 467.900 595.700 471.220 596.820 ;
        RECT 472.380 595.700 475.700 596.820 ;
        RECT 476.860 595.700 480.180 596.820 ;
        RECT 481.340 595.700 484.660 596.820 ;
        RECT 485.820 595.700 489.140 596.820 ;
        RECT 490.300 595.700 493.620 596.820 ;
        RECT 494.780 595.700 498.100 596.820 ;
        RECT 499.260 595.700 502.580 596.820 ;
        RECT 503.740 595.700 507.060 596.820 ;
        RECT 508.220 595.700 511.540 596.820 ;
        RECT 512.700 595.700 516.020 596.820 ;
        RECT 517.180 595.700 520.500 596.820 ;
        RECT 521.660 595.700 524.980 596.820 ;
        RECT 526.140 595.700 529.460 596.820 ;
        RECT 530.620 595.700 533.940 596.820 ;
        RECT 535.100 595.700 538.420 596.820 ;
        RECT 539.580 595.700 542.900 596.820 ;
        RECT 544.060 595.700 547.380 596.820 ;
        RECT 548.540 595.700 551.860 596.820 ;
        RECT 553.020 595.700 556.340 596.820 ;
        RECT 557.500 595.700 560.820 596.820 ;
        RECT 561.980 595.700 565.300 596.820 ;
        RECT 566.460 595.700 569.780 596.820 ;
        RECT 570.940 595.700 574.260 596.820 ;
        RECT 575.420 595.700 578.740 596.820 ;
        RECT 579.900 595.700 583.220 596.820 ;
        RECT 584.380 595.700 587.700 596.820 ;
        RECT 588.860 595.700 592.180 596.820 ;
        RECT 593.340 595.700 596.660 596.820 ;
        RECT 597.820 595.700 601.140 596.820 ;
        RECT 602.300 595.700 605.620 596.820 ;
        RECT 606.780 595.700 644.420 596.820 ;
        RECT 5.740 4.300 644.420 595.700 ;
        RECT 5.740 3.500 25.460 4.300 ;
        RECT 26.620 3.500 29.940 4.300 ;
        RECT 31.100 3.500 34.420 4.300 ;
        RECT 35.580 3.500 38.900 4.300 ;
        RECT 40.060 3.500 43.380 4.300 ;
        RECT 44.540 3.500 47.860 4.300 ;
        RECT 49.020 3.500 52.340 4.300 ;
        RECT 53.500 3.500 56.820 4.300 ;
        RECT 57.980 3.500 61.300 4.300 ;
        RECT 62.460 3.500 65.780 4.300 ;
        RECT 66.940 3.500 70.260 4.300 ;
        RECT 71.420 3.500 74.740 4.300 ;
        RECT 75.900 3.500 79.220 4.300 ;
        RECT 80.380 3.500 83.700 4.300 ;
        RECT 84.860 3.500 88.180 4.300 ;
        RECT 89.340 3.500 92.660 4.300 ;
        RECT 93.820 3.500 97.140 4.300 ;
        RECT 98.300 3.500 101.620 4.300 ;
        RECT 102.780 3.500 106.100 4.300 ;
        RECT 107.260 3.500 110.580 4.300 ;
        RECT 111.740 3.500 115.060 4.300 ;
        RECT 116.220 3.500 119.540 4.300 ;
        RECT 120.700 3.500 124.020 4.300 ;
        RECT 125.180 3.500 128.500 4.300 ;
        RECT 129.660 3.500 132.980 4.300 ;
        RECT 134.140 3.500 137.460 4.300 ;
        RECT 138.620 3.500 141.940 4.300 ;
        RECT 143.100 3.500 146.420 4.300 ;
        RECT 147.580 3.500 150.900 4.300 ;
        RECT 152.060 3.500 155.380 4.300 ;
        RECT 156.540 3.500 159.860 4.300 ;
        RECT 161.020 3.500 164.340 4.300 ;
        RECT 165.500 3.500 168.820 4.300 ;
        RECT 169.980 3.500 173.300 4.300 ;
        RECT 174.460 3.500 177.780 4.300 ;
        RECT 178.940 3.500 182.260 4.300 ;
        RECT 183.420 3.500 186.740 4.300 ;
        RECT 187.900 3.500 191.220 4.300 ;
        RECT 192.380 3.500 195.700 4.300 ;
        RECT 196.860 3.500 200.180 4.300 ;
        RECT 201.340 3.500 204.660 4.300 ;
        RECT 205.820 3.500 209.140 4.300 ;
        RECT 210.300 3.500 213.620 4.300 ;
        RECT 214.780 3.500 218.100 4.300 ;
        RECT 219.260 3.500 222.580 4.300 ;
        RECT 223.740 3.500 227.060 4.300 ;
        RECT 228.220 3.500 231.540 4.300 ;
        RECT 232.700 3.500 236.020 4.300 ;
        RECT 237.180 3.500 240.500 4.300 ;
        RECT 241.660 3.500 244.980 4.300 ;
        RECT 246.140 3.500 249.460 4.300 ;
        RECT 250.620 3.500 253.940 4.300 ;
        RECT 255.100 3.500 258.420 4.300 ;
        RECT 259.580 3.500 262.900 4.300 ;
        RECT 264.060 3.500 267.380 4.300 ;
        RECT 268.540 3.500 271.860 4.300 ;
        RECT 273.020 3.500 276.340 4.300 ;
        RECT 277.500 3.500 280.820 4.300 ;
        RECT 281.980 3.500 285.300 4.300 ;
        RECT 286.460 3.500 289.780 4.300 ;
        RECT 290.940 3.500 294.260 4.300 ;
        RECT 295.420 3.500 298.740 4.300 ;
        RECT 299.900 3.500 303.220 4.300 ;
        RECT 304.380 3.500 307.700 4.300 ;
        RECT 308.860 3.500 312.180 4.300 ;
        RECT 313.340 3.500 316.660 4.300 ;
        RECT 317.820 3.500 321.140 4.300 ;
        RECT 322.300 3.500 325.620 4.300 ;
        RECT 326.780 3.500 330.100 4.300 ;
        RECT 331.260 3.500 334.580 4.300 ;
        RECT 335.740 3.500 339.060 4.300 ;
        RECT 340.220 3.500 343.540 4.300 ;
        RECT 344.700 3.500 348.020 4.300 ;
        RECT 349.180 3.500 352.500 4.300 ;
        RECT 353.660 3.500 356.980 4.300 ;
        RECT 358.140 3.500 361.460 4.300 ;
        RECT 362.620 3.500 365.940 4.300 ;
        RECT 367.100 3.500 370.420 4.300 ;
        RECT 371.580 3.500 374.900 4.300 ;
        RECT 376.060 3.500 379.380 4.300 ;
        RECT 380.540 3.500 383.860 4.300 ;
        RECT 385.020 3.500 388.340 4.300 ;
        RECT 389.500 3.500 392.820 4.300 ;
        RECT 393.980 3.500 397.300 4.300 ;
        RECT 398.460 3.500 401.780 4.300 ;
        RECT 402.940 3.500 406.260 4.300 ;
        RECT 407.420 3.500 410.740 4.300 ;
        RECT 411.900 3.500 415.220 4.300 ;
        RECT 416.380 3.500 419.700 4.300 ;
        RECT 420.860 3.500 424.180 4.300 ;
        RECT 425.340 3.500 428.660 4.300 ;
        RECT 429.820 3.500 433.140 4.300 ;
        RECT 434.300 3.500 437.620 4.300 ;
        RECT 438.780 3.500 442.100 4.300 ;
        RECT 443.260 3.500 446.580 4.300 ;
        RECT 447.740 3.500 451.060 4.300 ;
        RECT 452.220 3.500 455.540 4.300 ;
        RECT 456.700 3.500 460.020 4.300 ;
        RECT 461.180 3.500 464.500 4.300 ;
        RECT 465.660 3.500 468.980 4.300 ;
        RECT 470.140 3.500 473.460 4.300 ;
        RECT 474.620 3.500 477.940 4.300 ;
        RECT 479.100 3.500 482.420 4.300 ;
        RECT 483.580 3.500 486.900 4.300 ;
        RECT 488.060 3.500 491.380 4.300 ;
        RECT 492.540 3.500 495.860 4.300 ;
        RECT 497.020 3.500 500.340 4.300 ;
        RECT 501.500 3.500 504.820 4.300 ;
        RECT 505.980 3.500 509.300 4.300 ;
        RECT 510.460 3.500 513.780 4.300 ;
        RECT 514.940 3.500 518.260 4.300 ;
        RECT 519.420 3.500 522.740 4.300 ;
        RECT 523.900 3.500 527.220 4.300 ;
        RECT 528.380 3.500 531.700 4.300 ;
        RECT 532.860 3.500 536.180 4.300 ;
        RECT 537.340 3.500 540.660 4.300 ;
        RECT 541.820 3.500 545.140 4.300 ;
        RECT 546.300 3.500 549.620 4.300 ;
        RECT 550.780 3.500 554.100 4.300 ;
        RECT 555.260 3.500 558.580 4.300 ;
        RECT 559.740 3.500 563.060 4.300 ;
        RECT 564.220 3.500 567.540 4.300 ;
        RECT 568.700 3.500 572.020 4.300 ;
        RECT 573.180 3.500 576.500 4.300 ;
        RECT 577.660 3.500 580.980 4.300 ;
        RECT 582.140 3.500 585.460 4.300 ;
        RECT 586.620 3.500 589.940 4.300 ;
        RECT 591.100 3.500 594.420 4.300 ;
        RECT 595.580 3.500 598.900 4.300 ;
        RECT 600.060 3.500 603.380 4.300 ;
        RECT 604.540 3.500 607.860 4.300 ;
        RECT 609.020 3.500 612.340 4.300 ;
        RECT 613.500 3.500 616.820 4.300 ;
        RECT 617.980 3.500 621.300 4.300 ;
        RECT 622.460 3.500 644.420 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 566.460 646.660 590.660 ;
        RECT 4.300 565.300 646.660 566.460 ;
        RECT 4.000 561.980 646.660 565.300 ;
        RECT 4.000 560.860 645.700 561.980 ;
        RECT 4.300 560.820 645.700 560.860 ;
        RECT 4.300 559.700 646.660 560.820 ;
        RECT 4.000 557.500 646.660 559.700 ;
        RECT 4.000 556.340 645.700 557.500 ;
        RECT 4.000 555.260 646.660 556.340 ;
        RECT 4.300 554.100 646.660 555.260 ;
        RECT 4.000 553.020 646.660 554.100 ;
        RECT 4.000 551.860 645.700 553.020 ;
        RECT 4.000 549.660 646.660 551.860 ;
        RECT 4.300 548.540 646.660 549.660 ;
        RECT 4.300 548.500 645.700 548.540 ;
        RECT 4.000 547.380 645.700 548.500 ;
        RECT 4.000 544.060 646.660 547.380 ;
        RECT 4.300 542.900 645.700 544.060 ;
        RECT 4.000 539.580 646.660 542.900 ;
        RECT 4.000 538.460 645.700 539.580 ;
        RECT 4.300 538.420 645.700 538.460 ;
        RECT 4.300 537.300 646.660 538.420 ;
        RECT 4.000 535.100 646.660 537.300 ;
        RECT 4.000 533.940 645.700 535.100 ;
        RECT 4.000 532.860 646.660 533.940 ;
        RECT 4.300 531.700 646.660 532.860 ;
        RECT 4.000 530.620 646.660 531.700 ;
        RECT 4.000 529.460 645.700 530.620 ;
        RECT 4.000 527.260 646.660 529.460 ;
        RECT 4.300 526.140 646.660 527.260 ;
        RECT 4.300 526.100 645.700 526.140 ;
        RECT 4.000 524.980 645.700 526.100 ;
        RECT 4.000 521.660 646.660 524.980 ;
        RECT 4.300 520.500 645.700 521.660 ;
        RECT 4.000 517.180 646.660 520.500 ;
        RECT 4.000 516.060 645.700 517.180 ;
        RECT 4.300 516.020 645.700 516.060 ;
        RECT 4.300 514.900 646.660 516.020 ;
        RECT 4.000 512.700 646.660 514.900 ;
        RECT 4.000 511.540 645.700 512.700 ;
        RECT 4.000 510.460 646.660 511.540 ;
        RECT 4.300 509.300 646.660 510.460 ;
        RECT 4.000 508.220 646.660 509.300 ;
        RECT 4.000 507.060 645.700 508.220 ;
        RECT 4.000 504.860 646.660 507.060 ;
        RECT 4.300 503.740 646.660 504.860 ;
        RECT 4.300 503.700 645.700 503.740 ;
        RECT 4.000 502.580 645.700 503.700 ;
        RECT 4.000 499.260 646.660 502.580 ;
        RECT 4.300 498.100 645.700 499.260 ;
        RECT 4.000 494.780 646.660 498.100 ;
        RECT 4.000 493.660 645.700 494.780 ;
        RECT 4.300 493.620 645.700 493.660 ;
        RECT 4.300 492.500 646.660 493.620 ;
        RECT 4.000 490.300 646.660 492.500 ;
        RECT 4.000 489.140 645.700 490.300 ;
        RECT 4.000 488.060 646.660 489.140 ;
        RECT 4.300 486.900 646.660 488.060 ;
        RECT 4.000 485.820 646.660 486.900 ;
        RECT 4.000 484.660 645.700 485.820 ;
        RECT 4.000 482.460 646.660 484.660 ;
        RECT 4.300 481.340 646.660 482.460 ;
        RECT 4.300 481.300 645.700 481.340 ;
        RECT 4.000 480.180 645.700 481.300 ;
        RECT 4.000 476.860 646.660 480.180 ;
        RECT 4.300 475.700 645.700 476.860 ;
        RECT 4.000 472.380 646.660 475.700 ;
        RECT 4.000 471.260 645.700 472.380 ;
        RECT 4.300 471.220 645.700 471.260 ;
        RECT 4.300 470.100 646.660 471.220 ;
        RECT 4.000 467.900 646.660 470.100 ;
        RECT 4.000 466.740 645.700 467.900 ;
        RECT 4.000 465.660 646.660 466.740 ;
        RECT 4.300 464.500 646.660 465.660 ;
        RECT 4.000 463.420 646.660 464.500 ;
        RECT 4.000 462.260 645.700 463.420 ;
        RECT 4.000 460.060 646.660 462.260 ;
        RECT 4.300 458.940 646.660 460.060 ;
        RECT 4.300 458.900 645.700 458.940 ;
        RECT 4.000 457.780 645.700 458.900 ;
        RECT 4.000 454.460 646.660 457.780 ;
        RECT 4.300 453.300 645.700 454.460 ;
        RECT 4.000 449.980 646.660 453.300 ;
        RECT 4.000 448.860 645.700 449.980 ;
        RECT 4.300 448.820 645.700 448.860 ;
        RECT 4.300 447.700 646.660 448.820 ;
        RECT 4.000 445.500 646.660 447.700 ;
        RECT 4.000 444.340 645.700 445.500 ;
        RECT 4.000 443.260 646.660 444.340 ;
        RECT 4.300 442.100 646.660 443.260 ;
        RECT 4.000 441.020 646.660 442.100 ;
        RECT 4.000 439.860 645.700 441.020 ;
        RECT 4.000 437.660 646.660 439.860 ;
        RECT 4.300 436.540 646.660 437.660 ;
        RECT 4.300 436.500 645.700 436.540 ;
        RECT 4.000 435.380 645.700 436.500 ;
        RECT 4.000 432.060 646.660 435.380 ;
        RECT 4.300 430.900 645.700 432.060 ;
        RECT 4.000 427.580 646.660 430.900 ;
        RECT 4.000 426.460 645.700 427.580 ;
        RECT 4.300 426.420 645.700 426.460 ;
        RECT 4.300 425.300 646.660 426.420 ;
        RECT 4.000 423.100 646.660 425.300 ;
        RECT 4.000 421.940 645.700 423.100 ;
        RECT 4.000 420.860 646.660 421.940 ;
        RECT 4.300 419.700 646.660 420.860 ;
        RECT 4.000 418.620 646.660 419.700 ;
        RECT 4.000 417.460 645.700 418.620 ;
        RECT 4.000 415.260 646.660 417.460 ;
        RECT 4.300 414.140 646.660 415.260 ;
        RECT 4.300 414.100 645.700 414.140 ;
        RECT 4.000 412.980 645.700 414.100 ;
        RECT 4.000 409.660 646.660 412.980 ;
        RECT 4.300 408.500 645.700 409.660 ;
        RECT 4.000 405.180 646.660 408.500 ;
        RECT 4.000 404.060 645.700 405.180 ;
        RECT 4.300 404.020 645.700 404.060 ;
        RECT 4.300 402.900 646.660 404.020 ;
        RECT 4.000 400.700 646.660 402.900 ;
        RECT 4.000 399.540 645.700 400.700 ;
        RECT 4.000 398.460 646.660 399.540 ;
        RECT 4.300 397.300 646.660 398.460 ;
        RECT 4.000 396.220 646.660 397.300 ;
        RECT 4.000 395.060 645.700 396.220 ;
        RECT 4.000 392.860 646.660 395.060 ;
        RECT 4.300 391.740 646.660 392.860 ;
        RECT 4.300 391.700 645.700 391.740 ;
        RECT 4.000 390.580 645.700 391.700 ;
        RECT 4.000 387.260 646.660 390.580 ;
        RECT 4.300 386.100 645.700 387.260 ;
        RECT 4.000 382.780 646.660 386.100 ;
        RECT 4.000 381.660 645.700 382.780 ;
        RECT 4.300 381.620 645.700 381.660 ;
        RECT 4.300 380.500 646.660 381.620 ;
        RECT 4.000 378.300 646.660 380.500 ;
        RECT 4.000 377.140 645.700 378.300 ;
        RECT 4.000 376.060 646.660 377.140 ;
        RECT 4.300 374.900 646.660 376.060 ;
        RECT 4.000 373.820 646.660 374.900 ;
        RECT 4.000 372.660 645.700 373.820 ;
        RECT 4.000 370.460 646.660 372.660 ;
        RECT 4.300 369.340 646.660 370.460 ;
        RECT 4.300 369.300 645.700 369.340 ;
        RECT 4.000 368.180 645.700 369.300 ;
        RECT 4.000 364.860 646.660 368.180 ;
        RECT 4.300 363.700 645.700 364.860 ;
        RECT 4.000 360.380 646.660 363.700 ;
        RECT 4.000 359.260 645.700 360.380 ;
        RECT 4.300 359.220 645.700 359.260 ;
        RECT 4.300 358.100 646.660 359.220 ;
        RECT 4.000 355.900 646.660 358.100 ;
        RECT 4.000 354.740 645.700 355.900 ;
        RECT 4.000 353.660 646.660 354.740 ;
        RECT 4.300 352.500 646.660 353.660 ;
        RECT 4.000 351.420 646.660 352.500 ;
        RECT 4.000 350.260 645.700 351.420 ;
        RECT 4.000 348.060 646.660 350.260 ;
        RECT 4.300 346.940 646.660 348.060 ;
        RECT 4.300 346.900 645.700 346.940 ;
        RECT 4.000 345.780 645.700 346.900 ;
        RECT 4.000 342.460 646.660 345.780 ;
        RECT 4.300 341.300 645.700 342.460 ;
        RECT 4.000 337.980 646.660 341.300 ;
        RECT 4.000 336.860 645.700 337.980 ;
        RECT 4.300 336.820 645.700 336.860 ;
        RECT 4.300 335.700 646.660 336.820 ;
        RECT 4.000 333.500 646.660 335.700 ;
        RECT 4.000 332.340 645.700 333.500 ;
        RECT 4.000 331.260 646.660 332.340 ;
        RECT 4.300 330.100 646.660 331.260 ;
        RECT 4.000 329.020 646.660 330.100 ;
        RECT 4.000 327.860 645.700 329.020 ;
        RECT 4.000 325.660 646.660 327.860 ;
        RECT 4.300 324.540 646.660 325.660 ;
        RECT 4.300 324.500 645.700 324.540 ;
        RECT 4.000 323.380 645.700 324.500 ;
        RECT 4.000 320.060 646.660 323.380 ;
        RECT 4.300 318.900 645.700 320.060 ;
        RECT 4.000 315.580 646.660 318.900 ;
        RECT 4.000 314.460 645.700 315.580 ;
        RECT 4.300 314.420 645.700 314.460 ;
        RECT 4.300 313.300 646.660 314.420 ;
        RECT 4.000 311.100 646.660 313.300 ;
        RECT 4.000 309.940 645.700 311.100 ;
        RECT 4.000 308.860 646.660 309.940 ;
        RECT 4.300 307.700 646.660 308.860 ;
        RECT 4.000 306.620 646.660 307.700 ;
        RECT 4.000 305.460 645.700 306.620 ;
        RECT 4.000 303.260 646.660 305.460 ;
        RECT 4.300 302.140 646.660 303.260 ;
        RECT 4.300 302.100 645.700 302.140 ;
        RECT 4.000 300.980 645.700 302.100 ;
        RECT 4.000 297.660 646.660 300.980 ;
        RECT 4.300 296.500 645.700 297.660 ;
        RECT 4.000 293.180 646.660 296.500 ;
        RECT 4.000 292.060 645.700 293.180 ;
        RECT 4.300 292.020 645.700 292.060 ;
        RECT 4.300 290.900 646.660 292.020 ;
        RECT 4.000 288.700 646.660 290.900 ;
        RECT 4.000 287.540 645.700 288.700 ;
        RECT 4.000 286.460 646.660 287.540 ;
        RECT 4.300 285.300 646.660 286.460 ;
        RECT 4.000 284.220 646.660 285.300 ;
        RECT 4.000 283.060 645.700 284.220 ;
        RECT 4.000 280.860 646.660 283.060 ;
        RECT 4.300 279.740 646.660 280.860 ;
        RECT 4.300 279.700 645.700 279.740 ;
        RECT 4.000 278.580 645.700 279.700 ;
        RECT 4.000 275.260 646.660 278.580 ;
        RECT 4.300 274.100 645.700 275.260 ;
        RECT 4.000 270.780 646.660 274.100 ;
        RECT 4.000 269.660 645.700 270.780 ;
        RECT 4.300 269.620 645.700 269.660 ;
        RECT 4.300 268.500 646.660 269.620 ;
        RECT 4.000 266.300 646.660 268.500 ;
        RECT 4.000 265.140 645.700 266.300 ;
        RECT 4.000 264.060 646.660 265.140 ;
        RECT 4.300 262.900 646.660 264.060 ;
        RECT 4.000 261.820 646.660 262.900 ;
        RECT 4.000 260.660 645.700 261.820 ;
        RECT 4.000 258.460 646.660 260.660 ;
        RECT 4.300 257.340 646.660 258.460 ;
        RECT 4.300 257.300 645.700 257.340 ;
        RECT 4.000 256.180 645.700 257.300 ;
        RECT 4.000 252.860 646.660 256.180 ;
        RECT 4.300 251.700 645.700 252.860 ;
        RECT 4.000 248.380 646.660 251.700 ;
        RECT 4.000 247.260 645.700 248.380 ;
        RECT 4.300 247.220 645.700 247.260 ;
        RECT 4.300 246.100 646.660 247.220 ;
        RECT 4.000 243.900 646.660 246.100 ;
        RECT 4.000 242.740 645.700 243.900 ;
        RECT 4.000 241.660 646.660 242.740 ;
        RECT 4.300 240.500 646.660 241.660 ;
        RECT 4.000 239.420 646.660 240.500 ;
        RECT 4.000 238.260 645.700 239.420 ;
        RECT 4.000 236.060 646.660 238.260 ;
        RECT 4.300 234.940 646.660 236.060 ;
        RECT 4.300 234.900 645.700 234.940 ;
        RECT 4.000 233.780 645.700 234.900 ;
        RECT 4.000 230.460 646.660 233.780 ;
        RECT 4.300 229.300 645.700 230.460 ;
        RECT 4.000 225.980 646.660 229.300 ;
        RECT 4.000 224.860 645.700 225.980 ;
        RECT 4.300 224.820 645.700 224.860 ;
        RECT 4.300 223.700 646.660 224.820 ;
        RECT 4.000 221.500 646.660 223.700 ;
        RECT 4.000 220.340 645.700 221.500 ;
        RECT 4.000 219.260 646.660 220.340 ;
        RECT 4.300 218.100 646.660 219.260 ;
        RECT 4.000 217.020 646.660 218.100 ;
        RECT 4.000 215.860 645.700 217.020 ;
        RECT 4.000 213.660 646.660 215.860 ;
        RECT 4.300 212.540 646.660 213.660 ;
        RECT 4.300 212.500 645.700 212.540 ;
        RECT 4.000 211.380 645.700 212.500 ;
        RECT 4.000 208.060 646.660 211.380 ;
        RECT 4.300 206.900 645.700 208.060 ;
        RECT 4.000 203.580 646.660 206.900 ;
        RECT 4.000 202.460 645.700 203.580 ;
        RECT 4.300 202.420 645.700 202.460 ;
        RECT 4.300 201.300 646.660 202.420 ;
        RECT 4.000 199.100 646.660 201.300 ;
        RECT 4.000 197.940 645.700 199.100 ;
        RECT 4.000 196.860 646.660 197.940 ;
        RECT 4.300 195.700 646.660 196.860 ;
        RECT 4.000 194.620 646.660 195.700 ;
        RECT 4.000 193.460 645.700 194.620 ;
        RECT 4.000 191.260 646.660 193.460 ;
        RECT 4.300 190.140 646.660 191.260 ;
        RECT 4.300 190.100 645.700 190.140 ;
        RECT 4.000 188.980 645.700 190.100 ;
        RECT 4.000 185.660 646.660 188.980 ;
        RECT 4.300 184.500 645.700 185.660 ;
        RECT 4.000 181.180 646.660 184.500 ;
        RECT 4.000 180.060 645.700 181.180 ;
        RECT 4.300 180.020 645.700 180.060 ;
        RECT 4.300 178.900 646.660 180.020 ;
        RECT 4.000 176.700 646.660 178.900 ;
        RECT 4.000 175.540 645.700 176.700 ;
        RECT 4.000 174.460 646.660 175.540 ;
        RECT 4.300 173.300 646.660 174.460 ;
        RECT 4.000 172.220 646.660 173.300 ;
        RECT 4.000 171.060 645.700 172.220 ;
        RECT 4.000 168.860 646.660 171.060 ;
        RECT 4.300 167.740 646.660 168.860 ;
        RECT 4.300 167.700 645.700 167.740 ;
        RECT 4.000 166.580 645.700 167.700 ;
        RECT 4.000 163.260 646.660 166.580 ;
        RECT 4.300 162.100 645.700 163.260 ;
        RECT 4.000 158.780 646.660 162.100 ;
        RECT 4.000 157.660 645.700 158.780 ;
        RECT 4.300 157.620 645.700 157.660 ;
        RECT 4.300 156.500 646.660 157.620 ;
        RECT 4.000 154.300 646.660 156.500 ;
        RECT 4.000 153.140 645.700 154.300 ;
        RECT 4.000 152.060 646.660 153.140 ;
        RECT 4.300 150.900 646.660 152.060 ;
        RECT 4.000 149.820 646.660 150.900 ;
        RECT 4.000 148.660 645.700 149.820 ;
        RECT 4.000 146.460 646.660 148.660 ;
        RECT 4.300 145.340 646.660 146.460 ;
        RECT 4.300 145.300 645.700 145.340 ;
        RECT 4.000 144.180 645.700 145.300 ;
        RECT 4.000 140.860 646.660 144.180 ;
        RECT 4.300 139.700 645.700 140.860 ;
        RECT 4.000 136.380 646.660 139.700 ;
        RECT 4.000 135.260 645.700 136.380 ;
        RECT 4.300 135.220 645.700 135.260 ;
        RECT 4.300 134.100 646.660 135.220 ;
        RECT 4.000 131.900 646.660 134.100 ;
        RECT 4.000 130.740 645.700 131.900 ;
        RECT 4.000 129.660 646.660 130.740 ;
        RECT 4.300 128.500 646.660 129.660 ;
        RECT 4.000 127.420 646.660 128.500 ;
        RECT 4.000 126.260 645.700 127.420 ;
        RECT 4.000 124.060 646.660 126.260 ;
        RECT 4.300 122.940 646.660 124.060 ;
        RECT 4.300 122.900 645.700 122.940 ;
        RECT 4.000 121.780 645.700 122.900 ;
        RECT 4.000 118.460 646.660 121.780 ;
        RECT 4.300 117.300 645.700 118.460 ;
        RECT 4.000 113.980 646.660 117.300 ;
        RECT 4.000 112.860 645.700 113.980 ;
        RECT 4.300 112.820 645.700 112.860 ;
        RECT 4.300 111.700 646.660 112.820 ;
        RECT 4.000 109.500 646.660 111.700 ;
        RECT 4.000 108.340 645.700 109.500 ;
        RECT 4.000 107.260 646.660 108.340 ;
        RECT 4.300 106.100 646.660 107.260 ;
        RECT 4.000 105.020 646.660 106.100 ;
        RECT 4.000 103.860 645.700 105.020 ;
        RECT 4.000 101.660 646.660 103.860 ;
        RECT 4.300 100.540 646.660 101.660 ;
        RECT 4.300 100.500 645.700 100.540 ;
        RECT 4.000 99.380 645.700 100.500 ;
        RECT 4.000 96.060 646.660 99.380 ;
        RECT 4.300 94.900 645.700 96.060 ;
        RECT 4.000 91.580 646.660 94.900 ;
        RECT 4.000 90.460 645.700 91.580 ;
        RECT 4.300 90.420 645.700 90.460 ;
        RECT 4.300 89.300 646.660 90.420 ;
        RECT 4.000 87.100 646.660 89.300 ;
        RECT 4.000 85.940 645.700 87.100 ;
        RECT 4.000 84.860 646.660 85.940 ;
        RECT 4.300 83.700 646.660 84.860 ;
        RECT 4.000 82.620 646.660 83.700 ;
        RECT 4.000 81.460 645.700 82.620 ;
        RECT 4.000 79.260 646.660 81.460 ;
        RECT 4.300 78.140 646.660 79.260 ;
        RECT 4.300 78.100 645.700 78.140 ;
        RECT 4.000 76.980 645.700 78.100 ;
        RECT 4.000 73.660 646.660 76.980 ;
        RECT 4.300 72.500 645.700 73.660 ;
        RECT 4.000 69.180 646.660 72.500 ;
        RECT 4.000 68.060 645.700 69.180 ;
        RECT 4.300 68.020 645.700 68.060 ;
        RECT 4.300 66.900 646.660 68.020 ;
        RECT 4.000 64.700 646.660 66.900 ;
        RECT 4.000 63.540 645.700 64.700 ;
        RECT 4.000 62.460 646.660 63.540 ;
        RECT 4.300 61.300 646.660 62.460 ;
        RECT 4.000 60.220 646.660 61.300 ;
        RECT 4.000 59.060 645.700 60.220 ;
        RECT 4.000 56.860 646.660 59.060 ;
        RECT 4.300 55.740 646.660 56.860 ;
        RECT 4.300 55.700 645.700 55.740 ;
        RECT 4.000 54.580 645.700 55.700 ;
        RECT 4.000 51.260 646.660 54.580 ;
        RECT 4.300 50.100 645.700 51.260 ;
        RECT 4.000 46.780 646.660 50.100 ;
        RECT 4.000 45.660 645.700 46.780 ;
        RECT 4.300 45.620 645.700 45.660 ;
        RECT 4.300 44.500 646.660 45.620 ;
        RECT 4.000 42.300 646.660 44.500 ;
        RECT 4.000 41.140 645.700 42.300 ;
        RECT 4.000 40.060 646.660 41.140 ;
        RECT 4.300 38.900 646.660 40.060 ;
        RECT 4.000 37.820 646.660 38.900 ;
        RECT 4.000 36.660 645.700 37.820 ;
        RECT 4.000 34.460 646.660 36.660 ;
        RECT 4.300 33.300 646.660 34.460 ;
        RECT 4.000 6.860 646.660 33.300 ;
      LAYER Metal4 ;
        RECT 18.620 15.080 21.940 581.750 ;
        RECT 24.140 15.080 98.740 581.750 ;
        RECT 100.940 15.080 175.540 581.750 ;
        RECT 177.740 15.080 252.340 581.750 ;
        RECT 254.540 15.080 329.140 581.750 ;
        RECT 331.340 15.080 405.940 581.750 ;
        RECT 408.140 15.080 482.740 581.750 ;
        RECT 484.940 15.080 559.540 581.750 ;
        RECT 561.740 15.080 636.340 581.750 ;
        RECT 638.540 15.080 638.820 581.750 ;
        RECT 18.620 13.530 638.820 15.080 ;
  END
END multiplexer
END LIBRARY

