VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_sid
  CLASS BLOCK ;
  FOREIGN wrapped_sid ;
  ORIGIN 0.000 0.000 ;
  SIZE 1150.000 BY 750.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 17.920 1150.000 18.480 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 152.320 1150.000 152.880 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 165.760 1150.000 166.320 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 179.200 1150.000 179.760 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 192.640 1150.000 193.200 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 206.080 1150.000 206.640 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 219.520 1150.000 220.080 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 232.960 1150.000 233.520 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 246.400 1150.000 246.960 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 259.840 1150.000 260.400 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 273.280 1150.000 273.840 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 31.360 1150.000 31.920 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 286.720 1150.000 287.280 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 300.160 1150.000 300.720 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 313.600 1150.000 314.160 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 327.040 1150.000 327.600 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 340.480 1150.000 341.040 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 353.920 1150.000 354.480 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 367.360 1150.000 367.920 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 380.800 1150.000 381.360 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 394.240 1150.000 394.800 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 407.680 1150.000 408.240 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 44.800 1150.000 45.360 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 421.120 1150.000 421.680 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 434.560 1150.000 435.120 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 448.000 1150.000 448.560 ;
    END
  END io_in[32]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 58.240 1150.000 58.800 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 71.680 1150.000 72.240 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 85.120 1150.000 85.680 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 98.560 1150.000 99.120 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 112.000 1150.000 112.560 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 125.440 1150.000 126.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 138.880 1150.000 139.440 ;
    END
  END io_in[9]
  PIN io_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 574.560 746.000 575.120 750.000 ;
    END
  END io_oeb
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 461.440 1150.000 462.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 595.840 1150.000 596.400 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 609.280 1150.000 609.840 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 622.720 1150.000 623.280 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 636.160 1150.000 636.720 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 649.600 1150.000 650.160 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 663.040 1150.000 663.600 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 676.480 1150.000 677.040 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 689.920 1150.000 690.480 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 703.360 1150.000 703.920 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 716.800 1150.000 717.360 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 474.880 1150.000 475.440 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 730.240 1150.000 730.800 ;
    END
  END io_out[20]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 488.320 1150.000 488.880 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 501.760 1150.000 502.320 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 515.200 1150.000 515.760 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 528.640 1150.000 529.200 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 542.080 1150.000 542.640 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 555.520 1150.000 556.080 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 568.960 1150.000 569.520 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 582.400 1150.000 582.960 ;
    END
  END io_out[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 861.280 0.000 861.840 4.000 ;
    END
  END rst_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 733.340 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 733.340 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 286.720 0.000 287.280 4.000 ;
    END
  END wb_clk_i
  OBS
      LAYER Nwell ;
        RECT 6.290 730.880 1143.390 733.470 ;
      LAYER Pwell ;
        RECT 6.290 727.360 1143.390 730.880 ;
      LAYER Nwell ;
        RECT 6.290 727.235 99.550 727.360 ;
        RECT 6.290 723.165 1143.390 727.235 ;
        RECT 6.290 723.040 88.630 723.165 ;
      LAYER Pwell ;
        RECT 6.290 719.520 1143.390 723.040 ;
      LAYER Nwell ;
        RECT 6.290 719.395 151.630 719.520 ;
        RECT 6.290 715.325 1143.390 719.395 ;
        RECT 6.290 715.200 132.030 715.325 ;
      LAYER Pwell ;
        RECT 6.290 711.680 1143.390 715.200 ;
      LAYER Nwell ;
        RECT 6.290 711.555 62.585 711.680 ;
        RECT 6.290 707.485 1143.390 711.555 ;
        RECT 6.290 707.360 148.355 707.485 ;
      LAYER Pwell ;
        RECT 6.290 703.840 1143.390 707.360 ;
      LAYER Nwell ;
        RECT 6.290 703.715 57.830 703.840 ;
        RECT 6.290 699.645 1143.390 703.715 ;
        RECT 6.290 699.520 134.315 699.645 ;
      LAYER Pwell ;
        RECT 6.290 696.000 1143.390 699.520 ;
      LAYER Nwell ;
        RECT 6.290 695.875 69.870 696.000 ;
        RECT 6.290 691.805 1143.390 695.875 ;
        RECT 6.290 691.680 49.710 691.805 ;
      LAYER Pwell ;
        RECT 6.290 688.160 1143.390 691.680 ;
      LAYER Nwell ;
        RECT 6.290 688.035 283.790 688.160 ;
        RECT 6.290 683.965 1143.390 688.035 ;
        RECT 6.290 683.840 43.270 683.965 ;
      LAYER Pwell ;
        RECT 6.290 680.320 1143.390 683.840 ;
      LAYER Nwell ;
        RECT 6.290 680.195 126.990 680.320 ;
        RECT 6.290 676.125 1143.390 680.195 ;
        RECT 6.290 676.000 156.110 676.125 ;
      LAYER Pwell ;
        RECT 6.290 672.480 1143.390 676.000 ;
      LAYER Nwell ;
        RECT 6.290 672.355 48.590 672.480 ;
        RECT 6.290 668.285 1143.390 672.355 ;
        RECT 6.290 668.160 364.005 668.285 ;
      LAYER Pwell ;
        RECT 6.290 664.640 1143.390 668.160 ;
      LAYER Nwell ;
        RECT 6.290 664.515 205.435 664.640 ;
        RECT 6.290 660.445 1143.390 664.515 ;
        RECT 6.290 660.320 37.435 660.445 ;
      LAYER Pwell ;
        RECT 6.290 656.800 1143.390 660.320 ;
      LAYER Nwell ;
        RECT 6.290 656.675 48.635 656.800 ;
        RECT 6.290 652.605 1143.390 656.675 ;
        RECT 6.290 652.480 79.390 652.605 ;
      LAYER Pwell ;
        RECT 6.290 648.960 1143.390 652.480 ;
      LAYER Nwell ;
        RECT 6.290 648.835 60.910 648.960 ;
        RECT 6.290 644.765 1143.390 648.835 ;
        RECT 6.290 644.640 53.130 644.765 ;
      LAYER Pwell ;
        RECT 6.290 641.120 1143.390 644.640 ;
      LAYER Nwell ;
        RECT 6.290 640.995 48.590 641.120 ;
        RECT 6.290 636.925 1143.390 640.995 ;
        RECT 6.290 636.800 179.795 636.925 ;
      LAYER Pwell ;
        RECT 6.290 633.280 1143.390 636.800 ;
      LAYER Nwell ;
        RECT 6.290 633.155 62.310 633.280 ;
        RECT 6.290 629.085 1143.390 633.155 ;
        RECT 6.290 628.960 37.390 629.085 ;
      LAYER Pwell ;
        RECT 6.290 625.440 1143.390 628.960 ;
      LAYER Nwell ;
        RECT 6.290 625.315 56.430 625.440 ;
        RECT 6.290 621.245 1143.390 625.315 ;
        RECT 6.290 621.120 47.470 621.245 ;
      LAYER Pwell ;
        RECT 6.290 617.600 1143.390 621.120 ;
      LAYER Nwell ;
        RECT 6.290 617.475 182.710 617.600 ;
        RECT 6.290 613.405 1143.390 617.475 ;
        RECT 6.290 613.280 56.990 613.405 ;
      LAYER Pwell ;
        RECT 6.290 609.760 1143.390 613.280 ;
      LAYER Nwell ;
        RECT 6.290 609.635 40.810 609.760 ;
        RECT 6.290 605.565 1143.390 609.635 ;
        RECT 6.290 605.440 39.070 605.565 ;
      LAYER Pwell ;
        RECT 6.290 601.920 1143.390 605.440 ;
      LAYER Nwell ;
        RECT 6.290 601.795 87.790 601.920 ;
        RECT 6.290 597.725 1143.390 601.795 ;
        RECT 6.290 597.600 39.910 597.725 ;
      LAYER Pwell ;
        RECT 6.290 594.080 1143.390 597.600 ;
      LAYER Nwell ;
        RECT 6.290 593.955 50.875 594.080 ;
        RECT 6.290 589.885 1143.390 593.955 ;
        RECT 6.290 589.760 109.070 589.885 ;
      LAYER Pwell ;
        RECT 6.290 586.240 1143.390 589.760 ;
      LAYER Nwell ;
        RECT 6.290 586.115 77.150 586.240 ;
        RECT 6.290 582.045 1143.390 586.115 ;
        RECT 6.290 581.920 123.630 582.045 ;
      LAYER Pwell ;
        RECT 6.290 578.400 1143.390 581.920 ;
      LAYER Nwell ;
        RECT 6.290 578.275 92.875 578.400 ;
        RECT 6.290 574.205 1143.390 578.275 ;
        RECT 6.290 574.080 77.710 574.205 ;
      LAYER Pwell ;
        RECT 6.290 570.560 1143.390 574.080 ;
      LAYER Nwell ;
        RECT 6.290 570.435 69.590 570.560 ;
        RECT 6.290 566.365 1143.390 570.435 ;
        RECT 6.290 566.240 114.670 566.365 ;
      LAYER Pwell ;
        RECT 6.290 562.720 1143.390 566.240 ;
      LAYER Nwell ;
        RECT 6.290 562.595 41.030 562.720 ;
        RECT 6.290 558.525 1143.390 562.595 ;
        RECT 6.290 558.400 73.875 558.525 ;
      LAYER Pwell ;
        RECT 6.290 554.880 1143.390 558.400 ;
      LAYER Nwell ;
        RECT 6.290 554.755 49.760 554.880 ;
        RECT 6.290 550.685 1143.390 554.755 ;
        RECT 6.290 550.560 110.540 550.685 ;
      LAYER Pwell ;
        RECT 6.290 547.040 1143.390 550.560 ;
      LAYER Nwell ;
        RECT 6.290 546.915 219.110 547.040 ;
        RECT 6.290 542.845 1143.390 546.915 ;
        RECT 6.290 542.720 90.545 542.845 ;
      LAYER Pwell ;
        RECT 6.290 539.200 1143.390 542.720 ;
      LAYER Nwell ;
        RECT 6.290 539.075 32.305 539.200 ;
        RECT 6.290 535.005 1143.390 539.075 ;
        RECT 6.290 534.880 49.665 535.005 ;
      LAYER Pwell ;
        RECT 6.290 531.360 1143.390 534.880 ;
      LAYER Nwell ;
        RECT 6.290 531.235 17.185 531.360 ;
        RECT 6.290 527.165 1143.390 531.235 ;
        RECT 6.290 527.040 120.785 527.165 ;
      LAYER Pwell ;
        RECT 6.290 523.520 1143.390 527.040 ;
      LAYER Nwell ;
        RECT 6.290 523.395 12.705 523.520 ;
        RECT 6.290 519.325 1143.390 523.395 ;
        RECT 6.290 519.200 172.630 519.325 ;
      LAYER Pwell ;
        RECT 6.290 515.680 1143.390 519.200 ;
      LAYER Nwell ;
        RECT 6.290 515.555 13.825 515.680 ;
        RECT 6.290 511.485 1143.390 515.555 ;
        RECT 6.290 511.360 49.865 511.485 ;
      LAYER Pwell ;
        RECT 6.290 507.840 1143.390 511.360 ;
      LAYER Nwell ;
        RECT 6.290 507.715 50.305 507.840 ;
        RECT 6.290 503.645 1143.390 507.715 ;
        RECT 6.290 503.520 12.705 503.645 ;
      LAYER Pwell ;
        RECT 6.290 500.000 1143.390 503.520 ;
      LAYER Nwell ;
        RECT 6.290 499.875 36.830 500.000 ;
        RECT 6.290 495.805 1143.390 499.875 ;
        RECT 6.290 495.680 161.665 495.805 ;
      LAYER Pwell ;
        RECT 6.290 492.160 1143.390 495.680 ;
      LAYER Nwell ;
        RECT 6.290 492.035 102.700 492.160 ;
        RECT 6.290 487.965 1143.390 492.035 ;
        RECT 6.290 487.840 51.390 487.965 ;
      LAYER Pwell ;
        RECT 6.290 484.320 1143.390 487.840 ;
      LAYER Nwell ;
        RECT 6.290 484.195 48.635 484.320 ;
        RECT 6.290 480.125 1143.390 484.195 ;
        RECT 6.290 480.000 34.180 480.125 ;
      LAYER Pwell ;
        RECT 6.290 476.480 1143.390 480.000 ;
      LAYER Nwell ;
        RECT 6.290 476.355 12.705 476.480 ;
        RECT 6.290 472.285 1143.390 476.355 ;
        RECT 6.290 472.160 91.260 472.285 ;
      LAYER Pwell ;
        RECT 6.290 468.640 1143.390 472.160 ;
      LAYER Nwell ;
        RECT 6.290 468.515 101.900 468.640 ;
        RECT 6.290 464.445 1143.390 468.515 ;
        RECT 6.290 464.320 160.545 464.445 ;
      LAYER Pwell ;
        RECT 6.290 460.800 1143.390 464.320 ;
      LAYER Nwell ;
        RECT 6.290 460.675 12.705 460.800 ;
        RECT 6.290 456.605 1143.390 460.675 ;
        RECT 6.290 456.480 236.705 456.605 ;
      LAYER Pwell ;
        RECT 6.290 452.960 1143.390 456.480 ;
      LAYER Nwell ;
        RECT 6.290 452.835 138.705 452.960 ;
        RECT 6.290 448.765 1143.390 452.835 ;
        RECT 6.290 448.640 161.665 448.765 ;
      LAYER Pwell ;
        RECT 6.290 445.120 1143.390 448.640 ;
      LAYER Nwell ;
        RECT 6.290 444.995 230.545 445.120 ;
        RECT 6.290 440.925 1143.390 444.995 ;
        RECT 6.290 440.800 83.865 440.925 ;
      LAYER Pwell ;
        RECT 6.290 437.280 1143.390 440.800 ;
      LAYER Nwell ;
        RECT 6.290 437.155 12.705 437.280 ;
        RECT 6.290 433.085 1143.390 437.155 ;
        RECT 6.290 432.960 83.405 433.085 ;
      LAYER Pwell ;
        RECT 6.290 429.440 1143.390 432.960 ;
      LAYER Nwell ;
        RECT 6.290 429.315 13.825 429.440 ;
        RECT 6.290 425.245 1143.390 429.315 ;
        RECT 6.290 425.120 559.825 425.245 ;
      LAYER Pwell ;
        RECT 6.290 421.600 1143.390 425.120 ;
      LAYER Nwell ;
        RECT 6.290 421.475 99.830 421.600 ;
        RECT 6.290 417.405 1143.390 421.475 ;
        RECT 6.290 417.280 12.705 417.405 ;
      LAYER Pwell ;
        RECT 6.290 413.760 1143.390 417.280 ;
      LAYER Nwell ;
        RECT 6.290 413.635 87.835 413.760 ;
        RECT 6.290 409.565 1143.390 413.635 ;
        RECT 6.290 409.440 146.610 409.565 ;
      LAYER Pwell ;
        RECT 6.290 405.920 1143.390 409.440 ;
      LAYER Nwell ;
        RECT 6.290 405.795 89.505 405.920 ;
        RECT 6.290 401.725 1143.390 405.795 ;
        RECT 6.290 401.600 193.025 401.725 ;
      LAYER Pwell ;
        RECT 6.290 398.080 1143.390 401.600 ;
      LAYER Nwell ;
        RECT 6.290 397.955 96.360 398.080 ;
        RECT 6.290 393.885 1143.390 397.955 ;
        RECT 6.290 393.760 59.400 393.885 ;
      LAYER Pwell ;
        RECT 6.290 390.240 1143.390 393.760 ;
      LAYER Nwell ;
        RECT 6.290 390.115 73.745 390.240 ;
        RECT 6.290 386.045 1143.390 390.115 ;
        RECT 6.290 385.920 120.785 386.045 ;
      LAYER Pwell ;
        RECT 6.290 382.400 1143.390 385.920 ;
      LAYER Nwell ;
        RECT 6.290 382.275 101.275 382.400 ;
        RECT 6.290 378.205 1143.390 382.275 ;
        RECT 6.290 378.080 91.150 378.205 ;
      LAYER Pwell ;
        RECT 6.290 374.560 1143.390 378.080 ;
      LAYER Nwell ;
        RECT 6.290 374.435 62.030 374.560 ;
        RECT 6.290 370.365 1143.390 374.435 ;
        RECT 6.290 370.240 46.385 370.365 ;
      LAYER Pwell ;
        RECT 6.290 366.720 1143.390 370.240 ;
      LAYER Nwell ;
        RECT 6.290 366.595 16.715 366.720 ;
        RECT 6.290 362.525 1143.390 366.595 ;
        RECT 6.290 362.400 20.875 362.525 ;
      LAYER Pwell ;
        RECT 6.290 358.880 1143.390 362.400 ;
      LAYER Nwell ;
        RECT 6.290 358.755 97.590 358.880 ;
        RECT 6.290 354.685 1143.390 358.755 ;
        RECT 6.290 354.560 30.670 354.685 ;
      LAYER Pwell ;
        RECT 6.290 351.040 1143.390 354.560 ;
      LAYER Nwell ;
        RECT 6.290 350.915 49.710 351.040 ;
        RECT 6.290 346.845 1143.390 350.915 ;
        RECT 6.290 346.720 45.810 346.845 ;
      LAYER Pwell ;
        RECT 6.290 343.200 1143.390 346.720 ;
      LAYER Nwell ;
        RECT 6.290 343.075 68.470 343.200 ;
        RECT 6.290 339.005 1143.390 343.075 ;
        RECT 6.290 338.880 36.270 339.005 ;
      LAYER Pwell ;
        RECT 6.290 335.360 1143.390 338.880 ;
      LAYER Nwell ;
        RECT 6.290 335.235 16.715 335.360 ;
        RECT 6.290 331.165 1143.390 335.235 ;
        RECT 6.290 331.040 48.590 331.165 ;
      LAYER Pwell ;
        RECT 6.290 327.520 1143.390 331.040 ;
      LAYER Nwell ;
        RECT 6.290 327.395 13.030 327.520 ;
        RECT 6.290 323.325 1143.390 327.395 ;
        RECT 6.290 323.200 49.710 323.325 ;
      LAYER Pwell ;
        RECT 6.290 319.680 1143.390 323.200 ;
      LAYER Nwell ;
        RECT 6.290 319.555 69.590 319.680 ;
        RECT 6.290 315.485 1143.390 319.555 ;
        RECT 6.290 315.360 35.150 315.485 ;
      LAYER Pwell ;
        RECT 6.290 311.840 1143.390 315.360 ;
      LAYER Nwell ;
        RECT 6.290 311.715 25.070 311.840 ;
        RECT 6.290 307.645 1143.390 311.715 ;
        RECT 6.290 307.520 272.085 307.645 ;
      LAYER Pwell ;
        RECT 6.290 304.000 1143.390 307.520 ;
      LAYER Nwell ;
        RECT 6.290 303.875 87.835 304.000 ;
        RECT 6.290 299.805 1143.390 303.875 ;
        RECT 6.290 299.680 9.440 299.805 ;
      LAYER Pwell ;
        RECT 6.290 296.160 1143.390 299.680 ;
      LAYER Nwell ;
        RECT 6.290 296.035 133.795 296.160 ;
        RECT 6.290 291.965 1143.390 296.035 ;
        RECT 6.290 291.840 16.950 291.965 ;
      LAYER Pwell ;
        RECT 6.290 288.320 1143.390 291.840 ;
      LAYER Nwell ;
        RECT 6.290 288.195 89.580 288.320 ;
        RECT 6.290 284.125 1143.390 288.195 ;
        RECT 6.290 284.000 13.310 284.125 ;
      LAYER Pwell ;
        RECT 6.290 280.480 1143.390 284.000 ;
      LAYER Nwell ;
        RECT 6.290 280.355 100.780 280.480 ;
        RECT 6.290 276.285 1143.390 280.355 ;
        RECT 6.290 276.160 21.210 276.285 ;
      LAYER Pwell ;
        RECT 6.290 272.640 1143.390 276.160 ;
      LAYER Nwell ;
        RECT 6.290 272.515 79.390 272.640 ;
        RECT 6.290 268.445 1143.390 272.515 ;
        RECT 6.290 268.320 68.190 268.445 ;
      LAYER Pwell ;
        RECT 6.290 264.800 1143.390 268.320 ;
      LAYER Nwell ;
        RECT 6.290 264.675 91.260 264.800 ;
        RECT 6.290 260.605 1143.390 264.675 ;
        RECT 6.290 260.480 91.430 260.605 ;
      LAYER Pwell ;
        RECT 6.290 256.960 1143.390 260.480 ;
      LAYER Nwell ;
        RECT 6.290 256.835 140.385 256.960 ;
        RECT 6.290 252.765 1143.390 256.835 ;
        RECT 6.290 252.640 13.590 252.765 ;
      LAYER Pwell ;
        RECT 6.290 249.120 1143.390 252.640 ;
      LAYER Nwell ;
        RECT 6.290 248.995 17.835 249.120 ;
        RECT 6.290 244.925 1143.390 248.995 ;
        RECT 6.290 244.800 124.885 244.925 ;
      LAYER Pwell ;
        RECT 6.290 241.280 1143.390 244.800 ;
      LAYER Nwell ;
        RECT 6.290 241.155 50.305 241.280 ;
        RECT 6.290 237.085 1143.390 241.155 ;
        RECT 6.290 236.960 403.800 237.085 ;
      LAYER Pwell ;
        RECT 6.290 233.440 1143.390 236.960 ;
      LAYER Nwell ;
        RECT 6.290 233.315 31.275 233.440 ;
        RECT 6.290 229.245 1143.390 233.315 ;
        RECT 6.290 229.120 19.080 229.245 ;
      LAYER Pwell ;
        RECT 6.290 225.600 1143.390 229.120 ;
      LAYER Nwell ;
        RECT 6.290 225.475 33.425 225.600 ;
        RECT 6.290 221.405 1143.390 225.475 ;
        RECT 6.290 221.280 77.105 221.405 ;
      LAYER Pwell ;
        RECT 6.290 217.760 1143.390 221.280 ;
      LAYER Nwell ;
        RECT 6.290 217.635 17.960 217.760 ;
        RECT 6.290 213.565 1143.390 217.635 ;
        RECT 6.290 213.440 71.650 213.565 ;
      LAYER Pwell ;
        RECT 6.290 209.920 1143.390 213.440 ;
      LAYER Nwell ;
        RECT 6.290 209.795 53.735 209.920 ;
        RECT 6.290 205.725 1143.390 209.795 ;
        RECT 6.290 205.600 14.945 205.725 ;
      LAYER Pwell ;
        RECT 6.290 202.080 1143.390 205.600 ;
      LAYER Nwell ;
        RECT 6.290 201.955 23.345 202.080 ;
        RECT 6.290 197.885 1143.390 201.955 ;
        RECT 6.290 197.760 110.705 197.885 ;
      LAYER Pwell ;
        RECT 6.290 194.240 1143.390 197.760 ;
      LAYER Nwell ;
        RECT 6.290 194.115 12.705 194.240 ;
        RECT 6.290 190.045 1143.390 194.115 ;
        RECT 6.290 189.920 43.505 190.045 ;
      LAYER Pwell ;
        RECT 6.290 186.400 1143.390 189.920 ;
      LAYER Nwell ;
        RECT 6.290 186.275 12.705 186.400 ;
        RECT 6.290 182.205 1143.390 186.275 ;
        RECT 6.290 182.080 32.305 182.205 ;
      LAYER Pwell ;
        RECT 6.290 178.560 1143.390 182.080 ;
      LAYER Nwell ;
        RECT 6.290 178.435 34.545 178.560 ;
        RECT 6.290 174.365 1143.390 178.435 ;
        RECT 6.290 174.240 12.705 174.365 ;
      LAYER Pwell ;
        RECT 6.290 170.720 1143.390 174.240 ;
      LAYER Nwell ;
        RECT 6.290 170.595 65.560 170.720 ;
        RECT 6.290 166.525 1143.390 170.595 ;
        RECT 6.290 166.400 39.585 166.525 ;
      LAYER Pwell ;
        RECT 6.290 162.880 1143.390 166.400 ;
      LAYER Nwell ;
        RECT 6.290 162.755 12.705 162.880 ;
        RECT 6.290 158.685 1143.390 162.755 ;
        RECT 6.290 158.560 53.205 158.685 ;
      LAYER Pwell ;
        RECT 6.290 155.040 1143.390 158.560 ;
      LAYER Nwell ;
        RECT 6.290 154.915 33.425 155.040 ;
        RECT 6.290 150.845 1143.390 154.915 ;
        RECT 6.290 150.720 13.265 150.845 ;
      LAYER Pwell ;
        RECT 6.290 147.200 1143.390 150.720 ;
      LAYER Nwell ;
        RECT 6.290 147.075 61.985 147.200 ;
        RECT 6.290 143.005 1143.390 147.075 ;
        RECT 6.290 142.880 14.385 143.005 ;
      LAYER Pwell ;
        RECT 6.290 139.360 1143.390 142.880 ;
      LAYER Nwell ;
        RECT 6.290 139.235 56.580 139.360 ;
        RECT 6.290 135.165 1143.390 139.235 ;
        RECT 6.290 135.040 45.745 135.165 ;
      LAYER Pwell ;
        RECT 6.290 131.520 1143.390 135.040 ;
      LAYER Nwell ;
        RECT 6.290 131.395 28.385 131.520 ;
        RECT 6.290 127.325 1143.390 131.395 ;
        RECT 6.290 127.200 13.825 127.325 ;
      LAYER Pwell ;
        RECT 6.290 123.680 1143.390 127.200 ;
      LAYER Nwell ;
        RECT 6.290 123.555 34.695 123.680 ;
        RECT 6.290 119.485 1143.390 123.555 ;
        RECT 6.290 119.360 13.265 119.485 ;
      LAYER Pwell ;
        RECT 6.290 115.840 1143.390 119.360 ;
      LAYER Nwell ;
        RECT 6.290 115.715 32.865 115.840 ;
        RECT 6.290 111.645 1143.390 115.715 ;
        RECT 6.290 111.520 14.385 111.645 ;
      LAYER Pwell ;
        RECT 6.290 108.000 1143.390 111.520 ;
      LAYER Nwell ;
        RECT 6.290 107.875 110.705 108.000 ;
        RECT 6.290 103.805 1143.390 107.875 ;
        RECT 6.290 103.680 71.505 103.805 ;
      LAYER Pwell ;
        RECT 6.290 100.160 1143.390 103.680 ;
      LAYER Nwell ;
        RECT 6.290 100.035 13.265 100.160 ;
        RECT 6.290 95.965 1143.390 100.035 ;
        RECT 6.290 95.840 54.235 95.965 ;
      LAYER Pwell ;
        RECT 6.290 92.320 1143.390 95.840 ;
      LAYER Nwell ;
        RECT 6.290 92.195 73.745 92.320 ;
        RECT 6.290 88.125 1143.390 92.195 ;
        RECT 6.290 88.000 12.705 88.125 ;
      LAYER Pwell ;
        RECT 6.290 84.480 1143.390 88.000 ;
      LAYER Nwell ;
        RECT 6.290 84.355 26.145 84.480 ;
        RECT 6.290 80.285 1143.390 84.355 ;
        RECT 6.290 80.160 50.885 80.285 ;
      LAYER Pwell ;
        RECT 6.290 76.640 1143.390 80.160 ;
      LAYER Nwell ;
        RECT 6.290 76.515 26.705 76.640 ;
        RECT 6.290 72.445 1143.390 76.515 ;
        RECT 6.290 72.320 12.705 72.445 ;
      LAYER Pwell ;
        RECT 6.290 68.800 1143.390 72.320 ;
      LAYER Nwell ;
        RECT 6.290 68.675 178.565 68.800 ;
        RECT 6.290 64.605 1143.390 68.675 ;
        RECT 6.290 64.480 83.825 64.605 ;
      LAYER Pwell ;
        RECT 6.290 60.960 1143.390 64.480 ;
      LAYER Nwell ;
        RECT 6.290 60.835 20.545 60.960 ;
        RECT 6.290 56.765 1143.390 60.835 ;
        RECT 6.290 56.640 12.705 56.765 ;
      LAYER Pwell ;
        RECT 6.290 53.120 1143.390 56.640 ;
      LAYER Nwell ;
        RECT 6.290 52.995 18.305 53.120 ;
        RECT 6.290 48.925 1143.390 52.995 ;
        RECT 6.290 48.800 89.525 48.925 ;
      LAYER Pwell ;
        RECT 6.290 45.280 1143.390 48.800 ;
      LAYER Nwell ;
        RECT 6.290 45.155 30.065 45.280 ;
        RECT 6.290 41.085 1143.390 45.155 ;
        RECT 6.290 40.960 81.125 41.085 ;
      LAYER Pwell ;
        RECT 6.290 37.440 1143.390 40.960 ;
      LAYER Nwell ;
        RECT 6.290 37.315 134.225 37.440 ;
        RECT 6.290 33.245 1143.390 37.315 ;
        RECT 6.290 33.120 37.905 33.245 ;
      LAYER Pwell ;
        RECT 6.290 29.600 1143.390 33.120 ;
      LAYER Nwell ;
        RECT 6.290 29.475 68.145 29.600 ;
        RECT 6.290 25.405 1143.390 29.475 ;
        RECT 6.290 25.280 78.785 25.405 ;
      LAYER Pwell ;
        RECT 6.290 21.760 1143.390 25.280 ;
      LAYER Nwell ;
        RECT 6.290 21.635 58.625 21.760 ;
        RECT 6.290 17.565 1143.390 21.635 ;
        RECT 6.290 17.440 299.985 17.565 ;
      LAYER Pwell ;
        RECT 6.290 15.250 1143.390 17.440 ;
      LAYER Metal1 ;
        RECT 6.720 15.380 1142.960 734.010 ;
      LAYER Metal2 ;
        RECT 8.540 745.700 574.260 746.000 ;
        RECT 575.420 745.700 1142.260 746.000 ;
        RECT 8.540 4.300 1142.260 745.700 ;
        RECT 8.540 4.000 286.420 4.300 ;
        RECT 287.580 4.000 860.980 4.300 ;
        RECT 862.140 4.000 1142.260 4.300 ;
      LAYER Metal3 ;
        RECT 8.490 731.100 1146.000 744.100 ;
        RECT 8.490 729.940 1145.700 731.100 ;
        RECT 8.490 717.660 1146.000 729.940 ;
        RECT 8.490 716.500 1145.700 717.660 ;
        RECT 8.490 704.220 1146.000 716.500 ;
        RECT 8.490 703.060 1145.700 704.220 ;
        RECT 8.490 690.780 1146.000 703.060 ;
        RECT 8.490 689.620 1145.700 690.780 ;
        RECT 8.490 677.340 1146.000 689.620 ;
        RECT 8.490 676.180 1145.700 677.340 ;
        RECT 8.490 663.900 1146.000 676.180 ;
        RECT 8.490 662.740 1145.700 663.900 ;
        RECT 8.490 650.460 1146.000 662.740 ;
        RECT 8.490 649.300 1145.700 650.460 ;
        RECT 8.490 637.020 1146.000 649.300 ;
        RECT 8.490 635.860 1145.700 637.020 ;
        RECT 8.490 623.580 1146.000 635.860 ;
        RECT 8.490 622.420 1145.700 623.580 ;
        RECT 8.490 610.140 1146.000 622.420 ;
        RECT 8.490 608.980 1145.700 610.140 ;
        RECT 8.490 596.700 1146.000 608.980 ;
        RECT 8.490 595.540 1145.700 596.700 ;
        RECT 8.490 583.260 1146.000 595.540 ;
        RECT 8.490 582.100 1145.700 583.260 ;
        RECT 8.490 569.820 1146.000 582.100 ;
        RECT 8.490 568.660 1145.700 569.820 ;
        RECT 8.490 556.380 1146.000 568.660 ;
        RECT 8.490 555.220 1145.700 556.380 ;
        RECT 8.490 542.940 1146.000 555.220 ;
        RECT 8.490 541.780 1145.700 542.940 ;
        RECT 8.490 529.500 1146.000 541.780 ;
        RECT 8.490 528.340 1145.700 529.500 ;
        RECT 8.490 516.060 1146.000 528.340 ;
        RECT 8.490 514.900 1145.700 516.060 ;
        RECT 8.490 502.620 1146.000 514.900 ;
        RECT 8.490 501.460 1145.700 502.620 ;
        RECT 8.490 489.180 1146.000 501.460 ;
        RECT 8.490 488.020 1145.700 489.180 ;
        RECT 8.490 475.740 1146.000 488.020 ;
        RECT 8.490 474.580 1145.700 475.740 ;
        RECT 8.490 462.300 1146.000 474.580 ;
        RECT 8.490 461.140 1145.700 462.300 ;
        RECT 8.490 448.860 1146.000 461.140 ;
        RECT 8.490 447.700 1145.700 448.860 ;
        RECT 8.490 435.420 1146.000 447.700 ;
        RECT 8.490 434.260 1145.700 435.420 ;
        RECT 8.490 421.980 1146.000 434.260 ;
        RECT 8.490 420.820 1145.700 421.980 ;
        RECT 8.490 408.540 1146.000 420.820 ;
        RECT 8.490 407.380 1145.700 408.540 ;
        RECT 8.490 395.100 1146.000 407.380 ;
        RECT 8.490 393.940 1145.700 395.100 ;
        RECT 8.490 381.660 1146.000 393.940 ;
        RECT 8.490 380.500 1145.700 381.660 ;
        RECT 8.490 368.220 1146.000 380.500 ;
        RECT 8.490 367.060 1145.700 368.220 ;
        RECT 8.490 354.780 1146.000 367.060 ;
        RECT 8.490 353.620 1145.700 354.780 ;
        RECT 8.490 341.340 1146.000 353.620 ;
        RECT 8.490 340.180 1145.700 341.340 ;
        RECT 8.490 327.900 1146.000 340.180 ;
        RECT 8.490 326.740 1145.700 327.900 ;
        RECT 8.490 314.460 1146.000 326.740 ;
        RECT 8.490 313.300 1145.700 314.460 ;
        RECT 8.490 301.020 1146.000 313.300 ;
        RECT 8.490 299.860 1145.700 301.020 ;
        RECT 8.490 287.580 1146.000 299.860 ;
        RECT 8.490 286.420 1145.700 287.580 ;
        RECT 8.490 274.140 1146.000 286.420 ;
        RECT 8.490 272.980 1145.700 274.140 ;
        RECT 8.490 260.700 1146.000 272.980 ;
        RECT 8.490 259.540 1145.700 260.700 ;
        RECT 8.490 247.260 1146.000 259.540 ;
        RECT 8.490 246.100 1145.700 247.260 ;
        RECT 8.490 233.820 1146.000 246.100 ;
        RECT 8.490 232.660 1145.700 233.820 ;
        RECT 8.490 220.380 1146.000 232.660 ;
        RECT 8.490 219.220 1145.700 220.380 ;
        RECT 8.490 206.940 1146.000 219.220 ;
        RECT 8.490 205.780 1145.700 206.940 ;
        RECT 8.490 193.500 1146.000 205.780 ;
        RECT 8.490 192.340 1145.700 193.500 ;
        RECT 8.490 180.060 1146.000 192.340 ;
        RECT 8.490 178.900 1145.700 180.060 ;
        RECT 8.490 166.620 1146.000 178.900 ;
        RECT 8.490 165.460 1145.700 166.620 ;
        RECT 8.490 153.180 1146.000 165.460 ;
        RECT 8.490 152.020 1145.700 153.180 ;
        RECT 8.490 139.740 1146.000 152.020 ;
        RECT 8.490 138.580 1145.700 139.740 ;
        RECT 8.490 126.300 1146.000 138.580 ;
        RECT 8.490 125.140 1145.700 126.300 ;
        RECT 8.490 112.860 1146.000 125.140 ;
        RECT 8.490 111.700 1145.700 112.860 ;
        RECT 8.490 99.420 1146.000 111.700 ;
        RECT 8.490 98.260 1145.700 99.420 ;
        RECT 8.490 85.980 1146.000 98.260 ;
        RECT 8.490 84.820 1145.700 85.980 ;
        RECT 8.490 72.540 1146.000 84.820 ;
        RECT 8.490 71.380 1145.700 72.540 ;
        RECT 8.490 59.100 1146.000 71.380 ;
        RECT 8.490 57.940 1145.700 59.100 ;
        RECT 8.490 45.660 1146.000 57.940 ;
        RECT 8.490 44.500 1145.700 45.660 ;
        RECT 8.490 32.220 1146.000 44.500 ;
        RECT 8.490 31.060 1145.700 32.220 ;
        RECT 8.490 18.780 1146.000 31.060 ;
        RECT 8.490 17.620 1145.700 18.780 ;
        RECT 8.490 3.500 1146.000 17.620 ;
      LAYER Metal4 ;
        RECT 39.340 733.640 1130.500 744.150 ;
        RECT 39.340 15.080 98.740 733.640 ;
        RECT 100.940 15.080 175.540 733.640 ;
        RECT 177.740 15.080 252.340 733.640 ;
        RECT 254.540 15.080 329.140 733.640 ;
        RECT 331.340 15.080 405.940 733.640 ;
        RECT 408.140 15.080 482.740 733.640 ;
        RECT 484.940 15.080 559.540 733.640 ;
        RECT 561.740 15.080 636.340 733.640 ;
        RECT 638.540 15.080 713.140 733.640 ;
        RECT 715.340 15.080 789.940 733.640 ;
        RECT 792.140 15.080 866.740 733.640 ;
        RECT 868.940 15.080 943.540 733.640 ;
        RECT 945.740 15.080 1020.340 733.640 ;
        RECT 1022.540 15.080 1097.140 733.640 ;
        RECT 1099.340 15.080 1130.500 733.640 ;
        RECT 39.340 3.450 1130.500 15.080 ;
  END
END wrapped_sid
END LIBRARY

