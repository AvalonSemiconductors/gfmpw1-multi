* NGSPICE file created from blinker.ext - technology: gf180mcuD

.subckt blinker io_out[0] io_out[1] io_out[2] rst_n vdd vss wb_clk_i
.ends

