VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_mc14500
  CLASS BLOCK ;
  FOREIGN wrapped_mc14500 ;
  ORIGIN 0.000 0.000 ;
  SIZE 175.000 BY 175.000 ;
  PIN SDI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 171.000 140.000 175.000 140.560 ;
    END
  END SDI
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 171.000 5.600 175.000 6.160 ;
    END
  END clk_i
  PIN custom_setting
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 171.000 166.880 175.000 167.440 ;
    END
  END custom_setting
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 171.000 32.480 175.000 33.040 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 171.000 45.920 175.000 46.480 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 171.000 59.360 175.000 59.920 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 171.000 72.800 175.000 73.360 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 171.000 86.240 175.000 86.800 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 171.000 99.680 175.000 100.240 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 171.000 113.120 175.000 113.680 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 171.000 126.560 175.000 127.120 ;
    END
  END io_in[7]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2.240 171.000 2.800 175.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 58.240 171.000 58.800 175.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 171.000 64.400 175.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 69.440 171.000 70.000 175.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 75.040 171.000 75.600 175.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 171.000 81.200 175.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 86.240 171.000 86.800 175.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 91.840 171.000 92.400 175.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 171.000 98.000 175.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 103.040 171.000 103.600 175.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 108.640 171.000 109.200 175.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 7.840 171.000 8.400 175.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 171.000 114.800 175.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 119.840 171.000 120.400 175.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 125.440 171.000 126.000 175.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 171.000 131.600 175.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 136.640 171.000 137.200 175.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 142.240 171.000 142.800 175.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 171.000 148.400 175.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 153.440 171.000 154.000 175.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 159.040 171.000 159.600 175.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 171.000 165.200 175.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 171.000 14.000 175.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 170.240 171.000 170.800 175.000 ;
    END
  END io_out[30]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 19.040 171.000 19.600 175.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 24.640 171.000 25.200 175.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 171.000 30.800 175.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 35.840 171.000 36.400 175.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 41.440 171.000 42.000 175.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 171.000 47.600 175.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 52.640 171.000 53.200 175.000 ;
    END
  END io_out[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 171.000 19.040 175.000 19.600 ;
    END
  END rst_n
  PIN sram_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 4.480 0.000 5.040 4.000 ;
    END
  END sram_addr[0]
  PIN sram_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 12.320 0.000 12.880 4.000 ;
    END
  END sram_addr[1]
  PIN sram_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 20.160 0.000 20.720 4.000 ;
    END
  END sram_addr[2]
  PIN sram_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 28.000 0.000 28.560 4.000 ;
    END
  END sram_addr[3]
  PIN sram_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 35.840 0.000 36.400 4.000 ;
    END
  END sram_addr[4]
  PIN sram_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 0.000 44.240 4.000 ;
    END
  END sram_addr[5]
  PIN sram_gwe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 171.000 153.440 175.000 154.000 ;
    END
  END sram_gwe
  PIN sram_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 51.520 0.000 52.080 4.000 ;
    END
  END sram_in[0]
  PIN sram_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 59.360 0.000 59.920 4.000 ;
    END
  END sram_in[1]
  PIN sram_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 0.000 67.760 4.000 ;
    END
  END sram_in[2]
  PIN sram_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 75.040 0.000 75.600 4.000 ;
    END
  END sram_in[3]
  PIN sram_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 82.880 0.000 83.440 4.000 ;
    END
  END sram_in[4]
  PIN sram_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 0.000 91.280 4.000 ;
    END
  END sram_in[5]
  PIN sram_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 98.560 0.000 99.120 4.000 ;
    END
  END sram_in[6]
  PIN sram_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 106.400 0.000 106.960 4.000 ;
    END
  END sram_in[7]
  PIN sram_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 0.000 114.800 4.000 ;
    END
  END sram_out[0]
  PIN sram_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 122.080 0.000 122.640 4.000 ;
    END
  END sram_out[1]
  PIN sram_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 129.920 0.000 130.480 4.000 ;
    END
  END sram_out[2]
  PIN sram_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 0.000 138.320 4.000 ;
    END
  END sram_out[3]
  PIN sram_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 145.600 0.000 146.160 4.000 ;
    END
  END sram_out[4]
  PIN sram_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 153.440 0.000 154.000 4.000 ;
    END
  END sram_out[5]
  PIN sram_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 0.000 161.840 4.000 ;
    END
  END sram_out[6]
  PIN sram_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 169.120 0.000 169.680 4.000 ;
    END
  END sram_out[7]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 26.080 15.380 27.680 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 66.400 15.380 68.000 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 106.720 15.380 108.320 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 147.040 15.380 148.640 157.100 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 46.240 15.380 47.840 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 86.560 15.380 88.160 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 126.880 15.380 128.480 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 167.200 15.380 168.800 157.100 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 2.330 15.380 168.800 157.770 ;
      LAYER Metal2 ;
        RECT 3.100 170.700 7.540 171.780 ;
        RECT 8.700 170.700 13.140 171.780 ;
        RECT 14.300 170.700 18.740 171.780 ;
        RECT 19.900 170.700 24.340 171.780 ;
        RECT 25.500 170.700 29.940 171.780 ;
        RECT 31.100 170.700 35.540 171.780 ;
        RECT 36.700 170.700 41.140 171.780 ;
        RECT 42.300 170.700 46.740 171.780 ;
        RECT 47.900 170.700 52.340 171.780 ;
        RECT 53.500 170.700 57.940 171.780 ;
        RECT 59.100 170.700 63.540 171.780 ;
        RECT 64.700 170.700 69.140 171.780 ;
        RECT 70.300 170.700 74.740 171.780 ;
        RECT 75.900 170.700 80.340 171.780 ;
        RECT 81.500 170.700 85.940 171.780 ;
        RECT 87.100 170.700 91.540 171.780 ;
        RECT 92.700 170.700 97.140 171.780 ;
        RECT 98.300 170.700 102.740 171.780 ;
        RECT 103.900 170.700 108.340 171.780 ;
        RECT 109.500 170.700 113.940 171.780 ;
        RECT 115.100 170.700 119.540 171.780 ;
        RECT 120.700 170.700 125.140 171.780 ;
        RECT 126.300 170.700 130.740 171.780 ;
        RECT 131.900 170.700 136.340 171.780 ;
        RECT 137.500 170.700 141.940 171.780 ;
        RECT 143.100 170.700 147.540 171.780 ;
        RECT 148.700 170.700 153.140 171.780 ;
        RECT 154.300 170.700 158.740 171.780 ;
        RECT 159.900 170.700 164.340 171.780 ;
        RECT 165.500 170.700 169.940 171.780 ;
        RECT 2.380 4.300 170.660 170.700 ;
        RECT 2.380 3.500 4.180 4.300 ;
        RECT 5.340 3.500 12.020 4.300 ;
        RECT 13.180 3.500 19.860 4.300 ;
        RECT 21.020 3.500 27.700 4.300 ;
        RECT 28.860 3.500 35.540 4.300 ;
        RECT 36.700 3.500 43.380 4.300 ;
        RECT 44.540 3.500 51.220 4.300 ;
        RECT 52.380 3.500 59.060 4.300 ;
        RECT 60.220 3.500 66.900 4.300 ;
        RECT 68.060 3.500 74.740 4.300 ;
        RECT 75.900 3.500 82.580 4.300 ;
        RECT 83.740 3.500 90.420 4.300 ;
        RECT 91.580 3.500 98.260 4.300 ;
        RECT 99.420 3.500 106.100 4.300 ;
        RECT 107.260 3.500 113.940 4.300 ;
        RECT 115.100 3.500 121.780 4.300 ;
        RECT 122.940 3.500 129.620 4.300 ;
        RECT 130.780 3.500 137.460 4.300 ;
        RECT 138.620 3.500 145.300 4.300 ;
        RECT 146.460 3.500 153.140 4.300 ;
        RECT 154.300 3.500 160.980 4.300 ;
        RECT 162.140 3.500 168.820 4.300 ;
        RECT 169.980 3.500 170.660 4.300 ;
      LAYER Metal3 ;
        RECT 4.570 166.580 170.700 167.300 ;
        RECT 4.570 154.300 171.000 166.580 ;
        RECT 4.570 153.140 170.700 154.300 ;
        RECT 4.570 140.860 171.000 153.140 ;
        RECT 4.570 139.700 170.700 140.860 ;
        RECT 4.570 127.420 171.000 139.700 ;
        RECT 4.570 126.260 170.700 127.420 ;
        RECT 4.570 113.980 171.000 126.260 ;
        RECT 4.570 112.820 170.700 113.980 ;
        RECT 4.570 100.540 171.000 112.820 ;
        RECT 4.570 99.380 170.700 100.540 ;
        RECT 4.570 87.100 171.000 99.380 ;
        RECT 4.570 85.940 170.700 87.100 ;
        RECT 4.570 73.660 171.000 85.940 ;
        RECT 4.570 72.500 170.700 73.660 ;
        RECT 4.570 60.220 171.000 72.500 ;
        RECT 4.570 59.060 170.700 60.220 ;
        RECT 4.570 46.780 171.000 59.060 ;
        RECT 4.570 45.620 170.700 46.780 ;
        RECT 4.570 33.340 171.000 45.620 ;
        RECT 4.570 32.180 170.700 33.340 ;
        RECT 4.570 19.900 171.000 32.180 ;
        RECT 4.570 18.740 170.700 19.900 ;
        RECT 4.570 6.460 171.000 18.740 ;
        RECT 4.570 5.740 170.700 6.460 ;
      LAYER Metal4 ;
        RECT 25.340 157.400 154.980 165.670 ;
        RECT 25.340 16.330 25.780 157.400 ;
        RECT 27.980 16.330 45.940 157.400 ;
        RECT 48.140 16.330 66.100 157.400 ;
        RECT 68.300 16.330 86.260 157.400 ;
        RECT 88.460 16.330 106.420 157.400 ;
        RECT 108.620 16.330 126.580 157.400 ;
        RECT 128.780 16.330 146.740 157.400 ;
        RECT 148.940 16.330 154.980 157.400 ;
  END
END wrapped_mc14500
END LIBRARY

