magic
tech gf180mcuD
magscale 1 5
timestamp 1753968502
<< nwell >>
rect 629 1525 24347 23171
<< obsm1 >>
rect 672 1538 24304 23158
<< metal2 >>
rect 1792 24600 1848 25000
rect 2576 24600 2632 25000
rect 3360 24600 3416 25000
rect 4144 24600 4200 25000
rect 4928 24600 4984 25000
rect 5712 24600 5768 25000
rect 6496 24600 6552 25000
rect 7280 24600 7336 25000
rect 8064 24600 8120 25000
rect 8848 24600 8904 25000
rect 9632 24600 9688 25000
rect 10416 24600 10472 25000
rect 11200 24600 11256 25000
rect 11984 24600 12040 25000
rect 12768 24600 12824 25000
rect 13552 24600 13608 25000
rect 14336 24600 14392 25000
rect 15120 24600 15176 25000
rect 15904 24600 15960 25000
rect 16688 24600 16744 25000
rect 17472 24600 17528 25000
rect 18256 24600 18312 25000
rect 19040 24600 19096 25000
rect 19824 24600 19880 25000
rect 20608 24600 20664 25000
rect 21392 24600 21448 25000
rect 22176 24600 22232 25000
rect 22960 24600 23016 25000
<< obsm2 >>
rect 14 24570 1762 24682
rect 1878 24570 2546 24682
rect 2662 24570 3330 24682
rect 3446 24570 4114 24682
rect 4230 24570 4898 24682
rect 5014 24570 5682 24682
rect 5798 24570 6466 24682
rect 6582 24570 7250 24682
rect 7366 24570 8034 24682
rect 8150 24570 8818 24682
rect 8934 24570 9602 24682
rect 9718 24570 10386 24682
rect 10502 24570 11170 24682
rect 11286 24570 11954 24682
rect 12070 24570 12738 24682
rect 12854 24570 13522 24682
rect 13638 24570 14306 24682
rect 14422 24570 15090 24682
rect 15206 24570 15874 24682
rect 15990 24570 16658 24682
rect 16774 24570 17442 24682
rect 17558 24570 18226 24682
rect 18342 24570 19010 24682
rect 19126 24570 19794 24682
rect 19910 24570 20578 24682
rect 20694 24570 21362 24682
rect 21478 24570 22146 24682
rect 22262 24570 22930 24682
rect 23046 24570 24402 24682
rect 14 1353 24402 24570
<< metal3 >>
rect 24600 23520 25000 23576
rect 24600 21056 25000 21112
rect 0 20720 400 20776
rect 24600 18592 25000 18648
rect 24600 16128 25000 16184
rect 24600 13664 25000 13720
rect 0 12432 400 12488
rect 24600 11200 25000 11256
rect 24600 8736 25000 8792
rect 24600 6272 25000 6328
rect 0 4144 400 4200
rect 24600 3808 25000 3864
rect 24600 1344 25000 1400
<< obsm3 >>
rect 9 23490 24570 23562
rect 9 21142 24682 23490
rect 9 21026 24570 21142
rect 9 20806 24682 21026
rect 430 20690 24682 20806
rect 9 18678 24682 20690
rect 9 18562 24570 18678
rect 9 16214 24682 18562
rect 9 16098 24570 16214
rect 9 13750 24682 16098
rect 9 13634 24570 13750
rect 9 12518 24682 13634
rect 430 12402 24682 12518
rect 9 11286 24682 12402
rect 9 11170 24570 11286
rect 9 8822 24682 11170
rect 9 8706 24570 8822
rect 9 6358 24682 8706
rect 9 6242 24570 6358
rect 9 4230 24682 6242
rect 430 4114 24682 4230
rect 9 3894 24682 4114
rect 9 3778 24570 3894
rect 9 1430 24682 3778
rect 9 1358 24570 1430
<< metal4 >>
rect 2224 1538 2384 23158
rect 9904 1538 10064 23158
rect 17584 1538 17744 23158
<< obsm4 >>
rect 3206 1633 9874 22783
rect 10094 1633 17554 22783
rect 17774 1633 23450 22783
<< labels >>
rlabel metal3 s 24600 21056 25000 21112 6 custom_settings[0]
port 1 nsew signal input
rlabel metal3 s 24600 23520 25000 23576 6 custom_settings[1]
port 2 nsew signal input
rlabel metal3 s 24600 1344 25000 1400 6 io_in_1[0]
port 3 nsew signal input
rlabel metal3 s 24600 3808 25000 3864 6 io_in_1[1]
port 4 nsew signal input
rlabel metal3 s 24600 6272 25000 6328 6 io_in_1[2]
port 5 nsew signal input
rlabel metal3 s 24600 8736 25000 8792 6 io_in_1[3]
port 6 nsew signal input
rlabel metal3 s 24600 11200 25000 11256 6 io_in_1[4]
port 7 nsew signal input
rlabel metal3 s 24600 13664 25000 13720 6 io_in_1[5]
port 8 nsew signal input
rlabel metal3 s 24600 16128 25000 16184 6 io_in_1[6]
port 9 nsew signal input
rlabel metal3 s 24600 18592 25000 18648 6 io_in_1[7]
port 10 nsew signal input
rlabel metal3 s 0 20720 400 20776 6 io_in_2
port 11 nsew signal input
rlabel metal2 s 1792 24600 1848 25000 6 io_out[0]
port 12 nsew signal output
rlabel metal2 s 9632 24600 9688 25000 6 io_out[10]
port 13 nsew signal output
rlabel metal2 s 10416 24600 10472 25000 6 io_out[11]
port 14 nsew signal output
rlabel metal2 s 11200 24600 11256 25000 6 io_out[12]
port 15 nsew signal output
rlabel metal2 s 11984 24600 12040 25000 6 io_out[13]
port 16 nsew signal output
rlabel metal2 s 12768 24600 12824 25000 6 io_out[14]
port 17 nsew signal output
rlabel metal2 s 13552 24600 13608 25000 6 io_out[15]
port 18 nsew signal output
rlabel metal2 s 14336 24600 14392 25000 6 io_out[16]
port 19 nsew signal output
rlabel metal2 s 15120 24600 15176 25000 6 io_out[17]
port 20 nsew signal output
rlabel metal2 s 15904 24600 15960 25000 6 io_out[18]
port 21 nsew signal output
rlabel metal2 s 16688 24600 16744 25000 6 io_out[19]
port 22 nsew signal output
rlabel metal2 s 2576 24600 2632 25000 6 io_out[1]
port 23 nsew signal output
rlabel metal2 s 17472 24600 17528 25000 6 io_out[20]
port 24 nsew signal output
rlabel metal2 s 18256 24600 18312 25000 6 io_out[21]
port 25 nsew signal output
rlabel metal2 s 19040 24600 19096 25000 6 io_out[22]
port 26 nsew signal output
rlabel metal2 s 19824 24600 19880 25000 6 io_out[23]
port 27 nsew signal output
rlabel metal2 s 20608 24600 20664 25000 6 io_out[24]
port 28 nsew signal output
rlabel metal2 s 21392 24600 21448 25000 6 io_out[25]
port 29 nsew signal output
rlabel metal2 s 22176 24600 22232 25000 6 io_out[26]
port 30 nsew signal output
rlabel metal2 s 22960 24600 23016 25000 6 io_out[27]
port 31 nsew signal output
rlabel metal2 s 3360 24600 3416 25000 6 io_out[2]
port 32 nsew signal output
rlabel metal2 s 4144 24600 4200 25000 6 io_out[3]
port 33 nsew signal output
rlabel metal2 s 4928 24600 4984 25000 6 io_out[4]
port 34 nsew signal output
rlabel metal2 s 5712 24600 5768 25000 6 io_out[5]
port 35 nsew signal output
rlabel metal2 s 6496 24600 6552 25000 6 io_out[6]
port 36 nsew signal output
rlabel metal2 s 7280 24600 7336 25000 6 io_out[7]
port 37 nsew signal output
rlabel metal2 s 8064 24600 8120 25000 6 io_out[8]
port 38 nsew signal output
rlabel metal2 s 8848 24600 8904 25000 6 io_out[9]
port 39 nsew signal output
rlabel metal3 s 0 12432 400 12488 6 rst_n
port 40 nsew signal input
rlabel metal4 s 2224 1538 2384 23158 6 vdd
port 41 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 23158 6 vdd
port 41 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 23158 6 vss
port 42 nsew ground bidirectional
rlabel metal3 s 0 4144 400 4200 6 wb_clk_i
port 43 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 25000 25000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2706390
string GDS_FILE /home/lucah/gfmpw1-multi/openlane/wrapped_sn76489/runs/25_07_31_15_25/results/signoff/wrapped_sn76489.magic.gds
string GDS_START 228656
<< end >>

