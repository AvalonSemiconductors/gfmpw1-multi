magic
tech gf180mcuD
magscale 1 5
timestamp 1702459010
<< metal1 >>
rect 672 10205 11392 10222
rect 672 10179 3267 10205
rect 3293 10179 3319 10205
rect 3345 10179 3371 10205
rect 3397 10179 5927 10205
rect 5953 10179 5979 10205
rect 6005 10179 6031 10205
rect 6057 10179 8587 10205
rect 8613 10179 8639 10205
rect 8665 10179 8691 10205
rect 8717 10179 11247 10205
rect 11273 10179 11299 10205
rect 11325 10179 11351 10205
rect 11377 10179 11392 10205
rect 672 10162 11392 10179
rect 1017 10039 1023 10065
rect 1049 10039 1055 10065
rect 2137 10039 2143 10065
rect 2169 10039 2175 10065
rect 3257 10039 3263 10065
rect 3289 10039 3295 10065
rect 4657 10039 4663 10065
rect 4689 10039 4695 10065
rect 5497 10039 5503 10065
rect 5529 10039 5535 10065
rect 6617 10039 6623 10065
rect 6649 10039 6655 10065
rect 7737 10039 7743 10065
rect 7769 10039 7775 10065
rect 8857 10039 8863 10065
rect 8889 10039 8895 10065
rect 10089 10039 10095 10065
rect 10121 10039 10127 10065
rect 10369 10039 10375 10065
rect 10401 10039 10407 10065
rect 11097 10039 11103 10065
rect 11129 10039 11135 10065
rect 2311 10009 2337 10015
rect 1129 9983 1135 10009
rect 1161 9983 1167 10009
rect 2311 9977 2337 9983
rect 3431 10009 3457 10015
rect 6791 10009 6817 10015
rect 9927 10009 9953 10015
rect 10935 10009 10961 10015
rect 4769 9983 4775 10009
rect 4801 9983 4807 10009
rect 5609 9983 5615 10009
rect 5641 9983 5647 10009
rect 7849 9983 7855 10009
rect 7881 9983 7887 10009
rect 8969 9983 8975 10009
rect 9001 9983 9007 10009
rect 10481 9983 10487 10009
rect 10513 9983 10519 10009
rect 3431 9977 3457 9983
rect 6791 9977 6817 9983
rect 9927 9977 9953 9983
rect 10935 9977 10961 9983
rect 672 9813 11312 9830
rect 672 9787 1937 9813
rect 1963 9787 1989 9813
rect 2015 9787 2041 9813
rect 2067 9787 4597 9813
rect 4623 9787 4649 9813
rect 4675 9787 4701 9813
rect 4727 9787 7257 9813
rect 7283 9787 7309 9813
rect 7335 9787 7361 9813
rect 7387 9787 9917 9813
rect 9943 9787 9969 9813
rect 9995 9787 10021 9813
rect 10047 9787 11312 9813
rect 672 9770 11312 9787
rect 2479 9729 2505 9735
rect 2479 9697 2505 9703
rect 8303 9729 8329 9735
rect 8303 9697 8329 9703
rect 2305 9647 2311 9673
rect 2337 9647 2343 9673
rect 8135 9617 8161 9623
rect 8471 9617 8497 9623
rect 5497 9591 5503 9617
rect 5529 9591 5535 9617
rect 7401 9591 7407 9617
rect 7433 9591 7439 9617
rect 8297 9591 8303 9617
rect 8329 9591 8335 9617
rect 8135 9585 8161 9591
rect 8471 9585 8497 9591
rect 8919 9617 8945 9623
rect 8919 9585 8945 9591
rect 9199 9617 9225 9623
rect 9199 9585 9225 9591
rect 2143 9561 2169 9567
rect 2143 9529 2169 9535
rect 2535 9561 2561 9567
rect 2535 9529 2561 9535
rect 3879 9561 3905 9567
rect 3879 9529 3905 9535
rect 4159 9561 4185 9567
rect 8079 9561 8105 9567
rect 5609 9535 5615 9561
rect 5641 9535 5647 9561
rect 7513 9535 7519 9561
rect 7545 9535 7551 9561
rect 4159 9529 4185 9535
rect 8079 9529 8105 9535
rect 10039 9561 10065 9567
rect 10039 9529 10065 9535
rect 10823 9561 10849 9567
rect 10823 9529 10849 9535
rect 11103 9561 11129 9567
rect 11103 9529 11129 9535
rect 2255 9505 2281 9511
rect 2255 9473 2281 9479
rect 3935 9505 3961 9511
rect 3935 9473 3961 9479
rect 4047 9505 4073 9511
rect 4047 9473 4073 9479
rect 8751 9505 8777 9511
rect 8751 9473 8777 9479
rect 8863 9505 8889 9511
rect 8863 9473 8889 9479
rect 8975 9505 9001 9511
rect 8975 9473 9001 9479
rect 9143 9505 9169 9511
rect 9143 9473 9169 9479
rect 9871 9505 9897 9511
rect 9871 9473 9897 9479
rect 10935 9505 10961 9511
rect 10935 9473 10961 9479
rect 672 9421 11392 9438
rect 672 9395 3267 9421
rect 3293 9395 3319 9421
rect 3345 9395 3371 9421
rect 3397 9395 5927 9421
rect 5953 9395 5979 9421
rect 6005 9395 6031 9421
rect 6057 9395 8587 9421
rect 8613 9395 8639 9421
rect 8665 9395 8691 9421
rect 8717 9395 11247 9421
rect 11273 9395 11299 9421
rect 11325 9395 11351 9421
rect 11377 9395 11392 9421
rect 672 9378 11392 9395
rect 2423 9337 2449 9343
rect 2423 9305 2449 9311
rect 5503 9337 5529 9343
rect 9143 9337 9169 9343
rect 8017 9311 8023 9337
rect 8049 9311 8055 9337
rect 5503 9305 5529 9311
rect 9143 9305 9169 9311
rect 10543 9337 10569 9343
rect 10543 9305 10569 9311
rect 2871 9281 2897 9287
rect 1633 9255 1639 9281
rect 1665 9255 1671 9281
rect 2871 9249 2897 9255
rect 2927 9281 2953 9287
rect 2927 9249 2953 9255
rect 4327 9281 4353 9287
rect 6343 9281 6369 9287
rect 7407 9281 7433 9287
rect 4769 9255 4775 9281
rect 4801 9255 4807 9281
rect 6673 9255 6679 9281
rect 6705 9255 6711 9281
rect 4327 9249 4353 9255
rect 6343 9249 6369 9255
rect 7407 9249 7433 9255
rect 7855 9281 7881 9287
rect 7855 9249 7881 9255
rect 9759 9281 9785 9287
rect 9759 9249 9785 9255
rect 2031 9225 2057 9231
rect 1521 9199 1527 9225
rect 1553 9199 1559 9225
rect 1801 9199 1807 9225
rect 1833 9199 1839 9225
rect 2031 9193 2057 9199
rect 2087 9225 2113 9231
rect 2087 9193 2113 9199
rect 2143 9225 2169 9231
rect 2759 9225 2785 9231
rect 2361 9199 2367 9225
rect 2393 9199 2399 9225
rect 2143 9193 2169 9199
rect 2759 9193 2785 9199
rect 4943 9225 4969 9231
rect 4943 9193 4969 9199
rect 5559 9225 5585 9231
rect 6175 9225 6201 9231
rect 5777 9199 5783 9225
rect 5809 9199 5815 9225
rect 5945 9199 5951 9225
rect 5977 9199 5983 9225
rect 5559 9193 5585 9199
rect 6175 9193 6201 9199
rect 6287 9225 6313 9231
rect 6287 9193 6313 9199
rect 6511 9225 6537 9231
rect 10599 9225 10625 9231
rect 9249 9199 9255 9225
rect 9281 9199 9287 9225
rect 10313 9199 10319 9225
rect 10345 9199 10351 9225
rect 10481 9199 10487 9225
rect 10513 9199 10519 9225
rect 6511 9193 6537 9199
rect 10599 9193 10625 9199
rect 2479 9169 2505 9175
rect 2479 9137 2505 9143
rect 3151 9169 3177 9175
rect 3151 9137 3177 9143
rect 4103 9169 4129 9175
rect 4103 9137 4129 9143
rect 10039 9169 10065 9175
rect 10039 9137 10065 9143
rect 2591 9113 2617 9119
rect 2591 9081 2617 9087
rect 3095 9113 3121 9119
rect 3095 9081 3121 9087
rect 4159 9113 4185 9119
rect 4159 9081 4185 9087
rect 4271 9113 4297 9119
rect 4271 9081 4297 9087
rect 5447 9113 5473 9119
rect 5447 9081 5473 9087
rect 5671 9113 5697 9119
rect 5671 9081 5697 9087
rect 6063 9113 6089 9119
rect 6063 9081 6089 9087
rect 7071 9113 7097 9119
rect 7071 9081 7097 9087
rect 7127 9113 7153 9119
rect 7127 9081 7153 9087
rect 7239 9113 7265 9119
rect 7239 9081 7265 9087
rect 7351 9113 7377 9119
rect 7351 9081 7377 9087
rect 9087 9113 9113 9119
rect 9087 9081 9113 9087
rect 9703 9113 9729 9119
rect 9703 9081 9729 9087
rect 9871 9113 9897 9119
rect 9871 9081 9897 9087
rect 10095 9113 10121 9119
rect 10095 9081 10121 9087
rect 10207 9113 10233 9119
rect 10207 9081 10233 9087
rect 10711 9113 10737 9119
rect 10711 9081 10737 9087
rect 672 9029 11312 9046
rect 672 9003 1937 9029
rect 1963 9003 1989 9029
rect 2015 9003 2041 9029
rect 2067 9003 4597 9029
rect 4623 9003 4649 9029
rect 4675 9003 4701 9029
rect 4727 9003 7257 9029
rect 7283 9003 7309 9029
rect 7335 9003 7361 9029
rect 7387 9003 9917 9029
rect 9943 9003 9969 9029
rect 9995 9003 10021 9029
rect 10047 9003 11312 9029
rect 672 8986 11312 9003
rect 2311 8945 2337 8951
rect 2311 8913 2337 8919
rect 2479 8945 2505 8951
rect 2479 8913 2505 8919
rect 4271 8945 4297 8951
rect 4271 8913 4297 8919
rect 5447 8945 5473 8951
rect 5447 8913 5473 8919
rect 5671 8945 5697 8951
rect 5671 8913 5697 8919
rect 6063 8945 6089 8951
rect 6063 8913 6089 8919
rect 7687 8945 7713 8951
rect 7687 8913 7713 8919
rect 10263 8945 10289 8951
rect 10263 8913 10289 8919
rect 1919 8889 1945 8895
rect 1919 8857 1945 8863
rect 5503 8889 5529 8895
rect 5503 8857 5529 8863
rect 5951 8889 5977 8895
rect 10145 8863 10151 8889
rect 10177 8863 10183 8889
rect 5951 8857 5977 8863
rect 1975 8833 2001 8839
rect 3991 8833 4017 8839
rect 2305 8807 2311 8833
rect 2337 8807 2343 8833
rect 1975 8801 2001 8807
rect 3991 8801 4017 8807
rect 4047 8833 4073 8839
rect 4047 8801 4073 8807
rect 4159 8833 4185 8839
rect 4159 8801 4185 8807
rect 5615 8833 5641 8839
rect 6169 8807 6175 8833
rect 6201 8807 6207 8833
rect 7513 8807 7519 8833
rect 7545 8807 7551 8833
rect 10089 8807 10095 8833
rect 10121 8807 10127 8833
rect 5615 8801 5641 8807
rect 2087 8777 2113 8783
rect 2087 8745 2113 8751
rect 1863 8721 1889 8727
rect 1863 8689 1889 8695
rect 3991 8721 4017 8727
rect 3991 8689 4017 8695
rect 6119 8721 6145 8727
rect 6119 8689 6145 8695
rect 7631 8721 7657 8727
rect 7631 8689 7657 8695
rect 672 8637 11392 8654
rect 672 8611 3267 8637
rect 3293 8611 3319 8637
rect 3345 8611 3371 8637
rect 3397 8611 5927 8637
rect 5953 8611 5979 8637
rect 6005 8611 6031 8637
rect 6057 8611 8587 8637
rect 8613 8611 8639 8637
rect 8665 8611 8691 8637
rect 8717 8611 11247 8637
rect 11273 8611 11299 8637
rect 11325 8611 11351 8637
rect 11377 8611 11392 8637
rect 672 8594 11392 8611
rect 2983 8553 3009 8559
rect 6175 8553 6201 8559
rect 2641 8527 2647 8553
rect 2673 8527 2679 8553
rect 4097 8527 4103 8553
rect 4129 8527 4135 8553
rect 2983 8521 3009 8527
rect 6175 8521 6201 8527
rect 10935 8497 10961 8503
rect 2809 8471 2815 8497
rect 2841 8471 2847 8497
rect 6001 8471 6007 8497
rect 6033 8471 6039 8497
rect 10935 8465 10961 8471
rect 3207 8441 3233 8447
rect 10823 8441 10849 8447
rect 2529 8415 2535 8441
rect 2561 8415 2567 8441
rect 4209 8415 4215 8441
rect 4241 8415 4247 8441
rect 10033 8415 10039 8441
rect 10065 8415 10071 8441
rect 3207 8409 3233 8415
rect 10823 8409 10849 8415
rect 11103 8441 11129 8447
rect 11103 8409 11129 8415
rect 9871 8329 9897 8335
rect 9871 8297 9897 8303
rect 10039 8329 10065 8335
rect 10039 8297 10065 8303
rect 672 8245 11312 8262
rect 672 8219 1937 8245
rect 1963 8219 1989 8245
rect 2015 8219 2041 8245
rect 2067 8219 4597 8245
rect 4623 8219 4649 8245
rect 4675 8219 4701 8245
rect 4727 8219 7257 8245
rect 7283 8219 7309 8245
rect 7335 8219 7361 8245
rect 7387 8219 9917 8245
rect 9943 8219 9969 8245
rect 9995 8219 10021 8245
rect 10047 8219 11312 8245
rect 672 8202 11312 8219
rect 6791 8161 6817 8167
rect 6791 8129 6817 8135
rect 9087 8161 9113 8167
rect 9087 8129 9113 8135
rect 9983 8105 10009 8111
rect 9529 8079 9535 8105
rect 9561 8079 9567 8105
rect 9983 8073 10009 8079
rect 6903 8049 6929 8055
rect 9031 8049 9057 8055
rect 9871 8049 9897 8055
rect 7009 8023 7015 8049
rect 7041 8023 7047 8049
rect 9193 8023 9199 8049
rect 9225 8023 9231 8049
rect 9585 8023 9591 8049
rect 9617 8023 9623 8049
rect 9753 8023 9759 8049
rect 9785 8023 9791 8049
rect 6903 8017 6929 8023
rect 9031 8017 9057 8023
rect 9871 8017 9897 8023
rect 10207 8049 10233 8055
rect 10207 8017 10233 8023
rect 1695 7993 1721 7999
rect 1695 7961 1721 7967
rect 1751 7993 1777 7999
rect 1751 7961 1777 7967
rect 1919 7993 1945 7999
rect 1919 7961 1945 7967
rect 8863 7993 8889 7999
rect 8863 7961 8889 7967
rect 9423 7993 9449 7999
rect 9423 7961 9449 7967
rect 10319 7993 10345 7999
rect 10319 7961 10345 7967
rect 1639 7937 1665 7943
rect 1639 7905 1665 7911
rect 1975 7937 2001 7943
rect 1975 7905 2001 7911
rect 2031 7937 2057 7943
rect 4719 7937 4745 7943
rect 4545 7911 4551 7937
rect 4577 7911 4583 7937
rect 2031 7905 2057 7911
rect 4719 7905 4745 7911
rect 6959 7937 6985 7943
rect 6959 7905 6985 7911
rect 9255 7937 9281 7943
rect 9255 7905 9281 7911
rect 9815 7937 9841 7943
rect 9815 7905 9841 7911
rect 10263 7937 10289 7943
rect 10263 7905 10289 7911
rect 672 7853 11392 7870
rect 672 7827 3267 7853
rect 3293 7827 3319 7853
rect 3345 7827 3371 7853
rect 3397 7827 5927 7853
rect 5953 7827 5979 7853
rect 6005 7827 6031 7853
rect 6057 7827 8587 7853
rect 8613 7827 8639 7853
rect 8665 7827 8691 7853
rect 8717 7827 11247 7853
rect 11273 7827 11299 7853
rect 11325 7827 11351 7853
rect 11377 7827 11392 7853
rect 672 7810 11392 7827
rect 7407 7769 7433 7775
rect 3985 7743 3991 7769
rect 4017 7743 4023 7769
rect 7407 7737 7433 7743
rect 10375 7769 10401 7775
rect 10375 7737 10401 7743
rect 1135 7713 1161 7719
rect 1135 7681 1161 7687
rect 1247 7713 1273 7719
rect 1247 7681 1273 7687
rect 1695 7713 1721 7719
rect 1695 7681 1721 7687
rect 2143 7713 2169 7719
rect 9871 7713 9897 7719
rect 6057 7687 6063 7713
rect 6089 7687 6095 7713
rect 7233 7687 7239 7713
rect 7265 7687 7271 7713
rect 2143 7681 2169 7687
rect 9871 7681 9897 7687
rect 10319 7713 10345 7719
rect 10319 7681 10345 7687
rect 10431 7713 10457 7719
rect 10431 7681 10457 7687
rect 1527 7657 1553 7663
rect 1975 7657 2001 7663
rect 1857 7631 1863 7657
rect 1889 7631 1895 7657
rect 1527 7625 1553 7631
rect 1975 7625 2001 7631
rect 4831 7657 4857 7663
rect 4831 7625 4857 7631
rect 6231 7657 6257 7663
rect 6231 7625 6257 7631
rect 10039 7657 10065 7663
rect 10039 7625 10065 7631
rect 10095 7657 10121 7663
rect 10095 7625 10121 7631
rect 1191 7601 1217 7607
rect 1191 7569 1217 7575
rect 1471 7601 1497 7607
rect 1471 7569 1497 7575
rect 1639 7601 1665 7607
rect 1639 7569 1665 7575
rect 2087 7601 2113 7607
rect 2087 7569 2113 7575
rect 2367 7601 2393 7607
rect 2367 7569 2393 7575
rect 4271 7601 4297 7607
rect 4271 7569 4297 7575
rect 4775 7601 4801 7607
rect 4775 7569 4801 7575
rect 4943 7601 4969 7607
rect 4943 7569 4969 7575
rect 4999 7601 5025 7607
rect 4999 7569 5025 7575
rect 9703 7601 9729 7607
rect 9703 7569 9729 7575
rect 9927 7601 9953 7607
rect 9927 7569 9953 7575
rect 4159 7545 4185 7551
rect 4159 7513 4185 7519
rect 672 7461 11312 7478
rect 672 7435 1937 7461
rect 1963 7435 1989 7461
rect 2015 7435 2041 7461
rect 2067 7435 4597 7461
rect 4623 7435 4649 7461
rect 4675 7435 4701 7461
rect 4727 7435 7257 7461
rect 7283 7435 7309 7461
rect 7335 7435 7361 7461
rect 7387 7435 9917 7461
rect 9943 7435 9969 7461
rect 9995 7435 10021 7461
rect 10047 7435 11312 7461
rect 672 7418 11312 7435
rect 1751 7377 1777 7383
rect 1751 7345 1777 7351
rect 2199 7377 2225 7383
rect 2199 7345 2225 7351
rect 3823 7377 3849 7383
rect 3823 7345 3849 7351
rect 3935 7377 3961 7383
rect 3935 7345 3961 7351
rect 4271 7377 4297 7383
rect 4271 7345 4297 7351
rect 4383 7377 4409 7383
rect 4383 7345 4409 7351
rect 5783 7377 5809 7383
rect 5783 7345 5809 7351
rect 7575 7377 7601 7383
rect 7575 7345 7601 7351
rect 9983 7321 10009 7327
rect 1857 7295 1863 7321
rect 1889 7295 1895 7321
rect 7793 7295 7799 7321
rect 7825 7295 7831 7321
rect 9809 7295 9815 7321
rect 9841 7295 9847 7321
rect 9983 7289 10009 7295
rect 5671 7265 5697 7271
rect 1913 7239 1919 7265
rect 1945 7239 1951 7265
rect 4041 7239 4047 7265
rect 4073 7239 4079 7265
rect 4489 7239 4495 7265
rect 4521 7239 4527 7265
rect 5385 7239 5391 7265
rect 5417 7239 5423 7265
rect 5671 7233 5697 7239
rect 5895 7265 5921 7271
rect 7015 7265 7041 7271
rect 7463 7265 7489 7271
rect 6337 7239 6343 7265
rect 6369 7239 6375 7265
rect 6897 7239 6903 7265
rect 6929 7239 6935 7265
rect 7177 7239 7183 7265
rect 7209 7239 7215 7265
rect 7345 7239 7351 7265
rect 7377 7239 7383 7265
rect 10145 7239 10151 7265
rect 10177 7239 10183 7265
rect 5895 7233 5921 7239
rect 7015 7233 7041 7239
rect 7463 7233 7489 7239
rect 2255 7209 2281 7215
rect 2255 7177 2281 7183
rect 3767 7209 3793 7215
rect 3767 7177 3793 7183
rect 4215 7209 4241 7215
rect 6791 7209 6817 7215
rect 5497 7183 5503 7209
rect 5529 7183 5535 7209
rect 4215 7177 4241 7183
rect 6791 7177 6817 7183
rect 7631 7209 7657 7215
rect 7631 7177 7657 7183
rect 7855 7209 7881 7215
rect 7855 7177 7881 7183
rect 7967 7209 7993 7215
rect 7967 7177 7993 7183
rect 9647 7209 9673 7215
rect 9647 7177 9673 7183
rect 2199 7153 2225 7159
rect 2199 7121 2225 7127
rect 6119 7153 6145 7159
rect 7183 7153 7209 7159
rect 6225 7127 6231 7153
rect 6257 7127 6263 7153
rect 6119 7121 6145 7127
rect 7183 7121 7209 7127
rect 9759 7153 9785 7159
rect 9759 7121 9785 7127
rect 10039 7153 10065 7159
rect 10039 7121 10065 7127
rect 672 7069 11392 7086
rect 672 7043 3267 7069
rect 3293 7043 3319 7069
rect 3345 7043 3371 7069
rect 3397 7043 5927 7069
rect 5953 7043 5979 7069
rect 6005 7043 6031 7069
rect 6057 7043 8587 7069
rect 8613 7043 8639 7069
rect 8665 7043 8691 7069
rect 8717 7043 11247 7069
rect 11273 7043 11299 7069
rect 11325 7043 11351 7069
rect 11377 7043 11392 7069
rect 672 7026 11392 7043
rect 7295 6985 7321 6991
rect 7121 6959 7127 6985
rect 7153 6959 7159 6985
rect 7295 6953 7321 6959
rect 7967 6985 7993 6991
rect 7967 6953 7993 6959
rect 9591 6985 9617 6991
rect 9591 6953 9617 6959
rect 7519 6929 7545 6935
rect 7519 6897 7545 6903
rect 7855 6929 7881 6935
rect 7855 6897 7881 6903
rect 9143 6929 9169 6935
rect 9143 6897 9169 6903
rect 9983 6929 10009 6935
rect 9983 6897 10009 6903
rect 10263 6929 10289 6935
rect 10263 6897 10289 6903
rect 10935 6929 10961 6935
rect 10935 6897 10961 6903
rect 1919 6873 1945 6879
rect 1919 6841 1945 6847
rect 4999 6873 5025 6879
rect 4999 6841 5025 6847
rect 5111 6873 5137 6879
rect 5111 6841 5137 6847
rect 5223 6873 5249 6879
rect 5223 6841 5249 6847
rect 5503 6873 5529 6879
rect 5503 6841 5529 6847
rect 5615 6873 5641 6879
rect 5615 6841 5641 6847
rect 5727 6873 5753 6879
rect 7799 6873 7825 6879
rect 5833 6847 5839 6873
rect 5865 6847 5871 6873
rect 5727 6841 5753 6847
rect 7799 6841 7825 6847
rect 9199 6873 9225 6879
rect 9199 6841 9225 6847
rect 9311 6873 9337 6879
rect 9759 6873 9785 6879
rect 9417 6847 9423 6873
rect 9449 6847 9455 6873
rect 9585 6847 9591 6873
rect 9617 6847 9623 6873
rect 9311 6841 9337 6847
rect 9759 6841 9785 6847
rect 9815 6873 9841 6879
rect 9815 6841 9841 6847
rect 11103 6873 11129 6879
rect 11103 6841 11129 6847
rect 4943 6817 4969 6823
rect 10207 6817 10233 6823
rect 7457 6791 7463 6817
rect 7489 6791 7495 6817
rect 4943 6785 4969 6791
rect 10207 6785 10233 6791
rect 10823 6817 10849 6823
rect 10823 6785 10849 6791
rect 1807 6761 1833 6767
rect 1633 6735 1639 6761
rect 1665 6735 1671 6761
rect 1807 6729 1833 6735
rect 5279 6761 5305 6767
rect 5279 6729 5305 6735
rect 5447 6761 5473 6767
rect 5447 6729 5473 6735
rect 7631 6761 7657 6767
rect 7631 6729 7657 6735
rect 10151 6761 10177 6767
rect 10151 6729 10177 6735
rect 672 6677 11312 6694
rect 672 6651 1937 6677
rect 1963 6651 1989 6677
rect 2015 6651 2041 6677
rect 2067 6651 4597 6677
rect 4623 6651 4649 6677
rect 4675 6651 4701 6677
rect 4727 6651 7257 6677
rect 7283 6651 7309 6677
rect 7335 6651 7361 6677
rect 7387 6651 9917 6677
rect 9943 6651 9969 6677
rect 9995 6651 10021 6677
rect 10047 6651 11312 6677
rect 672 6634 11312 6651
rect 9591 6593 9617 6599
rect 9591 6561 9617 6567
rect 9647 6593 9673 6599
rect 9647 6561 9673 6567
rect 2815 6537 2841 6543
rect 4377 6511 4383 6537
rect 4409 6511 4415 6537
rect 10145 6511 10151 6537
rect 10177 6511 10183 6537
rect 2815 6505 2841 6511
rect 1751 6481 1777 6487
rect 1751 6449 1777 6455
rect 4215 6481 4241 6487
rect 9759 6481 9785 6487
rect 7289 6455 7295 6481
rect 7321 6455 7327 6481
rect 4215 6449 4241 6455
rect 9759 6449 9785 6455
rect 9815 6481 9841 6487
rect 9815 6449 9841 6455
rect 10039 6481 10065 6487
rect 10201 6455 10207 6481
rect 10233 6455 10239 6481
rect 10039 6449 10065 6455
rect 4103 6425 4129 6431
rect 4103 6393 4129 6399
rect 2871 6369 2897 6375
rect 1913 6343 1919 6369
rect 1945 6343 1951 6369
rect 2871 6337 2897 6343
rect 4327 6369 4353 6375
rect 4327 6337 4353 6343
rect 4383 6369 4409 6375
rect 7177 6343 7183 6369
rect 7209 6343 7215 6369
rect 4383 6337 4409 6343
rect 672 6285 11392 6302
rect 672 6259 3267 6285
rect 3293 6259 3319 6285
rect 3345 6259 3371 6285
rect 3397 6259 5927 6285
rect 5953 6259 5979 6285
rect 6005 6259 6031 6285
rect 6057 6259 8587 6285
rect 8613 6259 8639 6285
rect 8665 6259 8691 6285
rect 8717 6259 11247 6285
rect 11273 6259 11299 6285
rect 11325 6259 11351 6285
rect 11377 6259 11392 6285
rect 672 6242 11392 6259
rect 3319 6201 3345 6207
rect 3319 6169 3345 6175
rect 4775 6201 4801 6207
rect 4775 6169 4801 6175
rect 4831 6201 4857 6207
rect 9753 6175 9759 6201
rect 9785 6175 9791 6201
rect 4831 6169 4857 6175
rect 2703 6145 2729 6151
rect 3929 6119 3935 6145
rect 3961 6119 3967 6145
rect 2703 6113 2729 6119
rect 2759 6089 2785 6095
rect 1969 6063 1975 6089
rect 2001 6063 2007 6089
rect 2759 6057 2785 6063
rect 2983 6089 3009 6095
rect 2983 6057 3009 6063
rect 3207 6089 3233 6095
rect 4887 6089 4913 6095
rect 9815 6089 9841 6095
rect 3817 6063 3823 6089
rect 3849 6063 3855 6089
rect 5049 6063 5055 6089
rect 5081 6063 5087 6089
rect 9585 6063 9591 6089
rect 9617 6063 9623 6089
rect 3207 6057 3233 6063
rect 4887 6057 4913 6063
rect 9815 6057 9841 6063
rect 9983 6089 10009 6095
rect 9983 6057 10009 6063
rect 1639 6033 1665 6039
rect 3263 6033 3289 6039
rect 2025 6007 2031 6033
rect 2057 6007 2063 6033
rect 1639 6001 1665 6007
rect 3263 6001 3289 6007
rect 9759 5977 9785 5983
rect 9759 5945 9785 5951
rect 672 5893 11312 5910
rect 672 5867 1937 5893
rect 1963 5867 1989 5893
rect 2015 5867 2041 5893
rect 2067 5867 4597 5893
rect 4623 5867 4649 5893
rect 4675 5867 4701 5893
rect 4727 5867 7257 5893
rect 7283 5867 7309 5893
rect 7335 5867 7361 5893
rect 7387 5867 9917 5893
rect 9943 5867 9969 5893
rect 9995 5867 10021 5893
rect 10047 5867 11312 5893
rect 672 5850 11312 5867
rect 4383 5809 4409 5815
rect 4383 5777 4409 5783
rect 2311 5753 2337 5759
rect 7513 5727 7519 5753
rect 7545 5727 7551 5753
rect 2311 5721 2337 5727
rect 2367 5697 2393 5703
rect 2367 5665 2393 5671
rect 4887 5697 4913 5703
rect 4887 5665 4913 5671
rect 5111 5697 5137 5703
rect 5111 5665 5137 5671
rect 5223 5697 5249 5703
rect 5223 5665 5249 5671
rect 9983 5697 10009 5703
rect 9983 5665 10009 5671
rect 4439 5641 4465 5647
rect 4439 5609 4465 5615
rect 4551 5641 4577 5647
rect 7575 5641 7601 5647
rect 7177 5615 7183 5641
rect 7209 5615 7215 5641
rect 4551 5609 4577 5615
rect 7575 5609 7601 5615
rect 7687 5641 7713 5647
rect 7687 5609 7713 5615
rect 5167 5585 5193 5591
rect 5167 5553 5193 5559
rect 7351 5585 7377 5591
rect 10145 5559 10151 5585
rect 10177 5559 10183 5585
rect 7351 5553 7377 5559
rect 672 5501 11392 5518
rect 672 5475 3267 5501
rect 3293 5475 3319 5501
rect 3345 5475 3371 5501
rect 3397 5475 5927 5501
rect 5953 5475 5979 5501
rect 6005 5475 6031 5501
rect 6057 5475 8587 5501
rect 8613 5475 8639 5501
rect 8665 5475 8691 5501
rect 8717 5475 11247 5501
rect 11273 5475 11299 5501
rect 11325 5475 11351 5501
rect 11377 5475 11392 5501
rect 672 5458 11392 5475
rect 1135 5417 1161 5423
rect 1135 5385 1161 5391
rect 7127 5417 7153 5423
rect 7127 5385 7153 5391
rect 7239 5417 7265 5423
rect 7239 5385 7265 5391
rect 7967 5417 7993 5423
rect 7967 5385 7993 5391
rect 9647 5417 9673 5423
rect 10935 5417 10961 5423
rect 10201 5391 10207 5417
rect 10233 5391 10239 5417
rect 9647 5385 9673 5391
rect 10935 5385 10961 5391
rect 6455 5361 6481 5367
rect 1297 5335 1303 5361
rect 1329 5335 1335 5361
rect 6455 5329 6481 5335
rect 9199 5361 9225 5367
rect 9199 5329 9225 5335
rect 10039 5361 10065 5367
rect 10039 5329 10065 5335
rect 6567 5305 6593 5311
rect 1633 5279 1639 5305
rect 1665 5279 1671 5305
rect 6567 5273 6593 5279
rect 6735 5305 6761 5311
rect 7463 5305 7489 5311
rect 7289 5279 7295 5305
rect 7321 5279 7327 5305
rect 6735 5273 6761 5279
rect 7463 5273 7489 5279
rect 7911 5305 7937 5311
rect 9871 5305 9897 5311
rect 11103 5305 11129 5311
rect 9473 5279 9479 5305
rect 9505 5279 9511 5305
rect 9641 5279 9647 5305
rect 9673 5279 9679 5305
rect 10313 5279 10319 5305
rect 10345 5279 10351 5305
rect 7911 5273 7937 5279
rect 9871 5273 9897 5279
rect 11103 5273 11129 5279
rect 1975 5249 2001 5255
rect 9367 5249 9393 5255
rect 1577 5223 1583 5249
rect 1609 5223 1615 5249
rect 7177 5223 7183 5249
rect 7209 5223 7215 5249
rect 1975 5217 2001 5223
rect 9367 5217 9393 5223
rect 10823 5249 10849 5255
rect 10823 5217 10849 5223
rect 6511 5193 6537 5199
rect 6511 5161 6537 5167
rect 6847 5193 6873 5199
rect 6847 5161 6873 5167
rect 7575 5193 7601 5199
rect 7575 5161 7601 5167
rect 7799 5193 7825 5199
rect 7799 5161 7825 5167
rect 7967 5193 7993 5199
rect 7967 5161 7993 5167
rect 9255 5193 9281 5199
rect 9753 5167 9759 5193
rect 9785 5167 9791 5193
rect 9255 5161 9281 5167
rect 672 5109 11312 5126
rect 672 5083 1937 5109
rect 1963 5083 1989 5109
rect 2015 5083 2041 5109
rect 2067 5083 4597 5109
rect 4623 5083 4649 5109
rect 4675 5083 4701 5109
rect 4727 5083 7257 5109
rect 7283 5083 7309 5109
rect 7335 5083 7361 5109
rect 7387 5083 9917 5109
rect 9943 5083 9969 5109
rect 9995 5083 10021 5109
rect 10047 5083 11312 5109
rect 672 5066 11312 5083
rect 2031 5025 2057 5031
rect 2031 4993 2057 4999
rect 4999 5025 5025 5031
rect 4999 4993 5025 4999
rect 9759 5025 9785 5031
rect 9759 4993 9785 4999
rect 4271 4969 4297 4975
rect 4271 4937 4297 4943
rect 4495 4969 4521 4975
rect 4495 4937 4521 4943
rect 4607 4969 4633 4975
rect 4607 4937 4633 4943
rect 7015 4969 7041 4975
rect 7015 4937 7041 4943
rect 7575 4969 7601 4975
rect 7575 4937 7601 4943
rect 9703 4969 9729 4975
rect 9703 4937 9729 4943
rect 9927 4969 9953 4975
rect 9927 4937 9953 4943
rect 2143 4913 2169 4919
rect 2143 4881 2169 4887
rect 4943 4913 4969 4919
rect 7687 4913 7713 4919
rect 9983 4913 10009 4919
rect 5441 4887 5447 4913
rect 5473 4887 5479 4913
rect 9361 4887 9367 4913
rect 9393 4887 9399 4913
rect 10089 4887 10095 4913
rect 10121 4887 10127 4913
rect 4943 4881 4969 4887
rect 7687 4881 7713 4887
rect 9983 4881 10009 4887
rect 4215 4857 4241 4863
rect 4215 4825 4241 4831
rect 4327 4857 4353 4863
rect 4327 4825 4353 4831
rect 5167 4857 5193 4863
rect 6959 4857 6985 4863
rect 5273 4831 5279 4857
rect 5305 4831 5311 4857
rect 5167 4825 5193 4831
rect 6959 4825 6985 4831
rect 7351 4857 7377 4863
rect 7351 4825 7377 4831
rect 7463 4857 7489 4863
rect 9647 4857 9673 4863
rect 9249 4831 9255 4857
rect 9281 4831 9287 4857
rect 7463 4825 7489 4831
rect 9647 4825 9673 4831
rect 5335 4801 5361 4807
rect 1857 4775 1863 4801
rect 1889 4775 1895 4801
rect 4769 4775 4775 4801
rect 4801 4775 4807 4801
rect 5335 4769 5361 4775
rect 672 4717 11392 4734
rect 672 4691 3267 4717
rect 3293 4691 3319 4717
rect 3345 4691 3371 4717
rect 3397 4691 5927 4717
rect 5953 4691 5979 4717
rect 6005 4691 6031 4717
rect 6057 4691 8587 4717
rect 8613 4691 8639 4717
rect 8665 4691 8691 4717
rect 8717 4691 11247 4717
rect 11273 4691 11299 4717
rect 11325 4691 11351 4717
rect 11377 4691 11392 4717
rect 672 4674 11392 4691
rect 5391 4633 5417 4639
rect 5391 4601 5417 4607
rect 7407 4633 7433 4639
rect 7407 4601 7433 4607
rect 9927 4633 9953 4639
rect 9927 4601 9953 4607
rect 5447 4577 5473 4583
rect 5447 4545 5473 4551
rect 7351 4577 7377 4583
rect 9753 4551 9759 4577
rect 9785 4551 9791 4577
rect 7351 4545 7377 4551
rect 1807 4521 1833 4527
rect 1807 4489 1833 4495
rect 1919 4521 1945 4527
rect 1919 4489 1945 4495
rect 2087 4521 2113 4527
rect 2087 4489 2113 4495
rect 2255 4521 2281 4527
rect 5167 4521 5193 4527
rect 2473 4495 2479 4521
rect 2505 4495 2511 4521
rect 4993 4495 4999 4521
rect 5025 4495 5031 4521
rect 9641 4495 9647 4521
rect 9673 4495 9679 4521
rect 10033 4495 10039 4521
rect 10065 4495 10071 4521
rect 2255 4489 2281 4495
rect 5167 4489 5193 4495
rect 1975 4465 2001 4471
rect 1975 4433 2001 4439
rect 2703 4465 2729 4471
rect 2703 4433 2729 4439
rect 5111 4465 5137 4471
rect 5111 4433 5137 4439
rect 5391 4409 5417 4415
rect 5391 4377 5417 4383
rect 672 4325 11312 4342
rect 672 4299 1937 4325
rect 1963 4299 1989 4325
rect 2015 4299 2041 4325
rect 2067 4299 4597 4325
rect 4623 4299 4649 4325
rect 4675 4299 4701 4325
rect 4727 4299 7257 4325
rect 7283 4299 7309 4325
rect 7335 4299 7361 4325
rect 7387 4299 9917 4325
rect 9943 4299 9969 4325
rect 9995 4299 10021 4325
rect 10047 4299 11312 4325
rect 672 4282 11312 4299
rect 9759 4241 9785 4247
rect 9759 4209 9785 4215
rect 2871 4185 2897 4191
rect 2871 4153 2897 4159
rect 4439 4185 4465 4191
rect 4439 4153 4465 4159
rect 4551 4185 4577 4191
rect 4551 4153 4577 4159
rect 4663 4185 4689 4191
rect 4663 4153 4689 4159
rect 5671 4185 5697 4191
rect 5671 4153 5697 4159
rect 7575 4185 7601 4191
rect 7575 4153 7601 4159
rect 1919 4129 1945 4135
rect 1577 4103 1583 4129
rect 1609 4103 1615 4129
rect 1919 4097 1945 4103
rect 2087 4129 2113 4135
rect 2983 4129 3009 4135
rect 2473 4103 2479 4129
rect 2505 4103 2511 4129
rect 2087 4097 2113 4103
rect 2983 4097 3009 4103
rect 3655 4129 3681 4135
rect 3655 4097 3681 4103
rect 3823 4129 3849 4135
rect 3823 4097 3849 4103
rect 4999 4129 5025 4135
rect 4999 4097 5025 4103
rect 5391 4129 5417 4135
rect 5391 4097 5417 4103
rect 7407 4129 7433 4135
rect 7407 4097 7433 4103
rect 7687 4129 7713 4135
rect 7687 4097 7713 4103
rect 9927 4129 9953 4135
rect 9927 4097 9953 4103
rect 10207 4129 10233 4135
rect 10207 4097 10233 4103
rect 3151 4073 3177 4079
rect 1689 4047 1695 4073
rect 1721 4047 1727 4073
rect 2361 4047 2367 4073
rect 2393 4047 2399 4073
rect 3151 4041 3177 4047
rect 3263 4073 3289 4079
rect 3263 4041 3289 4047
rect 3711 4073 3737 4079
rect 5615 4073 5641 4079
rect 5049 4047 5055 4073
rect 5081 4047 5087 4073
rect 5217 4047 5223 4073
rect 5249 4047 5255 4073
rect 3711 4041 3737 4047
rect 5615 4041 5641 4047
rect 5727 4073 5753 4079
rect 5727 4041 5753 4047
rect 7463 4073 7489 4079
rect 9815 4073 9841 4079
rect 9529 4047 9535 4073
rect 9561 4047 9567 4073
rect 7463 4041 7489 4047
rect 9815 4041 9841 4047
rect 10095 4073 10121 4079
rect 10095 4041 10121 4047
rect 10375 4073 10401 4079
rect 10375 4041 10401 4047
rect 10935 4073 10961 4079
rect 10935 4041 10961 4047
rect 11103 4073 11129 4079
rect 11103 4041 11129 4047
rect 2815 4017 2841 4023
rect 2815 3985 2841 3991
rect 4887 4017 4913 4023
rect 4887 3985 4913 3991
rect 5503 4017 5529 4023
rect 5503 3985 5529 3991
rect 7911 4017 7937 4023
rect 7911 3985 7937 3991
rect 9367 4017 9393 4023
rect 9367 3985 9393 3991
rect 10039 4017 10065 4023
rect 10039 3985 10065 3991
rect 10319 4017 10345 4023
rect 10319 3985 10345 3991
rect 10767 4017 10793 4023
rect 10767 3985 10793 3991
rect 672 3933 11392 3950
rect 672 3907 3267 3933
rect 3293 3907 3319 3933
rect 3345 3907 3371 3933
rect 3397 3907 5927 3933
rect 5953 3907 5979 3933
rect 6005 3907 6031 3933
rect 6057 3907 8587 3933
rect 8613 3907 8639 3933
rect 8665 3907 8691 3933
rect 8717 3907 11247 3933
rect 11273 3907 11299 3933
rect 11325 3907 11351 3933
rect 11377 3907 11392 3933
rect 672 3890 11392 3907
rect 2535 3849 2561 3855
rect 2535 3817 2561 3823
rect 4943 3849 4969 3855
rect 4943 3817 4969 3823
rect 5055 3849 5081 3855
rect 5055 3817 5081 3823
rect 7183 3849 7209 3855
rect 7183 3817 7209 3823
rect 2423 3793 2449 3799
rect 2423 3761 2449 3767
rect 5111 3793 5137 3799
rect 5559 3793 5585 3799
rect 5217 3767 5223 3793
rect 5249 3767 5255 3793
rect 5111 3761 5137 3767
rect 5559 3761 5585 3767
rect 7015 3793 7041 3799
rect 7015 3761 7041 3767
rect 7071 3793 7097 3799
rect 7071 3761 7097 3767
rect 7407 3793 7433 3799
rect 7407 3761 7433 3767
rect 7463 3793 7489 3799
rect 9977 3767 9983 3793
rect 10009 3767 10015 3793
rect 7463 3761 7489 3767
rect 2367 3737 2393 3743
rect 2367 3705 2393 3711
rect 2647 3737 2673 3743
rect 2647 3705 2673 3711
rect 7295 3737 7321 3743
rect 10151 3737 10177 3743
rect 7681 3711 7687 3737
rect 7713 3711 7719 3737
rect 7295 3705 7321 3711
rect 10151 3705 10177 3711
rect 11103 3737 11129 3743
rect 11103 3705 11129 3711
rect 2871 3681 2897 3687
rect 5329 3655 5335 3681
rect 5361 3655 5367 3681
rect 7457 3655 7463 3681
rect 7489 3655 7495 3681
rect 2871 3649 2897 3655
rect 672 3541 11312 3558
rect 672 3515 1937 3541
rect 1963 3515 1989 3541
rect 2015 3515 2041 3541
rect 2067 3515 4597 3541
rect 4623 3515 4649 3541
rect 4675 3515 4701 3541
rect 4727 3515 7257 3541
rect 7283 3515 7309 3541
rect 7335 3515 7361 3541
rect 7387 3515 9917 3541
rect 9943 3515 9969 3541
rect 9995 3515 10021 3541
rect 10047 3515 11312 3541
rect 672 3498 11312 3515
rect 7351 3457 7377 3463
rect 7351 3425 7377 3431
rect 7407 3401 7433 3407
rect 7407 3369 7433 3375
rect 7631 3401 7657 3407
rect 7631 3369 7657 3375
rect 672 3149 11392 3166
rect 672 3123 3267 3149
rect 3293 3123 3319 3149
rect 3345 3123 3371 3149
rect 3397 3123 5927 3149
rect 5953 3123 5979 3149
rect 6005 3123 6031 3149
rect 6057 3123 8587 3149
rect 8613 3123 8639 3149
rect 8665 3123 8691 3149
rect 8717 3123 11247 3149
rect 11273 3123 11299 3149
rect 11325 3123 11351 3149
rect 11377 3123 11392 3149
rect 672 3106 11392 3123
rect 672 2757 11312 2774
rect 672 2731 1937 2757
rect 1963 2731 1989 2757
rect 2015 2731 2041 2757
rect 2067 2731 4597 2757
rect 4623 2731 4649 2757
rect 4675 2731 4701 2757
rect 4727 2731 7257 2757
rect 7283 2731 7309 2757
rect 7335 2731 7361 2757
rect 7387 2731 9917 2757
rect 9943 2731 9969 2757
rect 9995 2731 10021 2757
rect 10047 2731 11312 2757
rect 672 2714 11312 2731
rect 10823 2561 10849 2567
rect 10823 2529 10849 2535
rect 11103 2561 11129 2567
rect 11103 2529 11129 2535
rect 10935 2505 10961 2511
rect 10935 2473 10961 2479
rect 672 2365 11392 2382
rect 672 2339 3267 2365
rect 3293 2339 3319 2365
rect 3345 2339 3371 2365
rect 3397 2339 5927 2365
rect 5953 2339 5979 2365
rect 6005 2339 6031 2365
rect 6057 2339 8587 2365
rect 8613 2339 8639 2365
rect 8665 2339 8691 2365
rect 8717 2339 11247 2365
rect 11273 2339 11299 2365
rect 11325 2339 11351 2365
rect 11377 2339 11392 2365
rect 672 2322 11392 2339
rect 672 1973 11312 1990
rect 672 1947 1937 1973
rect 1963 1947 1989 1973
rect 2015 1947 2041 1973
rect 2067 1947 4597 1973
rect 4623 1947 4649 1973
rect 4675 1947 4701 1973
rect 4727 1947 7257 1973
rect 7283 1947 7309 1973
rect 7335 1947 7361 1973
rect 7387 1947 9917 1973
rect 9943 1947 9969 1973
rect 9995 1947 10021 1973
rect 10047 1947 11312 1973
rect 672 1930 11312 1947
rect 672 1581 11392 1598
rect 672 1555 3267 1581
rect 3293 1555 3319 1581
rect 3345 1555 3371 1581
rect 3397 1555 5927 1581
rect 5953 1555 5979 1581
rect 6005 1555 6031 1581
rect 6057 1555 8587 1581
rect 8613 1555 8639 1581
rect 8665 1555 8691 1581
rect 8717 1555 11247 1581
rect 11273 1555 11299 1581
rect 11325 1555 11351 1581
rect 11377 1555 11392 1581
rect 672 1538 11392 1555
<< via1 >>
rect 3267 10179 3293 10205
rect 3319 10179 3345 10205
rect 3371 10179 3397 10205
rect 5927 10179 5953 10205
rect 5979 10179 6005 10205
rect 6031 10179 6057 10205
rect 8587 10179 8613 10205
rect 8639 10179 8665 10205
rect 8691 10179 8717 10205
rect 11247 10179 11273 10205
rect 11299 10179 11325 10205
rect 11351 10179 11377 10205
rect 1023 10039 1049 10065
rect 2143 10039 2169 10065
rect 3263 10039 3289 10065
rect 4663 10039 4689 10065
rect 5503 10039 5529 10065
rect 6623 10039 6649 10065
rect 7743 10039 7769 10065
rect 8863 10039 8889 10065
rect 10095 10039 10121 10065
rect 10375 10039 10401 10065
rect 11103 10039 11129 10065
rect 1135 9983 1161 10009
rect 2311 9983 2337 10009
rect 3431 9983 3457 10009
rect 4775 9983 4801 10009
rect 5615 9983 5641 10009
rect 6791 9983 6817 10009
rect 7855 9983 7881 10009
rect 8975 9983 9001 10009
rect 9927 9983 9953 10009
rect 10487 9983 10513 10009
rect 10935 9983 10961 10009
rect 1937 9787 1963 9813
rect 1989 9787 2015 9813
rect 2041 9787 2067 9813
rect 4597 9787 4623 9813
rect 4649 9787 4675 9813
rect 4701 9787 4727 9813
rect 7257 9787 7283 9813
rect 7309 9787 7335 9813
rect 7361 9787 7387 9813
rect 9917 9787 9943 9813
rect 9969 9787 9995 9813
rect 10021 9787 10047 9813
rect 2479 9703 2505 9729
rect 8303 9703 8329 9729
rect 2311 9647 2337 9673
rect 5503 9591 5529 9617
rect 7407 9591 7433 9617
rect 8135 9591 8161 9617
rect 8303 9591 8329 9617
rect 8471 9591 8497 9617
rect 8919 9591 8945 9617
rect 9199 9591 9225 9617
rect 2143 9535 2169 9561
rect 2535 9535 2561 9561
rect 3879 9535 3905 9561
rect 4159 9535 4185 9561
rect 5615 9535 5641 9561
rect 7519 9535 7545 9561
rect 8079 9535 8105 9561
rect 10039 9535 10065 9561
rect 10823 9535 10849 9561
rect 11103 9535 11129 9561
rect 2255 9479 2281 9505
rect 3935 9479 3961 9505
rect 4047 9479 4073 9505
rect 8751 9479 8777 9505
rect 8863 9479 8889 9505
rect 8975 9479 9001 9505
rect 9143 9479 9169 9505
rect 9871 9479 9897 9505
rect 10935 9479 10961 9505
rect 3267 9395 3293 9421
rect 3319 9395 3345 9421
rect 3371 9395 3397 9421
rect 5927 9395 5953 9421
rect 5979 9395 6005 9421
rect 6031 9395 6057 9421
rect 8587 9395 8613 9421
rect 8639 9395 8665 9421
rect 8691 9395 8717 9421
rect 11247 9395 11273 9421
rect 11299 9395 11325 9421
rect 11351 9395 11377 9421
rect 2423 9311 2449 9337
rect 5503 9311 5529 9337
rect 8023 9311 8049 9337
rect 9143 9311 9169 9337
rect 10543 9311 10569 9337
rect 1639 9255 1665 9281
rect 2871 9255 2897 9281
rect 2927 9255 2953 9281
rect 4327 9255 4353 9281
rect 4775 9255 4801 9281
rect 6343 9255 6369 9281
rect 6679 9255 6705 9281
rect 7407 9255 7433 9281
rect 7855 9255 7881 9281
rect 9759 9255 9785 9281
rect 1527 9199 1553 9225
rect 1807 9199 1833 9225
rect 2031 9199 2057 9225
rect 2087 9199 2113 9225
rect 2143 9199 2169 9225
rect 2367 9199 2393 9225
rect 2759 9199 2785 9225
rect 4943 9199 4969 9225
rect 5559 9199 5585 9225
rect 5783 9199 5809 9225
rect 5951 9199 5977 9225
rect 6175 9199 6201 9225
rect 6287 9199 6313 9225
rect 6511 9199 6537 9225
rect 9255 9199 9281 9225
rect 10319 9199 10345 9225
rect 10487 9199 10513 9225
rect 10599 9199 10625 9225
rect 2479 9143 2505 9169
rect 3151 9143 3177 9169
rect 4103 9143 4129 9169
rect 10039 9143 10065 9169
rect 2591 9087 2617 9113
rect 3095 9087 3121 9113
rect 4159 9087 4185 9113
rect 4271 9087 4297 9113
rect 5447 9087 5473 9113
rect 5671 9087 5697 9113
rect 6063 9087 6089 9113
rect 7071 9087 7097 9113
rect 7127 9087 7153 9113
rect 7239 9087 7265 9113
rect 7351 9087 7377 9113
rect 9087 9087 9113 9113
rect 9703 9087 9729 9113
rect 9871 9087 9897 9113
rect 10095 9087 10121 9113
rect 10207 9087 10233 9113
rect 10711 9087 10737 9113
rect 1937 9003 1963 9029
rect 1989 9003 2015 9029
rect 2041 9003 2067 9029
rect 4597 9003 4623 9029
rect 4649 9003 4675 9029
rect 4701 9003 4727 9029
rect 7257 9003 7283 9029
rect 7309 9003 7335 9029
rect 7361 9003 7387 9029
rect 9917 9003 9943 9029
rect 9969 9003 9995 9029
rect 10021 9003 10047 9029
rect 2311 8919 2337 8945
rect 2479 8919 2505 8945
rect 4271 8919 4297 8945
rect 5447 8919 5473 8945
rect 5671 8919 5697 8945
rect 6063 8919 6089 8945
rect 7687 8919 7713 8945
rect 10263 8919 10289 8945
rect 1919 8863 1945 8889
rect 5503 8863 5529 8889
rect 5951 8863 5977 8889
rect 10151 8863 10177 8889
rect 1975 8807 2001 8833
rect 2311 8807 2337 8833
rect 3991 8807 4017 8833
rect 4047 8807 4073 8833
rect 4159 8807 4185 8833
rect 5615 8807 5641 8833
rect 6175 8807 6201 8833
rect 7519 8807 7545 8833
rect 10095 8807 10121 8833
rect 2087 8751 2113 8777
rect 1863 8695 1889 8721
rect 3991 8695 4017 8721
rect 6119 8695 6145 8721
rect 7631 8695 7657 8721
rect 3267 8611 3293 8637
rect 3319 8611 3345 8637
rect 3371 8611 3397 8637
rect 5927 8611 5953 8637
rect 5979 8611 6005 8637
rect 6031 8611 6057 8637
rect 8587 8611 8613 8637
rect 8639 8611 8665 8637
rect 8691 8611 8717 8637
rect 11247 8611 11273 8637
rect 11299 8611 11325 8637
rect 11351 8611 11377 8637
rect 2647 8527 2673 8553
rect 2983 8527 3009 8553
rect 4103 8527 4129 8553
rect 6175 8527 6201 8553
rect 2815 8471 2841 8497
rect 6007 8471 6033 8497
rect 10935 8471 10961 8497
rect 2535 8415 2561 8441
rect 3207 8415 3233 8441
rect 4215 8415 4241 8441
rect 10039 8415 10065 8441
rect 10823 8415 10849 8441
rect 11103 8415 11129 8441
rect 9871 8303 9897 8329
rect 10039 8303 10065 8329
rect 1937 8219 1963 8245
rect 1989 8219 2015 8245
rect 2041 8219 2067 8245
rect 4597 8219 4623 8245
rect 4649 8219 4675 8245
rect 4701 8219 4727 8245
rect 7257 8219 7283 8245
rect 7309 8219 7335 8245
rect 7361 8219 7387 8245
rect 9917 8219 9943 8245
rect 9969 8219 9995 8245
rect 10021 8219 10047 8245
rect 6791 8135 6817 8161
rect 9087 8135 9113 8161
rect 9535 8079 9561 8105
rect 9983 8079 10009 8105
rect 6903 8023 6929 8049
rect 7015 8023 7041 8049
rect 9031 8023 9057 8049
rect 9199 8023 9225 8049
rect 9591 8023 9617 8049
rect 9759 8023 9785 8049
rect 9871 8023 9897 8049
rect 10207 8023 10233 8049
rect 1695 7967 1721 7993
rect 1751 7967 1777 7993
rect 1919 7967 1945 7993
rect 8863 7967 8889 7993
rect 9423 7967 9449 7993
rect 10319 7967 10345 7993
rect 1639 7911 1665 7937
rect 1975 7911 2001 7937
rect 2031 7911 2057 7937
rect 4551 7911 4577 7937
rect 4719 7911 4745 7937
rect 6959 7911 6985 7937
rect 9255 7911 9281 7937
rect 9815 7911 9841 7937
rect 10263 7911 10289 7937
rect 3267 7827 3293 7853
rect 3319 7827 3345 7853
rect 3371 7827 3397 7853
rect 5927 7827 5953 7853
rect 5979 7827 6005 7853
rect 6031 7827 6057 7853
rect 8587 7827 8613 7853
rect 8639 7827 8665 7853
rect 8691 7827 8717 7853
rect 11247 7827 11273 7853
rect 11299 7827 11325 7853
rect 11351 7827 11377 7853
rect 3991 7743 4017 7769
rect 7407 7743 7433 7769
rect 10375 7743 10401 7769
rect 1135 7687 1161 7713
rect 1247 7687 1273 7713
rect 1695 7687 1721 7713
rect 2143 7687 2169 7713
rect 6063 7687 6089 7713
rect 7239 7687 7265 7713
rect 9871 7687 9897 7713
rect 10319 7687 10345 7713
rect 10431 7687 10457 7713
rect 1527 7631 1553 7657
rect 1863 7631 1889 7657
rect 1975 7631 2001 7657
rect 4831 7631 4857 7657
rect 6231 7631 6257 7657
rect 10039 7631 10065 7657
rect 10095 7631 10121 7657
rect 1191 7575 1217 7601
rect 1471 7575 1497 7601
rect 1639 7575 1665 7601
rect 2087 7575 2113 7601
rect 2367 7575 2393 7601
rect 4271 7575 4297 7601
rect 4775 7575 4801 7601
rect 4943 7575 4969 7601
rect 4999 7575 5025 7601
rect 9703 7575 9729 7601
rect 9927 7575 9953 7601
rect 4159 7519 4185 7545
rect 1937 7435 1963 7461
rect 1989 7435 2015 7461
rect 2041 7435 2067 7461
rect 4597 7435 4623 7461
rect 4649 7435 4675 7461
rect 4701 7435 4727 7461
rect 7257 7435 7283 7461
rect 7309 7435 7335 7461
rect 7361 7435 7387 7461
rect 9917 7435 9943 7461
rect 9969 7435 9995 7461
rect 10021 7435 10047 7461
rect 1751 7351 1777 7377
rect 2199 7351 2225 7377
rect 3823 7351 3849 7377
rect 3935 7351 3961 7377
rect 4271 7351 4297 7377
rect 4383 7351 4409 7377
rect 5783 7351 5809 7377
rect 7575 7351 7601 7377
rect 1863 7295 1889 7321
rect 7799 7295 7825 7321
rect 9815 7295 9841 7321
rect 9983 7295 10009 7321
rect 1919 7239 1945 7265
rect 4047 7239 4073 7265
rect 4495 7239 4521 7265
rect 5391 7239 5417 7265
rect 5671 7239 5697 7265
rect 5895 7239 5921 7265
rect 6343 7239 6369 7265
rect 6903 7239 6929 7265
rect 7015 7239 7041 7265
rect 7183 7239 7209 7265
rect 7351 7239 7377 7265
rect 7463 7239 7489 7265
rect 10151 7239 10177 7265
rect 2255 7183 2281 7209
rect 3767 7183 3793 7209
rect 4215 7183 4241 7209
rect 5503 7183 5529 7209
rect 6791 7183 6817 7209
rect 7631 7183 7657 7209
rect 7855 7183 7881 7209
rect 7967 7183 7993 7209
rect 9647 7183 9673 7209
rect 2199 7127 2225 7153
rect 6119 7127 6145 7153
rect 6231 7127 6257 7153
rect 7183 7127 7209 7153
rect 9759 7127 9785 7153
rect 10039 7127 10065 7153
rect 3267 7043 3293 7069
rect 3319 7043 3345 7069
rect 3371 7043 3397 7069
rect 5927 7043 5953 7069
rect 5979 7043 6005 7069
rect 6031 7043 6057 7069
rect 8587 7043 8613 7069
rect 8639 7043 8665 7069
rect 8691 7043 8717 7069
rect 11247 7043 11273 7069
rect 11299 7043 11325 7069
rect 11351 7043 11377 7069
rect 7127 6959 7153 6985
rect 7295 6959 7321 6985
rect 7967 6959 7993 6985
rect 9591 6959 9617 6985
rect 7519 6903 7545 6929
rect 7855 6903 7881 6929
rect 9143 6903 9169 6929
rect 9983 6903 10009 6929
rect 10263 6903 10289 6929
rect 10935 6903 10961 6929
rect 1919 6847 1945 6873
rect 4999 6847 5025 6873
rect 5111 6847 5137 6873
rect 5223 6847 5249 6873
rect 5503 6847 5529 6873
rect 5615 6847 5641 6873
rect 5727 6847 5753 6873
rect 5839 6847 5865 6873
rect 7799 6847 7825 6873
rect 9199 6847 9225 6873
rect 9311 6847 9337 6873
rect 9423 6847 9449 6873
rect 9591 6847 9617 6873
rect 9759 6847 9785 6873
rect 9815 6847 9841 6873
rect 11103 6847 11129 6873
rect 4943 6791 4969 6817
rect 7463 6791 7489 6817
rect 10207 6791 10233 6817
rect 10823 6791 10849 6817
rect 1639 6735 1665 6761
rect 1807 6735 1833 6761
rect 5279 6735 5305 6761
rect 5447 6735 5473 6761
rect 7631 6735 7657 6761
rect 10151 6735 10177 6761
rect 1937 6651 1963 6677
rect 1989 6651 2015 6677
rect 2041 6651 2067 6677
rect 4597 6651 4623 6677
rect 4649 6651 4675 6677
rect 4701 6651 4727 6677
rect 7257 6651 7283 6677
rect 7309 6651 7335 6677
rect 7361 6651 7387 6677
rect 9917 6651 9943 6677
rect 9969 6651 9995 6677
rect 10021 6651 10047 6677
rect 9591 6567 9617 6593
rect 9647 6567 9673 6593
rect 2815 6511 2841 6537
rect 4383 6511 4409 6537
rect 10151 6511 10177 6537
rect 1751 6455 1777 6481
rect 4215 6455 4241 6481
rect 7295 6455 7321 6481
rect 9759 6455 9785 6481
rect 9815 6455 9841 6481
rect 10039 6455 10065 6481
rect 10207 6455 10233 6481
rect 4103 6399 4129 6425
rect 1919 6343 1945 6369
rect 2871 6343 2897 6369
rect 4327 6343 4353 6369
rect 4383 6343 4409 6369
rect 7183 6343 7209 6369
rect 3267 6259 3293 6285
rect 3319 6259 3345 6285
rect 3371 6259 3397 6285
rect 5927 6259 5953 6285
rect 5979 6259 6005 6285
rect 6031 6259 6057 6285
rect 8587 6259 8613 6285
rect 8639 6259 8665 6285
rect 8691 6259 8717 6285
rect 11247 6259 11273 6285
rect 11299 6259 11325 6285
rect 11351 6259 11377 6285
rect 3319 6175 3345 6201
rect 4775 6175 4801 6201
rect 4831 6175 4857 6201
rect 9759 6175 9785 6201
rect 2703 6119 2729 6145
rect 3935 6119 3961 6145
rect 1975 6063 2001 6089
rect 2759 6063 2785 6089
rect 2983 6063 3009 6089
rect 3207 6063 3233 6089
rect 3823 6063 3849 6089
rect 4887 6063 4913 6089
rect 5055 6063 5081 6089
rect 9591 6063 9617 6089
rect 9815 6063 9841 6089
rect 9983 6063 10009 6089
rect 1639 6007 1665 6033
rect 2031 6007 2057 6033
rect 3263 6007 3289 6033
rect 9759 5951 9785 5977
rect 1937 5867 1963 5893
rect 1989 5867 2015 5893
rect 2041 5867 2067 5893
rect 4597 5867 4623 5893
rect 4649 5867 4675 5893
rect 4701 5867 4727 5893
rect 7257 5867 7283 5893
rect 7309 5867 7335 5893
rect 7361 5867 7387 5893
rect 9917 5867 9943 5893
rect 9969 5867 9995 5893
rect 10021 5867 10047 5893
rect 4383 5783 4409 5809
rect 2311 5727 2337 5753
rect 7519 5727 7545 5753
rect 2367 5671 2393 5697
rect 4887 5671 4913 5697
rect 5111 5671 5137 5697
rect 5223 5671 5249 5697
rect 9983 5671 10009 5697
rect 4439 5615 4465 5641
rect 4551 5615 4577 5641
rect 7183 5615 7209 5641
rect 7575 5615 7601 5641
rect 7687 5615 7713 5641
rect 5167 5559 5193 5585
rect 7351 5559 7377 5585
rect 10151 5559 10177 5585
rect 3267 5475 3293 5501
rect 3319 5475 3345 5501
rect 3371 5475 3397 5501
rect 5927 5475 5953 5501
rect 5979 5475 6005 5501
rect 6031 5475 6057 5501
rect 8587 5475 8613 5501
rect 8639 5475 8665 5501
rect 8691 5475 8717 5501
rect 11247 5475 11273 5501
rect 11299 5475 11325 5501
rect 11351 5475 11377 5501
rect 1135 5391 1161 5417
rect 7127 5391 7153 5417
rect 7239 5391 7265 5417
rect 7967 5391 7993 5417
rect 9647 5391 9673 5417
rect 10207 5391 10233 5417
rect 10935 5391 10961 5417
rect 1303 5335 1329 5361
rect 6455 5335 6481 5361
rect 9199 5335 9225 5361
rect 10039 5335 10065 5361
rect 1639 5279 1665 5305
rect 6567 5279 6593 5305
rect 6735 5279 6761 5305
rect 7295 5279 7321 5305
rect 7463 5279 7489 5305
rect 7911 5279 7937 5305
rect 9479 5279 9505 5305
rect 9647 5279 9673 5305
rect 9871 5279 9897 5305
rect 10319 5279 10345 5305
rect 11103 5279 11129 5305
rect 1583 5223 1609 5249
rect 1975 5223 2001 5249
rect 7183 5223 7209 5249
rect 9367 5223 9393 5249
rect 10823 5223 10849 5249
rect 6511 5167 6537 5193
rect 6847 5167 6873 5193
rect 7575 5167 7601 5193
rect 7799 5167 7825 5193
rect 7967 5167 7993 5193
rect 9255 5167 9281 5193
rect 9759 5167 9785 5193
rect 1937 5083 1963 5109
rect 1989 5083 2015 5109
rect 2041 5083 2067 5109
rect 4597 5083 4623 5109
rect 4649 5083 4675 5109
rect 4701 5083 4727 5109
rect 7257 5083 7283 5109
rect 7309 5083 7335 5109
rect 7361 5083 7387 5109
rect 9917 5083 9943 5109
rect 9969 5083 9995 5109
rect 10021 5083 10047 5109
rect 2031 4999 2057 5025
rect 4999 4999 5025 5025
rect 9759 4999 9785 5025
rect 4271 4943 4297 4969
rect 4495 4943 4521 4969
rect 4607 4943 4633 4969
rect 7015 4943 7041 4969
rect 7575 4943 7601 4969
rect 9703 4943 9729 4969
rect 9927 4943 9953 4969
rect 2143 4887 2169 4913
rect 4943 4887 4969 4913
rect 5447 4887 5473 4913
rect 7687 4887 7713 4913
rect 9367 4887 9393 4913
rect 9983 4887 10009 4913
rect 10095 4887 10121 4913
rect 4215 4831 4241 4857
rect 4327 4831 4353 4857
rect 5167 4831 5193 4857
rect 5279 4831 5305 4857
rect 6959 4831 6985 4857
rect 7351 4831 7377 4857
rect 7463 4831 7489 4857
rect 9255 4831 9281 4857
rect 9647 4831 9673 4857
rect 1863 4775 1889 4801
rect 4775 4775 4801 4801
rect 5335 4775 5361 4801
rect 3267 4691 3293 4717
rect 3319 4691 3345 4717
rect 3371 4691 3397 4717
rect 5927 4691 5953 4717
rect 5979 4691 6005 4717
rect 6031 4691 6057 4717
rect 8587 4691 8613 4717
rect 8639 4691 8665 4717
rect 8691 4691 8717 4717
rect 11247 4691 11273 4717
rect 11299 4691 11325 4717
rect 11351 4691 11377 4717
rect 5391 4607 5417 4633
rect 7407 4607 7433 4633
rect 9927 4607 9953 4633
rect 5447 4551 5473 4577
rect 7351 4551 7377 4577
rect 9759 4551 9785 4577
rect 1807 4495 1833 4521
rect 1919 4495 1945 4521
rect 2087 4495 2113 4521
rect 2255 4495 2281 4521
rect 2479 4495 2505 4521
rect 4999 4495 5025 4521
rect 5167 4495 5193 4521
rect 9647 4495 9673 4521
rect 10039 4495 10065 4521
rect 1975 4439 2001 4465
rect 2703 4439 2729 4465
rect 5111 4439 5137 4465
rect 5391 4383 5417 4409
rect 1937 4299 1963 4325
rect 1989 4299 2015 4325
rect 2041 4299 2067 4325
rect 4597 4299 4623 4325
rect 4649 4299 4675 4325
rect 4701 4299 4727 4325
rect 7257 4299 7283 4325
rect 7309 4299 7335 4325
rect 7361 4299 7387 4325
rect 9917 4299 9943 4325
rect 9969 4299 9995 4325
rect 10021 4299 10047 4325
rect 9759 4215 9785 4241
rect 2871 4159 2897 4185
rect 4439 4159 4465 4185
rect 4551 4159 4577 4185
rect 4663 4159 4689 4185
rect 5671 4159 5697 4185
rect 7575 4159 7601 4185
rect 1583 4103 1609 4129
rect 1919 4103 1945 4129
rect 2087 4103 2113 4129
rect 2479 4103 2505 4129
rect 2983 4103 3009 4129
rect 3655 4103 3681 4129
rect 3823 4103 3849 4129
rect 4999 4103 5025 4129
rect 5391 4103 5417 4129
rect 7407 4103 7433 4129
rect 7687 4103 7713 4129
rect 9927 4103 9953 4129
rect 10207 4103 10233 4129
rect 1695 4047 1721 4073
rect 2367 4047 2393 4073
rect 3151 4047 3177 4073
rect 3263 4047 3289 4073
rect 3711 4047 3737 4073
rect 5055 4047 5081 4073
rect 5223 4047 5249 4073
rect 5615 4047 5641 4073
rect 5727 4047 5753 4073
rect 7463 4047 7489 4073
rect 9535 4047 9561 4073
rect 9815 4047 9841 4073
rect 10095 4047 10121 4073
rect 10375 4047 10401 4073
rect 10935 4047 10961 4073
rect 11103 4047 11129 4073
rect 2815 3991 2841 4017
rect 4887 3991 4913 4017
rect 5503 3991 5529 4017
rect 7911 3991 7937 4017
rect 9367 3991 9393 4017
rect 10039 3991 10065 4017
rect 10319 3991 10345 4017
rect 10767 3991 10793 4017
rect 3267 3907 3293 3933
rect 3319 3907 3345 3933
rect 3371 3907 3397 3933
rect 5927 3907 5953 3933
rect 5979 3907 6005 3933
rect 6031 3907 6057 3933
rect 8587 3907 8613 3933
rect 8639 3907 8665 3933
rect 8691 3907 8717 3933
rect 11247 3907 11273 3933
rect 11299 3907 11325 3933
rect 11351 3907 11377 3933
rect 2535 3823 2561 3849
rect 4943 3823 4969 3849
rect 5055 3823 5081 3849
rect 7183 3823 7209 3849
rect 2423 3767 2449 3793
rect 5111 3767 5137 3793
rect 5223 3767 5249 3793
rect 5559 3767 5585 3793
rect 7015 3767 7041 3793
rect 7071 3767 7097 3793
rect 7407 3767 7433 3793
rect 7463 3767 7489 3793
rect 9983 3767 10009 3793
rect 2367 3711 2393 3737
rect 2647 3711 2673 3737
rect 7295 3711 7321 3737
rect 7687 3711 7713 3737
rect 10151 3711 10177 3737
rect 11103 3711 11129 3737
rect 2871 3655 2897 3681
rect 5335 3655 5361 3681
rect 7463 3655 7489 3681
rect 1937 3515 1963 3541
rect 1989 3515 2015 3541
rect 2041 3515 2067 3541
rect 4597 3515 4623 3541
rect 4649 3515 4675 3541
rect 4701 3515 4727 3541
rect 7257 3515 7283 3541
rect 7309 3515 7335 3541
rect 7361 3515 7387 3541
rect 9917 3515 9943 3541
rect 9969 3515 9995 3541
rect 10021 3515 10047 3541
rect 7351 3431 7377 3457
rect 7407 3375 7433 3401
rect 7631 3375 7657 3401
rect 3267 3123 3293 3149
rect 3319 3123 3345 3149
rect 3371 3123 3397 3149
rect 5927 3123 5953 3149
rect 5979 3123 6005 3149
rect 6031 3123 6057 3149
rect 8587 3123 8613 3149
rect 8639 3123 8665 3149
rect 8691 3123 8717 3149
rect 11247 3123 11273 3149
rect 11299 3123 11325 3149
rect 11351 3123 11377 3149
rect 1937 2731 1963 2757
rect 1989 2731 2015 2757
rect 2041 2731 2067 2757
rect 4597 2731 4623 2757
rect 4649 2731 4675 2757
rect 4701 2731 4727 2757
rect 7257 2731 7283 2757
rect 7309 2731 7335 2757
rect 7361 2731 7387 2757
rect 9917 2731 9943 2757
rect 9969 2731 9995 2757
rect 10021 2731 10047 2757
rect 10823 2535 10849 2561
rect 11103 2535 11129 2561
rect 10935 2479 10961 2505
rect 3267 2339 3293 2365
rect 3319 2339 3345 2365
rect 3371 2339 3397 2365
rect 5927 2339 5953 2365
rect 5979 2339 6005 2365
rect 6031 2339 6057 2365
rect 8587 2339 8613 2365
rect 8639 2339 8665 2365
rect 8691 2339 8717 2365
rect 11247 2339 11273 2365
rect 11299 2339 11325 2365
rect 11351 2339 11377 2365
rect 1937 1947 1963 1973
rect 1989 1947 2015 1973
rect 2041 1947 2067 1973
rect 4597 1947 4623 1973
rect 4649 1947 4675 1973
rect 4701 1947 4727 1973
rect 7257 1947 7283 1973
rect 7309 1947 7335 1973
rect 7361 1947 7387 1973
rect 9917 1947 9943 1973
rect 9969 1947 9995 1973
rect 10021 1947 10047 1973
rect 3267 1555 3293 1581
rect 3319 1555 3345 1581
rect 3371 1555 3397 1581
rect 5927 1555 5953 1581
rect 5979 1555 6005 1581
rect 6031 1555 6057 1581
rect 8587 1555 8613 1581
rect 8639 1555 8665 1581
rect 8691 1555 8717 1581
rect 11247 1555 11273 1581
rect 11299 1555 11325 1581
rect 11351 1555 11377 1581
<< metal2 >>
rect 896 11600 952 12000
rect 2016 11600 2072 12000
rect 3136 11600 3192 12000
rect 4256 11600 4312 12000
rect 4438 11606 4690 11634
rect 910 10094 938 11600
rect 2030 10094 2058 11600
rect 3150 10094 3178 11600
rect 4270 11522 4298 11600
rect 4438 11522 4466 11606
rect 4270 11494 4466 11522
rect 3266 10206 3398 10211
rect 3294 10178 3318 10206
rect 3346 10178 3370 10206
rect 3266 10173 3398 10178
rect 910 10066 1050 10094
rect 2030 10066 2170 10094
rect 3150 10066 3290 10094
rect 1022 10065 1050 10066
rect 1022 10039 1023 10065
rect 1049 10039 1050 10065
rect 1022 10033 1050 10039
rect 2142 10065 2170 10066
rect 2142 10039 2143 10065
rect 2169 10039 2170 10065
rect 2142 10033 2170 10039
rect 3262 10065 3290 10066
rect 3262 10039 3263 10065
rect 3289 10039 3290 10065
rect 3262 10033 3290 10039
rect 4662 10065 4690 11606
rect 5376 11600 5432 12000
rect 6496 11600 6552 12000
rect 7616 11600 7672 12000
rect 8736 11600 8792 12000
rect 9856 11600 9912 12000
rect 10976 11600 11032 12000
rect 5390 10094 5418 11600
rect 5926 10206 6058 10211
rect 5954 10178 5978 10206
rect 6006 10178 6030 10206
rect 5926 10173 6058 10178
rect 6510 10094 6538 11600
rect 5390 10066 5530 10094
rect 6510 10066 6650 10094
rect 4662 10039 4663 10065
rect 4689 10039 4690 10065
rect 4662 10033 4690 10039
rect 5502 10065 5530 10066
rect 5502 10039 5503 10065
rect 5529 10039 5530 10065
rect 5502 10033 5530 10039
rect 6622 10065 6650 10066
rect 6622 10039 6623 10065
rect 6649 10039 6650 10065
rect 6622 10033 6650 10039
rect 7630 10066 7658 11600
rect 8586 10206 8718 10211
rect 8614 10178 8638 10206
rect 8666 10178 8690 10206
rect 8586 10173 8718 10178
rect 7742 10066 7770 10071
rect 7630 10065 7770 10066
rect 7630 10039 7743 10065
rect 7769 10039 7770 10065
rect 7630 10038 7770 10039
rect 8750 10066 8778 11600
rect 8862 10066 8890 10071
rect 8750 10065 8890 10066
rect 8750 10039 8863 10065
rect 8889 10039 8890 10065
rect 8750 10038 8890 10039
rect 7742 10033 7770 10038
rect 8862 10033 8890 10038
rect 9870 10066 9898 11600
rect 10038 11018 10066 11023
rect 10038 10066 10066 10990
rect 10094 10066 10122 10071
rect 10038 10065 10122 10066
rect 10038 10039 10095 10065
rect 10121 10039 10122 10065
rect 10038 10038 10122 10039
rect 9870 10033 9898 10038
rect 10094 10033 10122 10038
rect 10374 10066 10402 10071
rect 10990 10066 11018 11600
rect 11246 10206 11378 10211
rect 11274 10178 11298 10206
rect 11326 10178 11350 10206
rect 11246 10173 11378 10178
rect 11102 10066 11130 10071
rect 10990 10065 11130 10066
rect 10990 10039 11103 10065
rect 11129 10039 11130 10065
rect 10990 10038 11130 10039
rect 10374 10019 10402 10038
rect 11102 10033 11130 10038
rect 1134 10010 1162 10015
rect 1078 10009 1162 10010
rect 1078 9983 1135 10009
rect 1161 9983 1162 10009
rect 1078 9982 1162 9983
rect 1078 5418 1106 9982
rect 1134 9977 1162 9982
rect 2310 10010 2338 10015
rect 2310 10009 2506 10010
rect 2310 9983 2311 10009
rect 2337 9983 2506 10009
rect 2310 9982 2506 9983
rect 2310 9977 2338 9982
rect 1936 9814 2068 9819
rect 1964 9786 1988 9814
rect 2016 9786 2040 9814
rect 1936 9781 2068 9786
rect 2478 9729 2506 9982
rect 2478 9703 2479 9729
rect 2505 9703 2506 9729
rect 2478 9697 2506 9703
rect 3430 10009 3458 10015
rect 3430 9983 3431 10009
rect 3457 9983 3458 10009
rect 2310 9674 2338 9679
rect 2310 9673 2394 9674
rect 2310 9647 2311 9673
rect 2337 9647 2394 9673
rect 2310 9646 2394 9647
rect 2310 9641 2338 9646
rect 2142 9562 2170 9567
rect 2142 9561 2226 9562
rect 2142 9535 2143 9561
rect 2169 9535 2226 9561
rect 2142 9534 2226 9535
rect 2142 9529 2170 9534
rect 1638 9281 1666 9287
rect 1638 9255 1639 9281
rect 1665 9255 1666 9281
rect 1526 9226 1554 9231
rect 1526 9179 1554 9198
rect 1638 9170 1666 9255
rect 2086 9282 2114 9287
rect 1806 9226 1834 9231
rect 2030 9226 2058 9231
rect 1806 9179 1834 9198
rect 1862 9225 2058 9226
rect 1862 9199 2031 9225
rect 2057 9199 2058 9225
rect 1862 9198 2058 9199
rect 1638 9137 1666 9142
rect 1862 8890 1890 9198
rect 2030 9193 2058 9198
rect 2086 9225 2114 9254
rect 2086 9199 2087 9225
rect 2113 9199 2114 9225
rect 2086 9193 2114 9199
rect 2142 9226 2170 9231
rect 2142 9179 2170 9198
rect 2198 9114 2226 9534
rect 2254 9506 2282 9511
rect 2254 9505 2338 9506
rect 2254 9479 2255 9505
rect 2281 9479 2338 9505
rect 2254 9478 2338 9479
rect 2254 9473 2282 9478
rect 2310 9338 2338 9478
rect 2310 9305 2338 9310
rect 2366 9225 2394 9646
rect 2534 9562 2562 9567
rect 2534 9515 2562 9534
rect 3266 9422 3398 9427
rect 3294 9394 3318 9422
rect 3346 9394 3370 9422
rect 3266 9389 3398 9394
rect 2422 9338 2450 9343
rect 2422 9291 2450 9310
rect 2870 9281 2898 9287
rect 2870 9255 2871 9281
rect 2897 9255 2898 9281
rect 2758 9226 2786 9231
rect 2366 9199 2367 9225
rect 2393 9199 2394 9225
rect 2366 9193 2394 9199
rect 2534 9225 2786 9226
rect 2534 9199 2759 9225
rect 2785 9199 2786 9225
rect 2534 9198 2786 9199
rect 2478 9170 2506 9175
rect 2478 9123 2506 9142
rect 2198 9086 2282 9114
rect 1936 9030 2068 9035
rect 1964 9002 1988 9030
rect 2016 9002 2040 9030
rect 1936 8997 2068 9002
rect 2254 8946 2282 9086
rect 2310 8946 2338 8951
rect 1974 8945 2338 8946
rect 1974 8919 2311 8945
rect 2337 8919 2338 8945
rect 1974 8918 2338 8919
rect 1918 8890 1946 8895
rect 1862 8889 1946 8890
rect 1862 8863 1919 8889
rect 1945 8863 1946 8889
rect 1862 8862 1946 8863
rect 1862 8721 1890 8727
rect 1862 8695 1863 8721
rect 1889 8695 1890 8721
rect 1526 7994 1554 7999
rect 1246 7938 1274 7943
rect 1134 7713 1162 7719
rect 1134 7687 1135 7713
rect 1161 7687 1162 7713
rect 1134 7378 1162 7687
rect 1246 7713 1274 7910
rect 1246 7687 1247 7713
rect 1273 7687 1274 7713
rect 1246 7681 1274 7687
rect 1526 7657 1554 7966
rect 1694 7994 1722 7999
rect 1694 7947 1722 7966
rect 1750 7994 1778 7999
rect 1862 7994 1890 8695
rect 1918 8666 1946 8862
rect 1974 8833 2002 8918
rect 2310 8913 2338 8918
rect 2478 8946 2506 8951
rect 2534 8946 2562 9198
rect 2758 9193 2786 9198
rect 2870 9226 2898 9255
rect 2926 9282 2954 9287
rect 2926 9235 2954 9254
rect 2870 9193 2898 9198
rect 3150 9170 3178 9175
rect 3150 9123 3178 9142
rect 2590 9114 2618 9119
rect 2590 9113 2674 9114
rect 2590 9087 2591 9113
rect 2617 9087 2674 9113
rect 2590 9086 2674 9087
rect 2590 9081 2618 9086
rect 2478 8945 2562 8946
rect 2478 8919 2479 8945
rect 2505 8919 2562 8945
rect 2478 8918 2562 8919
rect 2478 8913 2506 8918
rect 2646 8890 2674 9086
rect 1974 8807 1975 8833
rect 2001 8807 2002 8833
rect 1974 8801 2002 8807
rect 2310 8833 2338 8839
rect 2310 8807 2311 8833
rect 2337 8807 2338 8833
rect 2086 8778 2114 8783
rect 2086 8731 2114 8750
rect 2310 8666 2338 8807
rect 1918 8638 2338 8666
rect 2646 8553 2674 8862
rect 3094 9113 3122 9119
rect 3094 9087 3095 9113
rect 3121 9087 3122 9113
rect 3094 8778 3122 9087
rect 3094 8745 3122 8750
rect 2646 8527 2647 8553
rect 2673 8527 2674 8553
rect 2646 8521 2674 8527
rect 2982 8722 3010 8727
rect 2982 8553 3010 8694
rect 3266 8638 3398 8643
rect 3294 8610 3318 8638
rect 3346 8610 3370 8638
rect 3266 8605 3398 8610
rect 2982 8527 2983 8553
rect 3009 8527 3010 8553
rect 2982 8521 3010 8527
rect 2814 8497 2842 8503
rect 2814 8471 2815 8497
rect 2841 8471 2842 8497
rect 2534 8441 2562 8447
rect 2534 8415 2535 8441
rect 2561 8415 2562 8441
rect 2534 8386 2562 8415
rect 1936 8246 2068 8251
rect 1964 8218 1988 8246
rect 2016 8218 2040 8246
rect 1936 8213 2068 8218
rect 1750 7993 1890 7994
rect 1750 7967 1751 7993
rect 1777 7967 1890 7993
rect 1750 7966 1890 7967
rect 1918 7994 1946 7999
rect 1750 7961 1778 7966
rect 1638 7937 1666 7943
rect 1638 7911 1639 7937
rect 1665 7911 1666 7937
rect 1638 7714 1666 7911
rect 1694 7714 1722 7719
rect 1638 7713 1778 7714
rect 1638 7687 1695 7713
rect 1721 7687 1778 7713
rect 1638 7686 1778 7687
rect 1694 7681 1722 7686
rect 1526 7631 1527 7657
rect 1553 7631 1554 7657
rect 1526 7625 1554 7631
rect 1190 7602 1218 7607
rect 1190 7555 1218 7574
rect 1470 7601 1498 7607
rect 1470 7575 1471 7601
rect 1497 7575 1498 7601
rect 1134 7345 1162 7350
rect 1470 7378 1498 7575
rect 1638 7602 1666 7607
rect 1638 7555 1666 7574
rect 1470 7345 1498 7350
rect 1750 7377 1778 7686
rect 1750 7351 1751 7377
rect 1777 7351 1778 7377
rect 1750 7345 1778 7351
rect 1638 6761 1666 6767
rect 1638 6735 1639 6761
rect 1665 6735 1666 6761
rect 1638 6538 1666 6735
rect 1806 6762 1834 7966
rect 1918 7947 1946 7966
rect 1974 7938 2002 7943
rect 1974 7891 2002 7910
rect 2030 7937 2058 7943
rect 2030 7911 2031 7937
rect 2057 7911 2058 7937
rect 1862 7657 1890 7663
rect 1862 7631 1863 7657
rect 1889 7631 1890 7657
rect 1862 7321 1890 7631
rect 1974 7658 2002 7663
rect 2030 7658 2058 7911
rect 1974 7657 2058 7658
rect 1974 7631 1975 7657
rect 2001 7631 2058 7657
rect 1974 7630 2058 7631
rect 2142 7770 2170 7775
rect 2142 7713 2170 7742
rect 2142 7687 2143 7713
rect 2169 7687 2170 7713
rect 1974 7602 2002 7630
rect 1974 7569 2002 7574
rect 2086 7602 2114 7607
rect 2086 7555 2114 7574
rect 1936 7462 2068 7467
rect 1964 7434 1988 7462
rect 2016 7434 2040 7462
rect 1936 7429 2068 7434
rect 2142 7322 2170 7687
rect 2310 7602 2338 7607
rect 2366 7602 2394 7607
rect 2338 7601 2394 7602
rect 2338 7575 2367 7601
rect 2393 7575 2394 7601
rect 2338 7574 2394 7575
rect 2198 7378 2226 7383
rect 2198 7331 2226 7350
rect 1862 7295 1863 7321
rect 1889 7295 1890 7321
rect 1862 7289 1890 7295
rect 1918 7294 2170 7322
rect 1918 7265 1946 7294
rect 1918 7239 1919 7265
rect 1945 7239 1946 7265
rect 1918 6873 1946 7239
rect 2254 7210 2282 7215
rect 2254 7163 2282 7182
rect 1918 6847 1919 6873
rect 1945 6847 1946 6873
rect 1918 6841 1946 6847
rect 2198 7154 2226 7159
rect 1806 6715 1834 6734
rect 1936 6678 2068 6683
rect 1964 6650 1988 6678
rect 2016 6650 2040 6678
rect 1936 6645 2068 6650
rect 1638 6510 1778 6538
rect 1750 6481 1778 6510
rect 1750 6455 1751 6481
rect 1777 6455 1778 6481
rect 1750 6449 1778 6455
rect 1918 6369 1946 6375
rect 1918 6343 1919 6369
rect 1945 6343 1946 6369
rect 1918 6146 1946 6343
rect 2198 6202 2226 7126
rect 2198 6169 2226 6174
rect 2310 6146 2338 7574
rect 2366 7569 2394 7574
rect 2478 7602 2506 7607
rect 2534 7602 2562 8358
rect 2506 7574 2562 7602
rect 2814 7574 2842 8471
rect 3206 8441 3234 8447
rect 3206 8415 3207 8441
rect 3233 8415 3234 8441
rect 3206 8386 3234 8415
rect 3206 8353 3234 8358
rect 3266 7854 3398 7859
rect 3294 7826 3318 7854
rect 3346 7826 3370 7854
rect 3266 7821 3398 7826
rect 2478 7569 2506 7574
rect 2702 7546 2842 7574
rect 1918 6118 2114 6146
rect 2310 6118 2450 6146
rect 1974 6089 2002 6118
rect 1974 6063 1975 6089
rect 2001 6063 2002 6089
rect 1974 6057 2002 6063
rect 2086 6090 2114 6118
rect 2086 6062 2338 6090
rect 1638 6033 1666 6039
rect 1638 6007 1639 6033
rect 1665 6007 1666 6033
rect 1134 5418 1162 5423
rect 1638 5418 1666 6007
rect 2030 6034 2058 6039
rect 2030 5987 2058 6006
rect 1936 5894 2068 5899
rect 1964 5866 1988 5894
rect 2016 5866 2040 5894
rect 1936 5861 2068 5866
rect 2310 5753 2338 6062
rect 2310 5727 2311 5753
rect 2337 5727 2338 5753
rect 2310 5721 2338 5727
rect 2366 5698 2394 5703
rect 2366 5651 2394 5670
rect 2422 5586 2450 6118
rect 2702 6145 2730 7546
rect 2814 7210 2842 7215
rect 2814 6537 2842 7182
rect 3266 7070 3398 7075
rect 3294 7042 3318 7070
rect 3346 7042 3370 7070
rect 3266 7037 3398 7042
rect 2814 6511 2815 6537
rect 2841 6511 2842 6537
rect 2814 6505 2842 6511
rect 2870 6370 2898 6375
rect 2870 6369 3234 6370
rect 2870 6343 2871 6369
rect 2897 6343 3234 6369
rect 2870 6342 3234 6343
rect 2870 6337 2898 6342
rect 2702 6119 2703 6145
rect 2729 6119 2730 6145
rect 2702 6034 2730 6119
rect 3150 6202 3178 6207
rect 3206 6202 3234 6342
rect 3266 6286 3398 6291
rect 3294 6258 3318 6286
rect 3346 6258 3370 6286
rect 3266 6253 3398 6258
rect 3318 6202 3346 6207
rect 3206 6201 3346 6202
rect 3206 6175 3319 6201
rect 3345 6175 3346 6201
rect 3206 6174 3346 6175
rect 2758 6090 2786 6095
rect 2982 6090 3010 6095
rect 2758 6089 3010 6090
rect 2758 6063 2759 6089
rect 2785 6063 2983 6089
rect 3009 6063 3010 6089
rect 2758 6062 3010 6063
rect 3150 6090 3178 6174
rect 3318 6169 3346 6174
rect 3206 6090 3234 6095
rect 3150 6089 3234 6090
rect 3150 6063 3207 6089
rect 3233 6063 3234 6089
rect 3150 6062 3234 6063
rect 2758 6057 2786 6062
rect 2982 6057 3010 6062
rect 3206 6057 3234 6062
rect 2702 6001 2730 6006
rect 3262 6033 3290 6039
rect 3262 6007 3263 6033
rect 3289 6007 3290 6033
rect 3262 5586 3290 6007
rect 2310 5558 2450 5586
rect 3206 5558 3290 5586
rect 1078 5417 1162 5418
rect 1078 5391 1135 5417
rect 1161 5391 1162 5417
rect 1078 5390 1162 5391
rect 1134 5306 1162 5390
rect 1582 5390 1890 5418
rect 1134 5273 1162 5278
rect 1302 5361 1330 5367
rect 1302 5335 1303 5361
rect 1329 5335 1330 5361
rect 1302 5026 1330 5335
rect 1582 5249 1610 5390
rect 1638 5306 1666 5311
rect 1638 5259 1666 5278
rect 1582 5223 1583 5249
rect 1609 5223 1610 5249
rect 1582 5217 1610 5223
rect 1862 5026 1890 5390
rect 1974 5249 2002 5255
rect 1974 5223 1975 5249
rect 2001 5223 2002 5249
rect 1974 5194 2002 5223
rect 1974 5166 2226 5194
rect 1936 5110 2068 5115
rect 1964 5082 1988 5110
rect 2016 5082 2040 5110
rect 1936 5077 2068 5082
rect 2030 5026 2058 5031
rect 1862 5025 2058 5026
rect 1862 4999 2031 5025
rect 2057 4999 2058 5025
rect 1862 4998 2058 4999
rect 1302 4993 1330 4998
rect 2030 4993 2058 4998
rect 2142 4914 2170 4919
rect 2142 4867 2170 4886
rect 1862 4802 1890 4807
rect 1806 4801 1890 4802
rect 1806 4775 1863 4801
rect 1889 4775 1890 4801
rect 1806 4774 1890 4775
rect 1694 4522 1722 4527
rect 1582 4130 1610 4135
rect 1582 4083 1610 4102
rect 1694 4073 1722 4494
rect 1806 4521 1834 4774
rect 1862 4769 1890 4774
rect 1806 4495 1807 4521
rect 1833 4495 1834 4521
rect 1806 4489 1834 4495
rect 1918 4522 1946 4527
rect 1918 4475 1946 4494
rect 2086 4522 2114 4527
rect 2198 4522 2226 5166
rect 2254 4522 2282 4527
rect 2086 4521 2282 4522
rect 2086 4495 2087 4521
rect 2113 4495 2255 4521
rect 2281 4495 2282 4521
rect 2086 4494 2282 4495
rect 2086 4489 2114 4494
rect 2254 4489 2282 4494
rect 1974 4465 2002 4471
rect 1974 4439 1975 4465
rect 2001 4439 2002 4465
rect 1974 4410 2002 4439
rect 1974 4382 2170 4410
rect 1936 4326 2068 4331
rect 1964 4298 1988 4326
rect 2016 4298 2040 4326
rect 1936 4293 2068 4298
rect 2142 4186 2170 4382
rect 2142 4153 2170 4158
rect 1918 4130 1946 4135
rect 1918 4083 1946 4102
rect 2086 4129 2114 4135
rect 2086 4103 2087 4129
rect 2113 4103 2114 4129
rect 1694 4047 1695 4073
rect 1721 4047 1722 4073
rect 1694 4041 1722 4047
rect 2086 4018 2114 4103
rect 2086 3985 2114 3990
rect 2310 3738 2338 5558
rect 2478 4522 2506 4527
rect 2366 4494 2478 4522
rect 2366 4073 2394 4494
rect 2478 4475 2506 4494
rect 2702 4465 2730 4471
rect 2702 4439 2703 4465
rect 2729 4439 2730 4465
rect 2366 4047 2367 4073
rect 2393 4047 2394 4073
rect 2366 4041 2394 4047
rect 2478 4129 2506 4135
rect 2478 4103 2479 4129
rect 2505 4103 2506 4129
rect 2422 4018 2450 4023
rect 2422 3793 2450 3990
rect 2422 3767 2423 3793
rect 2449 3767 2450 3793
rect 2422 3761 2450 3767
rect 2366 3738 2394 3743
rect 2310 3737 2394 3738
rect 2310 3711 2367 3737
rect 2393 3711 2394 3737
rect 2310 3710 2394 3711
rect 2478 3738 2506 4103
rect 2702 4130 2730 4439
rect 2870 4186 2898 4191
rect 2870 4139 2898 4158
rect 3206 4186 3234 5558
rect 3266 5502 3398 5507
rect 3294 5474 3318 5502
rect 3346 5474 3370 5502
rect 3266 5469 3398 5474
rect 3266 4718 3398 4723
rect 3294 4690 3318 4718
rect 3346 4690 3370 4718
rect 3266 4685 3398 4690
rect 3430 4522 3458 9983
rect 4774 10010 4802 10015
rect 4774 10009 4858 10010
rect 4774 9983 4775 10009
rect 4801 9983 4858 10009
rect 4774 9982 4858 9983
rect 4774 9977 4802 9982
rect 4596 9814 4728 9819
rect 4624 9786 4648 9814
rect 4676 9786 4700 9814
rect 4596 9781 4728 9786
rect 3878 9562 3906 9567
rect 3990 9562 4018 9567
rect 3878 9515 3906 9534
rect 3934 9534 3990 9562
rect 3934 9505 3962 9534
rect 3990 9529 4018 9534
rect 4158 9561 4186 9567
rect 4158 9535 4159 9561
rect 4185 9535 4186 9561
rect 3934 9479 3935 9505
rect 3961 9479 3962 9505
rect 3934 9338 3962 9479
rect 3934 9305 3962 9310
rect 4046 9505 4074 9511
rect 4046 9479 4047 9505
rect 4073 9479 4074 9505
rect 4046 8946 4074 9479
rect 4158 9226 4186 9535
rect 4326 9282 4354 9287
rect 4326 9235 4354 9254
rect 4774 9281 4802 9287
rect 4774 9255 4775 9281
rect 4801 9255 4802 9281
rect 4158 9193 4186 9198
rect 3934 8918 4074 8946
rect 4102 9170 4130 9175
rect 3878 8778 3906 8783
rect 3822 7378 3850 7383
rect 3822 7331 3850 7350
rect 3766 7210 3794 7215
rect 3766 7163 3794 7182
rect 3822 6202 3850 6207
rect 3822 6089 3850 6174
rect 3878 6146 3906 8750
rect 3934 7770 3962 8918
rect 3990 8834 4018 8839
rect 3990 8787 4018 8806
rect 4046 8834 4074 8839
rect 4102 8834 4130 9142
rect 4046 8833 4130 8834
rect 4046 8807 4047 8833
rect 4073 8807 4130 8833
rect 4046 8806 4130 8807
rect 4046 8801 4074 8806
rect 3990 8722 4018 8727
rect 3990 8675 4018 8694
rect 4102 8553 4130 8806
rect 4102 8527 4103 8553
rect 4129 8527 4130 8553
rect 4102 8521 4130 8527
rect 4158 9113 4186 9119
rect 4158 9087 4159 9113
rect 4185 9087 4186 9113
rect 4158 8833 4186 9087
rect 4270 9114 4298 9119
rect 4270 8945 4298 9086
rect 4774 9114 4802 9255
rect 4774 9081 4802 9086
rect 4596 9030 4728 9035
rect 4624 9002 4648 9030
rect 4676 9002 4700 9030
rect 4596 8997 4728 9002
rect 4270 8919 4271 8945
rect 4297 8919 4298 8945
rect 4270 8913 4298 8919
rect 4158 8807 4159 8833
rect 4185 8807 4186 8833
rect 4158 7938 4186 8807
rect 4158 7905 4186 7910
rect 4214 8441 4242 8447
rect 4214 8415 4215 8441
rect 4241 8415 4242 8441
rect 3990 7770 4018 7775
rect 3934 7769 4018 7770
rect 3934 7743 3991 7769
rect 4017 7743 4018 7769
rect 3934 7742 4018 7743
rect 3990 7737 4018 7742
rect 4158 7545 4186 7551
rect 4158 7519 4159 7545
rect 4185 7519 4186 7545
rect 3934 7434 3962 7439
rect 3934 7377 3962 7406
rect 3934 7351 3935 7377
rect 3961 7351 3962 7377
rect 3934 7098 3962 7351
rect 4046 7322 4074 7327
rect 4046 7265 4074 7294
rect 4046 7239 4047 7265
rect 4073 7239 4074 7265
rect 4046 7233 4074 7239
rect 4158 7210 4186 7519
rect 4214 7434 4242 8415
rect 4596 8246 4728 8251
rect 4624 8218 4648 8246
rect 4676 8218 4700 8246
rect 4596 8213 4728 8218
rect 4550 7938 4578 7943
rect 4550 7891 4578 7910
rect 4718 7937 4746 7943
rect 4718 7911 4719 7937
rect 4745 7911 4746 7937
rect 4326 7658 4354 7663
rect 4270 7602 4298 7607
rect 4326 7602 4354 7630
rect 4270 7601 4354 7602
rect 4270 7575 4271 7601
rect 4297 7575 4354 7601
rect 4270 7574 4354 7575
rect 4382 7602 4410 7607
rect 4270 7569 4298 7574
rect 4214 7401 4242 7406
rect 4270 7378 4298 7383
rect 4270 7331 4298 7350
rect 4382 7377 4410 7574
rect 4718 7546 4746 7911
rect 4830 7770 4858 9982
rect 5614 10009 5642 10015
rect 5614 9983 5615 10009
rect 5641 9983 5642 10009
rect 5502 9617 5530 9623
rect 5502 9591 5503 9617
rect 5529 9591 5530 9617
rect 5502 9337 5530 9591
rect 5614 9561 5642 9983
rect 6790 10009 6818 10015
rect 6790 9983 6791 10009
rect 6817 9983 6818 10009
rect 6790 9730 6818 9983
rect 7518 10010 7546 10015
rect 7256 9814 7388 9819
rect 7284 9786 7308 9814
rect 7336 9786 7360 9814
rect 7256 9781 7388 9786
rect 6790 9697 6818 9702
rect 5614 9535 5615 9561
rect 5641 9535 5642 9561
rect 5614 9529 5642 9535
rect 7406 9617 7434 9623
rect 7406 9591 7407 9617
rect 7433 9591 7434 9617
rect 5926 9422 6058 9427
rect 5954 9394 5978 9422
rect 6006 9394 6030 9422
rect 5926 9389 6058 9394
rect 5502 9311 5503 9337
rect 5529 9311 5530 9337
rect 5502 9305 5530 9311
rect 5558 9282 5586 9287
rect 4942 9225 4970 9231
rect 4942 9199 4943 9225
rect 4969 9199 4970 9225
rect 4942 8946 4970 9199
rect 5558 9225 5586 9254
rect 6062 9282 6090 9287
rect 5558 9199 5559 9225
rect 5585 9199 5586 9225
rect 5558 9193 5586 9199
rect 5614 9226 5642 9231
rect 5446 9114 5474 9119
rect 5446 9113 5530 9114
rect 5446 9087 5447 9113
rect 5473 9087 5530 9113
rect 5446 9086 5530 9087
rect 5446 9081 5474 9086
rect 4830 7737 4858 7742
rect 4886 8918 4942 8946
rect 4718 7513 4746 7518
rect 4774 7658 4802 7663
rect 4774 7601 4802 7630
rect 4774 7575 4775 7601
rect 4801 7575 4802 7601
rect 4596 7462 4728 7467
rect 4624 7434 4648 7462
rect 4676 7434 4700 7462
rect 4596 7429 4728 7434
rect 4382 7351 4383 7377
rect 4409 7351 4410 7377
rect 4382 7345 4410 7351
rect 4494 7322 4522 7327
rect 4494 7265 4522 7294
rect 4494 7239 4495 7265
rect 4521 7239 4522 7265
rect 4494 7233 4522 7239
rect 4214 7210 4242 7215
rect 4158 7209 4242 7210
rect 4158 7183 4215 7209
rect 4241 7183 4242 7209
rect 4158 7182 4242 7183
rect 3934 7065 3962 7070
rect 4214 6481 4242 7182
rect 4596 6678 4728 6683
rect 4624 6650 4648 6678
rect 4676 6650 4700 6678
rect 4596 6645 4728 6650
rect 4382 6538 4410 6543
rect 4382 6537 4466 6538
rect 4382 6511 4383 6537
rect 4409 6511 4466 6537
rect 4382 6510 4466 6511
rect 4382 6505 4410 6510
rect 4214 6455 4215 6481
rect 4241 6455 4242 6481
rect 4214 6449 4242 6455
rect 4102 6425 4130 6431
rect 4102 6399 4103 6425
rect 4129 6399 4130 6425
rect 3934 6146 3962 6151
rect 3878 6118 3934 6146
rect 3934 6099 3962 6118
rect 3822 6063 3823 6089
rect 3849 6063 3850 6089
rect 3822 6057 3850 6063
rect 4102 5306 4130 6399
rect 4438 6426 4466 6510
rect 4774 6426 4802 7575
rect 4830 7658 4858 7663
rect 4886 7658 4914 8918
rect 4942 8913 4970 8918
rect 5110 9058 5138 9063
rect 4830 7657 4914 7658
rect 4830 7631 4831 7657
rect 4857 7631 4914 7657
rect 4830 7630 4914 7631
rect 4830 7378 4858 7630
rect 4830 7345 4858 7350
rect 4942 7601 4970 7607
rect 4942 7575 4943 7601
rect 4969 7575 4970 7601
rect 4942 7546 4970 7575
rect 4998 7602 5026 7607
rect 4998 7555 5026 7574
rect 4942 7378 4970 7518
rect 4942 7345 4970 7350
rect 4998 7322 5026 7327
rect 4998 6873 5026 7294
rect 4998 6847 4999 6873
rect 5025 6847 5026 6873
rect 4998 6841 5026 6847
rect 5110 6873 5138 9030
rect 5502 9002 5530 9086
rect 5614 9002 5642 9198
rect 5782 9225 5810 9231
rect 5782 9199 5783 9225
rect 5809 9199 5810 9225
rect 5670 9113 5698 9119
rect 5670 9087 5671 9113
rect 5697 9087 5698 9113
rect 5670 9058 5698 9087
rect 5782 9058 5810 9199
rect 5950 9225 5978 9231
rect 5950 9199 5951 9225
rect 5977 9199 5978 9225
rect 5950 9170 5978 9199
rect 6062 9226 6090 9254
rect 6342 9282 6370 9287
rect 6342 9235 6370 9254
rect 6678 9281 6706 9287
rect 6678 9255 6679 9281
rect 6705 9255 6706 9281
rect 6174 9226 6202 9231
rect 6062 9225 6202 9226
rect 6062 9199 6175 9225
rect 6201 9199 6202 9225
rect 6062 9198 6202 9199
rect 6174 9170 6202 9198
rect 6286 9226 6314 9231
rect 6286 9179 6314 9198
rect 6510 9225 6538 9231
rect 6510 9199 6511 9225
rect 6537 9199 6538 9225
rect 5978 9142 6034 9170
rect 5950 9137 5978 9142
rect 5670 9025 5698 9030
rect 5726 9030 5782 9058
rect 5502 8974 5642 9002
rect 5446 8946 5474 8951
rect 5446 8899 5474 8918
rect 5502 8890 5530 8895
rect 5502 8843 5530 8862
rect 5614 8833 5642 8974
rect 5670 8946 5698 8951
rect 5670 8899 5698 8918
rect 5614 8807 5615 8833
rect 5641 8807 5642 8833
rect 5614 8442 5642 8807
rect 5614 8409 5642 8414
rect 5726 7826 5754 9030
rect 5782 9025 5810 9030
rect 6006 8946 6034 9142
rect 6174 9137 6202 9142
rect 6062 9113 6090 9119
rect 6062 9087 6063 9113
rect 6089 9087 6090 9113
rect 6062 9058 6090 9087
rect 6062 9030 6370 9058
rect 6062 8946 6090 8951
rect 6006 8945 6090 8946
rect 6006 8919 6063 8945
rect 6089 8919 6090 8945
rect 6006 8918 6090 8919
rect 6062 8913 6090 8918
rect 5950 8890 5978 8895
rect 5950 8843 5978 8862
rect 6174 8834 6202 8839
rect 6174 8833 6314 8834
rect 6174 8807 6175 8833
rect 6201 8807 6314 8833
rect 6174 8806 6314 8807
rect 6174 8801 6202 8806
rect 6118 8722 6146 8727
rect 6230 8722 6258 8727
rect 6118 8721 6230 8722
rect 6118 8695 6119 8721
rect 6145 8695 6230 8721
rect 6118 8694 6230 8695
rect 6118 8689 6146 8694
rect 5926 8638 6058 8643
rect 5954 8610 5978 8638
rect 6006 8610 6030 8638
rect 5926 8605 6058 8610
rect 6174 8553 6202 8694
rect 6230 8689 6258 8694
rect 6174 8527 6175 8553
rect 6201 8527 6202 8553
rect 6174 8521 6202 8527
rect 6006 8497 6034 8503
rect 6006 8471 6007 8497
rect 6033 8471 6034 8497
rect 6006 7938 6034 8471
rect 6174 8442 6202 8447
rect 6006 7910 6146 7938
rect 5502 7798 5754 7826
rect 5926 7854 6058 7859
rect 5954 7826 5978 7854
rect 6006 7826 6030 7854
rect 5926 7821 6058 7826
rect 5390 7322 5418 7327
rect 5390 7265 5418 7294
rect 5390 7239 5391 7265
rect 5417 7239 5418 7265
rect 5390 7233 5418 7239
rect 5110 6847 5111 6873
rect 5137 6847 5138 6873
rect 5110 6841 5138 6847
rect 5222 7210 5250 7215
rect 5222 6873 5250 7182
rect 5502 7209 5530 7798
rect 5502 7183 5503 7209
rect 5529 7183 5530 7209
rect 5502 7177 5530 7183
rect 5670 7265 5698 7271
rect 5670 7239 5671 7265
rect 5697 7239 5698 7265
rect 5670 7210 5698 7239
rect 5670 7177 5698 7182
rect 5614 7098 5642 7103
rect 5614 6986 5642 7070
rect 5222 6847 5223 6873
rect 5249 6847 5250 6873
rect 5222 6841 5250 6847
rect 5502 6874 5530 6879
rect 5502 6827 5530 6846
rect 5614 6873 5642 6958
rect 5614 6847 5615 6873
rect 5641 6847 5642 6873
rect 5614 6841 5642 6847
rect 5726 6930 5754 7798
rect 6062 7713 6090 7719
rect 6062 7687 6063 7713
rect 6089 7687 6090 7713
rect 5894 7602 5922 7607
rect 5782 7378 5810 7383
rect 5782 7331 5810 7350
rect 5894 7266 5922 7574
rect 6062 7322 6090 7687
rect 6118 7602 6146 7910
rect 6118 7569 6146 7574
rect 6174 7574 6202 8414
rect 6230 7658 6258 7663
rect 6230 7611 6258 7630
rect 6174 7546 6258 7574
rect 6062 7289 6090 7294
rect 5894 7219 5922 7238
rect 6118 7154 6146 7159
rect 5926 7070 6058 7075
rect 5954 7042 5978 7070
rect 6006 7042 6030 7070
rect 5926 7037 6058 7042
rect 5726 6873 5754 6902
rect 5726 6847 5727 6873
rect 5753 6847 5754 6873
rect 5726 6841 5754 6847
rect 5838 6873 5866 6879
rect 5838 6847 5839 6873
rect 5865 6847 5866 6873
rect 4942 6818 4970 6823
rect 4438 6398 4634 6426
rect 4326 6369 4354 6375
rect 4326 6343 4327 6369
rect 4353 6343 4354 6369
rect 4326 5894 4354 6343
rect 4382 6370 4410 6375
rect 4382 6314 4410 6342
rect 4382 6286 4522 6314
rect 4102 5273 4130 5278
rect 4214 5866 4354 5894
rect 4382 6090 4410 6095
rect 4214 4970 4242 5866
rect 4382 5809 4410 6062
rect 4382 5783 4383 5809
rect 4409 5783 4410 5809
rect 4382 5777 4410 5783
rect 4438 5754 4466 5759
rect 4438 5641 4466 5726
rect 4438 5615 4439 5641
rect 4465 5615 4466 5641
rect 4438 5609 4466 5615
rect 4494 5362 4522 6286
rect 4606 6258 4634 6398
rect 4662 6398 4802 6426
rect 4830 6762 4858 6767
rect 4662 6370 4690 6398
rect 4662 6337 4690 6342
rect 4606 6230 4802 6258
rect 4774 6201 4802 6230
rect 4774 6175 4775 6201
rect 4801 6175 4802 6201
rect 4774 6169 4802 6175
rect 4830 6201 4858 6734
rect 4830 6175 4831 6201
rect 4857 6175 4858 6201
rect 4830 6169 4858 6175
rect 4942 6202 4970 6790
rect 5838 6818 5866 6847
rect 5838 6785 5866 6790
rect 4942 6169 4970 6174
rect 5278 6761 5306 6767
rect 5278 6735 5279 6761
rect 5305 6735 5306 6761
rect 5110 6146 5138 6151
rect 4886 6090 4914 6095
rect 5054 6090 5082 6095
rect 4886 6089 4970 6090
rect 4886 6063 4887 6089
rect 4913 6063 4970 6089
rect 4886 6062 4970 6063
rect 4886 6057 4914 6062
rect 4596 5894 4728 5899
rect 4624 5866 4648 5894
rect 4676 5866 4700 5894
rect 4596 5861 4728 5866
rect 4942 5754 4970 6062
rect 5054 6043 5082 6062
rect 4606 5698 4634 5703
rect 4550 5642 4578 5647
rect 4550 5595 4578 5614
rect 4550 5362 4578 5367
rect 4494 5334 4550 5362
rect 4550 5329 4578 5334
rect 4214 4857 4242 4942
rect 4270 5306 4298 5311
rect 4270 4969 4298 5278
rect 4606 5194 4634 5670
rect 4270 4943 4271 4969
rect 4297 4943 4298 4969
rect 4270 4937 4298 4943
rect 4494 5166 4634 5194
rect 4886 5698 4914 5703
rect 4494 4969 4522 5166
rect 4596 5110 4728 5115
rect 4624 5082 4648 5110
rect 4676 5082 4700 5110
rect 4596 5077 4728 5082
rect 4494 4943 4495 4969
rect 4521 4943 4522 4969
rect 4494 4937 4522 4943
rect 4606 4970 4634 4975
rect 4606 4923 4634 4942
rect 4214 4831 4215 4857
rect 4241 4831 4242 4857
rect 4214 4825 4242 4831
rect 4326 4857 4354 4863
rect 4550 4858 4578 4863
rect 4326 4831 4327 4857
rect 4353 4831 4354 4857
rect 4326 4634 4354 4831
rect 4326 4601 4354 4606
rect 4494 4830 4550 4858
rect 3430 4489 3458 4494
rect 3206 4153 3234 4158
rect 3710 4186 3738 4191
rect 2702 4097 2730 4102
rect 2982 4129 3010 4135
rect 2982 4103 2983 4129
rect 3009 4103 3010 4129
rect 2814 4018 2842 4023
rect 2814 3971 2842 3990
rect 2982 4018 3010 4103
rect 3654 4130 3682 4135
rect 3654 4083 3682 4102
rect 3150 4074 3178 4079
rect 3262 4074 3290 4079
rect 3150 4027 3178 4046
rect 3206 4073 3290 4074
rect 3206 4047 3263 4073
rect 3289 4047 3290 4073
rect 3206 4046 3290 4047
rect 2982 3985 3010 3990
rect 3206 3906 3234 4046
rect 3262 4041 3290 4046
rect 3710 4073 3738 4158
rect 4438 4186 4466 4191
rect 4494 4186 4522 4830
rect 4550 4825 4578 4830
rect 4774 4802 4802 4807
rect 4886 4802 4914 5670
rect 4942 5642 4970 5726
rect 5110 5754 5138 6118
rect 5110 5697 5138 5726
rect 5110 5671 5111 5697
rect 5137 5671 5138 5697
rect 5110 5665 5138 5671
rect 5222 5698 5250 5703
rect 5222 5651 5250 5670
rect 4998 5642 5026 5647
rect 4942 5614 4998 5642
rect 4998 5609 5026 5614
rect 5166 5585 5194 5591
rect 5166 5559 5167 5585
rect 5193 5559 5194 5585
rect 5166 5250 5194 5559
rect 4998 5222 5194 5250
rect 4998 5025 5026 5222
rect 4998 4999 4999 5025
rect 5025 4999 5026 5025
rect 4998 4993 5026 4999
rect 5278 4970 5306 6735
rect 5054 4942 5306 4970
rect 5446 6761 5474 6767
rect 5446 6735 5447 6761
rect 5473 6735 5474 6761
rect 4942 4914 4970 4919
rect 4942 4867 4970 4886
rect 4886 4774 5026 4802
rect 4774 4755 4802 4774
rect 4998 4521 5026 4774
rect 4998 4495 4999 4521
rect 5025 4495 5026 4521
rect 4998 4489 5026 4495
rect 4596 4326 4728 4331
rect 4624 4298 4648 4326
rect 4676 4298 4700 4326
rect 4596 4293 4728 4298
rect 4662 4242 4690 4247
rect 5054 4242 5082 4942
rect 5390 4914 5418 4919
rect 5166 4858 5194 4863
rect 5166 4811 5194 4830
rect 5278 4857 5306 4863
rect 5278 4831 5279 4857
rect 5305 4831 5306 4857
rect 5278 4802 5306 4831
rect 5278 4769 5306 4774
rect 5334 4801 5362 4807
rect 5334 4775 5335 4801
rect 5361 4775 5362 4801
rect 5222 4578 5250 4583
rect 5166 4550 5222 4578
rect 5166 4521 5194 4550
rect 5222 4545 5250 4550
rect 5166 4495 5167 4521
rect 5193 4495 5194 4521
rect 5166 4489 5194 4495
rect 4550 4186 4578 4191
rect 4494 4185 4578 4186
rect 4494 4159 4551 4185
rect 4577 4159 4578 4185
rect 4494 4158 4578 4159
rect 3822 4130 3850 4135
rect 3822 4083 3850 4102
rect 3710 4047 3711 4073
rect 3737 4047 3738 4073
rect 3710 4041 3738 4047
rect 2534 3878 3234 3906
rect 3266 3934 3398 3939
rect 3294 3906 3318 3934
rect 3346 3906 3370 3934
rect 3266 3901 3398 3906
rect 2534 3849 2562 3878
rect 2534 3823 2535 3849
rect 2561 3823 2562 3849
rect 2534 3817 2562 3823
rect 4438 3850 4466 4158
rect 4550 4153 4578 4158
rect 4662 4185 4690 4214
rect 4662 4159 4663 4185
rect 4689 4159 4690 4185
rect 4662 4153 4690 4159
rect 4942 4214 5082 4242
rect 4942 4130 4970 4214
rect 5054 4186 5082 4214
rect 5054 4153 5082 4158
rect 5110 4465 5138 4471
rect 5110 4439 5111 4465
rect 5137 4439 5138 4465
rect 4830 4102 4970 4130
rect 4830 4074 4858 4102
rect 4830 4041 4858 4046
rect 4886 4017 4914 4023
rect 4886 3991 4887 4017
rect 4913 3991 4914 4017
rect 4886 3962 4914 3991
rect 4886 3929 4914 3934
rect 4438 3817 4466 3822
rect 4942 3849 4970 4102
rect 4998 4130 5026 4135
rect 4998 4083 5026 4102
rect 5054 4073 5082 4079
rect 5054 4047 5055 4073
rect 5081 4047 5082 4073
rect 5054 3962 5082 4047
rect 5110 4074 5138 4439
rect 5334 4410 5362 4775
rect 5390 4802 5418 4886
rect 5446 4913 5474 6735
rect 5926 6286 6058 6291
rect 5954 6258 5978 6286
rect 6006 6258 6030 6286
rect 5926 6253 6058 6258
rect 6118 5698 6146 7126
rect 6230 7153 6258 7546
rect 6286 7546 6314 8806
rect 6342 7938 6370 9030
rect 6510 8722 6538 9199
rect 6510 8689 6538 8694
rect 6622 9170 6650 9175
rect 6622 8386 6650 9142
rect 6678 9002 6706 9255
rect 7406 9281 7434 9591
rect 7518 9561 7546 9982
rect 7854 10010 7882 10015
rect 7854 9963 7882 9982
rect 8974 10009 9002 10015
rect 8974 9983 8975 10009
rect 9001 9983 9002 10009
rect 8974 9786 9002 9983
rect 8974 9753 9002 9758
rect 9254 10010 9282 10015
rect 8302 9730 8330 9735
rect 8302 9683 8330 9702
rect 8134 9618 8162 9623
rect 8302 9618 8330 9623
rect 8134 9617 8330 9618
rect 8134 9591 8135 9617
rect 8161 9591 8303 9617
rect 8329 9591 8330 9617
rect 8134 9590 8330 9591
rect 8134 9585 8162 9590
rect 8302 9585 8330 9590
rect 8470 9618 8498 9623
rect 8918 9618 8946 9623
rect 9198 9618 9226 9623
rect 8470 9617 8834 9618
rect 8470 9591 8471 9617
rect 8497 9591 8834 9617
rect 8470 9590 8834 9591
rect 8470 9585 8498 9590
rect 7518 9535 7519 9561
rect 7545 9535 7546 9561
rect 7518 9529 7546 9535
rect 8078 9561 8106 9567
rect 8078 9535 8079 9561
rect 8105 9535 8106 9561
rect 8078 9506 8106 9535
rect 8022 9478 8078 9506
rect 8022 9337 8050 9478
rect 8078 9473 8106 9478
rect 8750 9506 8778 9511
rect 8750 9459 8778 9478
rect 8586 9422 8718 9427
rect 8614 9394 8638 9422
rect 8666 9394 8690 9422
rect 8586 9389 8718 9394
rect 8806 9394 8834 9590
rect 8918 9617 9226 9618
rect 8918 9591 8919 9617
rect 8945 9591 9199 9617
rect 9225 9591 9226 9617
rect 8918 9590 9226 9591
rect 8918 9585 8946 9590
rect 9198 9585 9226 9590
rect 8862 9506 8890 9511
rect 8862 9459 8890 9478
rect 8974 9506 9002 9511
rect 9142 9506 9170 9511
rect 8974 9505 9170 9506
rect 8974 9479 8975 9505
rect 9001 9479 9143 9505
rect 9169 9479 9170 9505
rect 8974 9478 9170 9479
rect 8974 9394 9002 9478
rect 9142 9473 9170 9478
rect 8806 9366 9002 9394
rect 8022 9311 8023 9337
rect 8049 9311 8050 9337
rect 8022 9305 8050 9311
rect 9142 9338 9170 9343
rect 9254 9338 9282 9982
rect 9926 10009 9954 10015
rect 9926 9983 9927 10009
rect 9953 9983 9954 10009
rect 9926 9898 9954 9983
rect 10486 10010 10514 10015
rect 10486 9963 10514 9982
rect 10934 10010 10962 10015
rect 10934 10009 11018 10010
rect 10934 9983 10935 10009
rect 10961 9983 11018 10009
rect 10934 9982 11018 9983
rect 10934 9977 10962 9982
rect 9814 9870 9954 9898
rect 9142 9337 9282 9338
rect 9142 9311 9143 9337
rect 9169 9311 9282 9337
rect 9142 9310 9282 9311
rect 9478 9506 9506 9511
rect 9142 9305 9170 9310
rect 7406 9255 7407 9281
rect 7433 9255 7434 9281
rect 7406 9249 7434 9255
rect 7854 9282 7882 9287
rect 7854 9235 7882 9254
rect 9254 9226 9282 9231
rect 9254 9225 9338 9226
rect 9254 9199 9255 9225
rect 9281 9199 9338 9225
rect 9254 9198 9338 9199
rect 9254 9193 9282 9198
rect 7686 9170 7714 9175
rect 6678 8969 6706 8974
rect 7070 9113 7098 9119
rect 7070 9087 7071 9113
rect 7097 9087 7098 9113
rect 6622 8353 6650 8358
rect 6790 8890 6818 8895
rect 6790 8161 6818 8862
rect 7070 8778 7098 9087
rect 7126 9113 7154 9119
rect 7238 9114 7266 9119
rect 7126 9087 7127 9113
rect 7153 9087 7154 9113
rect 7126 9058 7154 9087
rect 7126 9025 7154 9030
rect 7182 9113 7266 9114
rect 7182 9087 7239 9113
rect 7265 9087 7266 9113
rect 7182 9086 7266 9087
rect 7070 8745 7098 8750
rect 7182 9002 7210 9086
rect 7238 9081 7266 9086
rect 7350 9114 7378 9133
rect 7378 9086 7490 9114
rect 7350 9081 7378 9086
rect 7256 9030 7388 9035
rect 7284 9002 7308 9030
rect 7336 9002 7360 9030
rect 7256 8997 7388 9002
rect 7182 8442 7210 8974
rect 7462 8834 7490 9086
rect 7686 8945 7714 9142
rect 9086 9114 9114 9119
rect 7686 8919 7687 8945
rect 7713 8919 7714 8945
rect 7686 8913 7714 8919
rect 9030 9113 9114 9114
rect 9030 9087 9087 9113
rect 9113 9087 9114 9113
rect 9030 9086 9114 9087
rect 7518 8834 7546 8839
rect 7462 8833 7546 8834
rect 7462 8807 7519 8833
rect 7545 8807 7546 8833
rect 7462 8806 7546 8807
rect 7518 8801 7546 8806
rect 7182 8409 7210 8414
rect 7630 8721 7658 8727
rect 7630 8695 7631 8721
rect 7657 8695 7658 8721
rect 6902 8386 6930 8391
rect 6790 8135 6791 8161
rect 6817 8135 6818 8161
rect 6790 8129 6818 8135
rect 6846 8358 6902 8386
rect 6342 7905 6370 7910
rect 6286 7513 6314 7518
rect 6342 7265 6370 7271
rect 6342 7239 6343 7265
rect 6369 7239 6370 7265
rect 6342 7210 6370 7239
rect 6342 7177 6370 7182
rect 6790 7209 6818 7215
rect 6790 7183 6791 7209
rect 6817 7183 6818 7209
rect 6230 7127 6231 7153
rect 6257 7127 6258 7153
rect 6230 6874 6258 7127
rect 6790 6986 6818 7183
rect 6790 6953 6818 6958
rect 6230 6841 6258 6846
rect 6846 6818 6874 8358
rect 6902 8353 6930 8358
rect 7256 8246 7388 8251
rect 7284 8218 7308 8246
rect 7336 8218 7360 8246
rect 7256 8213 7388 8218
rect 6902 8049 6930 8055
rect 6902 8023 6903 8049
rect 6929 8023 6930 8049
rect 6902 7938 6930 8023
rect 7014 8049 7042 8055
rect 7014 8023 7015 8049
rect 7041 8023 7042 8049
rect 6902 7905 6930 7910
rect 6958 7937 6986 7943
rect 6958 7911 6959 7937
rect 6985 7911 6986 7937
rect 6958 7658 6986 7911
rect 7014 7714 7042 8023
rect 7630 7882 7658 8695
rect 8586 8638 8718 8643
rect 8614 8610 8638 8638
rect 8666 8610 8690 8638
rect 8586 8605 8718 8610
rect 7406 7854 7658 7882
rect 7854 8442 7882 8447
rect 7406 7769 7434 7854
rect 7406 7743 7407 7769
rect 7433 7743 7434 7769
rect 7406 7737 7434 7743
rect 7238 7714 7266 7719
rect 7014 7681 7042 7686
rect 7182 7713 7266 7714
rect 7182 7687 7239 7713
rect 7265 7687 7266 7713
rect 7182 7686 7266 7687
rect 6958 7602 6986 7630
rect 6958 7574 7154 7602
rect 7014 7490 7042 7495
rect 6902 7266 6930 7271
rect 6902 7219 6930 7238
rect 7014 7265 7042 7462
rect 7126 7378 7154 7574
rect 7182 7490 7210 7686
rect 7238 7681 7266 7686
rect 7182 7457 7210 7462
rect 7256 7462 7388 7467
rect 7284 7434 7308 7462
rect 7336 7434 7360 7462
rect 7256 7429 7388 7434
rect 7126 7350 7378 7378
rect 7014 7239 7015 7265
rect 7041 7239 7042 7265
rect 7014 7210 7042 7239
rect 7182 7266 7210 7285
rect 7210 7238 7266 7266
rect 7182 7233 7210 7238
rect 7014 7177 7042 7182
rect 7182 7153 7210 7159
rect 7182 7127 7183 7153
rect 7209 7127 7210 7153
rect 7126 6986 7154 6991
rect 7126 6939 7154 6958
rect 6846 6790 7098 6818
rect 7070 6370 7098 6790
rect 7182 6482 7210 7127
rect 7238 6818 7266 7238
rect 7350 7265 7378 7350
rect 7574 7377 7602 7854
rect 7574 7351 7575 7377
rect 7601 7351 7602 7377
rect 7574 7345 7602 7351
rect 7798 7322 7826 7327
rect 7798 7275 7826 7294
rect 7350 7239 7351 7265
rect 7377 7239 7378 7265
rect 7350 7233 7378 7239
rect 7462 7266 7490 7271
rect 7294 6986 7322 6991
rect 7462 6986 7490 7238
rect 7294 6985 7490 6986
rect 7294 6959 7295 6985
rect 7321 6959 7490 6985
rect 7294 6958 7490 6959
rect 7630 7209 7658 7215
rect 7630 7183 7631 7209
rect 7657 7183 7658 7209
rect 7294 6953 7322 6958
rect 7518 6930 7546 6935
rect 7518 6883 7546 6902
rect 7630 6874 7658 7183
rect 7854 7209 7882 8414
rect 9030 8049 9058 9086
rect 9086 9081 9114 9086
rect 9086 8386 9114 8391
rect 9310 8386 9338 9198
rect 9114 8358 9338 8386
rect 9086 8161 9114 8358
rect 9254 8162 9282 8167
rect 9086 8135 9087 8161
rect 9113 8135 9114 8161
rect 9086 8129 9114 8135
rect 9198 8134 9254 8162
rect 9030 8023 9031 8049
rect 9057 8023 9058 8049
rect 8022 7994 8050 7999
rect 7854 7183 7855 7209
rect 7881 7183 7882 7209
rect 7854 7177 7882 7183
rect 7966 7210 7994 7215
rect 7966 7163 7994 7182
rect 7966 6986 7994 6991
rect 8022 6986 8050 7966
rect 8862 7994 8890 7999
rect 8862 7947 8890 7966
rect 8586 7854 8718 7859
rect 8614 7826 8638 7854
rect 8666 7826 8690 7854
rect 8586 7821 8718 7826
rect 9030 7154 9058 8023
rect 9198 8049 9226 8134
rect 9254 8129 9282 8134
rect 9198 8023 9199 8049
rect 9225 8023 9226 8049
rect 9198 8017 9226 8023
rect 9422 7994 9450 7999
rect 9254 7993 9450 7994
rect 9254 7967 9423 7993
rect 9449 7967 9450 7993
rect 9254 7966 9450 7967
rect 9254 7937 9282 7966
rect 9422 7961 9450 7966
rect 9254 7911 9255 7937
rect 9281 7911 9282 7937
rect 9254 7905 9282 7911
rect 9422 7770 9450 7775
rect 9254 7602 9282 7607
rect 9198 7546 9226 7551
rect 9030 7121 9058 7126
rect 9142 7210 9170 7215
rect 8586 7070 8718 7075
rect 8614 7042 8638 7070
rect 8666 7042 8690 7070
rect 8586 7037 8718 7042
rect 7966 6985 8050 6986
rect 7966 6959 7967 6985
rect 7993 6959 8050 6985
rect 7966 6958 8050 6959
rect 7966 6953 7994 6958
rect 7854 6929 7882 6935
rect 7854 6903 7855 6929
rect 7881 6903 7882 6929
rect 7798 6874 7826 6879
rect 7630 6873 7826 6874
rect 7630 6847 7799 6873
rect 7825 6847 7826 6873
rect 7630 6846 7826 6847
rect 7462 6818 7490 6823
rect 7238 6817 7490 6818
rect 7238 6791 7463 6817
rect 7489 6791 7490 6817
rect 7238 6790 7490 6791
rect 7462 6785 7490 6790
rect 7630 6761 7658 6767
rect 7630 6735 7631 6761
rect 7657 6735 7658 6761
rect 7256 6678 7388 6683
rect 7284 6650 7308 6678
rect 7336 6650 7360 6678
rect 7256 6645 7388 6650
rect 7630 6594 7658 6735
rect 7630 6561 7658 6566
rect 7182 6454 7266 6482
rect 7182 6370 7210 6375
rect 7070 6369 7210 6370
rect 7070 6343 7183 6369
rect 7209 6343 7210 6369
rect 7070 6342 7210 6343
rect 7182 6337 7210 6342
rect 7238 6202 7266 6454
rect 6118 5665 6146 5670
rect 7126 6174 7266 6202
rect 7294 6481 7322 6487
rect 7294 6455 7295 6481
rect 7321 6455 7322 6481
rect 6734 5642 6762 5647
rect 5926 5502 6058 5507
rect 5954 5474 5978 5502
rect 6006 5474 6030 5502
rect 5926 5469 6058 5474
rect 6454 5362 6482 5367
rect 6454 5315 6482 5334
rect 6566 5306 6594 5311
rect 6566 5259 6594 5278
rect 6734 5305 6762 5614
rect 7126 5417 7154 6174
rect 7294 5978 7322 6455
rect 7798 6426 7826 6846
rect 7182 5950 7322 5978
rect 7462 6398 7826 6426
rect 7182 5642 7210 5950
rect 7256 5894 7388 5899
rect 7284 5866 7308 5894
rect 7336 5866 7360 5894
rect 7256 5861 7388 5866
rect 7462 5810 7490 6398
rect 7182 5595 7210 5614
rect 7238 5782 7490 5810
rect 7126 5391 7127 5417
rect 7153 5391 7154 5417
rect 7126 5385 7154 5391
rect 7238 5417 7266 5782
rect 7518 5753 7546 5759
rect 7518 5727 7519 5753
rect 7545 5727 7546 5753
rect 7350 5586 7378 5591
rect 7518 5586 7546 5727
rect 7574 5642 7602 5647
rect 7574 5595 7602 5614
rect 7686 5642 7714 5647
rect 7686 5595 7714 5614
rect 7350 5585 7546 5586
rect 7350 5559 7351 5585
rect 7377 5559 7546 5585
rect 7350 5558 7546 5559
rect 7350 5553 7378 5558
rect 7238 5391 7239 5417
rect 7265 5391 7266 5417
rect 7238 5385 7266 5391
rect 6734 5279 6735 5305
rect 6761 5279 6762 5305
rect 6734 5273 6762 5279
rect 7294 5306 7322 5311
rect 7406 5306 7434 5558
rect 7686 5362 7714 5367
rect 7462 5306 7490 5311
rect 7322 5278 7378 5306
rect 7406 5278 7462 5306
rect 7294 5259 7322 5278
rect 7182 5249 7210 5255
rect 7182 5223 7183 5249
rect 7209 5223 7210 5249
rect 5446 4887 5447 4913
rect 5473 4887 5474 4913
rect 5446 4881 5474 4887
rect 5502 5194 5530 5199
rect 5390 4633 5418 4774
rect 5390 4607 5391 4633
rect 5417 4607 5418 4633
rect 5390 4601 5418 4607
rect 5446 4578 5474 4583
rect 5502 4578 5530 5166
rect 6510 5194 6538 5199
rect 6510 5147 6538 5166
rect 6846 5194 6874 5199
rect 6846 5147 6874 5166
rect 7182 5082 7210 5223
rect 7350 5194 7378 5278
rect 7462 5259 7490 5278
rect 7574 5194 7602 5199
rect 7350 5166 7490 5194
rect 7014 5054 7210 5082
rect 7256 5110 7388 5115
rect 7284 5082 7308 5110
rect 7336 5082 7360 5110
rect 7256 5077 7388 5082
rect 7462 5082 7490 5166
rect 7574 5147 7602 5166
rect 7014 4969 7042 5054
rect 7462 5049 7490 5054
rect 7014 4943 7015 4969
rect 7041 4943 7042 4969
rect 7014 4937 7042 4943
rect 7574 4970 7602 4975
rect 7574 4923 7602 4942
rect 7686 4913 7714 5334
rect 7798 5193 7826 5199
rect 7798 5167 7799 5193
rect 7825 5167 7826 5193
rect 7798 5082 7826 5167
rect 7798 5049 7826 5054
rect 7854 4970 7882 6903
rect 9142 6929 9170 7182
rect 9142 6903 9143 6929
rect 9169 6903 9170 6929
rect 7910 6874 7938 6879
rect 9142 6874 9170 6903
rect 7938 6846 7994 6874
rect 7910 6841 7938 6846
rect 7966 5417 7994 6846
rect 9142 6841 9170 6846
rect 9198 7154 9226 7518
rect 9198 6873 9226 7126
rect 9198 6847 9199 6873
rect 9225 6847 9226 6873
rect 9198 6841 9226 6847
rect 9254 6706 9282 7574
rect 9366 7210 9394 7215
rect 9310 6986 9338 6991
rect 9310 6873 9338 6958
rect 9310 6847 9311 6873
rect 9337 6847 9338 6873
rect 9310 6841 9338 6847
rect 9366 6762 9394 7182
rect 9422 6874 9450 7742
rect 9478 7098 9506 9478
rect 9814 9338 9842 9870
rect 9916 9814 10048 9819
rect 9944 9786 9968 9814
rect 9996 9786 10020 9814
rect 9916 9781 10048 9786
rect 10038 9561 10066 9567
rect 10038 9535 10039 9561
rect 10065 9535 10066 9561
rect 9870 9506 9898 9511
rect 9870 9459 9898 9478
rect 9814 9305 9842 9310
rect 9758 9281 9786 9287
rect 9758 9255 9759 9281
rect 9785 9255 9786 9281
rect 9758 9226 9786 9255
rect 10038 9282 10066 9535
rect 10822 9562 10850 9567
rect 10822 9515 10850 9534
rect 10934 9505 10962 9511
rect 10934 9479 10935 9505
rect 10961 9479 10962 9505
rect 10542 9338 10570 9343
rect 10038 9249 10066 9254
rect 10318 9337 10570 9338
rect 10318 9311 10543 9337
rect 10569 9311 10570 9337
rect 10318 9310 10570 9311
rect 9758 9193 9786 9198
rect 10206 9226 10234 9231
rect 10318 9226 10346 9310
rect 10542 9305 10570 9310
rect 10038 9170 10066 9175
rect 9702 9113 9730 9119
rect 9702 9087 9703 9113
rect 9729 9087 9730 9113
rect 9702 8946 9730 9087
rect 9870 9114 9898 9133
rect 10038 9123 10066 9142
rect 9870 9081 9898 9086
rect 10094 9113 10122 9119
rect 10094 9087 10095 9113
rect 10121 9087 10122 9113
rect 9916 9030 10048 9035
rect 9944 9002 9968 9030
rect 9996 9002 10020 9030
rect 9916 8997 10048 9002
rect 9702 8913 9730 8918
rect 10094 8946 10122 9087
rect 10094 8833 10122 8918
rect 10150 9114 10178 9119
rect 10150 8889 10178 9086
rect 10150 8863 10151 8889
rect 10177 8863 10178 8889
rect 10150 8857 10178 8863
rect 10206 9113 10234 9198
rect 10206 9087 10207 9113
rect 10233 9087 10234 9113
rect 10094 8807 10095 8833
rect 10121 8807 10122 8833
rect 10094 8801 10122 8807
rect 10038 8554 10066 8559
rect 10038 8442 10066 8526
rect 9982 8441 10066 8442
rect 9982 8415 10039 8441
rect 10065 8415 10066 8441
rect 9982 8414 10066 8415
rect 9870 8330 9898 8335
rect 9814 8329 9898 8330
rect 9814 8303 9871 8329
rect 9897 8303 9898 8329
rect 9814 8302 9898 8303
rect 9814 8162 9842 8302
rect 9870 8297 9898 8302
rect 9982 8330 10010 8414
rect 10038 8409 10066 8414
rect 10094 8442 10122 8447
rect 10206 8442 10234 9087
rect 10262 9225 10346 9226
rect 10262 9199 10319 9225
rect 10345 9199 10346 9225
rect 10262 9198 10346 9199
rect 10262 8945 10290 9198
rect 10318 9193 10346 9198
rect 10486 9225 10514 9231
rect 10486 9199 10487 9225
rect 10513 9199 10514 9225
rect 10486 9170 10514 9199
rect 10486 9137 10514 9142
rect 10598 9226 10626 9231
rect 10262 8919 10263 8945
rect 10289 8919 10290 8945
rect 10262 8913 10290 8919
rect 10598 8554 10626 9198
rect 10710 9114 10738 9119
rect 10710 9113 10906 9114
rect 10710 9087 10711 9113
rect 10737 9087 10906 9113
rect 10710 9086 10906 9087
rect 10710 9081 10738 9086
rect 10598 8521 10626 8526
rect 10878 8498 10906 9086
rect 10934 8610 10962 9479
rect 10990 9282 11018 9982
rect 11102 9562 11130 9567
rect 11102 9515 11130 9534
rect 11246 9422 11378 9427
rect 11274 9394 11298 9422
rect 11326 9394 11350 9422
rect 11246 9389 11378 9394
rect 10990 9249 11018 9254
rect 11246 8638 11378 8643
rect 11274 8610 11298 8638
rect 11326 8610 11350 8638
rect 10934 8582 11018 8610
rect 11246 8605 11378 8610
rect 10934 8498 10962 8503
rect 10878 8497 10962 8498
rect 10878 8471 10935 8497
rect 10961 8471 10962 8497
rect 10878 8470 10962 8471
rect 10934 8465 10962 8470
rect 10122 8414 10234 8442
rect 10822 8442 10850 8447
rect 10094 8409 10122 8414
rect 10822 8395 10850 8414
rect 9982 8297 10010 8302
rect 10038 8330 10066 8335
rect 10038 8329 10122 8330
rect 10038 8303 10039 8329
rect 10065 8303 10122 8329
rect 10038 8302 10122 8303
rect 10038 8297 10066 8302
rect 9916 8246 10048 8251
rect 9944 8218 9968 8246
rect 9996 8218 10020 8246
rect 9916 8213 10048 8218
rect 9590 8134 9842 8162
rect 9534 8105 9562 8111
rect 9534 8079 9535 8105
rect 9561 8079 9562 8105
rect 9534 8050 9562 8079
rect 9534 8017 9562 8022
rect 9590 8049 9618 8134
rect 9590 8023 9591 8049
rect 9617 8023 9618 8049
rect 9590 8017 9618 8023
rect 9758 8049 9786 8055
rect 9758 8023 9759 8049
rect 9785 8023 9786 8049
rect 9758 7770 9786 8023
rect 9814 7937 9842 8134
rect 9870 8162 9898 8167
rect 9898 8134 9954 8162
rect 9870 8129 9898 8134
rect 9870 8050 9898 8055
rect 9870 8003 9898 8022
rect 9814 7911 9815 7937
rect 9841 7911 9842 7937
rect 9814 7905 9842 7911
rect 9758 7737 9786 7742
rect 9870 7714 9898 7719
rect 9926 7714 9954 8134
rect 9982 8106 10010 8111
rect 10010 8078 10066 8106
rect 9982 8059 10010 8078
rect 9870 7713 9954 7714
rect 9870 7687 9871 7713
rect 9897 7687 9954 7713
rect 9870 7686 9954 7687
rect 9870 7681 9898 7686
rect 9702 7630 9842 7658
rect 9702 7601 9730 7630
rect 9702 7575 9703 7601
rect 9729 7575 9730 7601
rect 9702 7322 9730 7575
rect 9814 7602 9842 7630
rect 10038 7657 10066 8078
rect 10038 7631 10039 7657
rect 10065 7631 10066 7657
rect 10038 7625 10066 7631
rect 10094 7657 10122 8302
rect 10318 8106 10346 8111
rect 10206 8050 10234 8055
rect 10206 8003 10234 8022
rect 10318 7994 10346 8078
rect 10318 7993 10402 7994
rect 10318 7967 10319 7993
rect 10345 7967 10402 7993
rect 10318 7966 10402 7967
rect 10318 7961 10346 7966
rect 10262 7937 10290 7943
rect 10262 7911 10263 7937
rect 10289 7911 10290 7937
rect 10262 7714 10290 7911
rect 10374 7769 10402 7966
rect 10374 7743 10375 7769
rect 10401 7743 10402 7769
rect 10374 7737 10402 7743
rect 10318 7714 10346 7719
rect 10262 7713 10346 7714
rect 10262 7687 10319 7713
rect 10345 7687 10346 7713
rect 10262 7686 10346 7687
rect 10318 7681 10346 7686
rect 10430 7713 10458 7719
rect 10430 7687 10431 7713
rect 10457 7687 10458 7713
rect 10094 7631 10095 7657
rect 10121 7631 10122 7657
rect 10094 7625 10122 7631
rect 9926 7602 9954 7607
rect 9814 7601 9954 7602
rect 9814 7575 9927 7601
rect 9953 7575 9954 7601
rect 9814 7574 9954 7575
rect 10430 7574 10458 7687
rect 9926 7569 9954 7574
rect 9590 7294 9730 7322
rect 9758 7546 9786 7551
rect 9590 7210 9618 7294
rect 9758 7266 9786 7518
rect 10262 7546 10458 7574
rect 9916 7462 10048 7467
rect 9944 7434 9968 7462
rect 9996 7434 10020 7462
rect 9916 7429 10048 7434
rect 9814 7322 9842 7327
rect 9982 7322 10010 7327
rect 9814 7321 10010 7322
rect 9814 7295 9815 7321
rect 9841 7295 9983 7321
rect 10009 7295 10010 7321
rect 9814 7294 10010 7295
rect 9814 7289 9842 7294
rect 9982 7289 10010 7294
rect 9702 7238 9786 7266
rect 10150 7266 10178 7271
rect 10262 7266 10290 7546
rect 10150 7265 10290 7266
rect 10150 7239 10151 7265
rect 10177 7239 10290 7265
rect 10150 7238 10290 7239
rect 9590 7177 9618 7182
rect 9646 7209 9674 7215
rect 9646 7183 9647 7209
rect 9673 7183 9674 7209
rect 9478 7065 9506 7070
rect 9590 6986 9618 7005
rect 9646 6986 9674 7183
rect 9618 6958 9674 6986
rect 9590 6953 9618 6958
rect 9590 6874 9618 6879
rect 9422 6873 9506 6874
rect 9422 6847 9423 6873
rect 9449 6847 9506 6873
rect 9422 6846 9506 6847
rect 9422 6841 9450 6846
rect 9366 6734 9450 6762
rect 9254 6673 9282 6678
rect 8586 6286 8718 6291
rect 8614 6258 8638 6286
rect 8666 6258 8690 6286
rect 8586 6253 8718 6258
rect 9254 6090 9282 6095
rect 9282 6062 9338 6090
rect 9254 6057 9282 6062
rect 9198 5642 9226 5647
rect 8586 5502 8718 5507
rect 8614 5474 8638 5502
rect 8666 5474 8690 5502
rect 8586 5469 8718 5474
rect 7966 5391 7967 5417
rect 7993 5391 7994 5417
rect 7966 5385 7994 5391
rect 9198 5361 9226 5614
rect 9198 5335 9199 5361
rect 9225 5335 9226 5361
rect 7910 5306 7938 5311
rect 7910 5259 7938 5278
rect 9198 5306 9226 5335
rect 9198 5273 9226 5278
rect 7854 4937 7882 4942
rect 7966 5193 7994 5199
rect 7966 5167 7967 5193
rect 7993 5167 7994 5193
rect 7686 4887 7687 4913
rect 7713 4887 7714 4913
rect 7686 4881 7714 4887
rect 7966 4914 7994 5167
rect 7966 4881 7994 4886
rect 9254 5194 9282 5199
rect 6958 4858 6986 4863
rect 6958 4811 6986 4830
rect 7350 4857 7378 4863
rect 7350 4831 7351 4857
rect 7377 4831 7378 4857
rect 7350 4802 7378 4831
rect 7350 4769 7378 4774
rect 7462 4857 7490 4863
rect 7462 4831 7463 4857
rect 7489 4831 7490 4857
rect 5926 4718 6058 4723
rect 5954 4690 5978 4718
rect 6006 4690 6030 4718
rect 5926 4685 6058 4690
rect 5474 4550 5530 4578
rect 7350 4634 7378 4639
rect 7350 4577 7378 4606
rect 7406 4634 7434 4639
rect 7462 4634 7490 4831
rect 9254 4857 9282 5166
rect 9254 4831 9255 4857
rect 9281 4831 9282 4857
rect 9254 4825 9282 4831
rect 8586 4718 8718 4723
rect 8614 4690 8638 4718
rect 8666 4690 8690 4718
rect 8586 4685 8718 4690
rect 7406 4633 7490 4634
rect 7406 4607 7407 4633
rect 7433 4607 7490 4633
rect 7406 4606 7490 4607
rect 7406 4601 7434 4606
rect 7350 4551 7351 4577
rect 7377 4551 7378 4577
rect 5446 4531 5474 4550
rect 7350 4522 7378 4551
rect 7350 4494 7602 4522
rect 5110 4041 5138 4046
rect 5222 4382 5362 4410
rect 5390 4409 5418 4415
rect 5390 4383 5391 4409
rect 5417 4383 5418 4409
rect 5222 4073 5250 4382
rect 5334 4242 5362 4247
rect 5390 4242 5418 4383
rect 7256 4326 7388 4331
rect 7284 4298 7308 4326
rect 7336 4298 7360 4326
rect 7256 4293 7388 4298
rect 5362 4214 5418 4242
rect 5334 4209 5362 4214
rect 5670 4186 5698 4191
rect 5390 4185 5698 4186
rect 5390 4159 5671 4185
rect 5697 4159 5698 4185
rect 5390 4158 5698 4159
rect 5390 4129 5418 4158
rect 5670 4153 5698 4158
rect 5726 4186 5754 4191
rect 5390 4103 5391 4129
rect 5417 4103 5418 4129
rect 5390 4097 5418 4103
rect 5222 4047 5223 4073
rect 5249 4047 5250 4073
rect 5222 4041 5250 4047
rect 5614 4074 5642 4079
rect 5614 4027 5642 4046
rect 5726 4073 5754 4158
rect 7574 4185 7602 4494
rect 7574 4159 7575 4185
rect 7601 4159 7602 4185
rect 7574 4153 7602 4159
rect 5726 4047 5727 4073
rect 5753 4047 5754 4073
rect 5726 4041 5754 4047
rect 7406 4129 7434 4135
rect 7406 4103 7407 4129
rect 7433 4103 7434 4129
rect 5054 3929 5082 3934
rect 5334 4018 5362 4023
rect 4942 3823 4943 3849
rect 4969 3823 4970 3849
rect 4942 3817 4970 3823
rect 5054 3850 5082 3855
rect 5054 3803 5082 3822
rect 5222 3850 5250 3855
rect 2646 3794 2674 3799
rect 2646 3738 2674 3766
rect 5110 3794 5138 3799
rect 5110 3747 5138 3766
rect 5222 3793 5250 3822
rect 5222 3767 5223 3793
rect 5249 3767 5250 3793
rect 5222 3761 5250 3767
rect 2478 3737 2674 3738
rect 2478 3711 2647 3737
rect 2673 3711 2674 3737
rect 2478 3710 2674 3711
rect 2366 3626 2394 3710
rect 2646 3705 2674 3710
rect 2366 3593 2394 3598
rect 2870 3681 2898 3687
rect 2870 3655 2871 3681
rect 2897 3655 2898 3681
rect 2870 3626 2898 3655
rect 5334 3681 5362 3990
rect 5502 4017 5530 4023
rect 5502 3991 5503 4017
rect 5529 3991 5530 4017
rect 5502 3738 5530 3991
rect 7406 3962 7434 4103
rect 7686 4130 7714 4135
rect 7462 4074 7490 4079
rect 7462 4027 7490 4046
rect 5926 3934 6058 3939
rect 5954 3906 5978 3934
rect 6006 3906 6030 3934
rect 5926 3901 6058 3906
rect 7014 3934 7546 3962
rect 5502 3705 5530 3710
rect 5558 3794 5586 3799
rect 5334 3655 5335 3681
rect 5361 3655 5362 3681
rect 5334 3649 5362 3655
rect 2870 3593 2898 3598
rect 1936 3542 2068 3547
rect 1964 3514 1988 3542
rect 2016 3514 2040 3542
rect 1936 3509 2068 3514
rect 4596 3542 4728 3547
rect 4624 3514 4648 3542
rect 4676 3514 4700 3542
rect 4596 3509 4728 3514
rect 5558 3402 5586 3766
rect 7014 3793 7042 3934
rect 7182 3878 7490 3906
rect 7182 3849 7210 3878
rect 7182 3823 7183 3849
rect 7209 3823 7210 3849
rect 7182 3817 7210 3823
rect 7238 3822 7434 3850
rect 7014 3767 7015 3793
rect 7041 3767 7042 3793
rect 7014 3761 7042 3767
rect 7070 3793 7098 3799
rect 7070 3767 7071 3793
rect 7097 3767 7098 3793
rect 7070 3738 7098 3767
rect 7238 3738 7266 3822
rect 7406 3793 7434 3822
rect 7406 3767 7407 3793
rect 7433 3767 7434 3793
rect 7406 3761 7434 3767
rect 7462 3793 7490 3878
rect 7462 3767 7463 3793
rect 7489 3767 7490 3793
rect 7462 3761 7490 3767
rect 7070 3710 7266 3738
rect 7294 3738 7322 3743
rect 7182 3458 7210 3710
rect 7294 3691 7322 3710
rect 7462 3682 7490 3687
rect 7518 3682 7546 3934
rect 7686 3737 7714 4102
rect 9310 4074 9338 6062
rect 9366 5250 9394 5255
rect 9366 5203 9394 5222
rect 9366 4914 9394 4919
rect 9366 4867 9394 4886
rect 9422 4522 9450 6734
rect 9478 6426 9506 6846
rect 9590 6827 9618 6846
rect 9646 6706 9674 6711
rect 9478 5474 9506 6398
rect 9590 6594 9618 6599
rect 9478 5305 9506 5446
rect 9478 5279 9479 5305
rect 9505 5279 9506 5305
rect 9478 5273 9506 5279
rect 9534 6146 9562 6151
rect 9478 4522 9506 4527
rect 9422 4494 9478 4522
rect 9478 4489 9506 4494
rect 9310 4041 9338 4046
rect 9534 4130 9562 6118
rect 9590 6089 9618 6566
rect 9646 6593 9674 6678
rect 9646 6567 9647 6593
rect 9673 6567 9674 6593
rect 9646 6561 9674 6567
rect 9590 6063 9591 6089
rect 9617 6063 9618 6089
rect 9590 6057 9618 6063
rect 9646 5978 9674 5983
rect 9646 5698 9674 5950
rect 9702 5810 9730 7238
rect 10150 7233 10178 7238
rect 9758 7154 9786 7173
rect 9758 7121 9786 7126
rect 10038 7154 10066 7159
rect 10038 7107 10066 7126
rect 9758 7042 9786 7047
rect 9758 6873 9786 7014
rect 9982 6930 10010 6935
rect 9982 6883 10010 6902
rect 10262 6929 10290 7238
rect 10262 6903 10263 6929
rect 10289 6903 10290 6929
rect 9758 6847 9759 6873
rect 9785 6847 9786 6873
rect 9758 6841 9786 6847
rect 9814 6874 9842 6879
rect 9814 6827 9842 6846
rect 10206 6817 10234 6823
rect 10206 6791 10207 6817
rect 10233 6791 10234 6817
rect 10150 6761 10178 6767
rect 10150 6735 10151 6761
rect 10177 6735 10178 6761
rect 9916 6678 10048 6683
rect 9944 6650 9968 6678
rect 9996 6650 10020 6678
rect 9916 6645 10048 6650
rect 10150 6537 10178 6735
rect 10150 6511 10151 6537
rect 10177 6511 10178 6537
rect 10150 6505 10178 6511
rect 10206 6594 10234 6791
rect 9758 6482 9786 6487
rect 9758 6201 9786 6454
rect 9814 6481 9842 6487
rect 9814 6455 9815 6481
rect 9841 6455 9842 6481
rect 9814 6426 9842 6455
rect 10038 6482 10066 6487
rect 10038 6435 10066 6454
rect 10206 6481 10234 6566
rect 10206 6455 10207 6481
rect 10233 6455 10234 6481
rect 10206 6449 10234 6455
rect 9814 6393 9842 6398
rect 9758 6175 9759 6201
rect 9785 6175 9786 6201
rect 9758 6169 9786 6175
rect 9814 6146 9842 6151
rect 9814 6089 9842 6118
rect 9814 6063 9815 6089
rect 9841 6063 9842 6089
rect 9814 6057 9842 6063
rect 9982 6089 10010 6095
rect 9982 6063 9983 6089
rect 10009 6063 10010 6089
rect 9758 5978 9786 5983
rect 9982 5978 10010 6063
rect 9982 5950 10122 5978
rect 9758 5931 9786 5950
rect 9916 5894 10048 5899
rect 9944 5866 9968 5894
rect 9996 5866 10020 5894
rect 9916 5861 10048 5866
rect 10094 5866 10122 5950
rect 10094 5833 10122 5838
rect 10038 5810 10066 5815
rect 9702 5782 10010 5810
rect 9646 5670 9786 5698
rect 9646 5418 9674 5423
rect 9646 5417 9730 5418
rect 9646 5391 9647 5417
rect 9673 5391 9730 5417
rect 9646 5390 9730 5391
rect 9646 5385 9674 5390
rect 9646 5306 9674 5311
rect 9646 5259 9674 5278
rect 9702 5250 9730 5390
rect 9646 5194 9674 5199
rect 9590 5082 9618 5087
rect 9590 4746 9618 5054
rect 9646 4857 9674 5166
rect 9702 5082 9730 5222
rect 9758 5193 9786 5670
rect 9982 5697 10010 5782
rect 9982 5671 9983 5697
rect 10009 5671 10010 5697
rect 9870 5305 9898 5311
rect 9870 5279 9871 5305
rect 9897 5279 9898 5305
rect 9870 5194 9898 5279
rect 9982 5250 10010 5671
rect 10038 5361 10066 5782
rect 10150 5586 10178 5591
rect 10262 5586 10290 6903
rect 10934 6930 10962 6935
rect 10934 6883 10962 6902
rect 10822 6818 10850 6823
rect 10822 6771 10850 6790
rect 10934 5866 10962 5871
rect 10150 5585 10290 5586
rect 10150 5559 10151 5585
rect 10177 5559 10290 5585
rect 10150 5558 10290 5559
rect 10318 5586 10346 5591
rect 10038 5335 10039 5361
rect 10065 5335 10066 5361
rect 10038 5329 10066 5335
rect 10094 5362 10122 5367
rect 10150 5362 10178 5558
rect 10206 5474 10234 5479
rect 10206 5417 10234 5446
rect 10206 5391 10207 5417
rect 10233 5391 10234 5417
rect 10206 5385 10234 5391
rect 10122 5334 10178 5362
rect 10094 5329 10122 5334
rect 10318 5306 10346 5558
rect 10934 5417 10962 5838
rect 10990 5810 11018 8582
rect 11102 8442 11130 8447
rect 11102 8106 11130 8414
rect 11102 8073 11130 8078
rect 11246 7854 11378 7859
rect 11274 7826 11298 7854
rect 11326 7826 11350 7854
rect 11246 7821 11378 7826
rect 11246 7070 11378 7075
rect 11274 7042 11298 7070
rect 11326 7042 11350 7070
rect 11246 7037 11378 7042
rect 11102 6873 11130 6879
rect 11102 6847 11103 6873
rect 11129 6847 11130 6873
rect 11102 6818 11130 6847
rect 11102 6650 11130 6790
rect 11102 6617 11130 6622
rect 11246 6286 11378 6291
rect 11274 6258 11298 6286
rect 11326 6258 11350 6286
rect 11246 6253 11378 6258
rect 10990 5777 11018 5782
rect 11246 5502 11378 5507
rect 11274 5474 11298 5502
rect 11326 5474 11350 5502
rect 11246 5469 11378 5474
rect 10934 5391 10935 5417
rect 10961 5391 10962 5417
rect 10934 5385 10962 5391
rect 10150 5305 10346 5306
rect 10150 5279 10319 5305
rect 10345 5279 10346 5305
rect 10150 5278 10346 5279
rect 9982 5222 10066 5250
rect 9758 5167 9759 5193
rect 9785 5167 9786 5193
rect 9758 5161 9786 5167
rect 9814 5166 9898 5194
rect 10038 5194 10066 5222
rect 10038 5166 10122 5194
rect 9702 5054 9786 5082
rect 9758 5025 9786 5054
rect 9758 4999 9759 5025
rect 9785 4999 9786 5025
rect 9758 4993 9786 4999
rect 9702 4970 9730 4975
rect 9702 4923 9730 4942
rect 9646 4831 9647 4857
rect 9673 4831 9674 4857
rect 9646 4825 9674 4831
rect 9590 4718 9674 4746
rect 9646 4521 9674 4718
rect 9758 4578 9786 4583
rect 9646 4495 9647 4521
rect 9673 4495 9674 4521
rect 9534 4073 9562 4102
rect 9534 4047 9535 4073
rect 9561 4047 9562 4073
rect 9534 4041 9562 4047
rect 9590 4466 9618 4471
rect 7686 3711 7687 3737
rect 7713 3711 7714 3737
rect 7686 3705 7714 3711
rect 7910 4018 7938 4023
rect 7462 3681 7546 3682
rect 7462 3655 7463 3681
rect 7489 3655 7546 3681
rect 7462 3654 7546 3655
rect 7462 3649 7490 3654
rect 7256 3542 7388 3547
rect 7284 3514 7308 3542
rect 7336 3514 7360 3542
rect 7256 3509 7388 3514
rect 7350 3458 7378 3463
rect 7182 3457 7378 3458
rect 7182 3431 7351 3457
rect 7377 3431 7378 3457
rect 7182 3430 7378 3431
rect 7350 3425 7378 3430
rect 5558 3369 5586 3374
rect 7406 3402 7434 3407
rect 7406 3355 7434 3374
rect 7630 3402 7658 3407
rect 7630 3355 7658 3374
rect 7910 3402 7938 3990
rect 9366 4017 9394 4023
rect 9366 3991 9367 4017
rect 9393 3991 9394 4017
rect 8586 3934 8718 3939
rect 8614 3906 8638 3934
rect 8666 3906 8690 3934
rect 8586 3901 8718 3906
rect 9366 3794 9394 3991
rect 9366 3761 9394 3766
rect 9590 3626 9618 4438
rect 9646 4242 9674 4495
rect 9702 4577 9786 4578
rect 9702 4551 9759 4577
rect 9785 4551 9786 4577
rect 9702 4550 9786 4551
rect 9702 4522 9730 4550
rect 9758 4545 9786 4550
rect 9702 4489 9730 4494
rect 9758 4242 9786 4247
rect 9646 4241 9786 4242
rect 9646 4215 9759 4241
rect 9785 4215 9786 4241
rect 9646 4214 9786 4215
rect 9814 4242 9842 5166
rect 9916 5110 10048 5115
rect 9944 5082 9968 5110
rect 9996 5082 10020 5110
rect 9916 5077 10048 5082
rect 9926 4970 9954 4975
rect 9926 4923 9954 4942
rect 9982 4914 10010 4919
rect 10094 4914 10122 5166
rect 9982 4867 10010 4886
rect 10038 4913 10122 4914
rect 10038 4887 10095 4913
rect 10121 4887 10122 4913
rect 10038 4886 10122 4887
rect 10038 4802 10066 4886
rect 10094 4881 10122 4886
rect 9926 4774 10066 4802
rect 9926 4633 9954 4774
rect 9926 4607 9927 4633
rect 9953 4607 9954 4633
rect 9926 4601 9954 4607
rect 10038 4522 10066 4527
rect 10150 4522 10178 5278
rect 10318 5273 10346 5278
rect 11102 5305 11130 5311
rect 11102 5279 11103 5305
rect 11129 5279 11130 5305
rect 10822 5249 10850 5255
rect 10822 5223 10823 5249
rect 10849 5223 10850 5249
rect 10822 5194 10850 5223
rect 10822 5161 10850 5166
rect 11102 5194 11130 5279
rect 11102 5161 11130 5166
rect 11246 4718 11378 4723
rect 11274 4690 11298 4718
rect 11326 4690 11350 4718
rect 11246 4685 11378 4690
rect 10038 4521 10178 4522
rect 10038 4495 10039 4521
rect 10065 4495 10178 4521
rect 10038 4494 10178 4495
rect 10038 4489 10066 4494
rect 9916 4326 10048 4331
rect 9944 4298 9968 4326
rect 9996 4298 10020 4326
rect 9916 4293 10048 4298
rect 9814 4214 10066 4242
rect 9758 4209 9786 4214
rect 9926 4129 9954 4135
rect 9926 4103 9927 4129
rect 9953 4103 9954 4129
rect 9814 4073 9842 4079
rect 9814 4047 9815 4073
rect 9841 4047 9842 4073
rect 9814 3738 9842 4047
rect 9870 4074 9898 4079
rect 9926 4074 9954 4103
rect 9898 4046 9954 4074
rect 9870 4041 9898 4046
rect 10038 4017 10066 4214
rect 10150 4130 10178 4494
rect 10206 4130 10234 4135
rect 10150 4129 10234 4130
rect 10150 4103 10207 4129
rect 10233 4103 10234 4129
rect 10150 4102 10234 4103
rect 10206 4097 10234 4102
rect 10094 4074 10122 4079
rect 10094 4027 10122 4046
rect 10374 4073 10402 4079
rect 10374 4047 10375 4073
rect 10401 4047 10402 4073
rect 10038 3991 10039 4017
rect 10065 3991 10066 4017
rect 9982 3794 10010 3799
rect 10038 3794 10066 3991
rect 10010 3766 10066 3794
rect 10318 4018 10346 4023
rect 9982 3747 10010 3766
rect 9814 3705 9842 3710
rect 10150 3738 10178 3743
rect 10150 3691 10178 3710
rect 9590 3593 9618 3598
rect 9916 3542 10048 3547
rect 9944 3514 9968 3542
rect 9996 3514 10020 3542
rect 9916 3509 10048 3514
rect 7910 3369 7938 3374
rect 9814 3458 9842 3463
rect 3266 3150 3398 3155
rect 3294 3122 3318 3150
rect 3346 3122 3370 3150
rect 3266 3117 3398 3122
rect 5926 3150 6058 3155
rect 5954 3122 5978 3150
rect 6006 3122 6030 3150
rect 5926 3117 6058 3122
rect 8586 3150 8718 3155
rect 8614 3122 8638 3150
rect 8666 3122 8690 3150
rect 8586 3117 8718 3122
rect 1936 2758 2068 2763
rect 1964 2730 1988 2758
rect 2016 2730 2040 2758
rect 1936 2725 2068 2730
rect 4596 2758 4728 2763
rect 4624 2730 4648 2758
rect 4676 2730 4700 2758
rect 4596 2725 4728 2730
rect 7256 2758 7388 2763
rect 7284 2730 7308 2758
rect 7336 2730 7360 2758
rect 7256 2725 7388 2730
rect 3266 2366 3398 2371
rect 3294 2338 3318 2366
rect 3346 2338 3370 2366
rect 3266 2333 3398 2338
rect 5926 2366 6058 2371
rect 5954 2338 5978 2366
rect 6006 2338 6030 2366
rect 5926 2333 6058 2338
rect 8586 2366 8718 2371
rect 8614 2338 8638 2366
rect 8666 2338 8690 2366
rect 8586 2333 8718 2338
rect 1936 1974 2068 1979
rect 1964 1946 1988 1974
rect 2016 1946 2040 1974
rect 1936 1941 2068 1946
rect 4596 1974 4728 1979
rect 4624 1946 4648 1974
rect 4676 1946 4700 1974
rect 4596 1941 4728 1946
rect 7256 1974 7388 1979
rect 7284 1946 7308 1974
rect 7336 1946 7360 1974
rect 7256 1941 7388 1946
rect 3266 1582 3398 1587
rect 3294 1554 3318 1582
rect 3346 1554 3370 1582
rect 3266 1549 3398 1554
rect 5926 1582 6058 1587
rect 5954 1554 5978 1582
rect 6006 1554 6030 1582
rect 5926 1549 6058 1554
rect 8586 1582 8718 1587
rect 8614 1554 8638 1582
rect 8666 1554 8690 1582
rect 8586 1549 8718 1554
rect 9814 826 9842 3430
rect 10318 3458 10346 3990
rect 10374 3738 10402 4047
rect 10934 4074 10962 4079
rect 10934 4027 10962 4046
rect 11102 4073 11130 4079
rect 11102 4047 11103 4073
rect 11129 4047 11130 4073
rect 10766 4018 10794 4023
rect 10766 3971 10794 3990
rect 10374 3705 10402 3710
rect 10934 3738 10962 3743
rect 10318 3425 10346 3430
rect 9916 2758 10048 2763
rect 9944 2730 9968 2758
rect 9996 2730 10020 2758
rect 9916 2725 10048 2730
rect 10822 2562 10850 2567
rect 10822 2515 10850 2534
rect 10934 2505 10962 3710
rect 11102 3738 11130 4047
rect 11246 3934 11378 3939
rect 11274 3906 11298 3934
rect 11326 3906 11350 3934
rect 11246 3901 11378 3906
rect 11102 3691 11130 3710
rect 11246 3150 11378 3155
rect 11274 3122 11298 3150
rect 11326 3122 11350 3150
rect 11246 3117 11378 3122
rect 10934 2479 10935 2505
rect 10961 2479 10962 2505
rect 10934 2473 10962 2479
rect 11102 2562 11130 2567
rect 11102 2282 11130 2534
rect 11246 2366 11378 2371
rect 11274 2338 11298 2366
rect 11326 2338 11350 2366
rect 11246 2333 11378 2338
rect 11102 2249 11130 2254
rect 9916 1974 10048 1979
rect 9944 1946 9968 1974
rect 9996 1946 10020 1974
rect 9916 1941 10048 1946
rect 11246 1582 11378 1587
rect 11274 1554 11298 1582
rect 11326 1554 11350 1582
rect 11246 1549 11378 1554
rect 9814 793 9842 798
<< via2 >>
rect 3266 10205 3294 10206
rect 3266 10179 3267 10205
rect 3267 10179 3293 10205
rect 3293 10179 3294 10205
rect 3266 10178 3294 10179
rect 3318 10205 3346 10206
rect 3318 10179 3319 10205
rect 3319 10179 3345 10205
rect 3345 10179 3346 10205
rect 3318 10178 3346 10179
rect 3370 10205 3398 10206
rect 3370 10179 3371 10205
rect 3371 10179 3397 10205
rect 3397 10179 3398 10205
rect 3370 10178 3398 10179
rect 5926 10205 5954 10206
rect 5926 10179 5927 10205
rect 5927 10179 5953 10205
rect 5953 10179 5954 10205
rect 5926 10178 5954 10179
rect 5978 10205 6006 10206
rect 5978 10179 5979 10205
rect 5979 10179 6005 10205
rect 6005 10179 6006 10205
rect 5978 10178 6006 10179
rect 6030 10205 6058 10206
rect 6030 10179 6031 10205
rect 6031 10179 6057 10205
rect 6057 10179 6058 10205
rect 6030 10178 6058 10179
rect 8586 10205 8614 10206
rect 8586 10179 8587 10205
rect 8587 10179 8613 10205
rect 8613 10179 8614 10205
rect 8586 10178 8614 10179
rect 8638 10205 8666 10206
rect 8638 10179 8639 10205
rect 8639 10179 8665 10205
rect 8665 10179 8666 10205
rect 8638 10178 8666 10179
rect 8690 10205 8718 10206
rect 8690 10179 8691 10205
rect 8691 10179 8717 10205
rect 8717 10179 8718 10205
rect 8690 10178 8718 10179
rect 9870 10038 9898 10066
rect 10038 10990 10066 11018
rect 10374 10065 10402 10066
rect 10374 10039 10375 10065
rect 10375 10039 10401 10065
rect 10401 10039 10402 10065
rect 10374 10038 10402 10039
rect 11246 10205 11274 10206
rect 11246 10179 11247 10205
rect 11247 10179 11273 10205
rect 11273 10179 11274 10205
rect 11246 10178 11274 10179
rect 11298 10205 11326 10206
rect 11298 10179 11299 10205
rect 11299 10179 11325 10205
rect 11325 10179 11326 10205
rect 11298 10178 11326 10179
rect 11350 10205 11378 10206
rect 11350 10179 11351 10205
rect 11351 10179 11377 10205
rect 11377 10179 11378 10205
rect 11350 10178 11378 10179
rect 1936 9813 1964 9814
rect 1936 9787 1937 9813
rect 1937 9787 1963 9813
rect 1963 9787 1964 9813
rect 1936 9786 1964 9787
rect 1988 9813 2016 9814
rect 1988 9787 1989 9813
rect 1989 9787 2015 9813
rect 2015 9787 2016 9813
rect 1988 9786 2016 9787
rect 2040 9813 2068 9814
rect 2040 9787 2041 9813
rect 2041 9787 2067 9813
rect 2067 9787 2068 9813
rect 2040 9786 2068 9787
rect 1526 9225 1554 9226
rect 1526 9199 1527 9225
rect 1527 9199 1553 9225
rect 1553 9199 1554 9225
rect 1526 9198 1554 9199
rect 2086 9254 2114 9282
rect 1806 9225 1834 9226
rect 1806 9199 1807 9225
rect 1807 9199 1833 9225
rect 1833 9199 1834 9225
rect 1806 9198 1834 9199
rect 1638 9142 1666 9170
rect 2142 9225 2170 9226
rect 2142 9199 2143 9225
rect 2143 9199 2169 9225
rect 2169 9199 2170 9225
rect 2142 9198 2170 9199
rect 2310 9310 2338 9338
rect 2534 9561 2562 9562
rect 2534 9535 2535 9561
rect 2535 9535 2561 9561
rect 2561 9535 2562 9561
rect 2534 9534 2562 9535
rect 3266 9421 3294 9422
rect 3266 9395 3267 9421
rect 3267 9395 3293 9421
rect 3293 9395 3294 9421
rect 3266 9394 3294 9395
rect 3318 9421 3346 9422
rect 3318 9395 3319 9421
rect 3319 9395 3345 9421
rect 3345 9395 3346 9421
rect 3318 9394 3346 9395
rect 3370 9421 3398 9422
rect 3370 9395 3371 9421
rect 3371 9395 3397 9421
rect 3397 9395 3398 9421
rect 3370 9394 3398 9395
rect 2422 9337 2450 9338
rect 2422 9311 2423 9337
rect 2423 9311 2449 9337
rect 2449 9311 2450 9337
rect 2422 9310 2450 9311
rect 2478 9169 2506 9170
rect 2478 9143 2479 9169
rect 2479 9143 2505 9169
rect 2505 9143 2506 9169
rect 2478 9142 2506 9143
rect 1936 9029 1964 9030
rect 1936 9003 1937 9029
rect 1937 9003 1963 9029
rect 1963 9003 1964 9029
rect 1936 9002 1964 9003
rect 1988 9029 2016 9030
rect 1988 9003 1989 9029
rect 1989 9003 2015 9029
rect 2015 9003 2016 9029
rect 1988 9002 2016 9003
rect 2040 9029 2068 9030
rect 2040 9003 2041 9029
rect 2041 9003 2067 9029
rect 2067 9003 2068 9029
rect 2040 9002 2068 9003
rect 1526 7966 1554 7994
rect 1246 7910 1274 7938
rect 1694 7993 1722 7994
rect 1694 7967 1695 7993
rect 1695 7967 1721 7993
rect 1721 7967 1722 7993
rect 1694 7966 1722 7967
rect 2926 9281 2954 9282
rect 2926 9255 2927 9281
rect 2927 9255 2953 9281
rect 2953 9255 2954 9281
rect 2926 9254 2954 9255
rect 2870 9198 2898 9226
rect 3150 9169 3178 9170
rect 3150 9143 3151 9169
rect 3151 9143 3177 9169
rect 3177 9143 3178 9169
rect 3150 9142 3178 9143
rect 2646 8862 2674 8890
rect 2086 8777 2114 8778
rect 2086 8751 2087 8777
rect 2087 8751 2113 8777
rect 2113 8751 2114 8777
rect 2086 8750 2114 8751
rect 3094 8750 3122 8778
rect 2982 8694 3010 8722
rect 3266 8637 3294 8638
rect 3266 8611 3267 8637
rect 3267 8611 3293 8637
rect 3293 8611 3294 8637
rect 3266 8610 3294 8611
rect 3318 8637 3346 8638
rect 3318 8611 3319 8637
rect 3319 8611 3345 8637
rect 3345 8611 3346 8637
rect 3318 8610 3346 8611
rect 3370 8637 3398 8638
rect 3370 8611 3371 8637
rect 3371 8611 3397 8637
rect 3397 8611 3398 8637
rect 3370 8610 3398 8611
rect 2534 8358 2562 8386
rect 1936 8245 1964 8246
rect 1936 8219 1937 8245
rect 1937 8219 1963 8245
rect 1963 8219 1964 8245
rect 1936 8218 1964 8219
rect 1988 8245 2016 8246
rect 1988 8219 1989 8245
rect 1989 8219 2015 8245
rect 2015 8219 2016 8245
rect 1988 8218 2016 8219
rect 2040 8245 2068 8246
rect 2040 8219 2041 8245
rect 2041 8219 2067 8245
rect 2067 8219 2068 8245
rect 2040 8218 2068 8219
rect 1918 7993 1946 7994
rect 1918 7967 1919 7993
rect 1919 7967 1945 7993
rect 1945 7967 1946 7993
rect 1918 7966 1946 7967
rect 1190 7601 1218 7602
rect 1190 7575 1191 7601
rect 1191 7575 1217 7601
rect 1217 7575 1218 7601
rect 1190 7574 1218 7575
rect 1134 7350 1162 7378
rect 1638 7601 1666 7602
rect 1638 7575 1639 7601
rect 1639 7575 1665 7601
rect 1665 7575 1666 7601
rect 1638 7574 1666 7575
rect 1470 7350 1498 7378
rect 1974 7937 2002 7938
rect 1974 7911 1975 7937
rect 1975 7911 2001 7937
rect 2001 7911 2002 7937
rect 1974 7910 2002 7911
rect 2142 7742 2170 7770
rect 1974 7574 2002 7602
rect 2086 7601 2114 7602
rect 2086 7575 2087 7601
rect 2087 7575 2113 7601
rect 2113 7575 2114 7601
rect 2086 7574 2114 7575
rect 1936 7461 1964 7462
rect 1936 7435 1937 7461
rect 1937 7435 1963 7461
rect 1963 7435 1964 7461
rect 1936 7434 1964 7435
rect 1988 7461 2016 7462
rect 1988 7435 1989 7461
rect 1989 7435 2015 7461
rect 2015 7435 2016 7461
rect 1988 7434 2016 7435
rect 2040 7461 2068 7462
rect 2040 7435 2041 7461
rect 2041 7435 2067 7461
rect 2067 7435 2068 7461
rect 2040 7434 2068 7435
rect 2310 7574 2338 7602
rect 2198 7377 2226 7378
rect 2198 7351 2199 7377
rect 2199 7351 2225 7377
rect 2225 7351 2226 7377
rect 2198 7350 2226 7351
rect 2254 7209 2282 7210
rect 2254 7183 2255 7209
rect 2255 7183 2281 7209
rect 2281 7183 2282 7209
rect 2254 7182 2282 7183
rect 2198 7153 2226 7154
rect 2198 7127 2199 7153
rect 2199 7127 2225 7153
rect 2225 7127 2226 7153
rect 2198 7126 2226 7127
rect 1806 6761 1834 6762
rect 1806 6735 1807 6761
rect 1807 6735 1833 6761
rect 1833 6735 1834 6761
rect 1806 6734 1834 6735
rect 1936 6677 1964 6678
rect 1936 6651 1937 6677
rect 1937 6651 1963 6677
rect 1963 6651 1964 6677
rect 1936 6650 1964 6651
rect 1988 6677 2016 6678
rect 1988 6651 1989 6677
rect 1989 6651 2015 6677
rect 2015 6651 2016 6677
rect 1988 6650 2016 6651
rect 2040 6677 2068 6678
rect 2040 6651 2041 6677
rect 2041 6651 2067 6677
rect 2067 6651 2068 6677
rect 2040 6650 2068 6651
rect 2198 6174 2226 6202
rect 2478 7574 2506 7602
rect 3206 8358 3234 8386
rect 3266 7853 3294 7854
rect 3266 7827 3267 7853
rect 3267 7827 3293 7853
rect 3293 7827 3294 7853
rect 3266 7826 3294 7827
rect 3318 7853 3346 7854
rect 3318 7827 3319 7853
rect 3319 7827 3345 7853
rect 3345 7827 3346 7853
rect 3318 7826 3346 7827
rect 3370 7853 3398 7854
rect 3370 7827 3371 7853
rect 3371 7827 3397 7853
rect 3397 7827 3398 7853
rect 3370 7826 3398 7827
rect 2030 6033 2058 6034
rect 2030 6007 2031 6033
rect 2031 6007 2057 6033
rect 2057 6007 2058 6033
rect 2030 6006 2058 6007
rect 1936 5893 1964 5894
rect 1936 5867 1937 5893
rect 1937 5867 1963 5893
rect 1963 5867 1964 5893
rect 1936 5866 1964 5867
rect 1988 5893 2016 5894
rect 1988 5867 1989 5893
rect 1989 5867 2015 5893
rect 2015 5867 2016 5893
rect 1988 5866 2016 5867
rect 2040 5893 2068 5894
rect 2040 5867 2041 5893
rect 2041 5867 2067 5893
rect 2067 5867 2068 5893
rect 2040 5866 2068 5867
rect 2366 5697 2394 5698
rect 2366 5671 2367 5697
rect 2367 5671 2393 5697
rect 2393 5671 2394 5697
rect 2366 5670 2394 5671
rect 2814 7182 2842 7210
rect 3266 7069 3294 7070
rect 3266 7043 3267 7069
rect 3267 7043 3293 7069
rect 3293 7043 3294 7069
rect 3266 7042 3294 7043
rect 3318 7069 3346 7070
rect 3318 7043 3319 7069
rect 3319 7043 3345 7069
rect 3345 7043 3346 7069
rect 3318 7042 3346 7043
rect 3370 7069 3398 7070
rect 3370 7043 3371 7069
rect 3371 7043 3397 7069
rect 3397 7043 3398 7069
rect 3370 7042 3398 7043
rect 3150 6174 3178 6202
rect 3266 6285 3294 6286
rect 3266 6259 3267 6285
rect 3267 6259 3293 6285
rect 3293 6259 3294 6285
rect 3266 6258 3294 6259
rect 3318 6285 3346 6286
rect 3318 6259 3319 6285
rect 3319 6259 3345 6285
rect 3345 6259 3346 6285
rect 3318 6258 3346 6259
rect 3370 6285 3398 6286
rect 3370 6259 3371 6285
rect 3371 6259 3397 6285
rect 3397 6259 3398 6285
rect 3370 6258 3398 6259
rect 2702 6006 2730 6034
rect 1134 5278 1162 5306
rect 1638 5305 1666 5306
rect 1638 5279 1639 5305
rect 1639 5279 1665 5305
rect 1665 5279 1666 5305
rect 1638 5278 1666 5279
rect 1302 4998 1330 5026
rect 1936 5109 1964 5110
rect 1936 5083 1937 5109
rect 1937 5083 1963 5109
rect 1963 5083 1964 5109
rect 1936 5082 1964 5083
rect 1988 5109 2016 5110
rect 1988 5083 1989 5109
rect 1989 5083 2015 5109
rect 2015 5083 2016 5109
rect 1988 5082 2016 5083
rect 2040 5109 2068 5110
rect 2040 5083 2041 5109
rect 2041 5083 2067 5109
rect 2067 5083 2068 5109
rect 2040 5082 2068 5083
rect 2142 4913 2170 4914
rect 2142 4887 2143 4913
rect 2143 4887 2169 4913
rect 2169 4887 2170 4913
rect 2142 4886 2170 4887
rect 1694 4494 1722 4522
rect 1582 4129 1610 4130
rect 1582 4103 1583 4129
rect 1583 4103 1609 4129
rect 1609 4103 1610 4129
rect 1582 4102 1610 4103
rect 1918 4521 1946 4522
rect 1918 4495 1919 4521
rect 1919 4495 1945 4521
rect 1945 4495 1946 4521
rect 1918 4494 1946 4495
rect 1936 4325 1964 4326
rect 1936 4299 1937 4325
rect 1937 4299 1963 4325
rect 1963 4299 1964 4325
rect 1936 4298 1964 4299
rect 1988 4325 2016 4326
rect 1988 4299 1989 4325
rect 1989 4299 2015 4325
rect 2015 4299 2016 4325
rect 1988 4298 2016 4299
rect 2040 4325 2068 4326
rect 2040 4299 2041 4325
rect 2041 4299 2067 4325
rect 2067 4299 2068 4325
rect 2040 4298 2068 4299
rect 2142 4158 2170 4186
rect 1918 4129 1946 4130
rect 1918 4103 1919 4129
rect 1919 4103 1945 4129
rect 1945 4103 1946 4129
rect 1918 4102 1946 4103
rect 2086 3990 2114 4018
rect 2478 4521 2506 4522
rect 2478 4495 2479 4521
rect 2479 4495 2505 4521
rect 2505 4495 2506 4521
rect 2478 4494 2506 4495
rect 2422 3990 2450 4018
rect 2870 4185 2898 4186
rect 2870 4159 2871 4185
rect 2871 4159 2897 4185
rect 2897 4159 2898 4185
rect 2870 4158 2898 4159
rect 3266 5501 3294 5502
rect 3266 5475 3267 5501
rect 3267 5475 3293 5501
rect 3293 5475 3294 5501
rect 3266 5474 3294 5475
rect 3318 5501 3346 5502
rect 3318 5475 3319 5501
rect 3319 5475 3345 5501
rect 3345 5475 3346 5501
rect 3318 5474 3346 5475
rect 3370 5501 3398 5502
rect 3370 5475 3371 5501
rect 3371 5475 3397 5501
rect 3397 5475 3398 5501
rect 3370 5474 3398 5475
rect 3266 4717 3294 4718
rect 3266 4691 3267 4717
rect 3267 4691 3293 4717
rect 3293 4691 3294 4717
rect 3266 4690 3294 4691
rect 3318 4717 3346 4718
rect 3318 4691 3319 4717
rect 3319 4691 3345 4717
rect 3345 4691 3346 4717
rect 3318 4690 3346 4691
rect 3370 4717 3398 4718
rect 3370 4691 3371 4717
rect 3371 4691 3397 4717
rect 3397 4691 3398 4717
rect 3370 4690 3398 4691
rect 4596 9813 4624 9814
rect 4596 9787 4597 9813
rect 4597 9787 4623 9813
rect 4623 9787 4624 9813
rect 4596 9786 4624 9787
rect 4648 9813 4676 9814
rect 4648 9787 4649 9813
rect 4649 9787 4675 9813
rect 4675 9787 4676 9813
rect 4648 9786 4676 9787
rect 4700 9813 4728 9814
rect 4700 9787 4701 9813
rect 4701 9787 4727 9813
rect 4727 9787 4728 9813
rect 4700 9786 4728 9787
rect 3878 9561 3906 9562
rect 3878 9535 3879 9561
rect 3879 9535 3905 9561
rect 3905 9535 3906 9561
rect 3878 9534 3906 9535
rect 3990 9534 4018 9562
rect 3934 9310 3962 9338
rect 4326 9281 4354 9282
rect 4326 9255 4327 9281
rect 4327 9255 4353 9281
rect 4353 9255 4354 9281
rect 4326 9254 4354 9255
rect 4158 9198 4186 9226
rect 4102 9169 4130 9170
rect 4102 9143 4103 9169
rect 4103 9143 4129 9169
rect 4129 9143 4130 9169
rect 4102 9142 4130 9143
rect 3878 8750 3906 8778
rect 3822 7377 3850 7378
rect 3822 7351 3823 7377
rect 3823 7351 3849 7377
rect 3849 7351 3850 7377
rect 3822 7350 3850 7351
rect 3766 7209 3794 7210
rect 3766 7183 3767 7209
rect 3767 7183 3793 7209
rect 3793 7183 3794 7209
rect 3766 7182 3794 7183
rect 3822 6174 3850 6202
rect 3990 8833 4018 8834
rect 3990 8807 3991 8833
rect 3991 8807 4017 8833
rect 4017 8807 4018 8833
rect 3990 8806 4018 8807
rect 3990 8721 4018 8722
rect 3990 8695 3991 8721
rect 3991 8695 4017 8721
rect 4017 8695 4018 8721
rect 3990 8694 4018 8695
rect 4270 9113 4298 9114
rect 4270 9087 4271 9113
rect 4271 9087 4297 9113
rect 4297 9087 4298 9113
rect 4270 9086 4298 9087
rect 4774 9086 4802 9114
rect 4596 9029 4624 9030
rect 4596 9003 4597 9029
rect 4597 9003 4623 9029
rect 4623 9003 4624 9029
rect 4596 9002 4624 9003
rect 4648 9029 4676 9030
rect 4648 9003 4649 9029
rect 4649 9003 4675 9029
rect 4675 9003 4676 9029
rect 4648 9002 4676 9003
rect 4700 9029 4728 9030
rect 4700 9003 4701 9029
rect 4701 9003 4727 9029
rect 4727 9003 4728 9029
rect 4700 9002 4728 9003
rect 4158 7910 4186 7938
rect 3934 7406 3962 7434
rect 4046 7294 4074 7322
rect 4596 8245 4624 8246
rect 4596 8219 4597 8245
rect 4597 8219 4623 8245
rect 4623 8219 4624 8245
rect 4596 8218 4624 8219
rect 4648 8245 4676 8246
rect 4648 8219 4649 8245
rect 4649 8219 4675 8245
rect 4675 8219 4676 8245
rect 4648 8218 4676 8219
rect 4700 8245 4728 8246
rect 4700 8219 4701 8245
rect 4701 8219 4727 8245
rect 4727 8219 4728 8245
rect 4700 8218 4728 8219
rect 4550 7937 4578 7938
rect 4550 7911 4551 7937
rect 4551 7911 4577 7937
rect 4577 7911 4578 7937
rect 4550 7910 4578 7911
rect 4326 7630 4354 7658
rect 4382 7574 4410 7602
rect 4214 7406 4242 7434
rect 4270 7377 4298 7378
rect 4270 7351 4271 7377
rect 4271 7351 4297 7377
rect 4297 7351 4298 7377
rect 4270 7350 4298 7351
rect 7518 9982 7546 10010
rect 7256 9813 7284 9814
rect 7256 9787 7257 9813
rect 7257 9787 7283 9813
rect 7283 9787 7284 9813
rect 7256 9786 7284 9787
rect 7308 9813 7336 9814
rect 7308 9787 7309 9813
rect 7309 9787 7335 9813
rect 7335 9787 7336 9813
rect 7308 9786 7336 9787
rect 7360 9813 7388 9814
rect 7360 9787 7361 9813
rect 7361 9787 7387 9813
rect 7387 9787 7388 9813
rect 7360 9786 7388 9787
rect 6790 9702 6818 9730
rect 5926 9421 5954 9422
rect 5926 9395 5927 9421
rect 5927 9395 5953 9421
rect 5953 9395 5954 9421
rect 5926 9394 5954 9395
rect 5978 9421 6006 9422
rect 5978 9395 5979 9421
rect 5979 9395 6005 9421
rect 6005 9395 6006 9421
rect 5978 9394 6006 9395
rect 6030 9421 6058 9422
rect 6030 9395 6031 9421
rect 6031 9395 6057 9421
rect 6057 9395 6058 9421
rect 6030 9394 6058 9395
rect 5558 9254 5586 9282
rect 6062 9254 6090 9282
rect 5614 9198 5642 9226
rect 4830 7742 4858 7770
rect 4942 8918 4970 8946
rect 4718 7518 4746 7546
rect 4774 7630 4802 7658
rect 4596 7461 4624 7462
rect 4596 7435 4597 7461
rect 4597 7435 4623 7461
rect 4623 7435 4624 7461
rect 4596 7434 4624 7435
rect 4648 7461 4676 7462
rect 4648 7435 4649 7461
rect 4649 7435 4675 7461
rect 4675 7435 4676 7461
rect 4648 7434 4676 7435
rect 4700 7461 4728 7462
rect 4700 7435 4701 7461
rect 4701 7435 4727 7461
rect 4727 7435 4728 7461
rect 4700 7434 4728 7435
rect 4494 7294 4522 7322
rect 3934 7070 3962 7098
rect 4596 6677 4624 6678
rect 4596 6651 4597 6677
rect 4597 6651 4623 6677
rect 4623 6651 4624 6677
rect 4596 6650 4624 6651
rect 4648 6677 4676 6678
rect 4648 6651 4649 6677
rect 4649 6651 4675 6677
rect 4675 6651 4676 6677
rect 4648 6650 4676 6651
rect 4700 6677 4728 6678
rect 4700 6651 4701 6677
rect 4701 6651 4727 6677
rect 4727 6651 4728 6677
rect 4700 6650 4728 6651
rect 3934 6145 3962 6146
rect 3934 6119 3935 6145
rect 3935 6119 3961 6145
rect 3961 6119 3962 6145
rect 3934 6118 3962 6119
rect 5110 9030 5138 9058
rect 4830 7350 4858 7378
rect 4998 7601 5026 7602
rect 4998 7575 4999 7601
rect 4999 7575 5025 7601
rect 5025 7575 5026 7601
rect 4998 7574 5026 7575
rect 4942 7518 4970 7546
rect 4942 7350 4970 7378
rect 4998 7294 5026 7322
rect 6342 9281 6370 9282
rect 6342 9255 6343 9281
rect 6343 9255 6369 9281
rect 6369 9255 6370 9281
rect 6342 9254 6370 9255
rect 6286 9225 6314 9226
rect 6286 9199 6287 9225
rect 6287 9199 6313 9225
rect 6313 9199 6314 9225
rect 6286 9198 6314 9199
rect 5950 9142 5978 9170
rect 5670 9030 5698 9058
rect 5782 9030 5810 9058
rect 5446 8945 5474 8946
rect 5446 8919 5447 8945
rect 5447 8919 5473 8945
rect 5473 8919 5474 8945
rect 5446 8918 5474 8919
rect 5502 8889 5530 8890
rect 5502 8863 5503 8889
rect 5503 8863 5529 8889
rect 5529 8863 5530 8889
rect 5502 8862 5530 8863
rect 5670 8945 5698 8946
rect 5670 8919 5671 8945
rect 5671 8919 5697 8945
rect 5697 8919 5698 8945
rect 5670 8918 5698 8919
rect 5614 8414 5642 8442
rect 6174 9142 6202 9170
rect 5950 8889 5978 8890
rect 5950 8863 5951 8889
rect 5951 8863 5977 8889
rect 5977 8863 5978 8889
rect 5950 8862 5978 8863
rect 6230 8694 6258 8722
rect 5926 8637 5954 8638
rect 5926 8611 5927 8637
rect 5927 8611 5953 8637
rect 5953 8611 5954 8637
rect 5926 8610 5954 8611
rect 5978 8637 6006 8638
rect 5978 8611 5979 8637
rect 5979 8611 6005 8637
rect 6005 8611 6006 8637
rect 5978 8610 6006 8611
rect 6030 8637 6058 8638
rect 6030 8611 6031 8637
rect 6031 8611 6057 8637
rect 6057 8611 6058 8637
rect 6030 8610 6058 8611
rect 6174 8414 6202 8442
rect 5926 7853 5954 7854
rect 5926 7827 5927 7853
rect 5927 7827 5953 7853
rect 5953 7827 5954 7853
rect 5926 7826 5954 7827
rect 5978 7853 6006 7854
rect 5978 7827 5979 7853
rect 5979 7827 6005 7853
rect 6005 7827 6006 7853
rect 5978 7826 6006 7827
rect 6030 7853 6058 7854
rect 6030 7827 6031 7853
rect 6031 7827 6057 7853
rect 6057 7827 6058 7853
rect 6030 7826 6058 7827
rect 5390 7294 5418 7322
rect 5222 7182 5250 7210
rect 5670 7182 5698 7210
rect 5614 7070 5642 7098
rect 5614 6958 5642 6986
rect 5502 6873 5530 6874
rect 5502 6847 5503 6873
rect 5503 6847 5529 6873
rect 5529 6847 5530 6873
rect 5502 6846 5530 6847
rect 5894 7574 5922 7602
rect 5782 7377 5810 7378
rect 5782 7351 5783 7377
rect 5783 7351 5809 7377
rect 5809 7351 5810 7377
rect 5782 7350 5810 7351
rect 6118 7574 6146 7602
rect 6230 7657 6258 7658
rect 6230 7631 6231 7657
rect 6231 7631 6257 7657
rect 6257 7631 6258 7657
rect 6230 7630 6258 7631
rect 6062 7294 6090 7322
rect 5894 7265 5922 7266
rect 5894 7239 5895 7265
rect 5895 7239 5921 7265
rect 5921 7239 5922 7265
rect 5894 7238 5922 7239
rect 6118 7153 6146 7154
rect 6118 7127 6119 7153
rect 6119 7127 6145 7153
rect 6145 7127 6146 7153
rect 6118 7126 6146 7127
rect 5926 7069 5954 7070
rect 5926 7043 5927 7069
rect 5927 7043 5953 7069
rect 5953 7043 5954 7069
rect 5926 7042 5954 7043
rect 5978 7069 6006 7070
rect 5978 7043 5979 7069
rect 5979 7043 6005 7069
rect 6005 7043 6006 7069
rect 5978 7042 6006 7043
rect 6030 7069 6058 7070
rect 6030 7043 6031 7069
rect 6031 7043 6057 7069
rect 6057 7043 6058 7069
rect 6030 7042 6058 7043
rect 5726 6902 5754 6930
rect 4942 6817 4970 6818
rect 4942 6791 4943 6817
rect 4943 6791 4969 6817
rect 4969 6791 4970 6817
rect 4942 6790 4970 6791
rect 4382 6369 4410 6370
rect 4382 6343 4383 6369
rect 4383 6343 4409 6369
rect 4409 6343 4410 6369
rect 4382 6342 4410 6343
rect 4102 5278 4130 5306
rect 4382 6062 4410 6090
rect 4438 5726 4466 5754
rect 4830 6734 4858 6762
rect 4662 6342 4690 6370
rect 5838 6790 5866 6818
rect 4942 6174 4970 6202
rect 5110 6118 5138 6146
rect 4596 5893 4624 5894
rect 4596 5867 4597 5893
rect 4597 5867 4623 5893
rect 4623 5867 4624 5893
rect 4596 5866 4624 5867
rect 4648 5893 4676 5894
rect 4648 5867 4649 5893
rect 4649 5867 4675 5893
rect 4675 5867 4676 5893
rect 4648 5866 4676 5867
rect 4700 5893 4728 5894
rect 4700 5867 4701 5893
rect 4701 5867 4727 5893
rect 4727 5867 4728 5893
rect 4700 5866 4728 5867
rect 5054 6089 5082 6090
rect 5054 6063 5055 6089
rect 5055 6063 5081 6089
rect 5081 6063 5082 6089
rect 5054 6062 5082 6063
rect 4942 5726 4970 5754
rect 4606 5670 4634 5698
rect 4550 5641 4578 5642
rect 4550 5615 4551 5641
rect 4551 5615 4577 5641
rect 4577 5615 4578 5641
rect 4550 5614 4578 5615
rect 4550 5334 4578 5362
rect 4214 4942 4242 4970
rect 4270 5278 4298 5306
rect 4886 5697 4914 5698
rect 4886 5671 4887 5697
rect 4887 5671 4913 5697
rect 4913 5671 4914 5697
rect 4886 5670 4914 5671
rect 4596 5109 4624 5110
rect 4596 5083 4597 5109
rect 4597 5083 4623 5109
rect 4623 5083 4624 5109
rect 4596 5082 4624 5083
rect 4648 5109 4676 5110
rect 4648 5083 4649 5109
rect 4649 5083 4675 5109
rect 4675 5083 4676 5109
rect 4648 5082 4676 5083
rect 4700 5109 4728 5110
rect 4700 5083 4701 5109
rect 4701 5083 4727 5109
rect 4727 5083 4728 5109
rect 4700 5082 4728 5083
rect 4606 4969 4634 4970
rect 4606 4943 4607 4969
rect 4607 4943 4633 4969
rect 4633 4943 4634 4969
rect 4606 4942 4634 4943
rect 4326 4606 4354 4634
rect 4550 4830 4578 4858
rect 3430 4494 3458 4522
rect 3206 4158 3234 4186
rect 3710 4158 3738 4186
rect 2702 4102 2730 4130
rect 2814 4017 2842 4018
rect 2814 3991 2815 4017
rect 2815 3991 2841 4017
rect 2841 3991 2842 4017
rect 2814 3990 2842 3991
rect 3654 4129 3682 4130
rect 3654 4103 3655 4129
rect 3655 4103 3681 4129
rect 3681 4103 3682 4129
rect 3654 4102 3682 4103
rect 3150 4073 3178 4074
rect 3150 4047 3151 4073
rect 3151 4047 3177 4073
rect 3177 4047 3178 4073
rect 3150 4046 3178 4047
rect 2982 3990 3010 4018
rect 4438 4185 4466 4186
rect 4438 4159 4439 4185
rect 4439 4159 4465 4185
rect 4465 4159 4466 4185
rect 4438 4158 4466 4159
rect 4774 4801 4802 4802
rect 4774 4775 4775 4801
rect 4775 4775 4801 4801
rect 4801 4775 4802 4801
rect 4774 4774 4802 4775
rect 5110 5726 5138 5754
rect 5222 5697 5250 5698
rect 5222 5671 5223 5697
rect 5223 5671 5249 5697
rect 5249 5671 5250 5697
rect 5222 5670 5250 5671
rect 4998 5614 5026 5642
rect 4942 4913 4970 4914
rect 4942 4887 4943 4913
rect 4943 4887 4969 4913
rect 4969 4887 4970 4913
rect 4942 4886 4970 4887
rect 4596 4325 4624 4326
rect 4596 4299 4597 4325
rect 4597 4299 4623 4325
rect 4623 4299 4624 4325
rect 4596 4298 4624 4299
rect 4648 4325 4676 4326
rect 4648 4299 4649 4325
rect 4649 4299 4675 4325
rect 4675 4299 4676 4325
rect 4648 4298 4676 4299
rect 4700 4325 4728 4326
rect 4700 4299 4701 4325
rect 4701 4299 4727 4325
rect 4727 4299 4728 4325
rect 4700 4298 4728 4299
rect 5390 4886 5418 4914
rect 5166 4857 5194 4858
rect 5166 4831 5167 4857
rect 5167 4831 5193 4857
rect 5193 4831 5194 4857
rect 5166 4830 5194 4831
rect 5278 4774 5306 4802
rect 5222 4550 5250 4578
rect 4662 4214 4690 4242
rect 3822 4129 3850 4130
rect 3822 4103 3823 4129
rect 3823 4103 3849 4129
rect 3849 4103 3850 4129
rect 3822 4102 3850 4103
rect 3266 3933 3294 3934
rect 3266 3907 3267 3933
rect 3267 3907 3293 3933
rect 3293 3907 3294 3933
rect 3266 3906 3294 3907
rect 3318 3933 3346 3934
rect 3318 3907 3319 3933
rect 3319 3907 3345 3933
rect 3345 3907 3346 3933
rect 3318 3906 3346 3907
rect 3370 3933 3398 3934
rect 3370 3907 3371 3933
rect 3371 3907 3397 3933
rect 3397 3907 3398 3933
rect 3370 3906 3398 3907
rect 5054 4158 5082 4186
rect 4830 4046 4858 4074
rect 4886 3934 4914 3962
rect 4438 3822 4466 3850
rect 4998 4129 5026 4130
rect 4998 4103 4999 4129
rect 4999 4103 5025 4129
rect 5025 4103 5026 4129
rect 4998 4102 5026 4103
rect 5926 6285 5954 6286
rect 5926 6259 5927 6285
rect 5927 6259 5953 6285
rect 5953 6259 5954 6285
rect 5926 6258 5954 6259
rect 5978 6285 6006 6286
rect 5978 6259 5979 6285
rect 5979 6259 6005 6285
rect 6005 6259 6006 6285
rect 5978 6258 6006 6259
rect 6030 6285 6058 6286
rect 6030 6259 6031 6285
rect 6031 6259 6057 6285
rect 6057 6259 6058 6285
rect 6030 6258 6058 6259
rect 6510 8694 6538 8722
rect 6622 9142 6650 9170
rect 7854 10009 7882 10010
rect 7854 9983 7855 10009
rect 7855 9983 7881 10009
rect 7881 9983 7882 10009
rect 7854 9982 7882 9983
rect 8974 9758 9002 9786
rect 9254 9982 9282 10010
rect 8302 9729 8330 9730
rect 8302 9703 8303 9729
rect 8303 9703 8329 9729
rect 8329 9703 8330 9729
rect 8302 9702 8330 9703
rect 8078 9478 8106 9506
rect 8750 9505 8778 9506
rect 8750 9479 8751 9505
rect 8751 9479 8777 9505
rect 8777 9479 8778 9505
rect 8750 9478 8778 9479
rect 8586 9421 8614 9422
rect 8586 9395 8587 9421
rect 8587 9395 8613 9421
rect 8613 9395 8614 9421
rect 8586 9394 8614 9395
rect 8638 9421 8666 9422
rect 8638 9395 8639 9421
rect 8639 9395 8665 9421
rect 8665 9395 8666 9421
rect 8638 9394 8666 9395
rect 8690 9421 8718 9422
rect 8690 9395 8691 9421
rect 8691 9395 8717 9421
rect 8717 9395 8718 9421
rect 8690 9394 8718 9395
rect 8862 9505 8890 9506
rect 8862 9479 8863 9505
rect 8863 9479 8889 9505
rect 8889 9479 8890 9505
rect 8862 9478 8890 9479
rect 10486 10009 10514 10010
rect 10486 9983 10487 10009
rect 10487 9983 10513 10009
rect 10513 9983 10514 10009
rect 10486 9982 10514 9983
rect 9478 9478 9506 9506
rect 7854 9281 7882 9282
rect 7854 9255 7855 9281
rect 7855 9255 7881 9281
rect 7881 9255 7882 9281
rect 7854 9254 7882 9255
rect 7686 9142 7714 9170
rect 6678 8974 6706 9002
rect 6622 8358 6650 8386
rect 6790 8862 6818 8890
rect 7126 9030 7154 9058
rect 7070 8750 7098 8778
rect 7350 9113 7378 9114
rect 7350 9087 7351 9113
rect 7351 9087 7377 9113
rect 7377 9087 7378 9113
rect 7350 9086 7378 9087
rect 7182 8974 7210 9002
rect 7256 9029 7284 9030
rect 7256 9003 7257 9029
rect 7257 9003 7283 9029
rect 7283 9003 7284 9029
rect 7256 9002 7284 9003
rect 7308 9029 7336 9030
rect 7308 9003 7309 9029
rect 7309 9003 7335 9029
rect 7335 9003 7336 9029
rect 7308 9002 7336 9003
rect 7360 9029 7388 9030
rect 7360 9003 7361 9029
rect 7361 9003 7387 9029
rect 7387 9003 7388 9029
rect 7360 9002 7388 9003
rect 7182 8414 7210 8442
rect 6902 8358 6930 8386
rect 6342 7910 6370 7938
rect 6286 7518 6314 7546
rect 6342 7182 6370 7210
rect 6790 6958 6818 6986
rect 6230 6846 6258 6874
rect 7256 8245 7284 8246
rect 7256 8219 7257 8245
rect 7257 8219 7283 8245
rect 7283 8219 7284 8245
rect 7256 8218 7284 8219
rect 7308 8245 7336 8246
rect 7308 8219 7309 8245
rect 7309 8219 7335 8245
rect 7335 8219 7336 8245
rect 7308 8218 7336 8219
rect 7360 8245 7388 8246
rect 7360 8219 7361 8245
rect 7361 8219 7387 8245
rect 7387 8219 7388 8245
rect 7360 8218 7388 8219
rect 6902 7910 6930 7938
rect 8586 8637 8614 8638
rect 8586 8611 8587 8637
rect 8587 8611 8613 8637
rect 8613 8611 8614 8637
rect 8586 8610 8614 8611
rect 8638 8637 8666 8638
rect 8638 8611 8639 8637
rect 8639 8611 8665 8637
rect 8665 8611 8666 8637
rect 8638 8610 8666 8611
rect 8690 8637 8718 8638
rect 8690 8611 8691 8637
rect 8691 8611 8717 8637
rect 8717 8611 8718 8637
rect 8690 8610 8718 8611
rect 7854 8414 7882 8442
rect 7014 7686 7042 7714
rect 6958 7630 6986 7658
rect 7014 7462 7042 7490
rect 6902 7265 6930 7266
rect 6902 7239 6903 7265
rect 6903 7239 6929 7265
rect 6929 7239 6930 7265
rect 6902 7238 6930 7239
rect 7182 7462 7210 7490
rect 7256 7461 7284 7462
rect 7256 7435 7257 7461
rect 7257 7435 7283 7461
rect 7283 7435 7284 7461
rect 7256 7434 7284 7435
rect 7308 7461 7336 7462
rect 7308 7435 7309 7461
rect 7309 7435 7335 7461
rect 7335 7435 7336 7461
rect 7308 7434 7336 7435
rect 7360 7461 7388 7462
rect 7360 7435 7361 7461
rect 7361 7435 7387 7461
rect 7387 7435 7388 7461
rect 7360 7434 7388 7435
rect 7182 7265 7210 7266
rect 7182 7239 7183 7265
rect 7183 7239 7209 7265
rect 7209 7239 7210 7265
rect 7182 7238 7210 7239
rect 7014 7182 7042 7210
rect 7126 6985 7154 6986
rect 7126 6959 7127 6985
rect 7127 6959 7153 6985
rect 7153 6959 7154 6985
rect 7126 6958 7154 6959
rect 7798 7321 7826 7322
rect 7798 7295 7799 7321
rect 7799 7295 7825 7321
rect 7825 7295 7826 7321
rect 7798 7294 7826 7295
rect 7462 7265 7490 7266
rect 7462 7239 7463 7265
rect 7463 7239 7489 7265
rect 7489 7239 7490 7265
rect 7462 7238 7490 7239
rect 7518 6929 7546 6930
rect 7518 6903 7519 6929
rect 7519 6903 7545 6929
rect 7545 6903 7546 6929
rect 7518 6902 7546 6903
rect 9086 8358 9114 8386
rect 9254 8134 9282 8162
rect 8022 7966 8050 7994
rect 7966 7209 7994 7210
rect 7966 7183 7967 7209
rect 7967 7183 7993 7209
rect 7993 7183 7994 7209
rect 7966 7182 7994 7183
rect 8862 7993 8890 7994
rect 8862 7967 8863 7993
rect 8863 7967 8889 7993
rect 8889 7967 8890 7993
rect 8862 7966 8890 7967
rect 8586 7853 8614 7854
rect 8586 7827 8587 7853
rect 8587 7827 8613 7853
rect 8613 7827 8614 7853
rect 8586 7826 8614 7827
rect 8638 7853 8666 7854
rect 8638 7827 8639 7853
rect 8639 7827 8665 7853
rect 8665 7827 8666 7853
rect 8638 7826 8666 7827
rect 8690 7853 8718 7854
rect 8690 7827 8691 7853
rect 8691 7827 8717 7853
rect 8717 7827 8718 7853
rect 8690 7826 8718 7827
rect 9422 7742 9450 7770
rect 9254 7574 9282 7602
rect 9198 7518 9226 7546
rect 9030 7126 9058 7154
rect 9142 7182 9170 7210
rect 8586 7069 8614 7070
rect 8586 7043 8587 7069
rect 8587 7043 8613 7069
rect 8613 7043 8614 7069
rect 8586 7042 8614 7043
rect 8638 7069 8666 7070
rect 8638 7043 8639 7069
rect 8639 7043 8665 7069
rect 8665 7043 8666 7069
rect 8638 7042 8666 7043
rect 8690 7069 8718 7070
rect 8690 7043 8691 7069
rect 8691 7043 8717 7069
rect 8717 7043 8718 7069
rect 8690 7042 8718 7043
rect 7256 6677 7284 6678
rect 7256 6651 7257 6677
rect 7257 6651 7283 6677
rect 7283 6651 7284 6677
rect 7256 6650 7284 6651
rect 7308 6677 7336 6678
rect 7308 6651 7309 6677
rect 7309 6651 7335 6677
rect 7335 6651 7336 6677
rect 7308 6650 7336 6651
rect 7360 6677 7388 6678
rect 7360 6651 7361 6677
rect 7361 6651 7387 6677
rect 7387 6651 7388 6677
rect 7360 6650 7388 6651
rect 7630 6566 7658 6594
rect 6118 5670 6146 5698
rect 6734 5614 6762 5642
rect 5926 5501 5954 5502
rect 5926 5475 5927 5501
rect 5927 5475 5953 5501
rect 5953 5475 5954 5501
rect 5926 5474 5954 5475
rect 5978 5501 6006 5502
rect 5978 5475 5979 5501
rect 5979 5475 6005 5501
rect 6005 5475 6006 5501
rect 5978 5474 6006 5475
rect 6030 5501 6058 5502
rect 6030 5475 6031 5501
rect 6031 5475 6057 5501
rect 6057 5475 6058 5501
rect 6030 5474 6058 5475
rect 6454 5361 6482 5362
rect 6454 5335 6455 5361
rect 6455 5335 6481 5361
rect 6481 5335 6482 5361
rect 6454 5334 6482 5335
rect 6566 5305 6594 5306
rect 6566 5279 6567 5305
rect 6567 5279 6593 5305
rect 6593 5279 6594 5305
rect 6566 5278 6594 5279
rect 7256 5893 7284 5894
rect 7256 5867 7257 5893
rect 7257 5867 7283 5893
rect 7283 5867 7284 5893
rect 7256 5866 7284 5867
rect 7308 5893 7336 5894
rect 7308 5867 7309 5893
rect 7309 5867 7335 5893
rect 7335 5867 7336 5893
rect 7308 5866 7336 5867
rect 7360 5893 7388 5894
rect 7360 5867 7361 5893
rect 7361 5867 7387 5893
rect 7387 5867 7388 5893
rect 7360 5866 7388 5867
rect 7182 5641 7210 5642
rect 7182 5615 7183 5641
rect 7183 5615 7209 5641
rect 7209 5615 7210 5641
rect 7182 5614 7210 5615
rect 7574 5641 7602 5642
rect 7574 5615 7575 5641
rect 7575 5615 7601 5641
rect 7601 5615 7602 5641
rect 7574 5614 7602 5615
rect 7686 5641 7714 5642
rect 7686 5615 7687 5641
rect 7687 5615 7713 5641
rect 7713 5615 7714 5641
rect 7686 5614 7714 5615
rect 7686 5334 7714 5362
rect 7294 5305 7322 5306
rect 7294 5279 7295 5305
rect 7295 5279 7321 5305
rect 7321 5279 7322 5305
rect 7294 5278 7322 5279
rect 7462 5305 7490 5306
rect 7462 5279 7463 5305
rect 7463 5279 7489 5305
rect 7489 5279 7490 5305
rect 7462 5278 7490 5279
rect 5502 5166 5530 5194
rect 5390 4774 5418 4802
rect 6510 5193 6538 5194
rect 6510 5167 6511 5193
rect 6511 5167 6537 5193
rect 6537 5167 6538 5193
rect 6510 5166 6538 5167
rect 6846 5193 6874 5194
rect 6846 5167 6847 5193
rect 6847 5167 6873 5193
rect 6873 5167 6874 5193
rect 6846 5166 6874 5167
rect 7256 5109 7284 5110
rect 7256 5083 7257 5109
rect 7257 5083 7283 5109
rect 7283 5083 7284 5109
rect 7256 5082 7284 5083
rect 7308 5109 7336 5110
rect 7308 5083 7309 5109
rect 7309 5083 7335 5109
rect 7335 5083 7336 5109
rect 7308 5082 7336 5083
rect 7360 5109 7388 5110
rect 7360 5083 7361 5109
rect 7361 5083 7387 5109
rect 7387 5083 7388 5109
rect 7360 5082 7388 5083
rect 7574 5193 7602 5194
rect 7574 5167 7575 5193
rect 7575 5167 7601 5193
rect 7601 5167 7602 5193
rect 7574 5166 7602 5167
rect 7462 5054 7490 5082
rect 7574 4969 7602 4970
rect 7574 4943 7575 4969
rect 7575 4943 7601 4969
rect 7601 4943 7602 4969
rect 7574 4942 7602 4943
rect 7798 5054 7826 5082
rect 7910 6846 7938 6874
rect 9142 6846 9170 6874
rect 9198 7126 9226 7154
rect 9366 7182 9394 7210
rect 9310 6958 9338 6986
rect 9916 9813 9944 9814
rect 9916 9787 9917 9813
rect 9917 9787 9943 9813
rect 9943 9787 9944 9813
rect 9916 9786 9944 9787
rect 9968 9813 9996 9814
rect 9968 9787 9969 9813
rect 9969 9787 9995 9813
rect 9995 9787 9996 9813
rect 9968 9786 9996 9787
rect 10020 9813 10048 9814
rect 10020 9787 10021 9813
rect 10021 9787 10047 9813
rect 10047 9787 10048 9813
rect 10020 9786 10048 9787
rect 9870 9505 9898 9506
rect 9870 9479 9871 9505
rect 9871 9479 9897 9505
rect 9897 9479 9898 9505
rect 9870 9478 9898 9479
rect 9814 9310 9842 9338
rect 10822 9561 10850 9562
rect 10822 9535 10823 9561
rect 10823 9535 10849 9561
rect 10849 9535 10850 9561
rect 10822 9534 10850 9535
rect 10038 9254 10066 9282
rect 9758 9198 9786 9226
rect 10206 9198 10234 9226
rect 10038 9169 10066 9170
rect 10038 9143 10039 9169
rect 10039 9143 10065 9169
rect 10065 9143 10066 9169
rect 10038 9142 10066 9143
rect 9870 9113 9898 9114
rect 9870 9087 9871 9113
rect 9871 9087 9897 9113
rect 9897 9087 9898 9113
rect 9870 9086 9898 9087
rect 9916 9029 9944 9030
rect 9916 9003 9917 9029
rect 9917 9003 9943 9029
rect 9943 9003 9944 9029
rect 9916 9002 9944 9003
rect 9968 9029 9996 9030
rect 9968 9003 9969 9029
rect 9969 9003 9995 9029
rect 9995 9003 9996 9029
rect 9968 9002 9996 9003
rect 10020 9029 10048 9030
rect 10020 9003 10021 9029
rect 10021 9003 10047 9029
rect 10047 9003 10048 9029
rect 10020 9002 10048 9003
rect 9702 8918 9730 8946
rect 10094 8918 10122 8946
rect 10150 9086 10178 9114
rect 10038 8526 10066 8554
rect 10486 9142 10514 9170
rect 10598 9225 10626 9226
rect 10598 9199 10599 9225
rect 10599 9199 10625 9225
rect 10625 9199 10626 9225
rect 10598 9198 10626 9199
rect 10598 8526 10626 8554
rect 11102 9561 11130 9562
rect 11102 9535 11103 9561
rect 11103 9535 11129 9561
rect 11129 9535 11130 9561
rect 11102 9534 11130 9535
rect 11246 9421 11274 9422
rect 11246 9395 11247 9421
rect 11247 9395 11273 9421
rect 11273 9395 11274 9421
rect 11246 9394 11274 9395
rect 11298 9421 11326 9422
rect 11298 9395 11299 9421
rect 11299 9395 11325 9421
rect 11325 9395 11326 9421
rect 11298 9394 11326 9395
rect 11350 9421 11378 9422
rect 11350 9395 11351 9421
rect 11351 9395 11377 9421
rect 11377 9395 11378 9421
rect 11350 9394 11378 9395
rect 10990 9254 11018 9282
rect 11246 8637 11274 8638
rect 11246 8611 11247 8637
rect 11247 8611 11273 8637
rect 11273 8611 11274 8637
rect 11246 8610 11274 8611
rect 11298 8637 11326 8638
rect 11298 8611 11299 8637
rect 11299 8611 11325 8637
rect 11325 8611 11326 8637
rect 11298 8610 11326 8611
rect 11350 8637 11378 8638
rect 11350 8611 11351 8637
rect 11351 8611 11377 8637
rect 11377 8611 11378 8637
rect 11350 8610 11378 8611
rect 10094 8414 10122 8442
rect 10822 8441 10850 8442
rect 10822 8415 10823 8441
rect 10823 8415 10849 8441
rect 10849 8415 10850 8441
rect 10822 8414 10850 8415
rect 9982 8302 10010 8330
rect 9916 8245 9944 8246
rect 9916 8219 9917 8245
rect 9917 8219 9943 8245
rect 9943 8219 9944 8245
rect 9916 8218 9944 8219
rect 9968 8245 9996 8246
rect 9968 8219 9969 8245
rect 9969 8219 9995 8245
rect 9995 8219 9996 8245
rect 9968 8218 9996 8219
rect 10020 8245 10048 8246
rect 10020 8219 10021 8245
rect 10021 8219 10047 8245
rect 10047 8219 10048 8245
rect 10020 8218 10048 8219
rect 9534 8022 9562 8050
rect 9870 8134 9898 8162
rect 9870 8049 9898 8050
rect 9870 8023 9871 8049
rect 9871 8023 9897 8049
rect 9897 8023 9898 8049
rect 9870 8022 9898 8023
rect 9758 7742 9786 7770
rect 9982 8105 10010 8106
rect 9982 8079 9983 8105
rect 9983 8079 10009 8105
rect 10009 8079 10010 8105
rect 9982 8078 10010 8079
rect 10318 8078 10346 8106
rect 10206 8049 10234 8050
rect 10206 8023 10207 8049
rect 10207 8023 10233 8049
rect 10233 8023 10234 8049
rect 10206 8022 10234 8023
rect 9758 7518 9786 7546
rect 9916 7461 9944 7462
rect 9916 7435 9917 7461
rect 9917 7435 9943 7461
rect 9943 7435 9944 7461
rect 9916 7434 9944 7435
rect 9968 7461 9996 7462
rect 9968 7435 9969 7461
rect 9969 7435 9995 7461
rect 9995 7435 9996 7461
rect 9968 7434 9996 7435
rect 10020 7461 10048 7462
rect 10020 7435 10021 7461
rect 10021 7435 10047 7461
rect 10047 7435 10048 7461
rect 10020 7434 10048 7435
rect 9590 7182 9618 7210
rect 9478 7070 9506 7098
rect 9590 6985 9618 6986
rect 9590 6959 9591 6985
rect 9591 6959 9617 6985
rect 9617 6959 9618 6985
rect 9590 6958 9618 6959
rect 9254 6678 9282 6706
rect 8586 6285 8614 6286
rect 8586 6259 8587 6285
rect 8587 6259 8613 6285
rect 8613 6259 8614 6285
rect 8586 6258 8614 6259
rect 8638 6285 8666 6286
rect 8638 6259 8639 6285
rect 8639 6259 8665 6285
rect 8665 6259 8666 6285
rect 8638 6258 8666 6259
rect 8690 6285 8718 6286
rect 8690 6259 8691 6285
rect 8691 6259 8717 6285
rect 8717 6259 8718 6285
rect 8690 6258 8718 6259
rect 9254 6062 9282 6090
rect 9198 5614 9226 5642
rect 8586 5501 8614 5502
rect 8586 5475 8587 5501
rect 8587 5475 8613 5501
rect 8613 5475 8614 5501
rect 8586 5474 8614 5475
rect 8638 5501 8666 5502
rect 8638 5475 8639 5501
rect 8639 5475 8665 5501
rect 8665 5475 8666 5501
rect 8638 5474 8666 5475
rect 8690 5501 8718 5502
rect 8690 5475 8691 5501
rect 8691 5475 8717 5501
rect 8717 5475 8718 5501
rect 8690 5474 8718 5475
rect 7910 5305 7938 5306
rect 7910 5279 7911 5305
rect 7911 5279 7937 5305
rect 7937 5279 7938 5305
rect 7910 5278 7938 5279
rect 9198 5278 9226 5306
rect 7854 4942 7882 4970
rect 7966 4886 7994 4914
rect 9254 5193 9282 5194
rect 9254 5167 9255 5193
rect 9255 5167 9281 5193
rect 9281 5167 9282 5193
rect 9254 5166 9282 5167
rect 6958 4857 6986 4858
rect 6958 4831 6959 4857
rect 6959 4831 6985 4857
rect 6985 4831 6986 4857
rect 6958 4830 6986 4831
rect 7350 4774 7378 4802
rect 5926 4717 5954 4718
rect 5926 4691 5927 4717
rect 5927 4691 5953 4717
rect 5953 4691 5954 4717
rect 5926 4690 5954 4691
rect 5978 4717 6006 4718
rect 5978 4691 5979 4717
rect 5979 4691 6005 4717
rect 6005 4691 6006 4717
rect 5978 4690 6006 4691
rect 6030 4717 6058 4718
rect 6030 4691 6031 4717
rect 6031 4691 6057 4717
rect 6057 4691 6058 4717
rect 6030 4690 6058 4691
rect 5446 4577 5474 4578
rect 5446 4551 5447 4577
rect 5447 4551 5473 4577
rect 5473 4551 5474 4577
rect 5446 4550 5474 4551
rect 7350 4606 7378 4634
rect 8586 4717 8614 4718
rect 8586 4691 8587 4717
rect 8587 4691 8613 4717
rect 8613 4691 8614 4717
rect 8586 4690 8614 4691
rect 8638 4717 8666 4718
rect 8638 4691 8639 4717
rect 8639 4691 8665 4717
rect 8665 4691 8666 4717
rect 8638 4690 8666 4691
rect 8690 4717 8718 4718
rect 8690 4691 8691 4717
rect 8691 4691 8717 4717
rect 8717 4691 8718 4717
rect 8690 4690 8718 4691
rect 5110 4046 5138 4074
rect 7256 4325 7284 4326
rect 7256 4299 7257 4325
rect 7257 4299 7283 4325
rect 7283 4299 7284 4325
rect 7256 4298 7284 4299
rect 7308 4325 7336 4326
rect 7308 4299 7309 4325
rect 7309 4299 7335 4325
rect 7335 4299 7336 4325
rect 7308 4298 7336 4299
rect 7360 4325 7388 4326
rect 7360 4299 7361 4325
rect 7361 4299 7387 4325
rect 7387 4299 7388 4325
rect 7360 4298 7388 4299
rect 5334 4214 5362 4242
rect 5726 4158 5754 4186
rect 5614 4073 5642 4074
rect 5614 4047 5615 4073
rect 5615 4047 5641 4073
rect 5641 4047 5642 4073
rect 5614 4046 5642 4047
rect 5054 3934 5082 3962
rect 5334 3990 5362 4018
rect 5054 3849 5082 3850
rect 5054 3823 5055 3849
rect 5055 3823 5081 3849
rect 5081 3823 5082 3849
rect 5054 3822 5082 3823
rect 5222 3822 5250 3850
rect 2646 3766 2674 3794
rect 5110 3793 5138 3794
rect 5110 3767 5111 3793
rect 5111 3767 5137 3793
rect 5137 3767 5138 3793
rect 5110 3766 5138 3767
rect 2366 3598 2394 3626
rect 7686 4129 7714 4130
rect 7686 4103 7687 4129
rect 7687 4103 7713 4129
rect 7713 4103 7714 4129
rect 7686 4102 7714 4103
rect 7462 4073 7490 4074
rect 7462 4047 7463 4073
rect 7463 4047 7489 4073
rect 7489 4047 7490 4073
rect 7462 4046 7490 4047
rect 5926 3933 5954 3934
rect 5926 3907 5927 3933
rect 5927 3907 5953 3933
rect 5953 3907 5954 3933
rect 5926 3906 5954 3907
rect 5978 3933 6006 3934
rect 5978 3907 5979 3933
rect 5979 3907 6005 3933
rect 6005 3907 6006 3933
rect 5978 3906 6006 3907
rect 6030 3933 6058 3934
rect 6030 3907 6031 3933
rect 6031 3907 6057 3933
rect 6057 3907 6058 3933
rect 6030 3906 6058 3907
rect 5502 3710 5530 3738
rect 5558 3793 5586 3794
rect 5558 3767 5559 3793
rect 5559 3767 5585 3793
rect 5585 3767 5586 3793
rect 5558 3766 5586 3767
rect 2870 3598 2898 3626
rect 1936 3541 1964 3542
rect 1936 3515 1937 3541
rect 1937 3515 1963 3541
rect 1963 3515 1964 3541
rect 1936 3514 1964 3515
rect 1988 3541 2016 3542
rect 1988 3515 1989 3541
rect 1989 3515 2015 3541
rect 2015 3515 2016 3541
rect 1988 3514 2016 3515
rect 2040 3541 2068 3542
rect 2040 3515 2041 3541
rect 2041 3515 2067 3541
rect 2067 3515 2068 3541
rect 2040 3514 2068 3515
rect 4596 3541 4624 3542
rect 4596 3515 4597 3541
rect 4597 3515 4623 3541
rect 4623 3515 4624 3541
rect 4596 3514 4624 3515
rect 4648 3541 4676 3542
rect 4648 3515 4649 3541
rect 4649 3515 4675 3541
rect 4675 3515 4676 3541
rect 4648 3514 4676 3515
rect 4700 3541 4728 3542
rect 4700 3515 4701 3541
rect 4701 3515 4727 3541
rect 4727 3515 4728 3541
rect 4700 3514 4728 3515
rect 7294 3737 7322 3738
rect 7294 3711 7295 3737
rect 7295 3711 7321 3737
rect 7321 3711 7322 3737
rect 7294 3710 7322 3711
rect 9366 5249 9394 5250
rect 9366 5223 9367 5249
rect 9367 5223 9393 5249
rect 9393 5223 9394 5249
rect 9366 5222 9394 5223
rect 9366 4913 9394 4914
rect 9366 4887 9367 4913
rect 9367 4887 9393 4913
rect 9393 4887 9394 4913
rect 9366 4886 9394 4887
rect 9590 6873 9618 6874
rect 9590 6847 9591 6873
rect 9591 6847 9617 6873
rect 9617 6847 9618 6873
rect 9590 6846 9618 6847
rect 9646 6678 9674 6706
rect 9478 6398 9506 6426
rect 9590 6593 9618 6594
rect 9590 6567 9591 6593
rect 9591 6567 9617 6593
rect 9617 6567 9618 6593
rect 9590 6566 9618 6567
rect 9478 5446 9506 5474
rect 9534 6118 9562 6146
rect 9478 4494 9506 4522
rect 9310 4046 9338 4074
rect 9646 5950 9674 5978
rect 9758 7153 9786 7154
rect 9758 7127 9759 7153
rect 9759 7127 9785 7153
rect 9785 7127 9786 7153
rect 9758 7126 9786 7127
rect 10038 7153 10066 7154
rect 10038 7127 10039 7153
rect 10039 7127 10065 7153
rect 10065 7127 10066 7153
rect 10038 7126 10066 7127
rect 9758 7014 9786 7042
rect 9982 6929 10010 6930
rect 9982 6903 9983 6929
rect 9983 6903 10009 6929
rect 10009 6903 10010 6929
rect 9982 6902 10010 6903
rect 9814 6873 9842 6874
rect 9814 6847 9815 6873
rect 9815 6847 9841 6873
rect 9841 6847 9842 6873
rect 9814 6846 9842 6847
rect 9916 6677 9944 6678
rect 9916 6651 9917 6677
rect 9917 6651 9943 6677
rect 9943 6651 9944 6677
rect 9916 6650 9944 6651
rect 9968 6677 9996 6678
rect 9968 6651 9969 6677
rect 9969 6651 9995 6677
rect 9995 6651 9996 6677
rect 9968 6650 9996 6651
rect 10020 6677 10048 6678
rect 10020 6651 10021 6677
rect 10021 6651 10047 6677
rect 10047 6651 10048 6677
rect 10020 6650 10048 6651
rect 10206 6566 10234 6594
rect 9758 6481 9786 6482
rect 9758 6455 9759 6481
rect 9759 6455 9785 6481
rect 9785 6455 9786 6481
rect 9758 6454 9786 6455
rect 10038 6481 10066 6482
rect 10038 6455 10039 6481
rect 10039 6455 10065 6481
rect 10065 6455 10066 6481
rect 10038 6454 10066 6455
rect 9814 6398 9842 6426
rect 9814 6118 9842 6146
rect 9758 5977 9786 5978
rect 9758 5951 9759 5977
rect 9759 5951 9785 5977
rect 9785 5951 9786 5977
rect 9758 5950 9786 5951
rect 9916 5893 9944 5894
rect 9916 5867 9917 5893
rect 9917 5867 9943 5893
rect 9943 5867 9944 5893
rect 9916 5866 9944 5867
rect 9968 5893 9996 5894
rect 9968 5867 9969 5893
rect 9969 5867 9995 5893
rect 9995 5867 9996 5893
rect 9968 5866 9996 5867
rect 10020 5893 10048 5894
rect 10020 5867 10021 5893
rect 10021 5867 10047 5893
rect 10047 5867 10048 5893
rect 10020 5866 10048 5867
rect 10094 5838 10122 5866
rect 9646 5305 9674 5306
rect 9646 5279 9647 5305
rect 9647 5279 9673 5305
rect 9673 5279 9674 5305
rect 9646 5278 9674 5279
rect 9702 5222 9730 5250
rect 9646 5166 9674 5194
rect 9590 5054 9618 5082
rect 10038 5782 10066 5810
rect 10934 6929 10962 6930
rect 10934 6903 10935 6929
rect 10935 6903 10961 6929
rect 10961 6903 10962 6929
rect 10934 6902 10962 6903
rect 10822 6817 10850 6818
rect 10822 6791 10823 6817
rect 10823 6791 10849 6817
rect 10849 6791 10850 6817
rect 10822 6790 10850 6791
rect 10934 5838 10962 5866
rect 10318 5558 10346 5586
rect 10206 5446 10234 5474
rect 10094 5334 10122 5362
rect 11102 8441 11130 8442
rect 11102 8415 11103 8441
rect 11103 8415 11129 8441
rect 11129 8415 11130 8441
rect 11102 8414 11130 8415
rect 11102 8078 11130 8106
rect 11246 7853 11274 7854
rect 11246 7827 11247 7853
rect 11247 7827 11273 7853
rect 11273 7827 11274 7853
rect 11246 7826 11274 7827
rect 11298 7853 11326 7854
rect 11298 7827 11299 7853
rect 11299 7827 11325 7853
rect 11325 7827 11326 7853
rect 11298 7826 11326 7827
rect 11350 7853 11378 7854
rect 11350 7827 11351 7853
rect 11351 7827 11377 7853
rect 11377 7827 11378 7853
rect 11350 7826 11378 7827
rect 11246 7069 11274 7070
rect 11246 7043 11247 7069
rect 11247 7043 11273 7069
rect 11273 7043 11274 7069
rect 11246 7042 11274 7043
rect 11298 7069 11326 7070
rect 11298 7043 11299 7069
rect 11299 7043 11325 7069
rect 11325 7043 11326 7069
rect 11298 7042 11326 7043
rect 11350 7069 11378 7070
rect 11350 7043 11351 7069
rect 11351 7043 11377 7069
rect 11377 7043 11378 7069
rect 11350 7042 11378 7043
rect 11102 6790 11130 6818
rect 11102 6622 11130 6650
rect 11246 6285 11274 6286
rect 11246 6259 11247 6285
rect 11247 6259 11273 6285
rect 11273 6259 11274 6285
rect 11246 6258 11274 6259
rect 11298 6285 11326 6286
rect 11298 6259 11299 6285
rect 11299 6259 11325 6285
rect 11325 6259 11326 6285
rect 11298 6258 11326 6259
rect 11350 6285 11378 6286
rect 11350 6259 11351 6285
rect 11351 6259 11377 6285
rect 11377 6259 11378 6285
rect 11350 6258 11378 6259
rect 10990 5782 11018 5810
rect 11246 5501 11274 5502
rect 11246 5475 11247 5501
rect 11247 5475 11273 5501
rect 11273 5475 11274 5501
rect 11246 5474 11274 5475
rect 11298 5501 11326 5502
rect 11298 5475 11299 5501
rect 11299 5475 11325 5501
rect 11325 5475 11326 5501
rect 11298 5474 11326 5475
rect 11350 5501 11378 5502
rect 11350 5475 11351 5501
rect 11351 5475 11377 5501
rect 11377 5475 11378 5501
rect 11350 5474 11378 5475
rect 9702 4969 9730 4970
rect 9702 4943 9703 4969
rect 9703 4943 9729 4969
rect 9729 4943 9730 4969
rect 9702 4942 9730 4943
rect 9534 4102 9562 4130
rect 9590 4438 9618 4466
rect 7910 4017 7938 4018
rect 7910 3991 7911 4017
rect 7911 3991 7937 4017
rect 7937 3991 7938 4017
rect 7910 3990 7938 3991
rect 7256 3541 7284 3542
rect 7256 3515 7257 3541
rect 7257 3515 7283 3541
rect 7283 3515 7284 3541
rect 7256 3514 7284 3515
rect 7308 3541 7336 3542
rect 7308 3515 7309 3541
rect 7309 3515 7335 3541
rect 7335 3515 7336 3541
rect 7308 3514 7336 3515
rect 7360 3541 7388 3542
rect 7360 3515 7361 3541
rect 7361 3515 7387 3541
rect 7387 3515 7388 3541
rect 7360 3514 7388 3515
rect 5558 3374 5586 3402
rect 7406 3401 7434 3402
rect 7406 3375 7407 3401
rect 7407 3375 7433 3401
rect 7433 3375 7434 3401
rect 7406 3374 7434 3375
rect 7630 3401 7658 3402
rect 7630 3375 7631 3401
rect 7631 3375 7657 3401
rect 7657 3375 7658 3401
rect 7630 3374 7658 3375
rect 8586 3933 8614 3934
rect 8586 3907 8587 3933
rect 8587 3907 8613 3933
rect 8613 3907 8614 3933
rect 8586 3906 8614 3907
rect 8638 3933 8666 3934
rect 8638 3907 8639 3933
rect 8639 3907 8665 3933
rect 8665 3907 8666 3933
rect 8638 3906 8666 3907
rect 8690 3933 8718 3934
rect 8690 3907 8691 3933
rect 8691 3907 8717 3933
rect 8717 3907 8718 3933
rect 8690 3906 8718 3907
rect 9366 3766 9394 3794
rect 9702 4494 9730 4522
rect 9916 5109 9944 5110
rect 9916 5083 9917 5109
rect 9917 5083 9943 5109
rect 9943 5083 9944 5109
rect 9916 5082 9944 5083
rect 9968 5109 9996 5110
rect 9968 5083 9969 5109
rect 9969 5083 9995 5109
rect 9995 5083 9996 5109
rect 9968 5082 9996 5083
rect 10020 5109 10048 5110
rect 10020 5083 10021 5109
rect 10021 5083 10047 5109
rect 10047 5083 10048 5109
rect 10020 5082 10048 5083
rect 9926 4969 9954 4970
rect 9926 4943 9927 4969
rect 9927 4943 9953 4969
rect 9953 4943 9954 4969
rect 9926 4942 9954 4943
rect 9982 4913 10010 4914
rect 9982 4887 9983 4913
rect 9983 4887 10009 4913
rect 10009 4887 10010 4913
rect 9982 4886 10010 4887
rect 10822 5166 10850 5194
rect 11102 5166 11130 5194
rect 11246 4717 11274 4718
rect 11246 4691 11247 4717
rect 11247 4691 11273 4717
rect 11273 4691 11274 4717
rect 11246 4690 11274 4691
rect 11298 4717 11326 4718
rect 11298 4691 11299 4717
rect 11299 4691 11325 4717
rect 11325 4691 11326 4717
rect 11298 4690 11326 4691
rect 11350 4717 11378 4718
rect 11350 4691 11351 4717
rect 11351 4691 11377 4717
rect 11377 4691 11378 4717
rect 11350 4690 11378 4691
rect 9916 4325 9944 4326
rect 9916 4299 9917 4325
rect 9917 4299 9943 4325
rect 9943 4299 9944 4325
rect 9916 4298 9944 4299
rect 9968 4325 9996 4326
rect 9968 4299 9969 4325
rect 9969 4299 9995 4325
rect 9995 4299 9996 4325
rect 9968 4298 9996 4299
rect 10020 4325 10048 4326
rect 10020 4299 10021 4325
rect 10021 4299 10047 4325
rect 10047 4299 10048 4325
rect 10020 4298 10048 4299
rect 9870 4046 9898 4074
rect 10094 4073 10122 4074
rect 10094 4047 10095 4073
rect 10095 4047 10121 4073
rect 10121 4047 10122 4073
rect 10094 4046 10122 4047
rect 9982 3793 10010 3794
rect 9982 3767 9983 3793
rect 9983 3767 10009 3793
rect 10009 3767 10010 3793
rect 9982 3766 10010 3767
rect 10318 4017 10346 4018
rect 10318 3991 10319 4017
rect 10319 3991 10345 4017
rect 10345 3991 10346 4017
rect 10318 3990 10346 3991
rect 9814 3710 9842 3738
rect 10150 3737 10178 3738
rect 10150 3711 10151 3737
rect 10151 3711 10177 3737
rect 10177 3711 10178 3737
rect 10150 3710 10178 3711
rect 9590 3598 9618 3626
rect 9916 3541 9944 3542
rect 9916 3515 9917 3541
rect 9917 3515 9943 3541
rect 9943 3515 9944 3541
rect 9916 3514 9944 3515
rect 9968 3541 9996 3542
rect 9968 3515 9969 3541
rect 9969 3515 9995 3541
rect 9995 3515 9996 3541
rect 9968 3514 9996 3515
rect 10020 3541 10048 3542
rect 10020 3515 10021 3541
rect 10021 3515 10047 3541
rect 10047 3515 10048 3541
rect 10020 3514 10048 3515
rect 7910 3374 7938 3402
rect 9814 3430 9842 3458
rect 3266 3149 3294 3150
rect 3266 3123 3267 3149
rect 3267 3123 3293 3149
rect 3293 3123 3294 3149
rect 3266 3122 3294 3123
rect 3318 3149 3346 3150
rect 3318 3123 3319 3149
rect 3319 3123 3345 3149
rect 3345 3123 3346 3149
rect 3318 3122 3346 3123
rect 3370 3149 3398 3150
rect 3370 3123 3371 3149
rect 3371 3123 3397 3149
rect 3397 3123 3398 3149
rect 3370 3122 3398 3123
rect 5926 3149 5954 3150
rect 5926 3123 5927 3149
rect 5927 3123 5953 3149
rect 5953 3123 5954 3149
rect 5926 3122 5954 3123
rect 5978 3149 6006 3150
rect 5978 3123 5979 3149
rect 5979 3123 6005 3149
rect 6005 3123 6006 3149
rect 5978 3122 6006 3123
rect 6030 3149 6058 3150
rect 6030 3123 6031 3149
rect 6031 3123 6057 3149
rect 6057 3123 6058 3149
rect 6030 3122 6058 3123
rect 8586 3149 8614 3150
rect 8586 3123 8587 3149
rect 8587 3123 8613 3149
rect 8613 3123 8614 3149
rect 8586 3122 8614 3123
rect 8638 3149 8666 3150
rect 8638 3123 8639 3149
rect 8639 3123 8665 3149
rect 8665 3123 8666 3149
rect 8638 3122 8666 3123
rect 8690 3149 8718 3150
rect 8690 3123 8691 3149
rect 8691 3123 8717 3149
rect 8717 3123 8718 3149
rect 8690 3122 8718 3123
rect 1936 2757 1964 2758
rect 1936 2731 1937 2757
rect 1937 2731 1963 2757
rect 1963 2731 1964 2757
rect 1936 2730 1964 2731
rect 1988 2757 2016 2758
rect 1988 2731 1989 2757
rect 1989 2731 2015 2757
rect 2015 2731 2016 2757
rect 1988 2730 2016 2731
rect 2040 2757 2068 2758
rect 2040 2731 2041 2757
rect 2041 2731 2067 2757
rect 2067 2731 2068 2757
rect 2040 2730 2068 2731
rect 4596 2757 4624 2758
rect 4596 2731 4597 2757
rect 4597 2731 4623 2757
rect 4623 2731 4624 2757
rect 4596 2730 4624 2731
rect 4648 2757 4676 2758
rect 4648 2731 4649 2757
rect 4649 2731 4675 2757
rect 4675 2731 4676 2757
rect 4648 2730 4676 2731
rect 4700 2757 4728 2758
rect 4700 2731 4701 2757
rect 4701 2731 4727 2757
rect 4727 2731 4728 2757
rect 4700 2730 4728 2731
rect 7256 2757 7284 2758
rect 7256 2731 7257 2757
rect 7257 2731 7283 2757
rect 7283 2731 7284 2757
rect 7256 2730 7284 2731
rect 7308 2757 7336 2758
rect 7308 2731 7309 2757
rect 7309 2731 7335 2757
rect 7335 2731 7336 2757
rect 7308 2730 7336 2731
rect 7360 2757 7388 2758
rect 7360 2731 7361 2757
rect 7361 2731 7387 2757
rect 7387 2731 7388 2757
rect 7360 2730 7388 2731
rect 3266 2365 3294 2366
rect 3266 2339 3267 2365
rect 3267 2339 3293 2365
rect 3293 2339 3294 2365
rect 3266 2338 3294 2339
rect 3318 2365 3346 2366
rect 3318 2339 3319 2365
rect 3319 2339 3345 2365
rect 3345 2339 3346 2365
rect 3318 2338 3346 2339
rect 3370 2365 3398 2366
rect 3370 2339 3371 2365
rect 3371 2339 3397 2365
rect 3397 2339 3398 2365
rect 3370 2338 3398 2339
rect 5926 2365 5954 2366
rect 5926 2339 5927 2365
rect 5927 2339 5953 2365
rect 5953 2339 5954 2365
rect 5926 2338 5954 2339
rect 5978 2365 6006 2366
rect 5978 2339 5979 2365
rect 5979 2339 6005 2365
rect 6005 2339 6006 2365
rect 5978 2338 6006 2339
rect 6030 2365 6058 2366
rect 6030 2339 6031 2365
rect 6031 2339 6057 2365
rect 6057 2339 6058 2365
rect 6030 2338 6058 2339
rect 8586 2365 8614 2366
rect 8586 2339 8587 2365
rect 8587 2339 8613 2365
rect 8613 2339 8614 2365
rect 8586 2338 8614 2339
rect 8638 2365 8666 2366
rect 8638 2339 8639 2365
rect 8639 2339 8665 2365
rect 8665 2339 8666 2365
rect 8638 2338 8666 2339
rect 8690 2365 8718 2366
rect 8690 2339 8691 2365
rect 8691 2339 8717 2365
rect 8717 2339 8718 2365
rect 8690 2338 8718 2339
rect 1936 1973 1964 1974
rect 1936 1947 1937 1973
rect 1937 1947 1963 1973
rect 1963 1947 1964 1973
rect 1936 1946 1964 1947
rect 1988 1973 2016 1974
rect 1988 1947 1989 1973
rect 1989 1947 2015 1973
rect 2015 1947 2016 1973
rect 1988 1946 2016 1947
rect 2040 1973 2068 1974
rect 2040 1947 2041 1973
rect 2041 1947 2067 1973
rect 2067 1947 2068 1973
rect 2040 1946 2068 1947
rect 4596 1973 4624 1974
rect 4596 1947 4597 1973
rect 4597 1947 4623 1973
rect 4623 1947 4624 1973
rect 4596 1946 4624 1947
rect 4648 1973 4676 1974
rect 4648 1947 4649 1973
rect 4649 1947 4675 1973
rect 4675 1947 4676 1973
rect 4648 1946 4676 1947
rect 4700 1973 4728 1974
rect 4700 1947 4701 1973
rect 4701 1947 4727 1973
rect 4727 1947 4728 1973
rect 4700 1946 4728 1947
rect 7256 1973 7284 1974
rect 7256 1947 7257 1973
rect 7257 1947 7283 1973
rect 7283 1947 7284 1973
rect 7256 1946 7284 1947
rect 7308 1973 7336 1974
rect 7308 1947 7309 1973
rect 7309 1947 7335 1973
rect 7335 1947 7336 1973
rect 7308 1946 7336 1947
rect 7360 1973 7388 1974
rect 7360 1947 7361 1973
rect 7361 1947 7387 1973
rect 7387 1947 7388 1973
rect 7360 1946 7388 1947
rect 3266 1581 3294 1582
rect 3266 1555 3267 1581
rect 3267 1555 3293 1581
rect 3293 1555 3294 1581
rect 3266 1554 3294 1555
rect 3318 1581 3346 1582
rect 3318 1555 3319 1581
rect 3319 1555 3345 1581
rect 3345 1555 3346 1581
rect 3318 1554 3346 1555
rect 3370 1581 3398 1582
rect 3370 1555 3371 1581
rect 3371 1555 3397 1581
rect 3397 1555 3398 1581
rect 3370 1554 3398 1555
rect 5926 1581 5954 1582
rect 5926 1555 5927 1581
rect 5927 1555 5953 1581
rect 5953 1555 5954 1581
rect 5926 1554 5954 1555
rect 5978 1581 6006 1582
rect 5978 1555 5979 1581
rect 5979 1555 6005 1581
rect 6005 1555 6006 1581
rect 5978 1554 6006 1555
rect 6030 1581 6058 1582
rect 6030 1555 6031 1581
rect 6031 1555 6057 1581
rect 6057 1555 6058 1581
rect 6030 1554 6058 1555
rect 8586 1581 8614 1582
rect 8586 1555 8587 1581
rect 8587 1555 8613 1581
rect 8613 1555 8614 1581
rect 8586 1554 8614 1555
rect 8638 1581 8666 1582
rect 8638 1555 8639 1581
rect 8639 1555 8665 1581
rect 8665 1555 8666 1581
rect 8638 1554 8666 1555
rect 8690 1581 8718 1582
rect 8690 1555 8691 1581
rect 8691 1555 8717 1581
rect 8717 1555 8718 1581
rect 8690 1554 8718 1555
rect 10934 4073 10962 4074
rect 10934 4047 10935 4073
rect 10935 4047 10961 4073
rect 10961 4047 10962 4073
rect 10934 4046 10962 4047
rect 10766 4017 10794 4018
rect 10766 3991 10767 4017
rect 10767 3991 10793 4017
rect 10793 3991 10794 4017
rect 10766 3990 10794 3991
rect 10374 3710 10402 3738
rect 10934 3710 10962 3738
rect 10318 3430 10346 3458
rect 9916 2757 9944 2758
rect 9916 2731 9917 2757
rect 9917 2731 9943 2757
rect 9943 2731 9944 2757
rect 9916 2730 9944 2731
rect 9968 2757 9996 2758
rect 9968 2731 9969 2757
rect 9969 2731 9995 2757
rect 9995 2731 9996 2757
rect 9968 2730 9996 2731
rect 10020 2757 10048 2758
rect 10020 2731 10021 2757
rect 10021 2731 10047 2757
rect 10047 2731 10048 2757
rect 10020 2730 10048 2731
rect 10822 2561 10850 2562
rect 10822 2535 10823 2561
rect 10823 2535 10849 2561
rect 10849 2535 10850 2561
rect 10822 2534 10850 2535
rect 11246 3933 11274 3934
rect 11246 3907 11247 3933
rect 11247 3907 11273 3933
rect 11273 3907 11274 3933
rect 11246 3906 11274 3907
rect 11298 3933 11326 3934
rect 11298 3907 11299 3933
rect 11299 3907 11325 3933
rect 11325 3907 11326 3933
rect 11298 3906 11326 3907
rect 11350 3933 11378 3934
rect 11350 3907 11351 3933
rect 11351 3907 11377 3933
rect 11377 3907 11378 3933
rect 11350 3906 11378 3907
rect 11102 3737 11130 3738
rect 11102 3711 11103 3737
rect 11103 3711 11129 3737
rect 11129 3711 11130 3737
rect 11102 3710 11130 3711
rect 11246 3149 11274 3150
rect 11246 3123 11247 3149
rect 11247 3123 11273 3149
rect 11273 3123 11274 3149
rect 11246 3122 11274 3123
rect 11298 3149 11326 3150
rect 11298 3123 11299 3149
rect 11299 3123 11325 3149
rect 11325 3123 11326 3149
rect 11298 3122 11326 3123
rect 11350 3149 11378 3150
rect 11350 3123 11351 3149
rect 11351 3123 11377 3149
rect 11377 3123 11378 3149
rect 11350 3122 11378 3123
rect 11102 2561 11130 2562
rect 11102 2535 11103 2561
rect 11103 2535 11129 2561
rect 11129 2535 11130 2561
rect 11102 2534 11130 2535
rect 11246 2365 11274 2366
rect 11246 2339 11247 2365
rect 11247 2339 11273 2365
rect 11273 2339 11274 2365
rect 11246 2338 11274 2339
rect 11298 2365 11326 2366
rect 11298 2339 11299 2365
rect 11299 2339 11325 2365
rect 11325 2339 11326 2365
rect 11298 2338 11326 2339
rect 11350 2365 11378 2366
rect 11350 2339 11351 2365
rect 11351 2339 11377 2365
rect 11377 2339 11378 2365
rect 11350 2338 11378 2339
rect 11102 2254 11130 2282
rect 9916 1973 9944 1974
rect 9916 1947 9917 1973
rect 9917 1947 9943 1973
rect 9943 1947 9944 1973
rect 9916 1946 9944 1947
rect 9968 1973 9996 1974
rect 9968 1947 9969 1973
rect 9969 1947 9995 1973
rect 9995 1947 9996 1973
rect 9968 1946 9996 1947
rect 10020 1973 10048 1974
rect 10020 1947 10021 1973
rect 10021 1947 10047 1973
rect 10047 1947 10048 1973
rect 10020 1946 10048 1947
rect 11246 1581 11274 1582
rect 11246 1555 11247 1581
rect 11247 1555 11273 1581
rect 11273 1555 11274 1581
rect 11246 1554 11274 1555
rect 11298 1581 11326 1582
rect 11298 1555 11299 1581
rect 11299 1555 11325 1581
rect 11325 1555 11326 1581
rect 11298 1554 11326 1555
rect 11350 1581 11378 1582
rect 11350 1555 11351 1581
rect 11351 1555 11377 1581
rect 11377 1555 11378 1581
rect 11350 1554 11378 1555
rect 9814 798 9842 826
<< metal3 >>
rect 11600 11018 12000 11032
rect 10033 10990 10038 11018
rect 10066 10990 12000 11018
rect 11600 10976 12000 10990
rect 3261 10178 3266 10206
rect 3294 10178 3318 10206
rect 3346 10178 3370 10206
rect 3398 10178 3403 10206
rect 5921 10178 5926 10206
rect 5954 10178 5978 10206
rect 6006 10178 6030 10206
rect 6058 10178 6063 10206
rect 8581 10178 8586 10206
rect 8614 10178 8638 10206
rect 8666 10178 8690 10206
rect 8718 10178 8723 10206
rect 11241 10178 11246 10206
rect 11274 10178 11298 10206
rect 11326 10178 11350 10206
rect 11378 10178 11383 10206
rect 9865 10038 9870 10066
rect 9898 10038 10374 10066
rect 10402 10038 10407 10066
rect 7513 9982 7518 10010
rect 7546 9982 7854 10010
rect 7882 9982 7887 10010
rect 9249 9982 9254 10010
rect 9282 9982 10486 10010
rect 10514 9982 10519 10010
rect 1931 9786 1936 9814
rect 1964 9786 1988 9814
rect 2016 9786 2040 9814
rect 2068 9786 2073 9814
rect 4591 9786 4596 9814
rect 4624 9786 4648 9814
rect 4676 9786 4700 9814
rect 4728 9786 4733 9814
rect 7251 9786 7256 9814
rect 7284 9786 7308 9814
rect 7336 9786 7360 9814
rect 7388 9786 7393 9814
rect 9911 9786 9916 9814
rect 9944 9786 9968 9814
rect 9996 9786 10020 9814
rect 10048 9786 10053 9814
rect 8969 9758 8974 9786
rect 9002 9758 9007 9786
rect 6785 9702 6790 9730
rect 6818 9702 8302 9730
rect 8330 9702 8335 9730
rect 8974 9562 9002 9758
rect 11600 9562 12000 9576
rect 2529 9534 2534 9562
rect 2562 9534 3878 9562
rect 3906 9534 3911 9562
rect 3985 9534 3990 9562
rect 4018 9534 9002 9562
rect 10817 9534 10822 9562
rect 10850 9534 11102 9562
rect 11130 9534 12000 9562
rect 3878 9506 3906 9534
rect 11600 9520 12000 9534
rect 3878 9478 4214 9506
rect 8073 9478 8078 9506
rect 8106 9478 8750 9506
rect 8778 9478 8783 9506
rect 8857 9478 8862 9506
rect 8890 9478 9478 9506
rect 9506 9478 9870 9506
rect 9898 9478 9903 9506
rect 3261 9394 3266 9422
rect 3294 9394 3318 9422
rect 3346 9394 3370 9422
rect 3398 9394 3403 9422
rect 4186 9338 4214 9478
rect 5921 9394 5926 9422
rect 5954 9394 5978 9422
rect 6006 9394 6030 9422
rect 6058 9394 6063 9422
rect 8581 9394 8586 9422
rect 8614 9394 8638 9422
rect 8666 9394 8690 9422
rect 8718 9394 8723 9422
rect 11241 9394 11246 9422
rect 11274 9394 11298 9422
rect 11326 9394 11350 9422
rect 11378 9394 11383 9422
rect 2305 9310 2310 9338
rect 2338 9310 2422 9338
rect 2450 9310 3934 9338
rect 3962 9310 3967 9338
rect 4186 9310 9814 9338
rect 9842 9310 9847 9338
rect 2081 9254 2086 9282
rect 2114 9254 2926 9282
rect 2954 9254 4326 9282
rect 4354 9254 4359 9282
rect 5553 9254 5558 9282
rect 5586 9254 6062 9282
rect 6090 9254 6095 9282
rect 6337 9254 6342 9282
rect 6370 9254 7854 9282
rect 7882 9254 7887 9282
rect 10033 9254 10038 9282
rect 10066 9254 10990 9282
rect 11018 9254 11023 9282
rect 10598 9226 10626 9254
rect 1521 9198 1526 9226
rect 1554 9198 1806 9226
rect 1834 9198 1839 9226
rect 2137 9198 2142 9226
rect 2170 9198 2198 9226
rect 2226 9198 2870 9226
rect 2898 9198 4158 9226
rect 4186 9198 4191 9226
rect 5609 9198 5614 9226
rect 5642 9198 6286 9226
rect 6314 9198 6319 9226
rect 9753 9198 9758 9226
rect 9786 9198 10206 9226
rect 10234 9198 10239 9226
rect 10593 9198 10598 9226
rect 10626 9198 10631 9226
rect 1633 9142 1638 9170
rect 1666 9142 2478 9170
rect 2506 9142 3150 9170
rect 3178 9142 3183 9170
rect 4097 9142 4102 9170
rect 4130 9142 5950 9170
rect 5978 9142 5983 9170
rect 6169 9142 6174 9170
rect 6202 9142 6622 9170
rect 6650 9142 6655 9170
rect 7681 9142 7686 9170
rect 7714 9142 10038 9170
rect 10066 9142 10486 9170
rect 10514 9142 10519 9170
rect 4265 9086 4270 9114
rect 4298 9086 4774 9114
rect 4802 9086 7350 9114
rect 7378 9086 7383 9114
rect 9865 9086 9870 9114
rect 9898 9086 10150 9114
rect 10178 9086 10183 9114
rect 5105 9030 5110 9058
rect 5138 9030 5670 9058
rect 5698 9030 5703 9058
rect 5777 9030 5782 9058
rect 5810 9030 7126 9058
rect 7154 9030 7159 9058
rect 1931 9002 1936 9030
rect 1964 9002 1988 9030
rect 2016 9002 2040 9030
rect 2068 9002 2073 9030
rect 4591 9002 4596 9030
rect 4624 9002 4648 9030
rect 4676 9002 4700 9030
rect 4728 9002 4733 9030
rect 5670 9002 5698 9030
rect 7251 9002 7256 9030
rect 7284 9002 7308 9030
rect 7336 9002 7360 9030
rect 7388 9002 7393 9030
rect 9911 9002 9916 9030
rect 9944 9002 9968 9030
rect 9996 9002 10020 9030
rect 10048 9002 10053 9030
rect 5670 8974 6678 9002
rect 6706 8974 7182 9002
rect 7210 8974 7215 9002
rect 4937 8918 4942 8946
rect 4970 8918 5446 8946
rect 5474 8918 5479 8946
rect 5665 8918 5670 8946
rect 5698 8918 9702 8946
rect 9730 8918 10094 8946
rect 10122 8918 10127 8946
rect 2641 8862 2646 8890
rect 2674 8862 5502 8890
rect 5530 8862 5950 8890
rect 5978 8862 6790 8890
rect 6818 8862 6823 8890
rect 3985 8806 3990 8834
rect 4018 8806 4023 8834
rect 3990 8778 4018 8806
rect 2081 8750 2086 8778
rect 2114 8750 3094 8778
rect 3122 8750 3127 8778
rect 3873 8750 3878 8778
rect 3906 8750 7070 8778
rect 7098 8750 7103 8778
rect 2977 8694 2982 8722
rect 3010 8694 3990 8722
rect 4018 8694 4023 8722
rect 6225 8694 6230 8722
rect 6258 8694 6510 8722
rect 6538 8694 6543 8722
rect 3261 8610 3266 8638
rect 3294 8610 3318 8638
rect 3346 8610 3370 8638
rect 3398 8610 3403 8638
rect 5921 8610 5926 8638
rect 5954 8610 5978 8638
rect 6006 8610 6030 8638
rect 6058 8610 6063 8638
rect 8581 8610 8586 8638
rect 8614 8610 8638 8638
rect 8666 8610 8690 8638
rect 8718 8610 8723 8638
rect 11241 8610 11246 8638
rect 11274 8610 11298 8638
rect 11326 8610 11350 8638
rect 11378 8610 11383 8638
rect 10033 8526 10038 8554
rect 10066 8526 10598 8554
rect 10626 8526 10631 8554
rect 5609 8414 5614 8442
rect 5642 8414 6174 8442
rect 6202 8414 6207 8442
rect 7177 8414 7182 8442
rect 7210 8414 7854 8442
rect 7882 8414 7887 8442
rect 10075 8414 10094 8442
rect 10122 8414 10127 8442
rect 10817 8414 10822 8442
rect 10850 8414 11102 8442
rect 11130 8414 11135 8442
rect 2529 8358 2534 8386
rect 2562 8358 3206 8386
rect 3234 8358 3239 8386
rect 6617 8358 6622 8386
rect 6650 8358 6902 8386
rect 6930 8358 9086 8386
rect 9114 8358 9119 8386
rect 9814 8302 9982 8330
rect 10010 8302 10015 8330
rect 1931 8218 1936 8246
rect 1964 8218 1988 8246
rect 2016 8218 2040 8246
rect 2068 8218 2073 8246
rect 4591 8218 4596 8246
rect 4624 8218 4648 8246
rect 4676 8218 4700 8246
rect 4728 8218 4733 8246
rect 7251 8218 7256 8246
rect 7284 8218 7308 8246
rect 7336 8218 7360 8246
rect 7388 8218 7393 8246
rect 9814 8162 9842 8302
rect 9911 8218 9916 8246
rect 9944 8218 9968 8246
rect 9996 8218 10020 8246
rect 10048 8218 10053 8246
rect 9249 8134 9254 8162
rect 9282 8134 9870 8162
rect 9898 8134 9903 8162
rect 11600 8106 12000 8120
rect 9977 8078 9982 8106
rect 10010 8078 10318 8106
rect 10346 8078 10351 8106
rect 11097 8078 11102 8106
rect 11130 8078 12000 8106
rect 11600 8064 12000 8078
rect 9529 8022 9534 8050
rect 9562 8022 9870 8050
rect 9898 8022 10206 8050
rect 10234 8022 10239 8050
rect 1521 7966 1526 7994
rect 1554 7966 1694 7994
rect 1722 7966 1918 7994
rect 1946 7966 1951 7994
rect 8017 7966 8022 7994
rect 8050 7966 8862 7994
rect 8890 7966 8895 7994
rect 1241 7910 1246 7938
rect 1274 7910 1974 7938
rect 2002 7910 2007 7938
rect 4153 7910 4158 7938
rect 4186 7910 4550 7938
rect 4578 7910 6342 7938
rect 6370 7910 6902 7938
rect 6930 7910 6935 7938
rect 3261 7826 3266 7854
rect 3294 7826 3318 7854
rect 3346 7826 3370 7854
rect 3398 7826 3403 7854
rect 5921 7826 5926 7854
rect 5954 7826 5978 7854
rect 6006 7826 6030 7854
rect 6058 7826 6063 7854
rect 8581 7826 8586 7854
rect 8614 7826 8638 7854
rect 8666 7826 8690 7854
rect 8718 7826 8723 7854
rect 11241 7826 11246 7854
rect 11274 7826 11298 7854
rect 11326 7826 11350 7854
rect 11378 7826 11383 7854
rect 2137 7742 2142 7770
rect 2170 7742 4830 7770
rect 4858 7742 4863 7770
rect 9417 7742 9422 7770
rect 9450 7742 9758 7770
rect 9786 7742 9791 7770
rect 7009 7686 7014 7714
rect 7042 7686 7574 7714
rect 4321 7630 4326 7658
rect 4354 7630 4774 7658
rect 4802 7630 4807 7658
rect 6225 7630 6230 7658
rect 6258 7630 6958 7658
rect 6986 7630 6991 7658
rect 7546 7602 7574 7686
rect 1185 7574 1190 7602
rect 1218 7574 1638 7602
rect 1666 7574 1974 7602
rect 2002 7574 2007 7602
rect 2081 7574 2086 7602
rect 2114 7574 2310 7602
rect 2338 7574 2478 7602
rect 2506 7574 2511 7602
rect 4377 7574 4382 7602
rect 4410 7574 4998 7602
rect 5026 7574 5894 7602
rect 5922 7574 6118 7602
rect 6146 7574 6151 7602
rect 7546 7574 9254 7602
rect 9282 7574 9287 7602
rect 4713 7518 4718 7546
rect 4746 7518 4942 7546
rect 4970 7518 4975 7546
rect 6281 7518 6286 7546
rect 6314 7518 9198 7546
rect 9226 7518 9231 7546
rect 9753 7518 9758 7546
rect 9786 7518 10094 7546
rect 10122 7518 10127 7546
rect 7009 7462 7014 7490
rect 7042 7462 7182 7490
rect 7210 7462 7215 7490
rect 1931 7434 1936 7462
rect 1964 7434 1988 7462
rect 2016 7434 2040 7462
rect 2068 7434 2073 7462
rect 4591 7434 4596 7462
rect 4624 7434 4648 7462
rect 4676 7434 4700 7462
rect 4728 7434 4733 7462
rect 7251 7434 7256 7462
rect 7284 7434 7308 7462
rect 7336 7434 7360 7462
rect 7388 7434 7393 7462
rect 9911 7434 9916 7462
rect 9944 7434 9968 7462
rect 9996 7434 10020 7462
rect 10048 7434 10053 7462
rect 3929 7406 3934 7434
rect 3962 7406 4214 7434
rect 4242 7406 4247 7434
rect 1129 7350 1134 7378
rect 1162 7350 1470 7378
rect 1498 7350 2198 7378
rect 2226 7350 2231 7378
rect 3817 7350 3822 7378
rect 3850 7350 4270 7378
rect 4298 7350 4830 7378
rect 4858 7350 4863 7378
rect 4937 7350 4942 7378
rect 4970 7350 5782 7378
rect 5810 7350 7210 7378
rect 4041 7294 4046 7322
rect 4074 7294 4494 7322
rect 4522 7294 4998 7322
rect 5026 7294 5390 7322
rect 5418 7294 6062 7322
rect 6090 7294 6095 7322
rect 7182 7266 7210 7350
rect 7546 7294 7798 7322
rect 7826 7294 7831 7322
rect 7546 7266 7574 7294
rect 5889 7238 5894 7266
rect 5922 7238 6902 7266
rect 6930 7238 6935 7266
rect 7177 7238 7182 7266
rect 7210 7238 7215 7266
rect 7457 7238 7462 7266
rect 7490 7238 7574 7266
rect 2249 7182 2254 7210
rect 2282 7182 2814 7210
rect 2842 7182 3766 7210
rect 3794 7182 3799 7210
rect 5217 7182 5222 7210
rect 5250 7182 5670 7210
rect 5698 7182 6342 7210
rect 6370 7182 7014 7210
rect 7042 7182 7047 7210
rect 7961 7182 7966 7210
rect 7994 7182 9142 7210
rect 9170 7182 9175 7210
rect 9361 7182 9366 7210
rect 9394 7182 9590 7210
rect 9618 7182 9623 7210
rect 2179 7126 2198 7154
rect 2226 7126 2231 7154
rect 6113 7126 6118 7154
rect 6146 7126 9030 7154
rect 9058 7126 9063 7154
rect 9193 7126 9198 7154
rect 9226 7126 9758 7154
rect 9786 7126 10038 7154
rect 10066 7126 10071 7154
rect 3929 7070 3934 7098
rect 3962 7070 5614 7098
rect 5642 7070 5647 7098
rect 9473 7070 9478 7098
rect 9506 7070 9786 7098
rect 3261 7042 3266 7070
rect 3294 7042 3318 7070
rect 3346 7042 3370 7070
rect 3398 7042 3403 7070
rect 5921 7042 5926 7070
rect 5954 7042 5978 7070
rect 6006 7042 6030 7070
rect 6058 7042 6063 7070
rect 8581 7042 8586 7070
rect 8614 7042 8638 7070
rect 8666 7042 8690 7070
rect 8718 7042 8723 7070
rect 9758 7042 9786 7070
rect 11241 7042 11246 7070
rect 11274 7042 11298 7070
rect 11326 7042 11350 7070
rect 11378 7042 11383 7070
rect 9739 7014 9758 7042
rect 9786 7014 9791 7042
rect 5609 6958 5614 6986
rect 5642 6958 6790 6986
rect 6818 6958 7126 6986
rect 7154 6958 7159 6986
rect 9305 6958 9310 6986
rect 9338 6958 9590 6986
rect 9618 6958 9623 6986
rect 5721 6902 5726 6930
rect 5754 6902 7518 6930
rect 7546 6902 7551 6930
rect 9977 6902 9982 6930
rect 10010 6902 10934 6930
rect 10962 6902 10967 6930
rect 5497 6846 5502 6874
rect 5530 6846 6230 6874
rect 6258 6846 6263 6874
rect 7546 6846 7910 6874
rect 7938 6846 7943 6874
rect 9137 6846 9142 6874
rect 9170 6846 9590 6874
rect 9618 6846 9623 6874
rect 9795 6846 9814 6874
rect 9842 6846 9847 6874
rect 7546 6818 7574 6846
rect 4937 6790 4942 6818
rect 4970 6790 5838 6818
rect 5866 6790 7574 6818
rect 10817 6790 10822 6818
rect 10850 6790 11102 6818
rect 11130 6790 11135 6818
rect 1801 6734 1806 6762
rect 1834 6734 4830 6762
rect 4858 6734 4863 6762
rect 9249 6678 9254 6706
rect 9282 6678 9646 6706
rect 9674 6678 9842 6706
rect 1931 6650 1936 6678
rect 1964 6650 1988 6678
rect 2016 6650 2040 6678
rect 2068 6650 2073 6678
rect 4591 6650 4596 6678
rect 4624 6650 4648 6678
rect 4676 6650 4700 6678
rect 4728 6650 4733 6678
rect 7251 6650 7256 6678
rect 7284 6650 7308 6678
rect 7336 6650 7360 6678
rect 7388 6650 7393 6678
rect 9814 6594 9842 6678
rect 9911 6650 9916 6678
rect 9944 6650 9968 6678
rect 9996 6650 10020 6678
rect 10048 6650 10053 6678
rect 11600 6650 12000 6664
rect 11097 6622 11102 6650
rect 11130 6622 12000 6650
rect 11600 6608 12000 6622
rect 7625 6566 7630 6594
rect 7658 6566 9590 6594
rect 9618 6566 9623 6594
rect 9814 6566 10206 6594
rect 10234 6566 10239 6594
rect 9753 6454 9758 6482
rect 9786 6454 10038 6482
rect 10066 6454 10071 6482
rect 9473 6398 9478 6426
rect 9506 6398 9814 6426
rect 9842 6398 9847 6426
rect 4377 6342 4382 6370
rect 4410 6342 4662 6370
rect 4690 6342 4695 6370
rect 3261 6258 3266 6286
rect 3294 6258 3318 6286
rect 3346 6258 3370 6286
rect 3398 6258 3403 6286
rect 5921 6258 5926 6286
rect 5954 6258 5978 6286
rect 6006 6258 6030 6286
rect 6058 6258 6063 6286
rect 8581 6258 8586 6286
rect 8614 6258 8638 6286
rect 8666 6258 8690 6286
rect 8718 6258 8723 6286
rect 11241 6258 11246 6286
rect 11274 6258 11298 6286
rect 11326 6258 11350 6286
rect 11378 6258 11383 6286
rect 2193 6174 2198 6202
rect 2226 6174 2231 6202
rect 3145 6174 3150 6202
rect 3178 6174 3822 6202
rect 3850 6174 4942 6202
rect 4970 6174 4975 6202
rect 2198 6090 2226 6174
rect 3929 6118 3934 6146
rect 3962 6118 5110 6146
rect 5138 6118 5143 6146
rect 9529 6118 9534 6146
rect 9562 6118 9814 6146
rect 9842 6118 9847 6146
rect 2198 6062 4382 6090
rect 4410 6062 4415 6090
rect 5049 6062 5054 6090
rect 5082 6062 9254 6090
rect 9282 6062 9287 6090
rect 2025 6006 2030 6034
rect 2058 6006 2702 6034
rect 2730 6006 2735 6034
rect 9641 5950 9646 5978
rect 9674 5950 9758 5978
rect 9786 5950 9791 5978
rect 1931 5866 1936 5894
rect 1964 5866 1988 5894
rect 2016 5866 2040 5894
rect 2068 5866 2073 5894
rect 4591 5866 4596 5894
rect 4624 5866 4648 5894
rect 4676 5866 4700 5894
rect 4728 5866 4733 5894
rect 7251 5866 7256 5894
rect 7284 5866 7308 5894
rect 7336 5866 7360 5894
rect 7388 5866 7393 5894
rect 9911 5866 9916 5894
rect 9944 5866 9968 5894
rect 9996 5866 10020 5894
rect 10048 5866 10053 5894
rect 10089 5838 10094 5866
rect 10122 5838 10934 5866
rect 10962 5838 10967 5866
rect 10033 5782 10038 5810
rect 10066 5782 10990 5810
rect 11018 5782 11023 5810
rect 4433 5726 4438 5754
rect 4466 5726 4942 5754
rect 4970 5726 4975 5754
rect 5105 5726 5110 5754
rect 5138 5726 7574 5754
rect 2361 5670 2366 5698
rect 2394 5670 4606 5698
rect 4634 5670 4886 5698
rect 4914 5670 4919 5698
rect 5217 5670 5222 5698
rect 5250 5670 6118 5698
rect 6146 5670 6151 5698
rect 4545 5614 4550 5642
rect 4578 5614 4583 5642
rect 4993 5614 4998 5642
rect 5026 5614 6734 5642
rect 6762 5614 7182 5642
rect 7210 5614 7215 5642
rect 7546 5614 7574 5726
rect 7602 5614 7607 5642
rect 7681 5614 7686 5642
rect 7714 5614 9198 5642
rect 9226 5614 9231 5642
rect 4550 5586 4578 5614
rect 4550 5558 10318 5586
rect 10346 5558 10351 5586
rect 3261 5474 3266 5502
rect 3294 5474 3318 5502
rect 3346 5474 3370 5502
rect 3398 5474 3403 5502
rect 5921 5474 5926 5502
rect 5954 5474 5978 5502
rect 6006 5474 6030 5502
rect 6058 5474 6063 5502
rect 8581 5474 8586 5502
rect 8614 5474 8638 5502
rect 8666 5474 8690 5502
rect 8718 5474 8723 5502
rect 11241 5474 11246 5502
rect 11274 5474 11298 5502
rect 11326 5474 11350 5502
rect 11378 5474 11383 5502
rect 9473 5446 9478 5474
rect 9506 5446 10206 5474
rect 10234 5446 10239 5474
rect 4545 5334 4550 5362
rect 4578 5334 6454 5362
rect 6482 5334 6487 5362
rect 7681 5334 7686 5362
rect 7714 5334 10094 5362
rect 10122 5334 10127 5362
rect 1129 5278 1134 5306
rect 1162 5278 1638 5306
rect 1666 5278 4102 5306
rect 4130 5278 4270 5306
rect 4298 5278 4303 5306
rect 6561 5278 6566 5306
rect 6594 5278 7294 5306
rect 7322 5278 7327 5306
rect 7457 5278 7462 5306
rect 7490 5278 7910 5306
rect 7938 5278 7943 5306
rect 9193 5278 9198 5306
rect 9226 5278 9646 5306
rect 9674 5278 9679 5306
rect 9361 5222 9366 5250
rect 9394 5222 9702 5250
rect 9730 5222 9735 5250
rect 11600 5194 12000 5208
rect 5497 5166 5502 5194
rect 5530 5166 6510 5194
rect 6538 5166 6543 5194
rect 6841 5166 6846 5194
rect 6874 5166 7574 5194
rect 7602 5166 9254 5194
rect 9282 5166 9646 5194
rect 9674 5166 9679 5194
rect 10817 5166 10822 5194
rect 10850 5166 11102 5194
rect 11130 5166 12000 5194
rect 11600 5152 12000 5166
rect 1931 5082 1936 5110
rect 1964 5082 1988 5110
rect 2016 5082 2040 5110
rect 2068 5082 2073 5110
rect 4591 5082 4596 5110
rect 4624 5082 4648 5110
rect 4676 5082 4700 5110
rect 4728 5082 4733 5110
rect 7251 5082 7256 5110
rect 7284 5082 7308 5110
rect 7336 5082 7360 5110
rect 7388 5082 7393 5110
rect 9911 5082 9916 5110
rect 9944 5082 9968 5110
rect 9996 5082 10020 5110
rect 10048 5082 10053 5110
rect 7457 5054 7462 5082
rect 7490 5054 7798 5082
rect 7826 5054 9590 5082
rect 9618 5054 9623 5082
rect 1297 4998 1302 5026
rect 1330 4998 2170 5026
rect 2142 4914 2170 4998
rect 4209 4942 4214 4970
rect 4242 4942 4606 4970
rect 4634 4942 7574 4970
rect 7602 4942 7854 4970
rect 7882 4942 7887 4970
rect 9697 4942 9702 4970
rect 9730 4942 9926 4970
rect 9954 4942 9959 4970
rect 2137 4886 2142 4914
rect 2170 4886 4942 4914
rect 4970 4886 5390 4914
rect 5418 4886 5423 4914
rect 7961 4886 7966 4914
rect 7994 4886 9366 4914
rect 9394 4886 9982 4914
rect 10010 4886 10015 4914
rect 4545 4830 4550 4858
rect 4578 4830 5166 4858
rect 5194 4830 6958 4858
rect 6986 4830 6991 4858
rect 4769 4774 4774 4802
rect 4802 4774 5278 4802
rect 5306 4774 5311 4802
rect 5385 4774 5390 4802
rect 5418 4774 7350 4802
rect 7378 4774 7383 4802
rect 3261 4690 3266 4718
rect 3294 4690 3318 4718
rect 3346 4690 3370 4718
rect 3398 4690 3403 4718
rect 5921 4690 5926 4718
rect 5954 4690 5978 4718
rect 6006 4690 6030 4718
rect 6058 4690 6063 4718
rect 8581 4690 8586 4718
rect 8614 4690 8638 4718
rect 8666 4690 8690 4718
rect 8718 4690 8723 4718
rect 11241 4690 11246 4718
rect 11274 4690 11298 4718
rect 11326 4690 11350 4718
rect 11378 4690 11383 4718
rect 4321 4606 4326 4634
rect 4354 4606 7350 4634
rect 7378 4606 7383 4634
rect 5217 4550 5222 4578
rect 5250 4550 5446 4578
rect 5474 4550 5479 4578
rect 1689 4494 1694 4522
rect 1722 4494 1918 4522
rect 1946 4494 2478 4522
rect 2506 4494 3430 4522
rect 3458 4494 3463 4522
rect 9473 4494 9478 4522
rect 9506 4494 9702 4522
rect 9730 4494 9735 4522
rect 9590 4466 9618 4494
rect 9585 4438 9590 4466
rect 9618 4438 9623 4466
rect 1931 4298 1936 4326
rect 1964 4298 1988 4326
rect 2016 4298 2040 4326
rect 2068 4298 2073 4326
rect 4591 4298 4596 4326
rect 4624 4298 4648 4326
rect 4676 4298 4700 4326
rect 4728 4298 4733 4326
rect 7251 4298 7256 4326
rect 7284 4298 7308 4326
rect 7336 4298 7360 4326
rect 7388 4298 7393 4326
rect 9911 4298 9916 4326
rect 9944 4298 9968 4326
rect 9996 4298 10020 4326
rect 10048 4298 10053 4326
rect 4657 4214 4662 4242
rect 4690 4214 5334 4242
rect 5362 4214 5367 4242
rect 2137 4158 2142 4186
rect 2170 4158 2870 4186
rect 2898 4158 2903 4186
rect 3201 4158 3206 4186
rect 3234 4158 3710 4186
rect 3738 4158 4438 4186
rect 4466 4158 4471 4186
rect 5049 4158 5054 4186
rect 5082 4158 5726 4186
rect 5754 4158 5759 4186
rect 1577 4102 1582 4130
rect 1610 4102 1918 4130
rect 1946 4102 1951 4130
rect 2697 4102 2702 4130
rect 2730 4102 3654 4130
rect 3682 4102 3687 4130
rect 3817 4102 3822 4130
rect 3850 4102 4998 4130
rect 5026 4102 5031 4130
rect 7681 4102 7686 4130
rect 7714 4102 9534 4130
rect 9562 4102 9567 4130
rect 3145 4046 3150 4074
rect 3178 4046 4830 4074
rect 4858 4046 4863 4074
rect 5105 4046 5110 4074
rect 5138 4046 5614 4074
rect 5642 4046 5647 4074
rect 7457 4046 7462 4074
rect 7490 4046 7574 4074
rect 9305 4046 9310 4074
rect 9338 4046 9870 4074
rect 9898 4046 9903 4074
rect 10089 4046 10094 4074
rect 10122 4046 10934 4074
rect 10962 4046 10967 4074
rect 7546 4018 7574 4046
rect 2081 3990 2086 4018
rect 2114 3990 2422 4018
rect 2450 3990 2814 4018
rect 2842 3990 2847 4018
rect 2977 3990 2982 4018
rect 3010 3990 5334 4018
rect 5362 3990 5367 4018
rect 7546 3990 7910 4018
rect 7938 3990 10318 4018
rect 10346 3990 10766 4018
rect 10794 3990 10799 4018
rect 2982 3794 3010 3990
rect 4881 3934 4886 3962
rect 4914 3934 5054 3962
rect 5082 3934 5087 3962
rect 3261 3906 3266 3934
rect 3294 3906 3318 3934
rect 3346 3906 3370 3934
rect 3398 3906 3403 3934
rect 5921 3906 5926 3934
rect 5954 3906 5978 3934
rect 6006 3906 6030 3934
rect 6058 3906 6063 3934
rect 8581 3906 8586 3934
rect 8614 3906 8638 3934
rect 8666 3906 8690 3934
rect 8718 3906 8723 3934
rect 11241 3906 11246 3934
rect 11274 3906 11298 3934
rect 11326 3906 11350 3934
rect 11378 3906 11383 3934
rect 4433 3822 4438 3850
rect 4466 3822 5054 3850
rect 5082 3822 5087 3850
rect 5217 3822 5222 3850
rect 5250 3822 7574 3850
rect 7546 3794 7574 3822
rect 2641 3766 2646 3794
rect 2674 3766 3010 3794
rect 5105 3766 5110 3794
rect 5138 3766 5558 3794
rect 5586 3766 5591 3794
rect 7546 3766 9366 3794
rect 9394 3766 9982 3794
rect 10010 3766 10015 3794
rect 11600 3738 12000 3752
rect 5497 3710 5502 3738
rect 5530 3710 7294 3738
rect 7322 3710 7327 3738
rect 9809 3710 9814 3738
rect 9842 3710 10150 3738
rect 10178 3710 10374 3738
rect 10402 3710 10934 3738
rect 10962 3710 10967 3738
rect 11097 3710 11102 3738
rect 11130 3710 12000 3738
rect 11600 3696 12000 3710
rect 2361 3598 2366 3626
rect 2394 3598 2870 3626
rect 2898 3598 9590 3626
rect 9618 3598 9623 3626
rect 1931 3514 1936 3542
rect 1964 3514 1988 3542
rect 2016 3514 2040 3542
rect 2068 3514 2073 3542
rect 4591 3514 4596 3542
rect 4624 3514 4648 3542
rect 4676 3514 4700 3542
rect 4728 3514 4733 3542
rect 7251 3514 7256 3542
rect 7284 3514 7308 3542
rect 7336 3514 7360 3542
rect 7388 3514 7393 3542
rect 9911 3514 9916 3542
rect 9944 3514 9968 3542
rect 9996 3514 10020 3542
rect 10048 3514 10053 3542
rect 9809 3430 9814 3458
rect 9842 3430 10318 3458
rect 10346 3430 10351 3458
rect 5553 3374 5558 3402
rect 5586 3374 7406 3402
rect 7434 3374 7630 3402
rect 7658 3374 7910 3402
rect 7938 3374 7943 3402
rect 3261 3122 3266 3150
rect 3294 3122 3318 3150
rect 3346 3122 3370 3150
rect 3398 3122 3403 3150
rect 5921 3122 5926 3150
rect 5954 3122 5978 3150
rect 6006 3122 6030 3150
rect 6058 3122 6063 3150
rect 8581 3122 8586 3150
rect 8614 3122 8638 3150
rect 8666 3122 8690 3150
rect 8718 3122 8723 3150
rect 11241 3122 11246 3150
rect 11274 3122 11298 3150
rect 11326 3122 11350 3150
rect 11378 3122 11383 3150
rect 1931 2730 1936 2758
rect 1964 2730 1988 2758
rect 2016 2730 2040 2758
rect 2068 2730 2073 2758
rect 4591 2730 4596 2758
rect 4624 2730 4648 2758
rect 4676 2730 4700 2758
rect 4728 2730 4733 2758
rect 7251 2730 7256 2758
rect 7284 2730 7308 2758
rect 7336 2730 7360 2758
rect 7388 2730 7393 2758
rect 9911 2730 9916 2758
rect 9944 2730 9968 2758
rect 9996 2730 10020 2758
rect 10048 2730 10053 2758
rect 10817 2534 10822 2562
rect 10850 2534 11102 2562
rect 11130 2534 11135 2562
rect 3261 2338 3266 2366
rect 3294 2338 3318 2366
rect 3346 2338 3370 2366
rect 3398 2338 3403 2366
rect 5921 2338 5926 2366
rect 5954 2338 5978 2366
rect 6006 2338 6030 2366
rect 6058 2338 6063 2366
rect 8581 2338 8586 2366
rect 8614 2338 8638 2366
rect 8666 2338 8690 2366
rect 8718 2338 8723 2366
rect 11241 2338 11246 2366
rect 11274 2338 11298 2366
rect 11326 2338 11350 2366
rect 11378 2338 11383 2366
rect 11600 2282 12000 2296
rect 11097 2254 11102 2282
rect 11130 2254 12000 2282
rect 11600 2240 12000 2254
rect 1931 1946 1936 1974
rect 1964 1946 1988 1974
rect 2016 1946 2040 1974
rect 2068 1946 2073 1974
rect 4591 1946 4596 1974
rect 4624 1946 4648 1974
rect 4676 1946 4700 1974
rect 4728 1946 4733 1974
rect 7251 1946 7256 1974
rect 7284 1946 7308 1974
rect 7336 1946 7360 1974
rect 7388 1946 7393 1974
rect 9911 1946 9916 1974
rect 9944 1946 9968 1974
rect 9996 1946 10020 1974
rect 10048 1946 10053 1974
rect 3261 1554 3266 1582
rect 3294 1554 3318 1582
rect 3346 1554 3370 1582
rect 3398 1554 3403 1582
rect 5921 1554 5926 1582
rect 5954 1554 5978 1582
rect 6006 1554 6030 1582
rect 6058 1554 6063 1582
rect 8581 1554 8586 1582
rect 8614 1554 8638 1582
rect 8666 1554 8690 1582
rect 8718 1554 8723 1582
rect 11241 1554 11246 1582
rect 11274 1554 11298 1582
rect 11326 1554 11350 1582
rect 11378 1554 11383 1582
rect 11600 826 12000 840
rect 9809 798 9814 826
rect 9842 798 12000 826
rect 11600 784 12000 798
<< via3 >>
rect 3266 10178 3294 10206
rect 3318 10178 3346 10206
rect 3370 10178 3398 10206
rect 5926 10178 5954 10206
rect 5978 10178 6006 10206
rect 6030 10178 6058 10206
rect 8586 10178 8614 10206
rect 8638 10178 8666 10206
rect 8690 10178 8718 10206
rect 11246 10178 11274 10206
rect 11298 10178 11326 10206
rect 11350 10178 11378 10206
rect 1936 9786 1964 9814
rect 1988 9786 2016 9814
rect 2040 9786 2068 9814
rect 4596 9786 4624 9814
rect 4648 9786 4676 9814
rect 4700 9786 4728 9814
rect 7256 9786 7284 9814
rect 7308 9786 7336 9814
rect 7360 9786 7388 9814
rect 9916 9786 9944 9814
rect 9968 9786 9996 9814
rect 10020 9786 10048 9814
rect 3266 9394 3294 9422
rect 3318 9394 3346 9422
rect 3370 9394 3398 9422
rect 5926 9394 5954 9422
rect 5978 9394 6006 9422
rect 6030 9394 6058 9422
rect 8586 9394 8614 9422
rect 8638 9394 8666 9422
rect 8690 9394 8718 9422
rect 11246 9394 11274 9422
rect 11298 9394 11326 9422
rect 11350 9394 11378 9422
rect 2198 9198 2226 9226
rect 1936 9002 1964 9030
rect 1988 9002 2016 9030
rect 2040 9002 2068 9030
rect 4596 9002 4624 9030
rect 4648 9002 4676 9030
rect 4700 9002 4728 9030
rect 7256 9002 7284 9030
rect 7308 9002 7336 9030
rect 7360 9002 7388 9030
rect 9916 9002 9944 9030
rect 9968 9002 9996 9030
rect 10020 9002 10048 9030
rect 3266 8610 3294 8638
rect 3318 8610 3346 8638
rect 3370 8610 3398 8638
rect 5926 8610 5954 8638
rect 5978 8610 6006 8638
rect 6030 8610 6058 8638
rect 8586 8610 8614 8638
rect 8638 8610 8666 8638
rect 8690 8610 8718 8638
rect 11246 8610 11274 8638
rect 11298 8610 11326 8638
rect 11350 8610 11378 8638
rect 10094 8414 10122 8442
rect 1936 8218 1964 8246
rect 1988 8218 2016 8246
rect 2040 8218 2068 8246
rect 4596 8218 4624 8246
rect 4648 8218 4676 8246
rect 4700 8218 4728 8246
rect 7256 8218 7284 8246
rect 7308 8218 7336 8246
rect 7360 8218 7388 8246
rect 9916 8218 9944 8246
rect 9968 8218 9996 8246
rect 10020 8218 10048 8246
rect 3266 7826 3294 7854
rect 3318 7826 3346 7854
rect 3370 7826 3398 7854
rect 5926 7826 5954 7854
rect 5978 7826 6006 7854
rect 6030 7826 6058 7854
rect 8586 7826 8614 7854
rect 8638 7826 8666 7854
rect 8690 7826 8718 7854
rect 11246 7826 11274 7854
rect 11298 7826 11326 7854
rect 11350 7826 11378 7854
rect 10094 7518 10122 7546
rect 1936 7434 1964 7462
rect 1988 7434 2016 7462
rect 2040 7434 2068 7462
rect 4596 7434 4624 7462
rect 4648 7434 4676 7462
rect 4700 7434 4728 7462
rect 7256 7434 7284 7462
rect 7308 7434 7336 7462
rect 7360 7434 7388 7462
rect 9916 7434 9944 7462
rect 9968 7434 9996 7462
rect 10020 7434 10048 7462
rect 2198 7126 2226 7154
rect 3266 7042 3294 7070
rect 3318 7042 3346 7070
rect 3370 7042 3398 7070
rect 5926 7042 5954 7070
rect 5978 7042 6006 7070
rect 6030 7042 6058 7070
rect 8586 7042 8614 7070
rect 8638 7042 8666 7070
rect 8690 7042 8718 7070
rect 11246 7042 11274 7070
rect 11298 7042 11326 7070
rect 11350 7042 11378 7070
rect 9758 7014 9786 7042
rect 9814 6846 9842 6874
rect 1936 6650 1964 6678
rect 1988 6650 2016 6678
rect 2040 6650 2068 6678
rect 4596 6650 4624 6678
rect 4648 6650 4676 6678
rect 4700 6650 4728 6678
rect 7256 6650 7284 6678
rect 7308 6650 7336 6678
rect 7360 6650 7388 6678
rect 9916 6650 9944 6678
rect 9968 6650 9996 6678
rect 10020 6650 10048 6678
rect 3266 6258 3294 6286
rect 3318 6258 3346 6286
rect 3370 6258 3398 6286
rect 5926 6258 5954 6286
rect 5978 6258 6006 6286
rect 6030 6258 6058 6286
rect 8586 6258 8614 6286
rect 8638 6258 8666 6286
rect 8690 6258 8718 6286
rect 11246 6258 11274 6286
rect 11298 6258 11326 6286
rect 11350 6258 11378 6286
rect 9814 6118 9842 6146
rect 9758 5950 9786 5978
rect 1936 5866 1964 5894
rect 1988 5866 2016 5894
rect 2040 5866 2068 5894
rect 4596 5866 4624 5894
rect 4648 5866 4676 5894
rect 4700 5866 4728 5894
rect 7256 5866 7284 5894
rect 7308 5866 7336 5894
rect 7360 5866 7388 5894
rect 9916 5866 9944 5894
rect 9968 5866 9996 5894
rect 10020 5866 10048 5894
rect 3266 5474 3294 5502
rect 3318 5474 3346 5502
rect 3370 5474 3398 5502
rect 5926 5474 5954 5502
rect 5978 5474 6006 5502
rect 6030 5474 6058 5502
rect 8586 5474 8614 5502
rect 8638 5474 8666 5502
rect 8690 5474 8718 5502
rect 11246 5474 11274 5502
rect 11298 5474 11326 5502
rect 11350 5474 11378 5502
rect 1936 5082 1964 5110
rect 1988 5082 2016 5110
rect 2040 5082 2068 5110
rect 4596 5082 4624 5110
rect 4648 5082 4676 5110
rect 4700 5082 4728 5110
rect 7256 5082 7284 5110
rect 7308 5082 7336 5110
rect 7360 5082 7388 5110
rect 9916 5082 9944 5110
rect 9968 5082 9996 5110
rect 10020 5082 10048 5110
rect 3266 4690 3294 4718
rect 3318 4690 3346 4718
rect 3370 4690 3398 4718
rect 5926 4690 5954 4718
rect 5978 4690 6006 4718
rect 6030 4690 6058 4718
rect 8586 4690 8614 4718
rect 8638 4690 8666 4718
rect 8690 4690 8718 4718
rect 11246 4690 11274 4718
rect 11298 4690 11326 4718
rect 11350 4690 11378 4718
rect 1936 4298 1964 4326
rect 1988 4298 2016 4326
rect 2040 4298 2068 4326
rect 4596 4298 4624 4326
rect 4648 4298 4676 4326
rect 4700 4298 4728 4326
rect 7256 4298 7284 4326
rect 7308 4298 7336 4326
rect 7360 4298 7388 4326
rect 9916 4298 9944 4326
rect 9968 4298 9996 4326
rect 10020 4298 10048 4326
rect 3266 3906 3294 3934
rect 3318 3906 3346 3934
rect 3370 3906 3398 3934
rect 5926 3906 5954 3934
rect 5978 3906 6006 3934
rect 6030 3906 6058 3934
rect 8586 3906 8614 3934
rect 8638 3906 8666 3934
rect 8690 3906 8718 3934
rect 11246 3906 11274 3934
rect 11298 3906 11326 3934
rect 11350 3906 11378 3934
rect 1936 3514 1964 3542
rect 1988 3514 2016 3542
rect 2040 3514 2068 3542
rect 4596 3514 4624 3542
rect 4648 3514 4676 3542
rect 4700 3514 4728 3542
rect 7256 3514 7284 3542
rect 7308 3514 7336 3542
rect 7360 3514 7388 3542
rect 9916 3514 9944 3542
rect 9968 3514 9996 3542
rect 10020 3514 10048 3542
rect 3266 3122 3294 3150
rect 3318 3122 3346 3150
rect 3370 3122 3398 3150
rect 5926 3122 5954 3150
rect 5978 3122 6006 3150
rect 6030 3122 6058 3150
rect 8586 3122 8614 3150
rect 8638 3122 8666 3150
rect 8690 3122 8718 3150
rect 11246 3122 11274 3150
rect 11298 3122 11326 3150
rect 11350 3122 11378 3150
rect 1936 2730 1964 2758
rect 1988 2730 2016 2758
rect 2040 2730 2068 2758
rect 4596 2730 4624 2758
rect 4648 2730 4676 2758
rect 4700 2730 4728 2758
rect 7256 2730 7284 2758
rect 7308 2730 7336 2758
rect 7360 2730 7388 2758
rect 9916 2730 9944 2758
rect 9968 2730 9996 2758
rect 10020 2730 10048 2758
rect 3266 2338 3294 2366
rect 3318 2338 3346 2366
rect 3370 2338 3398 2366
rect 5926 2338 5954 2366
rect 5978 2338 6006 2366
rect 6030 2338 6058 2366
rect 8586 2338 8614 2366
rect 8638 2338 8666 2366
rect 8690 2338 8718 2366
rect 11246 2338 11274 2366
rect 11298 2338 11326 2366
rect 11350 2338 11378 2366
rect 1936 1946 1964 1974
rect 1988 1946 2016 1974
rect 2040 1946 2068 1974
rect 4596 1946 4624 1974
rect 4648 1946 4676 1974
rect 4700 1946 4728 1974
rect 7256 1946 7284 1974
rect 7308 1946 7336 1974
rect 7360 1946 7388 1974
rect 9916 1946 9944 1974
rect 9968 1946 9996 1974
rect 10020 1946 10048 1974
rect 3266 1554 3294 1582
rect 3318 1554 3346 1582
rect 3370 1554 3398 1582
rect 5926 1554 5954 1582
rect 5978 1554 6006 1582
rect 6030 1554 6058 1582
rect 8586 1554 8614 1582
rect 8638 1554 8666 1582
rect 8690 1554 8718 1582
rect 11246 1554 11274 1582
rect 11298 1554 11326 1582
rect 11350 1554 11378 1582
<< metal4 >>
rect 1922 9814 2082 10222
rect 1922 9786 1936 9814
rect 1964 9786 1988 9814
rect 2016 9786 2040 9814
rect 2068 9786 2082 9814
rect 1922 9030 2082 9786
rect 3252 10206 3412 10222
rect 3252 10178 3266 10206
rect 3294 10178 3318 10206
rect 3346 10178 3370 10206
rect 3398 10178 3412 10206
rect 3252 9422 3412 10178
rect 3252 9394 3266 9422
rect 3294 9394 3318 9422
rect 3346 9394 3370 9422
rect 3398 9394 3412 9422
rect 1922 9002 1936 9030
rect 1964 9002 1988 9030
rect 2016 9002 2040 9030
rect 2068 9002 2082 9030
rect 1922 8246 2082 9002
rect 1922 8218 1936 8246
rect 1964 8218 1988 8246
rect 2016 8218 2040 8246
rect 2068 8218 2082 8246
rect 1922 7462 2082 8218
rect 1922 7434 1936 7462
rect 1964 7434 1988 7462
rect 2016 7434 2040 7462
rect 2068 7434 2082 7462
rect 1922 6678 2082 7434
rect 2198 9226 2226 9231
rect 2198 7154 2226 9198
rect 2198 7121 2226 7126
rect 3252 8638 3412 9394
rect 3252 8610 3266 8638
rect 3294 8610 3318 8638
rect 3346 8610 3370 8638
rect 3398 8610 3412 8638
rect 3252 7854 3412 8610
rect 3252 7826 3266 7854
rect 3294 7826 3318 7854
rect 3346 7826 3370 7854
rect 3398 7826 3412 7854
rect 1922 6650 1936 6678
rect 1964 6650 1988 6678
rect 2016 6650 2040 6678
rect 2068 6650 2082 6678
rect 1922 5894 2082 6650
rect 1922 5866 1936 5894
rect 1964 5866 1988 5894
rect 2016 5866 2040 5894
rect 2068 5866 2082 5894
rect 1922 5110 2082 5866
rect 1922 5082 1936 5110
rect 1964 5082 1988 5110
rect 2016 5082 2040 5110
rect 2068 5082 2082 5110
rect 1922 4326 2082 5082
rect 1922 4298 1936 4326
rect 1964 4298 1988 4326
rect 2016 4298 2040 4326
rect 2068 4298 2082 4326
rect 1922 3542 2082 4298
rect 1922 3514 1936 3542
rect 1964 3514 1988 3542
rect 2016 3514 2040 3542
rect 2068 3514 2082 3542
rect 1922 2758 2082 3514
rect 1922 2730 1936 2758
rect 1964 2730 1988 2758
rect 2016 2730 2040 2758
rect 2068 2730 2082 2758
rect 1922 1974 2082 2730
rect 1922 1946 1936 1974
rect 1964 1946 1988 1974
rect 2016 1946 2040 1974
rect 2068 1946 2082 1974
rect 1922 1538 2082 1946
rect 3252 7070 3412 7826
rect 3252 7042 3266 7070
rect 3294 7042 3318 7070
rect 3346 7042 3370 7070
rect 3398 7042 3412 7070
rect 3252 6286 3412 7042
rect 3252 6258 3266 6286
rect 3294 6258 3318 6286
rect 3346 6258 3370 6286
rect 3398 6258 3412 6286
rect 3252 5502 3412 6258
rect 3252 5474 3266 5502
rect 3294 5474 3318 5502
rect 3346 5474 3370 5502
rect 3398 5474 3412 5502
rect 3252 4718 3412 5474
rect 3252 4690 3266 4718
rect 3294 4690 3318 4718
rect 3346 4690 3370 4718
rect 3398 4690 3412 4718
rect 3252 3934 3412 4690
rect 3252 3906 3266 3934
rect 3294 3906 3318 3934
rect 3346 3906 3370 3934
rect 3398 3906 3412 3934
rect 3252 3150 3412 3906
rect 3252 3122 3266 3150
rect 3294 3122 3318 3150
rect 3346 3122 3370 3150
rect 3398 3122 3412 3150
rect 3252 2366 3412 3122
rect 3252 2338 3266 2366
rect 3294 2338 3318 2366
rect 3346 2338 3370 2366
rect 3398 2338 3412 2366
rect 3252 1582 3412 2338
rect 3252 1554 3266 1582
rect 3294 1554 3318 1582
rect 3346 1554 3370 1582
rect 3398 1554 3412 1582
rect 3252 1538 3412 1554
rect 4582 9814 4742 10222
rect 4582 9786 4596 9814
rect 4624 9786 4648 9814
rect 4676 9786 4700 9814
rect 4728 9786 4742 9814
rect 4582 9030 4742 9786
rect 4582 9002 4596 9030
rect 4624 9002 4648 9030
rect 4676 9002 4700 9030
rect 4728 9002 4742 9030
rect 4582 8246 4742 9002
rect 4582 8218 4596 8246
rect 4624 8218 4648 8246
rect 4676 8218 4700 8246
rect 4728 8218 4742 8246
rect 4582 7462 4742 8218
rect 4582 7434 4596 7462
rect 4624 7434 4648 7462
rect 4676 7434 4700 7462
rect 4728 7434 4742 7462
rect 4582 6678 4742 7434
rect 4582 6650 4596 6678
rect 4624 6650 4648 6678
rect 4676 6650 4700 6678
rect 4728 6650 4742 6678
rect 4582 5894 4742 6650
rect 4582 5866 4596 5894
rect 4624 5866 4648 5894
rect 4676 5866 4700 5894
rect 4728 5866 4742 5894
rect 4582 5110 4742 5866
rect 4582 5082 4596 5110
rect 4624 5082 4648 5110
rect 4676 5082 4700 5110
rect 4728 5082 4742 5110
rect 4582 4326 4742 5082
rect 4582 4298 4596 4326
rect 4624 4298 4648 4326
rect 4676 4298 4700 4326
rect 4728 4298 4742 4326
rect 4582 3542 4742 4298
rect 4582 3514 4596 3542
rect 4624 3514 4648 3542
rect 4676 3514 4700 3542
rect 4728 3514 4742 3542
rect 4582 2758 4742 3514
rect 4582 2730 4596 2758
rect 4624 2730 4648 2758
rect 4676 2730 4700 2758
rect 4728 2730 4742 2758
rect 4582 1974 4742 2730
rect 4582 1946 4596 1974
rect 4624 1946 4648 1974
rect 4676 1946 4700 1974
rect 4728 1946 4742 1974
rect 4582 1538 4742 1946
rect 5912 10206 6072 10222
rect 5912 10178 5926 10206
rect 5954 10178 5978 10206
rect 6006 10178 6030 10206
rect 6058 10178 6072 10206
rect 5912 9422 6072 10178
rect 5912 9394 5926 9422
rect 5954 9394 5978 9422
rect 6006 9394 6030 9422
rect 6058 9394 6072 9422
rect 5912 8638 6072 9394
rect 5912 8610 5926 8638
rect 5954 8610 5978 8638
rect 6006 8610 6030 8638
rect 6058 8610 6072 8638
rect 5912 7854 6072 8610
rect 5912 7826 5926 7854
rect 5954 7826 5978 7854
rect 6006 7826 6030 7854
rect 6058 7826 6072 7854
rect 5912 7070 6072 7826
rect 5912 7042 5926 7070
rect 5954 7042 5978 7070
rect 6006 7042 6030 7070
rect 6058 7042 6072 7070
rect 5912 6286 6072 7042
rect 5912 6258 5926 6286
rect 5954 6258 5978 6286
rect 6006 6258 6030 6286
rect 6058 6258 6072 6286
rect 5912 5502 6072 6258
rect 5912 5474 5926 5502
rect 5954 5474 5978 5502
rect 6006 5474 6030 5502
rect 6058 5474 6072 5502
rect 5912 4718 6072 5474
rect 5912 4690 5926 4718
rect 5954 4690 5978 4718
rect 6006 4690 6030 4718
rect 6058 4690 6072 4718
rect 5912 3934 6072 4690
rect 5912 3906 5926 3934
rect 5954 3906 5978 3934
rect 6006 3906 6030 3934
rect 6058 3906 6072 3934
rect 5912 3150 6072 3906
rect 5912 3122 5926 3150
rect 5954 3122 5978 3150
rect 6006 3122 6030 3150
rect 6058 3122 6072 3150
rect 5912 2366 6072 3122
rect 5912 2338 5926 2366
rect 5954 2338 5978 2366
rect 6006 2338 6030 2366
rect 6058 2338 6072 2366
rect 5912 1582 6072 2338
rect 5912 1554 5926 1582
rect 5954 1554 5978 1582
rect 6006 1554 6030 1582
rect 6058 1554 6072 1582
rect 5912 1538 6072 1554
rect 7242 9814 7402 10222
rect 7242 9786 7256 9814
rect 7284 9786 7308 9814
rect 7336 9786 7360 9814
rect 7388 9786 7402 9814
rect 7242 9030 7402 9786
rect 7242 9002 7256 9030
rect 7284 9002 7308 9030
rect 7336 9002 7360 9030
rect 7388 9002 7402 9030
rect 7242 8246 7402 9002
rect 7242 8218 7256 8246
rect 7284 8218 7308 8246
rect 7336 8218 7360 8246
rect 7388 8218 7402 8246
rect 7242 7462 7402 8218
rect 7242 7434 7256 7462
rect 7284 7434 7308 7462
rect 7336 7434 7360 7462
rect 7388 7434 7402 7462
rect 7242 6678 7402 7434
rect 7242 6650 7256 6678
rect 7284 6650 7308 6678
rect 7336 6650 7360 6678
rect 7388 6650 7402 6678
rect 7242 5894 7402 6650
rect 7242 5866 7256 5894
rect 7284 5866 7308 5894
rect 7336 5866 7360 5894
rect 7388 5866 7402 5894
rect 7242 5110 7402 5866
rect 7242 5082 7256 5110
rect 7284 5082 7308 5110
rect 7336 5082 7360 5110
rect 7388 5082 7402 5110
rect 7242 4326 7402 5082
rect 7242 4298 7256 4326
rect 7284 4298 7308 4326
rect 7336 4298 7360 4326
rect 7388 4298 7402 4326
rect 7242 3542 7402 4298
rect 7242 3514 7256 3542
rect 7284 3514 7308 3542
rect 7336 3514 7360 3542
rect 7388 3514 7402 3542
rect 7242 2758 7402 3514
rect 7242 2730 7256 2758
rect 7284 2730 7308 2758
rect 7336 2730 7360 2758
rect 7388 2730 7402 2758
rect 7242 1974 7402 2730
rect 7242 1946 7256 1974
rect 7284 1946 7308 1974
rect 7336 1946 7360 1974
rect 7388 1946 7402 1974
rect 7242 1538 7402 1946
rect 8572 10206 8732 10222
rect 8572 10178 8586 10206
rect 8614 10178 8638 10206
rect 8666 10178 8690 10206
rect 8718 10178 8732 10206
rect 8572 9422 8732 10178
rect 8572 9394 8586 9422
rect 8614 9394 8638 9422
rect 8666 9394 8690 9422
rect 8718 9394 8732 9422
rect 8572 8638 8732 9394
rect 8572 8610 8586 8638
rect 8614 8610 8638 8638
rect 8666 8610 8690 8638
rect 8718 8610 8732 8638
rect 8572 7854 8732 8610
rect 8572 7826 8586 7854
rect 8614 7826 8638 7854
rect 8666 7826 8690 7854
rect 8718 7826 8732 7854
rect 8572 7070 8732 7826
rect 8572 7042 8586 7070
rect 8614 7042 8638 7070
rect 8666 7042 8690 7070
rect 8718 7042 8732 7070
rect 9902 9814 10062 10222
rect 9902 9786 9916 9814
rect 9944 9786 9968 9814
rect 9996 9786 10020 9814
rect 10048 9786 10062 9814
rect 9902 9030 10062 9786
rect 9902 9002 9916 9030
rect 9944 9002 9968 9030
rect 9996 9002 10020 9030
rect 10048 9002 10062 9030
rect 9902 8246 10062 9002
rect 11232 10206 11392 10222
rect 11232 10178 11246 10206
rect 11274 10178 11298 10206
rect 11326 10178 11350 10206
rect 11378 10178 11392 10206
rect 11232 9422 11392 10178
rect 11232 9394 11246 9422
rect 11274 9394 11298 9422
rect 11326 9394 11350 9422
rect 11378 9394 11392 9422
rect 11232 8638 11392 9394
rect 11232 8610 11246 8638
rect 11274 8610 11298 8638
rect 11326 8610 11350 8638
rect 11378 8610 11392 8638
rect 9902 8218 9916 8246
rect 9944 8218 9968 8246
rect 9996 8218 10020 8246
rect 10048 8218 10062 8246
rect 9902 7462 10062 8218
rect 10094 8442 10122 8447
rect 10094 7546 10122 8414
rect 10094 7513 10122 7518
rect 11232 7854 11392 8610
rect 11232 7826 11246 7854
rect 11274 7826 11298 7854
rect 11326 7826 11350 7854
rect 11378 7826 11392 7854
rect 9902 7434 9916 7462
rect 9944 7434 9968 7462
rect 9996 7434 10020 7462
rect 10048 7434 10062 7462
rect 8572 6286 8732 7042
rect 8572 6258 8586 6286
rect 8614 6258 8638 6286
rect 8666 6258 8690 6286
rect 8718 6258 8732 6286
rect 8572 5502 8732 6258
rect 9758 7042 9786 7047
rect 9758 5978 9786 7014
rect 9814 6874 9842 6879
rect 9814 6146 9842 6846
rect 9814 6113 9842 6118
rect 9902 6678 10062 7434
rect 9902 6650 9916 6678
rect 9944 6650 9968 6678
rect 9996 6650 10020 6678
rect 10048 6650 10062 6678
rect 9758 5945 9786 5950
rect 8572 5474 8586 5502
rect 8614 5474 8638 5502
rect 8666 5474 8690 5502
rect 8718 5474 8732 5502
rect 8572 4718 8732 5474
rect 8572 4690 8586 4718
rect 8614 4690 8638 4718
rect 8666 4690 8690 4718
rect 8718 4690 8732 4718
rect 8572 3934 8732 4690
rect 8572 3906 8586 3934
rect 8614 3906 8638 3934
rect 8666 3906 8690 3934
rect 8718 3906 8732 3934
rect 8572 3150 8732 3906
rect 8572 3122 8586 3150
rect 8614 3122 8638 3150
rect 8666 3122 8690 3150
rect 8718 3122 8732 3150
rect 8572 2366 8732 3122
rect 8572 2338 8586 2366
rect 8614 2338 8638 2366
rect 8666 2338 8690 2366
rect 8718 2338 8732 2366
rect 8572 1582 8732 2338
rect 8572 1554 8586 1582
rect 8614 1554 8638 1582
rect 8666 1554 8690 1582
rect 8718 1554 8732 1582
rect 8572 1538 8732 1554
rect 9902 5894 10062 6650
rect 9902 5866 9916 5894
rect 9944 5866 9968 5894
rect 9996 5866 10020 5894
rect 10048 5866 10062 5894
rect 9902 5110 10062 5866
rect 9902 5082 9916 5110
rect 9944 5082 9968 5110
rect 9996 5082 10020 5110
rect 10048 5082 10062 5110
rect 9902 4326 10062 5082
rect 9902 4298 9916 4326
rect 9944 4298 9968 4326
rect 9996 4298 10020 4326
rect 10048 4298 10062 4326
rect 9902 3542 10062 4298
rect 9902 3514 9916 3542
rect 9944 3514 9968 3542
rect 9996 3514 10020 3542
rect 10048 3514 10062 3542
rect 9902 2758 10062 3514
rect 9902 2730 9916 2758
rect 9944 2730 9968 2758
rect 9996 2730 10020 2758
rect 10048 2730 10062 2758
rect 9902 1974 10062 2730
rect 9902 1946 9916 1974
rect 9944 1946 9968 1974
rect 9996 1946 10020 1974
rect 10048 1946 10062 1974
rect 9902 1538 10062 1946
rect 11232 7070 11392 7826
rect 11232 7042 11246 7070
rect 11274 7042 11298 7070
rect 11326 7042 11350 7070
rect 11378 7042 11392 7070
rect 11232 6286 11392 7042
rect 11232 6258 11246 6286
rect 11274 6258 11298 6286
rect 11326 6258 11350 6286
rect 11378 6258 11392 6286
rect 11232 5502 11392 6258
rect 11232 5474 11246 5502
rect 11274 5474 11298 5502
rect 11326 5474 11350 5502
rect 11378 5474 11392 5502
rect 11232 4718 11392 5474
rect 11232 4690 11246 4718
rect 11274 4690 11298 4718
rect 11326 4690 11350 4718
rect 11378 4690 11392 4718
rect 11232 3934 11392 4690
rect 11232 3906 11246 3934
rect 11274 3906 11298 3934
rect 11326 3906 11350 3934
rect 11378 3906 11392 3934
rect 11232 3150 11392 3906
rect 11232 3122 11246 3150
rect 11274 3122 11298 3150
rect 11326 3122 11350 3150
rect 11378 3122 11392 3150
rect 11232 2366 11392 3122
rect 11232 2338 11246 2366
rect 11274 2338 11298 2366
rect 11326 2338 11350 2366
rect 11378 2338 11392 2366
rect 11232 1582 11392 2338
rect 11232 1554 11246 1582
rect 11274 1554 11298 1582
rect 11326 1554 11350 1582
rect 11378 1554 11392 1582
rect 11232 1538 11392 1554
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _096_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 9912 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _097_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9520 0 -1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _098_
timestamp 1698431365
transform 1 0 2408 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _099_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2072 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _100_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2296 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _101_
timestamp 1698431365
transform -1 0 7392 0 -1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _102_
timestamp 1698431365
transform -1 0 4368 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _103_
timestamp 1698431365
transform -1 0 6272 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _104_
timestamp 1698431365
transform -1 0 6328 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _105_
timestamp 1698431365
transform 1 0 5264 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _106_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10472 0 1 3920
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _107_
timestamp 1698431365
transform -1 0 10472 0 -1 5488
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _108_
timestamp 1698431365
transform -1 0 9968 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _109_
timestamp 1698431365
transform -1 0 7728 0 -1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _110_
timestamp 1698431365
transform -1 0 7504 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _111_
timestamp 1698431365
transform -1 0 6496 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _112_
timestamp 1698431365
transform -1 0 5824 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _113_
timestamp 1698431365
transform -1 0 8120 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _114_
timestamp 1698431365
transform 1 0 3696 0 -1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _115_
timestamp 1698431365
transform -1 0 9520 0 1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _116_
timestamp 1698431365
transform -1 0 9576 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _117_
timestamp 1698431365
transform -1 0 7784 0 1 5488
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _118_
timestamp 1698431365
transform -1 0 4816 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _119_
timestamp 1698431365
transform -1 0 7112 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _120_
timestamp 1698431365
transform -1 0 6272 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _121_
timestamp 1698431365
transform -1 0 5152 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _122_
timestamp 1698431365
transform -1 0 4592 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _123_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 4368 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _124_
timestamp 1698431365
transform -1 0 7448 0 1 5488
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _125_
timestamp 1698431365
transform -1 0 4648 0 1 5488
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _126_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 4256 0 1 9408
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _127_
timestamp 1698431365
transform -1 0 2632 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _128_
timestamp 1698431365
transform 1 0 6440 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _129_
timestamp 1698431365
transform -1 0 9520 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _130_
timestamp 1698431365
transform -1 0 8064 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _131_
timestamp 1698431365
transform -1 0 5040 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _132_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3864 0 1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _133_
timestamp 1698431365
transform -1 0 3080 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _134_
timestamp 1698431365
transform -1 0 10248 0 -1 3920
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _135_
timestamp 1698431365
transform 1 0 9296 0 1 3920
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _136_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10136 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _137_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10080 0 -1 6272
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _138_
timestamp 1698431365
transform -1 0 10192 0 -1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _139_
timestamp 1698431365
transform 1 0 9912 0 1 5488
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _140_
timestamp 1698431365
transform 1 0 9968 0 1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _141_
timestamp 1698431365
transform 1 0 10080 0 -1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _142_
timestamp 1698431365
transform -1 0 4424 0 1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _143_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7728 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _144_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7280 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _145_
timestamp 1698431365
transform 1 0 1064 0 -1 5488
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _146_
timestamp 1698431365
transform -1 0 7728 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _147_
timestamp 1698431365
transform -1 0 7784 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _148_
timestamp 1698431365
transform -1 0 7448 0 1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _149_
timestamp 1698431365
transform 1 0 5880 0 -1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _150_
timestamp 1698431365
transform 1 0 7784 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _151_
timestamp 1698431365
transform -1 0 4144 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _152_
timestamp 1698431365
transform -1 0 2352 0 1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _153_
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _154_
timestamp 1698431365
transform 1 0 1680 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _155_
timestamp 1698431365
transform 1 0 1792 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _156_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4032 0 1 6272
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _157_
timestamp 1698431365
transform -1 0 10192 0 1 3920
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _158_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4704 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _159_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 2016 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _160_
timestamp 1698431365
transform 1 0 1680 0 1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _161_
timestamp 1698431365
transform -1 0 7504 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _162_
timestamp 1698431365
transform 1 0 2744 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _163_
timestamp 1698431365
transform 1 0 2632 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _164_
timestamp 1698431365
transform -1 0 3416 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _165_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 2240 0 -1 6272
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _166_
timestamp 1698431365
transform 1 0 1400 0 -1 5488
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _167_
timestamp 1698431365
transform 1 0 2128 0 -1 4704
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _168_
timestamp 1698431365
transform 1 0 3584 0 1 3920
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _169_
timestamp 1698431365
transform 1 0 7280 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _170_
timestamp 1698431365
transform 1 0 6720 0 1 7056
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _171_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7672 0 -1 5488
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _172_
timestamp 1698431365
transform -1 0 7112 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _173_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6384 0 -1 5488
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _174_
timestamp 1698431365
transform -1 0 5544 0 -1 4704
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _175_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4368 0 1 3920
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _176_
timestamp 1698431365
transform -1 0 5936 0 -1 7056
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _177_
timestamp 1698431365
transform 1 0 2240 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _178_
timestamp 1698431365
transform 1 0 4424 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _179_
timestamp 1698431365
transform 1 0 5600 0 1 7056
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _180_
timestamp 1698431365
transform -1 0 5320 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _181_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4872 0 1 4704
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _182_
timestamp 1698431365
transform 1 0 4816 0 -1 7056
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _183_
timestamp 1698431365
transform -1 0 5264 0 -1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _184_
timestamp 1698431365
transform 1 0 5544 0 1 3920
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _185_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4928 0 1 3920
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _186_
timestamp 1698431365
transform 1 0 6944 0 -1 3920
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _187_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7224 0 -1 3920
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _188_
timestamp 1698431365
transform 1 0 9576 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _189_
timestamp 1698431365
transform 1 0 9912 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _190_
timestamp 1698431365
transform -1 0 10080 0 -1 7056
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _191_
timestamp 1698431365
transform 1 0 9688 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _192_
timestamp 1698431365
transform 1 0 9800 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _193_
timestamp 1698431365
transform -1 0 10248 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _194_
timestamp 1698431365
transform 1 0 10136 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _195_
timestamp 1698431365
transform 1 0 10248 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _196_
timestamp 1698431365
transform 1 0 7728 0 -1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _197_
timestamp 1698431365
transform 1 0 8792 0 1 7840
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _198_
timestamp 1698431365
transform 1 0 9352 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _199_
timestamp 1698431365
transform -1 0 10136 0 -1 5488
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _200_
timestamp 1698431365
transform -1 0 9856 0 1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _201_
timestamp 1698431365
transform 1 0 9856 0 1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _202_
timestamp 1698431365
transform -1 0 1848 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _203_
timestamp 1698431365
transform 1 0 1848 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _204_
timestamp 1698431365
transform -1 0 1344 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _205_
timestamp 1698431365
transform 1 0 6944 0 -1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _206_
timestamp 1698431365
transform 1 0 7280 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _207_
timestamp 1698431365
transform 1 0 3976 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _208_
timestamp 1698431365
transform -1 0 3248 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _209_
timestamp 1698431365
transform 1 0 1792 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _210_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 2296 0 -1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _211_
timestamp 1698431365
transform 1 0 1400 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _212_
timestamp 1698431365
transform -1 0 3024 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _213_
timestamp 1698431365
transform -1 0 2576 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _214_
timestamp 1698431365
transform 1 0 9016 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _215_
timestamp 1698431365
transform 1 0 4872 0 -1 3920
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _216_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1792 0 1 3920
box -43 -43 883 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _217_
timestamp 1698431365
transform 1 0 1456 0 1 3920
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _218_
timestamp 1698431365
transform -1 0 2240 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _219_
timestamp 1698431365
transform -1 0 2128 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _220_
timestamp 1698431365
transform -1 0 2688 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _221_
timestamp 1698431365
transform -1 0 3360 0 1 3920
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _222_
timestamp 1698431365
transform -1 0 9072 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _223_
timestamp 1698431365
transform -1 0 9296 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _224_
timestamp 1698431365
transform 1 0 10416 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _225_
timestamp 1698431365
transform -1 0 10360 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _226_
timestamp 1698431365
transform -1 0 9968 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _227_
timestamp 1698431365
transform -1 0 10416 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _228_
timestamp 1698431365
transform -1 0 5880 0 -1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _229_
timestamp 1698431365
transform 1 0 5376 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _230_
timestamp 1698431365
transform 1 0 8008 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _231_
timestamp 1698431365
transform -1 0 8568 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__098__I $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3192 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__106__A1
timestamp 1698431365
transform -1 0 10808 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__143__A1
timestamp 1698431365
transform -1 0 7952 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__155__A1
timestamp 1698431365
transform 1 0 2352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__161__I
timestamp 1698431365
transform 1 0 7616 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__193__A1
timestamp 1698431365
transform 1 0 9688 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__B
timestamp 1698431365
transform 1 0 5544 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__B
timestamp 1698431365
transform -1 0 2912 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 11088 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 10864 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 10864 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 10864 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 10864 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 10864 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698431365
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698431365
transform 1 0 8400 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_172 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10304 0 1 1568
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698431365
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_142
timestamp 1698431365
transform 1 0 8624 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_174 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10416 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_182
timestamp 1698431365
transform 1 0 10864 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_186 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11088 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698431365
transform 1 0 6664 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698431365
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_177
timestamp 1698431365
transform 1 0 10584 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_179
timestamp 1698431365
transform 1 0 10696 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698431365
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_142
timestamp 1698431365
transform 1 0 8624 0 -1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_174
timestamp 1698431365
transform 1 0 10416 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_182
timestamp 1698431365
transform 1 0 10864 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_186
timestamp 1698431365
transform 1 0 11088 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_107
timestamp 1698431365
transform 1 0 6664 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_115
timestamp 1698431365
transform 1 0 7112 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_117
timestamp 1698431365
transform 1 0 7224 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_122
timestamp 1698431365
transform 1 0 7504 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_126
timestamp 1698431365
transform 1 0 7728 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_158
timestamp 1698431365
transform 1 0 9520 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_174
timestamp 1698431365
transform 1 0 10416 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_177
timestamp 1698431365
transform 1 0 10584 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_185
timestamp 1698431365
transform 1 0 11032 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_187
timestamp 1698431365
transform 1 0 11144 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_2
timestamp 1698431365
transform 1 0 784 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_18
timestamp 1698431365
transform 1 0 1680 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_26
timestamp 1698431365
transform 1 0 2128 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_36
timestamp 1698431365
transform 1 0 2688 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_40
timestamp 1698431365
transform 1 0 2912 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_56
timestamp 1698431365
transform 1 0 3808 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_64
timestamp 1698431365
transform 1 0 4256 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_68
timestamp 1698431365
transform 1 0 4480 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_72
timestamp 1698431365
transform 1 0 4704 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_74
timestamp 1698431365
transform 1 0 4816 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_85
timestamp 1698431365
transform 1 0 5432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_89
timestamp 1698431365
transform 1 0 5656 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_105
timestamp 1698431365
transform 1 0 6552 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_109
timestamp 1698431365
transform 1 0 6776 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_111
timestamp 1698431365
transform 1 0 6888 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_127
timestamp 1698431365
transform 1 0 7784 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_135
timestamp 1698431365
transform 1 0 8232 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_139
timestamp 1698431365
transform 1 0 8456 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_142
timestamp 1698431365
transform 1 0 8624 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_158
timestamp 1698431365
transform 1 0 9520 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_162
timestamp 1698431365
transform 1 0 9744 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_164
timestamp 1698431365
transform 1 0 9856 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_171
timestamp 1698431365
transform 1 0 10248 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_179
timestamp 1698431365
transform 1 0 10696 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_183
timestamp 1698431365
transform 1 0 10920 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_185
timestamp 1698431365
transform 1 0 11032 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_2
timestamp 1698431365
transform 1 0 784 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_10
timestamp 1698431365
transform 1 0 1232 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_48
timestamp 1698431365
transform 1 0 3360 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_57
timestamp 1698431365
transform 1 0 3864 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_65
timestamp 1698431365
transform 1 0 4312 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_93
timestamp 1698431365
transform 1 0 5880 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698431365
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_107
timestamp 1698431365
transform 1 0 6664 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_115
timestamp 1698431365
transform 1 0 7112 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_117
timestamp 1698431365
transform 1 0 7224 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_126
timestamp 1698431365
transform 1 0 7728 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_130
timestamp 1698431365
transform 1 0 7952 0 1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_146
timestamp 1698431365
transform 1 0 8848 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_160
timestamp 1698431365
transform 1 0 9632 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_177
timestamp 1698431365
transform 1 0 10584 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_181
timestamp 1698431365
transform 1 0 10808 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_2
timestamp 1698431365
transform 1 0 784 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_38
timestamp 1698431365
transform 1 0 2800 0 -1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_72
timestamp 1698431365
transform 1 0 4704 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_87
timestamp 1698431365
transform 1 0 5544 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_103
timestamp 1698431365
transform 1 0 6440 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_111
timestamp 1698431365
transform 1 0 6888 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_115
timestamp 1698431365
transform 1 0 7112 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_117
timestamp 1698431365
transform 1 0 7224 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_122
timestamp 1698431365
transform 1 0 7504 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_138
timestamp 1698431365
transform 1 0 8400 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_142
timestamp 1698431365
transform 1 0 8624 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_170
timestamp 1698431365
transform 1 0 10192 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_186
timestamp 1698431365
transform 1 0 11088 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_2
timestamp 1698431365
transform 1 0 784 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_18
timestamp 1698431365
transform 1 0 1680 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_28
timestamp 1698431365
transform 1 0 2240 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_32
timestamp 1698431365
transform 1 0 2464 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_37
timestamp 1698431365
transform 1 0 2744 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_53
timestamp 1698431365
transform 1 0 3640 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_87
timestamp 1698431365
transform 1 0 5544 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_103
timestamp 1698431365
transform 1 0 6440 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_107
timestamp 1698431365
transform 1 0 6664 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_115
timestamp 1698431365
transform 1 0 7112 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_117
timestamp 1698431365
transform 1 0 7224 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_126
timestamp 1698431365
transform 1 0 7728 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_142
timestamp 1698431365
transform 1 0 8624 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_150
timestamp 1698431365
transform 1 0 9072 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_170
timestamp 1698431365
transform 1 0 10192 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_174
timestamp 1698431365
transform 1 0 10416 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_177
timestamp 1698431365
transform 1 0 10584 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_185
timestamp 1698431365
transform 1 0 11032 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_187
timestamp 1698431365
transform 1 0 11144 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_2
timestamp 1698431365
transform 1 0 784 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_6
timestamp 1698431365
transform 1 0 1008 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_25
timestamp 1698431365
transform 1 0 2072 0 -1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_57
timestamp 1698431365
transform 1 0 3864 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_65
timestamp 1698431365
transform 1 0 4312 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_69
timestamp 1698431365
transform 1 0 4536 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_72
timestamp 1698431365
transform 1 0 4704 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_88
timestamp 1698431365
transform 1 0 5600 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_96
timestamp 1698431365
transform 1 0 6048 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_100
timestamp 1698431365
transform 1 0 6272 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_133
timestamp 1698431365
transform 1 0 8120 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_137
timestamp 1698431365
transform 1 0 8344 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_139
timestamp 1698431365
transform 1 0 8456 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_142
timestamp 1698431365
transform 1 0 8624 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_150
timestamp 1698431365
transform 1 0 9072 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_175
timestamp 1698431365
transform 1 0 10472 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_179
timestamp 1698431365
transform 1 0 10696 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_2
timestamp 1698431365
transform 1 0 784 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_18
timestamp 1698431365
transform 1 0 1680 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_26
timestamp 1698431365
transform 1 0 2128 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_32
timestamp 1698431365
transform 1 0 2464 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_37
timestamp 1698431365
transform 1 0 2744 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_53
timestamp 1698431365
transform 1 0 3640 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_61
timestamp 1698431365
transform 1 0 4088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_71
timestamp 1698431365
transform 1 0 4648 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_83
timestamp 1698431365
transform 1 0 5320 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_99
timestamp 1698431365
transform 1 0 6216 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_103
timestamp 1698431365
transform 1 0 6440 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_107
timestamp 1698431365
transform 1 0 6664 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_127
timestamp 1698431365
transform 1 0 7784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_159
timestamp 1698431365
transform 1 0 9576 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_163
timestamp 1698431365
transform 1 0 9800 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698431365
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_177
timestamp 1698431365
transform 1 0 10584 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_185
timestamp 1698431365
transform 1 0 11032 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_187
timestamp 1698431365
transform 1 0 11144 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_2
timestamp 1698431365
transform 1 0 784 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_10
timestamp 1698431365
transform 1 0 1232 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_14
timestamp 1698431365
transform 1 0 1456 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_28
timestamp 1698431365
transform 1 0 2240 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_32
timestamp 1698431365
transform 1 0 2464 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_34
timestamp 1698431365
transform 1 0 2576 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_39
timestamp 1698431365
transform 1 0 2856 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_49
timestamp 1698431365
transform 1 0 3416 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_53
timestamp 1698431365
transform 1 0 3640 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_60
timestamp 1698431365
transform 1 0 4032 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_68
timestamp 1698431365
transform 1 0 4480 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_80
timestamp 1698431365
transform 1 0 5152 0 -1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_112
timestamp 1698431365
transform 1 0 6944 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_128
timestamp 1698431365
transform 1 0 7840 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698431365
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_142
timestamp 1698431365
transform 1 0 8624 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_168
timestamp 1698431365
transform 1 0 10080 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_184
timestamp 1698431365
transform 1 0 10976 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_2
timestamp 1698431365
transform 1 0 784 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_24
timestamp 1698431365
transform 1 0 2016 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_32
timestamp 1698431365
transform 1 0 2464 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_41
timestamp 1698431365
transform 1 0 2968 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_57
timestamp 1698431365
transform 1 0 3864 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_59
timestamp 1698431365
transform 1 0 3976 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_69
timestamp 1698431365
transform 1 0 4536 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698431365
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_107
timestamp 1698431365
transform 1 0 6664 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_121
timestamp 1698431365
transform 1 0 7448 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_153
timestamp 1698431365
transform 1 0 9240 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_157
timestamp 1698431365
transform 1 0 9464 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_172
timestamp 1698431365
transform 1 0 10304 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698431365
transform 1 0 10416 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_177
timestamp 1698431365
transform 1 0 10584 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_185
timestamp 1698431365
transform 1 0 11032 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_187
timestamp 1698431365
transform 1 0 11144 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_2
timestamp 1698431365
transform 1 0 784 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_10
timestamp 1698431365
transform 1 0 1232 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_14
timestamp 1698431365
transform 1 0 1456 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_24
timestamp 1698431365
transform 1 0 2016 0 -1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_56
timestamp 1698431365
transform 1 0 3808 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_64
timestamp 1698431365
transform 1 0 4256 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_68
timestamp 1698431365
transform 1 0 4480 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_72
timestamp 1698431365
transform 1 0 4704 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_94
timestamp 1698431365
transform 1 0 5936 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_110
timestamp 1698431365
transform 1 0 6832 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_131
timestamp 1698431365
transform 1 0 8008 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_139
timestamp 1698431365
transform 1 0 8456 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_142
timestamp 1698431365
transform 1 0 8624 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_174
timestamp 1698431365
transform 1 0 10416 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_178
timestamp 1698431365
transform 1 0 10640 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_2
timestamp 1698431365
transform 1 0 784 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_24
timestamp 1698431365
transform 1 0 2016 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_30
timestamp 1698431365
transform 1 0 2352 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_37
timestamp 1698431365
transform 1 0 2744 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_53
timestamp 1698431365
transform 1 0 3640 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_70
timestamp 1698431365
transform 1 0 4592 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_78
timestamp 1698431365
transform 1 0 5040 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_104
timestamp 1698431365
transform 1 0 6496 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_107
timestamp 1698431365
transform 1 0 6664 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_132
timestamp 1698431365
transform 1 0 8064 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_148
timestamp 1698431365
transform 1 0 8960 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_156
timestamp 1698431365
transform 1 0 9408 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_158
timestamp 1698431365
transform 1 0 9520 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_171
timestamp 1698431365
transform 1 0 10248 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_177
timestamp 1698431365
transform 1 0 10584 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_185
timestamp 1698431365
transform 1 0 11032 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_187
timestamp 1698431365
transform 1 0 11144 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_2
timestamp 1698431365
transform 1 0 784 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_28
timestamp 1698431365
transform 1 0 2240 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_32
timestamp 1698431365
transform 1 0 2464 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_48
timestamp 1698431365
transform 1 0 3360 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_56
timestamp 1698431365
transform 1 0 3808 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698431365
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_80
timestamp 1698431365
transform 1 0 5152 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_88
timestamp 1698431365
transform 1 0 5600 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_92
timestamp 1698431365
transform 1 0 5824 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_94
timestamp 1698431365
transform 1 0 5936 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_101
timestamp 1698431365
transform 1 0 6328 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_109
timestamp 1698431365
transform 1 0 6776 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_113
timestamp 1698431365
transform 1 0 7000 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_115
timestamp 1698431365
transform 1 0 7112 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_122
timestamp 1698431365
transform 1 0 7504 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_138
timestamp 1698431365
transform 1 0 8400 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_142
timestamp 1698431365
transform 1 0 8624 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_158
timestamp 1698431365
transform 1 0 9520 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_160
timestamp 1698431365
transform 1 0 9632 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_177
timestamp 1698431365
transform 1 0 10584 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_185
timestamp 1698431365
transform 1 0 11032 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_187
timestamp 1698431365
transform 1 0 11144 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_2
timestamp 1698431365
transform 1 0 784 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_10
timestamp 1698431365
transform 1 0 1232 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_14
timestamp 1698431365
transform 1 0 1456 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_27
timestamp 1698431365
transform 1 0 2184 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_37
timestamp 1698431365
transform 1 0 2744 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_53
timestamp 1698431365
transform 1 0 3640 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_61
timestamp 1698431365
transform 1 0 4088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_65
timestamp 1698431365
transform 1 0 4312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_67
timestamp 1698431365
transform 1 0 4424 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_74
timestamp 1698431365
transform 1 0 4816 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_90
timestamp 1698431365
transform 1 0 5712 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_98
timestamp 1698431365
transform 1 0 6160 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_102
timestamp 1698431365
transform 1 0 6384 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_104
timestamp 1698431365
transform 1 0 6496 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_115
timestamp 1698431365
transform 1 0 7112 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_131
timestamp 1698431365
transform 1 0 8008 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_139
timestamp 1698431365
transform 1 0 8456 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_143
timestamp 1698431365
transform 1 0 8680 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_177
timestamp 1698431365
transform 1 0 10584 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_185
timestamp 1698431365
transform 1 0 11032 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_187
timestamp 1698431365
transform 1 0 11144 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_2
timestamp 1698431365
transform 1 0 784 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_18
timestamp 1698431365
transform 1 0 1680 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_26
timestamp 1698431365
transform 1 0 2128 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_30
timestamp 1698431365
transform 1 0 2352 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_43
timestamp 1698431365
transform 1 0 3080 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_47
timestamp 1698431365
transform 1 0 3304 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_55
timestamp 1698431365
transform 1 0 3752 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_59
timestamp 1698431365
transform 1 0 3976 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698431365
transform 1 0 4368 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698431365
transform 1 0 4704 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_88
timestamp 1698431365
transform 1 0 5600 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_92
timestamp 1698431365
transform 1 0 5824 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_100
timestamp 1698431365
transform 1 0 6272 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_132
timestamp 1698431365
transform 1 0 8064 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_142
timestamp 1698431365
transform 1 0 8624 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_158
timestamp 1698431365
transform 1 0 9520 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_162
timestamp 1698431365
transform 1 0 9744 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_169
timestamp 1698431365
transform 1 0 10136 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_177
timestamp 1698431365
transform 1 0 10584 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_179
timestamp 1698431365
transform 1 0 10696 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_2
timestamp 1698431365
transform 1 0 784 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_18
timestamp 1698431365
transform 1 0 1680 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_37
timestamp 1698431365
transform 1 0 2744 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_53
timestamp 1698431365
transform 1 0 3640 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_67
timestamp 1698431365
transform 1 0 4424 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_83
timestamp 1698431365
transform 1 0 5320 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_100
timestamp 1698431365
transform 1 0 6272 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_104
timestamp 1698431365
transform 1 0 6496 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_107
timestamp 1698431365
transform 1 0 6664 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_115
timestamp 1698431365
transform 1 0 7112 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_119
timestamp 1698431365
transform 1 0 7336 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_127
timestamp 1698431365
transform 1 0 7784 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_159
timestamp 1698431365
transform 1 0 9576 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_173
timestamp 1698431365
transform 1 0 10360 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_177
timestamp 1698431365
transform 1 0 10584 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_185
timestamp 1698431365
transform 1 0 11032 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_187
timestamp 1698431365
transform 1 0 11144 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_2
timestamp 1698431365
transform 1 0 784 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_10
timestamp 1698431365
transform 1 0 1232 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_12
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_46
timestamp 1698431365
transform 1 0 3248 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_54
timestamp 1698431365
transform 1 0 3696 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_58
timestamp 1698431365
transform 1 0 3920 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_67
timestamp 1698431365
transform 1 0 4424 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_69
timestamp 1698431365
transform 1 0 4536 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_78
timestamp 1698431365
transform 1 0 5040 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_82
timestamp 1698431365
transform 1 0 5264 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_109
timestamp 1698431365
transform 1 0 6776 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_111
timestamp 1698431365
transform 1 0 6888 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_122
timestamp 1698431365
transform 1 0 7504 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_126
timestamp 1698431365
transform 1 0 7728 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_133
timestamp 1698431365
transform 1 0 8120 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_137
timestamp 1698431365
transform 1 0 8344 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698431365
transform 1 0 8456 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_142
timestamp 1698431365
transform 1 0 8624 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_146
timestamp 1698431365
transform 1 0 8848 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_148
timestamp 1698431365
transform 1 0 8960 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_155
timestamp 1698431365
transform 1 0 9352 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_159
timestamp 1698431365
transform 1 0 9576 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_182
timestamp 1698431365
transform 1 0 10864 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_186
timestamp 1698431365
transform 1 0 11088 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_2
timestamp 1698431365
transform 1 0 784 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_18
timestamp 1698431365
transform 1 0 1680 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_22
timestamp 1698431365
transform 1 0 1904 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_24
timestamp 1698431365
transform 1 0 2016 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_37
timestamp 1698431365
transform 1 0 2744 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_53
timestamp 1698431365
transform 1 0 3640 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_64
timestamp 1698431365
transform 1 0 4256 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_80
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_90
timestamp 1698431365
transform 1 0 5712 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_98
timestamp 1698431365
transform 1 0 6160 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_102
timestamp 1698431365
transform 1 0 6384 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_104
timestamp 1698431365
transform 1 0 6496 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_107
timestamp 1698431365
transform 1 0 6664 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_115
timestamp 1698431365
transform 1 0 7112 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_117
timestamp 1698431365
transform 1 0 7224 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_124
timestamp 1698431365
transform 1 0 7616 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_128
timestamp 1698431365
transform 1 0 7840 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_130
timestamp 1698431365
transform 1 0 7952 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_141
timestamp 1698431365
transform 1 0 8568 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_154
timestamp 1698431365
transform 1 0 9296 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_162
timestamp 1698431365
transform 1 0 9744 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_169
timestamp 1698431365
transform 1 0 10136 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_173
timestamp 1698431365
transform 1 0 10360 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_177
timestamp 1698431365
transform 1 0 10584 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_179
timestamp 1698431365
transform 1 0 10696 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_2
timestamp 1698431365
transform 1 0 784 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_4
timestamp 1698431365
transform 1 0 896 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_11
timestamp 1698431365
transform 1 0 1288 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_19
timestamp 1698431365
transform 1 0 1736 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_23
timestamp 1698431365
transform 1 0 1960 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_31
timestamp 1698431365
transform 1 0 2408 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_33
timestamp 1698431365
transform 1 0 2520 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_36
timestamp 1698431365
transform 1 0 2688 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_44
timestamp 1698431365
transform 1 0 3136 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_51
timestamp 1698431365
transform 1 0 3528 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_67
timestamp 1698431365
transform 1 0 4424 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_76
timestamp 1698431365
transform 1 0 4928 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_84
timestamp 1698431365
transform 1 0 5376 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_91
timestamp 1698431365
transform 1 0 5768 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_99
timestamp 1698431365
transform 1 0 6216 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_101
timestamp 1698431365
transform 1 0 6328 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_104
timestamp 1698431365
transform 1 0 6496 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_111
timestamp 1698431365
transform 1 0 6888 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_119
timestamp 1698431365
transform 1 0 7336 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_123
timestamp 1698431365
transform 1 0 7560 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_131
timestamp 1698431365
transform 1 0 8008 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_135
timestamp 1698431365
transform 1 0 8232 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_138
timestamp 1698431365
transform 1 0 8400 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698431365
transform 1 0 8624 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_144
timestamp 1698431365
transform 1 0 8736 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_151
timestamp 1698431365
transform 1 0 9128 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_159
timestamp 1698431365
transform 1 0 9576 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_163
timestamp 1698431365
transform 1 0 9800 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_178
timestamp 1698431365
transform 1 0 10640 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform -1 0 11200 0 1 3920
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform -1 0 11200 0 -1 5488
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform -1 0 11200 0 -1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform -1 0 11200 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform -1 0 11200 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform -1 0 11200 0 1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output7
timestamp 1698431365
transform 1 0 9856 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output8
timestamp 1698431365
transform -1 0 1288 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output9
timestamp 1698431365
transform -1 0 2408 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output10
timestamp 1698431365
transform -1 0 3528 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output11
timestamp 1698431365
transform -1 0 4928 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output12
timestamp 1698431365
transform -1 0 5768 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output13
timestamp 1698431365
transform -1 0 6888 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output14
timestamp 1698431365
transform -1 0 8008 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output15
timestamp 1698431365
transform -1 0 9128 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output16
timestamp 1698431365
transform -1 0 10640 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output17
timestamp 1698431365
transform 1 0 10864 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_22 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 11312 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_23
timestamp 1698431365
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 11312 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_24
timestamp 1698431365
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 11312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_25
timestamp 1698431365
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 11312 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_26
timestamp 1698431365
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 11312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_27
timestamp 1698431365
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 11312 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_28
timestamp 1698431365
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 11312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_29
timestamp 1698431365
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 11312 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_30
timestamp 1698431365
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 11312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_31
timestamp 1698431365
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 11312 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_32
timestamp 1698431365
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 11312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_33
timestamp 1698431365
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 11312 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_34
timestamp 1698431365
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 11312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_35
timestamp 1698431365
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 11312 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_36
timestamp 1698431365
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 11312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_37
timestamp 1698431365
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 11312 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_38
timestamp 1698431365
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 11312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_39
timestamp 1698431365
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 11312 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_40
timestamp 1698431365
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 11312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_41
timestamp 1698431365
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 11312 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_42
timestamp 1698431365
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 11312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_43
timestamp 1698431365
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 11312 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_44 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_45
timestamp 1698431365
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_46
timestamp 1698431365
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_47
timestamp 1698431365
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_48
timestamp 1698431365
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_49
timestamp 1698431365
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_50
timestamp 1698431365
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_51
timestamp 1698431365
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_52
timestamp 1698431365
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_53
timestamp 1698431365
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_54
timestamp 1698431365
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_55
timestamp 1698431365
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_56
timestamp 1698431365
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_57
timestamp 1698431365
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_58
timestamp 1698431365
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_59
timestamp 1698431365
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_60
timestamp 1698431365
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_61
timestamp 1698431365
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_62
timestamp 1698431365
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_63
timestamp 1698431365
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_64
timestamp 1698431365
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_65
timestamp 1698431365
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_66
timestamp 1698431365
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_67
timestamp 1698431365
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_68
timestamp 1698431365
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_69
timestamp 1698431365
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_70
timestamp 1698431365
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_71
timestamp 1698431365
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_72
timestamp 1698431365
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_73
timestamp 1698431365
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_74
timestamp 1698431365
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_75
timestamp 1698431365
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_76
timestamp 1698431365
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_77
timestamp 1698431365
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_78
timestamp 1698431365
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_79
timestamp 1698431365
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_80
timestamp 1698431365
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_81
timestamp 1698431365
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_82
timestamp 1698431365
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_83
timestamp 1698431365
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_84
timestamp 1698431365
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_85
timestamp 1698431365
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_86
timestamp 1698431365
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_87
timestamp 1698431365
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_88
timestamp 1698431365
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_89
timestamp 1698431365
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_90
timestamp 1698431365
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_91
timestamp 1698431365
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_92
timestamp 1698431365
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_93
timestamp 1698431365
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_94
timestamp 1698431365
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_95
timestamp 1698431365
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_96
timestamp 1698431365
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_97
timestamp 1698431365
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_98
timestamp 1698431365
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_99
timestamp 1698431365
transform 1 0 2576 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_100
timestamp 1698431365
transform 1 0 4480 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_101
timestamp 1698431365
transform 1 0 6384 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_102
timestamp 1698431365
transform 1 0 8288 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_103
timestamp 1698431365
transform 1 0 10192 0 -1 10192
box -43 -43 155 435
<< labels >>
flabel metal3 s 11600 784 12000 840 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 11600 3696 12000 3752 0 FreeSans 224 0 0 0 io_in[0]
port 1 nsew signal input
flabel metal3 s 11600 5152 12000 5208 0 FreeSans 224 0 0 0 io_in[1]
port 2 nsew signal input
flabel metal3 s 11600 6608 12000 6664 0 FreeSans 224 0 0 0 io_in[2]
port 3 nsew signal input
flabel metal3 s 11600 8064 12000 8120 0 FreeSans 224 0 0 0 io_in[3]
port 4 nsew signal input
flabel metal3 s 11600 9520 12000 9576 0 FreeSans 224 0 0 0 io_in[4]
port 5 nsew signal input
flabel metal3 s 11600 10976 12000 11032 0 FreeSans 224 0 0 0 io_oeb
port 6 nsew signal tristate
flabel metal2 s 896 11600 952 12000 0 FreeSans 224 90 0 0 io_out[0]
port 7 nsew signal tristate
flabel metal2 s 2016 11600 2072 12000 0 FreeSans 224 90 0 0 io_out[1]
port 8 nsew signal tristate
flabel metal2 s 3136 11600 3192 12000 0 FreeSans 224 90 0 0 io_out[2]
port 9 nsew signal tristate
flabel metal2 s 4256 11600 4312 12000 0 FreeSans 224 90 0 0 io_out[3]
port 10 nsew signal tristate
flabel metal2 s 5376 11600 5432 12000 0 FreeSans 224 90 0 0 io_out[4]
port 11 nsew signal tristate
flabel metal2 s 6496 11600 6552 12000 0 FreeSans 224 90 0 0 io_out[5]
port 12 nsew signal tristate
flabel metal2 s 7616 11600 7672 12000 0 FreeSans 224 90 0 0 io_out[6]
port 13 nsew signal tristate
flabel metal2 s 8736 11600 8792 12000 0 FreeSans 224 90 0 0 io_out[7]
port 14 nsew signal tristate
flabel metal2 s 9856 11600 9912 12000 0 FreeSans 224 90 0 0 io_out[8]
port 15 nsew signal tristate
flabel metal2 s 10976 11600 11032 12000 0 FreeSans 224 90 0 0 io_out[9]
port 16 nsew signal tristate
flabel metal3 s 11600 2240 12000 2296 0 FreeSans 224 0 0 0 rst_n
port 17 nsew signal input
flabel metal4 s 1922 1538 2082 10222 0 FreeSans 640 90 0 0 vdd
port 18 nsew power bidirectional
flabel metal4 s 4582 1538 4742 10222 0 FreeSans 640 90 0 0 vdd
port 18 nsew power bidirectional
flabel metal4 s 7242 1538 7402 10222 0 FreeSans 640 90 0 0 vdd
port 18 nsew power bidirectional
flabel metal4 s 9902 1538 10062 10222 0 FreeSans 640 90 0 0 vdd
port 18 nsew power bidirectional
flabel metal4 s 3252 1538 3412 10222 0 FreeSans 640 90 0 0 vss
port 19 nsew ground bidirectional
flabel metal4 s 5912 1538 6072 10222 0 FreeSans 640 90 0 0 vss
port 19 nsew ground bidirectional
flabel metal4 s 8572 1538 8732 10222 0 FreeSans 640 90 0 0 vss
port 19 nsew ground bidirectional
flabel metal4 s 11232 1538 11392 10222 0 FreeSans 640 90 0 0 vss
port 19 nsew ground bidirectional
rlabel metal1 5992 9800 5992 9800 0 vdd
rlabel via1 6032 10192 6032 10192 0 vss
rlabel metal3 4004 8792 4004 8792 0 _000_
rlabel metal3 8428 5180 8428 5180 0 _001_
rlabel metal2 9212 5488 9212 5488 0 _002_
rlabel metal2 4172 8372 4172 8372 0 _003_
rlabel metal3 5460 7588 5460 7588 0 _004_
rlabel metal2 4312 7588 4312 7588 0 _005_
rlabel metal2 4228 6832 4228 6832 0 _006_
rlabel metal2 3976 7756 3976 7756 0 _007_
rlabel metal2 7196 5796 7196 5796 0 _008_
rlabel metal2 2212 6664 2212 6664 0 _009_
rlabel metal2 5684 9072 5684 9072 0 _010_
rlabel metal2 9156 7056 9156 7056 0 _011_
rlabel metal2 7420 9100 7420 9100 0 _012_
rlabel metal3 3500 8708 3500 8708 0 _013_
rlabel metal2 9380 3892 9380 3892 0 _014_
rlabel metal3 8624 4116 8624 4116 0 _015_
rlabel metal3 9688 9492 9688 9492 0 _016_
rlabel metal2 10220 8764 10220 8764 0 _017_
rlabel metal2 10444 7630 10444 7630 0 _018_
rlabel metal2 10164 6636 10164 6636 0 _019_
rlabel metal2 7448 4620 7448 4620 0 _020_
rlabel metal2 1316 5180 1316 5180 0 _021_
rlabel metal2 6132 9212 6132 9212 0 _022_
rlabel metal3 7112 9268 7112 9268 0 _023_
rlabel metal3 3024 7196 3024 7196 0 _024_
rlabel metal2 1484 7476 1484 7476 0 _025_
rlabel metal2 1680 7700 1680 7700 0 _026_
rlabel metal2 1876 7476 1876 7476 0 _027_
rlabel metal2 4788 6216 4788 6216 0 _028_
rlabel metal2 9940 4088 9940 4088 0 _029_
rlabel metal2 1792 7980 1792 7980 0 _030_
rlabel metal2 1652 6636 1652 6636 0 _031_
rlabel metal2 7420 3808 7420 3808 0 _032_
rlabel metal2 3276 6188 3276 6188 0 _033_
rlabel metal2 2884 6076 2884 6076 0 _034_
rlabel metal2 3724 4116 3724 4116 0 _035_
rlabel metal2 1596 5320 1596 5320 0 _036_
rlabel metal2 2184 4508 2184 4508 0 _037_
rlabel metal3 3192 4116 3192 4116 0 _038_
rlabel metal3 4424 4116 4424 4116 0 _039_
rlabel metal2 7812 6636 7812 6636 0 _040_
rlabel metal2 7140 5796 7140 5796 0 _041_
rlabel metal2 7028 5012 7028 5012 0 _042_
rlabel metal3 6076 4844 6076 4844 0 _043_
rlabel metal2 5488 4564 5488 4564 0 _044_
rlabel metal2 4676 4200 4676 4200 0 _045_
rlabel metal2 5068 4004 5068 4004 0 _046_
rlabel metal2 5460 5824 5460 5824 0 _047_
rlabel metal3 3640 5684 3640 5684 0 _048_
rlabel metal2 5292 4816 5292 4816 0 _049_
rlabel metal2 9044 8568 9044 8568 0 _050_
rlabel metal2 5012 5124 5012 5124 0 _051_
rlabel metal2 5236 4228 5236 4228 0 _052_
rlabel metal2 4956 4032 4956 4032 0 _053_
rlabel metal3 5376 4060 5376 4060 0 _054_
rlabel metal2 5404 4144 5404 4144 0 _055_
rlabel metal3 6412 3724 6412 3724 0 _056_
rlabel metal2 7196 3864 7196 3864 0 _057_
rlabel metal2 9912 7308 9912 7308 0 _058_
rlabel metal2 9828 8120 9828 8120 0 _059_
rlabel metal2 10108 7980 10108 7980 0 _060_
rlabel metal2 10304 7700 10304 7700 0 _061_
rlabel metal3 8456 7980 8456 7980 0 _062_
rlabel metal2 9268 7952 9268 7952 0 _063_
rlabel metal3 9828 4956 9828 4956 0 _064_
rlabel metal2 1260 7812 1260 7812 0 _065_
rlabel metal2 7420 9436 7420 9436 0 _066_
rlabel metal2 2100 9240 2100 9240 0 _067_
rlabel metal3 2604 8764 2604 8764 0 _068_
rlabel metal2 1904 8876 1904 8876 0 _069_
rlabel metal3 1680 9212 1680 9212 0 _070_
rlabel metal2 2520 8932 2520 8932 0 _071_
rlabel metal2 2996 4060 2996 4060 0 _072_
rlabel metal3 1764 4116 1764 4116 0 _073_
rlabel metal2 1820 4648 1820 4648 0 _074_
rlabel metal3 2520 4172 2520 4172 0 _075_
rlabel metal2 2548 3864 2548 3864 0 _076_
rlabel metal2 9072 9604 9072 9604 0 _077_
rlabel metal2 10332 9268 10332 9268 0 _078_
rlabel metal2 10164 8988 10164 8988 0 _079_
rlabel metal2 5516 9464 5516 9464 0 _080_
rlabel metal2 8232 9604 8232 9604 0 _081_
rlabel metal2 9660 4368 9660 4368 0 _082_
rlabel metal2 2352 7588 2352 7588 0 _083_
rlabel metal2 2660 8708 2660 8708 0 _084_
rlabel metal2 2380 9436 2380 9436 0 _085_
rlabel metal2 3948 7392 3948 7392 0 _086_
rlabel metal2 4088 8820 4088 8820 0 _087_
rlabel metal2 5404 7280 5404 7280 0 _088_
rlabel metal2 5796 9128 5796 9128 0 _089_
rlabel metal2 10332 5432 10332 5432 0 _090_
rlabel metal2 10220 5432 10220 5432 0 _091_
rlabel metal3 8624 6580 8624 6580 0 _092_
rlabel metal2 7224 7700 7224 7700 0 _093_
rlabel metal2 5628 8624 5628 8624 0 _094_
rlabel metal2 7980 6132 7980 6132 0 _095_
rlabel metal3 10717 812 10717 812 0 clk
rlabel metal3 11361 3724 11361 3724 0 io_in[0]
rlabel metal2 11116 5236 11116 5236 0 io_in[1]
rlabel metal2 11116 6748 11116 6748 0 io_in[2]
rlabel metal2 11116 8260 11116 8260 0 io_in[3]
rlabel metal3 11361 9548 11361 9548 0 io_in[4]
rlabel metal2 10080 10052 10080 10052 0 io_oeb
rlabel metal2 924 10843 924 10843 0 io_out[0]
rlabel metal2 2044 10843 2044 10843 0 io_out[1]
rlabel metal2 3164 10843 3164 10843 0 io_out[2]
rlabel metal2 4564 11620 4564 11620 0 io_out[3]
rlabel metal2 5404 10843 5404 10843 0 io_out[4]
rlabel metal2 6524 10843 6524 10843 0 io_out[5]
rlabel metal2 7700 10052 7700 10052 0 io_out[6]
rlabel metal2 8820 10052 8820 10052 0 io_out[7]
rlabel metal3 10136 10052 10136 10052 0 io_out[8]
rlabel metal2 11060 10052 11060 10052 0 io_out[9]
rlabel metal2 8092 9520 8092 9520 0 main.GATES_100.input2
rlabel metal2 7224 7252 7224 7252 0 main.GATES_102.input1
rlabel metal2 6188 8708 6188 8708 0 main.GATES_102.input2
rlabel metal2 7420 7812 7420 7812 0 main.GATES_102.input3
rlabel metal2 2016 7644 2016 7644 0 main.GATES_103.input2
rlabel metal3 1820 7980 1820 7980 0 main.GATES_105.input3
rlabel metal3 2072 9156 2072 9156 0 main.GATES_106.input2
rlabel metal3 7686 7308 7686 7308 0 main.GATES_107.input2
rlabel metal2 7588 4340 7588 4340 0 main.GATES_108.input1
rlabel metal2 2296 8932 2296 8932 0 main.GATES_109.input2
rlabel metal2 7392 5572 7392 5572 0 main.GATES_11.input2
rlabel metal2 1988 6104 1988 6104 0 main.GATES_110.input1
rlabel metal2 7504 3668 7504 3668 0 main.GATES_113.input1
rlabel metal2 2828 8022 2828 8022 0 main.GATES_114.input2
rlabel metal2 6244 8820 6244 8820 0 main.GATES_115.input2
rlabel metal2 6972 7756 6972 7756 0 main.GATES_116.input1
rlabel metal2 4956 9072 4956 9072 0 main.GATES_116.input3
rlabel metal2 7868 5936 7868 5936 0 main.GATES_119.result
rlabel metal3 8680 4900 8680 4900 0 main.GATES_124.input2
rlabel metal2 7028 7868 7028 7868 0 main.GATES_127.result
rlabel metal2 2436 3892 2436 3892 0 main.GATES_132.input1
rlabel metal3 9912 6468 9912 6468 0 main.GATES_15.input3
rlabel metal2 8988 9436 8988 9436 0 main.GATES_16.input1
rlabel metal2 10332 8036 10332 8036 0 main.GATES_18.result
rlabel metal3 8876 9156 8876 9156 0 main.GATES_19.input1
rlabel metal2 9716 9016 9716 9016 0 main.GATES_20.result
rlabel metal2 9772 5040 9772 5040 0 main.GATES_26.input3
rlabel metal2 9660 7084 9660 7084 0 main.GATES_29.input3
rlabel metal3 10052 8036 10052 8036 0 main.GATES_46.input3
rlabel metal3 10528 4060 10528 4060 0 net1
rlabel metal3 2968 4508 2968 4508 0 net10
rlabel metal2 2156 7728 2156 7728 0 net11
rlabel metal2 5628 9772 5628 9772 0 net12
rlabel metal2 6804 9856 6804 9856 0 net13
rlabel metal2 7532 9772 7532 9772 0 net14
rlabel metal2 3948 9520 3948 9520 0 net15
rlabel metal2 9212 9324 9212 9324 0 net16
rlabel metal3 10612 9240 10612 9240 0 net17
rlabel metal2 10948 5628 10948 5628 0 net2
rlabel metal3 10472 6916 10472 6916 0 net3
rlabel metal2 10920 8484 10920 8484 0 net4
rlabel metal2 10976 8596 10976 8596 0 net5
rlabel metal3 10556 3724 10556 3724 0 net6
rlabel metal3 3220 9548 3220 9548 0 net7
rlabel metal2 1120 5404 1120 5404 0 net8
rlabel metal2 2492 9856 2492 9856 0 net9
rlabel metal2 11116 2408 11116 2408 0 rst_n
<< properties >>
string FIXED_BBOX 0 0 12000 12000
<< end >>
