magic
tech gf180mcuD
magscale 1 5
timestamp 1753965785
<< nwell >>
rect 629 15857 17347 16115
rect 629 15073 17347 15503
rect 629 14289 17347 14719
rect 629 13505 17347 13935
rect 629 12721 17347 13151
rect 629 11937 17347 12367
rect 629 11153 17347 11583
rect 629 10369 17347 10799
rect 629 9585 17347 10015
rect 629 8801 17347 9231
rect 629 8017 17347 8447
rect 629 7233 17347 7663
rect 629 6449 17347 6879
rect 629 5665 17347 6095
rect 629 4881 17347 5311
rect 629 4097 17347 4527
rect 629 3313 17347 3743
rect 629 2529 17347 2959
rect 629 1745 17347 2175
<< pwell >>
rect 629 15503 17347 15857
rect 629 14719 17347 15073
rect 629 13935 17347 14289
rect 629 13151 17347 13505
rect 629 12367 17347 12721
rect 629 11583 17347 11937
rect 629 10799 17347 11153
rect 629 10015 17347 10369
rect 629 9231 17347 9585
rect 629 8447 17347 8801
rect 629 7663 17347 8017
rect 629 6879 17347 7233
rect 629 6095 17347 6449
rect 629 5311 17347 5665
rect 629 4527 17347 4881
rect 629 3743 17347 4097
rect 629 2959 17347 3313
rect 629 2175 17347 2529
rect 629 1525 17347 1745
<< obsm1 >>
rect 672 1538 17384 16102
<< metal2 >>
rect 1792 0 1848 400
rect 5376 0 5432 400
rect 8960 0 9016 400
rect 12544 0 12600 400
rect 16128 0 16184 400
<< obsm2 >>
rect 798 430 17370 16091
rect 798 400 1762 430
rect 1878 400 5346 430
rect 5462 400 8930 430
rect 9046 400 12514 430
rect 12630 400 16098 430
rect 16214 400 17370 430
<< obsm3 >>
rect 793 1554 17375 16086
<< metal4 >>
rect 2671 1538 2831 16102
rect 4750 1538 4910 16102
rect 6829 1538 6989 16102
rect 8908 1538 9068 16102
rect 10987 1538 11147 16102
rect 13066 1538 13226 16102
rect 15145 1538 15305 16102
rect 17224 1538 17384 16102
<< obsm4 >>
rect 1694 2865 2641 12647
rect 2861 2865 4720 12647
rect 4940 2865 6799 12647
rect 7019 2865 8878 12647
rect 9098 2865 10957 12647
rect 11177 2865 11802 12647
<< labels >>
rlabel metal2 s 8960 0 9016 400 6 io_out[0]
port 1 nsew signal output
rlabel metal2 s 12544 0 12600 400 6 io_out[1]
port 2 nsew signal output
rlabel metal2 s 16128 0 16184 400 6 io_out[2]
port 3 nsew signal output
rlabel metal2 s 5376 0 5432 400 6 rst_n
port 4 nsew signal input
rlabel metal4 s 2671 1538 2831 16102 6 vdd
port 5 nsew power bidirectional
rlabel metal4 s 6829 1538 6989 16102 6 vdd
port 5 nsew power bidirectional
rlabel metal4 s 10987 1538 11147 16102 6 vdd
port 5 nsew power bidirectional
rlabel metal4 s 15145 1538 15305 16102 6 vdd
port 5 nsew power bidirectional
rlabel metal4 s 4750 1538 4910 16102 6 vss
port 6 nsew ground bidirectional
rlabel metal4 s 8908 1538 9068 16102 6 vss
port 6 nsew ground bidirectional
rlabel metal4 s 13066 1538 13226 16102 6 vss
port 6 nsew ground bidirectional
rlabel metal4 s 17224 1538 17384 16102 6 vss
port 6 nsew ground bidirectional
rlabel metal2 s 1792 0 1848 400 6 wb_clk_i
port 7 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 18000 18000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1068034
string GDS_FILE /home/lucah/gfmpw1-multi/openlane/blinker/runs/25_07_31_14_42/results/signoff/blinker.magic.gds
string GDS_START 173308
<< end >>

