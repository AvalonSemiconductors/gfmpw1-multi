VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO blinker
  CLASS BLOCK ;
  FOREIGN blinker ;
  ORIGIN 0.000 0.000 ;
  SIZE 180.000 BY 180.000 ;
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 89.600 0.000 90.160 4.000 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 125.440 0.000 126.000 4.000 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 0.000 161.840 4.000 ;
    END
  END io_out[2]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 0.000 54.320 4.000 ;
    END
  END rst_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 26.710 15.380 28.310 161.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 68.290 15.380 69.890 161.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 109.870 15.380 111.470 161.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 151.450 15.380 153.050 161.020 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 47.500 15.380 49.100 161.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 89.080 15.380 90.680 161.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 130.660 15.380 132.260 161.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 172.240 15.380 173.840 161.020 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.352000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 17.920 0.000 18.480 4.000 ;
    END
  END wb_clk_i
  OBS
      LAYER Nwell ;
        RECT 6.290 158.570 173.470 161.150 ;
      LAYER Pwell ;
        RECT 6.290 155.030 173.470 158.570 ;
      LAYER Nwell ;
        RECT 6.290 150.730 173.470 155.030 ;
      LAYER Pwell ;
        RECT 6.290 147.190 173.470 150.730 ;
      LAYER Nwell ;
        RECT 6.290 142.890 173.470 147.190 ;
      LAYER Pwell ;
        RECT 6.290 139.350 173.470 142.890 ;
      LAYER Nwell ;
        RECT 6.290 135.050 173.470 139.350 ;
      LAYER Pwell ;
        RECT 6.290 131.510 173.470 135.050 ;
      LAYER Nwell ;
        RECT 6.290 127.210 173.470 131.510 ;
      LAYER Pwell ;
        RECT 6.290 123.670 173.470 127.210 ;
      LAYER Nwell ;
        RECT 6.290 119.370 173.470 123.670 ;
      LAYER Pwell ;
        RECT 6.290 115.830 173.470 119.370 ;
      LAYER Nwell ;
        RECT 6.290 111.530 173.470 115.830 ;
      LAYER Pwell ;
        RECT 6.290 107.990 173.470 111.530 ;
      LAYER Nwell ;
        RECT 6.290 103.690 173.470 107.990 ;
      LAYER Pwell ;
        RECT 6.290 100.150 173.470 103.690 ;
      LAYER Nwell ;
        RECT 6.290 95.850 173.470 100.150 ;
      LAYER Pwell ;
        RECT 6.290 92.310 173.470 95.850 ;
      LAYER Nwell ;
        RECT 6.290 88.010 173.470 92.310 ;
      LAYER Pwell ;
        RECT 6.290 84.470 173.470 88.010 ;
      LAYER Nwell ;
        RECT 6.290 80.170 173.470 84.470 ;
      LAYER Pwell ;
        RECT 6.290 76.630 173.470 80.170 ;
      LAYER Nwell ;
        RECT 6.290 72.330 173.470 76.630 ;
      LAYER Pwell ;
        RECT 6.290 68.790 173.470 72.330 ;
      LAYER Nwell ;
        RECT 6.290 64.490 173.470 68.790 ;
      LAYER Pwell ;
        RECT 6.290 60.950 173.470 64.490 ;
      LAYER Nwell ;
        RECT 6.290 56.650 173.470 60.950 ;
      LAYER Pwell ;
        RECT 6.290 53.110 173.470 56.650 ;
      LAYER Nwell ;
        RECT 6.290 48.810 173.470 53.110 ;
      LAYER Pwell ;
        RECT 6.290 45.270 173.470 48.810 ;
      LAYER Nwell ;
        RECT 6.290 40.970 173.470 45.270 ;
      LAYER Pwell ;
        RECT 6.290 37.430 173.470 40.970 ;
      LAYER Nwell ;
        RECT 6.290 33.130 173.470 37.430 ;
      LAYER Pwell ;
        RECT 6.290 29.590 173.470 33.130 ;
      LAYER Nwell ;
        RECT 6.290 25.290 173.470 29.590 ;
      LAYER Pwell ;
        RECT 6.290 21.750 173.470 25.290 ;
      LAYER Nwell ;
        RECT 6.290 17.450 173.470 21.750 ;
      LAYER Pwell ;
        RECT 6.290 15.250 173.470 17.450 ;
      LAYER Metal1 ;
        RECT 6.720 15.380 173.840 161.020 ;
      LAYER Metal2 ;
        RECT 7.980 4.300 173.700 160.910 ;
        RECT 7.980 4.000 17.620 4.300 ;
        RECT 18.780 4.000 53.460 4.300 ;
        RECT 54.620 4.000 89.300 4.300 ;
        RECT 90.460 4.000 125.140 4.300 ;
        RECT 126.300 4.000 160.980 4.300 ;
        RECT 162.140 4.000 173.700 4.300 ;
      LAYER Metal3 ;
        RECT 7.930 15.540 173.750 160.860 ;
      LAYER Metal4 ;
        RECT 16.940 28.650 26.410 126.470 ;
        RECT 28.610 28.650 47.200 126.470 ;
        RECT 49.400 28.650 67.990 126.470 ;
        RECT 70.190 28.650 88.780 126.470 ;
        RECT 90.980 28.650 109.570 126.470 ;
        RECT 111.770 28.650 118.020 126.470 ;
  END
END blinker
END LIBRARY

