magic
tech gf180mcuD
magscale 1 10
timestamp 1702247292
<< metal1 >>
rect 30930 46398 30942 46450
rect 30994 46447 31006 46450
rect 32610 46447 32622 46450
rect 30994 46401 32622 46447
rect 30994 46398 31006 46401
rect 32610 46398 32622 46401
rect 32674 46447 32686 46450
rect 33170 46447 33182 46450
rect 32674 46401 33182 46447
rect 32674 46398 32686 46401
rect 33170 46398 33182 46401
rect 33234 46398 33246 46450
rect 40338 46398 40350 46450
rect 40402 46447 40414 46450
rect 41794 46447 41806 46450
rect 40402 46401 41806 46447
rect 40402 46398 40414 46401
rect 41794 46398 41806 46401
rect 41858 46398 41870 46450
rect 1344 46282 48608 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 48608 46282
rect 1344 46196 48608 46230
rect 18510 46002 18562 46014
rect 43150 46002 43202 46014
rect 21522 45950 21534 46002
rect 21586 45950 21598 46002
rect 23650 45950 23662 46002
rect 23714 45950 23726 46002
rect 24546 45950 24558 46002
rect 24610 45950 24622 46002
rect 18510 45938 18562 45950
rect 43150 45938 43202 45950
rect 44942 46002 44994 46014
rect 44942 45938 44994 45950
rect 11342 45890 11394 45902
rect 32174 45890 32226 45902
rect 18722 45838 18734 45890
rect 18786 45838 18798 45890
rect 19618 45838 19630 45890
rect 19682 45838 19694 45890
rect 20850 45838 20862 45890
rect 20914 45838 20926 45890
rect 27458 45838 27470 45890
rect 27522 45838 27534 45890
rect 28354 45838 28366 45890
rect 28418 45838 28430 45890
rect 32610 45838 32622 45890
rect 32674 45838 32686 45890
rect 38210 45838 38222 45890
rect 38274 45838 38286 45890
rect 43810 45838 43822 45890
rect 43874 45838 43886 45890
rect 45266 45838 45278 45890
rect 45330 45838 45342 45890
rect 11342 45826 11394 45838
rect 32174 45826 32226 45838
rect 10670 45778 10722 45790
rect 10670 45714 10722 45726
rect 10894 45778 10946 45790
rect 33070 45778 33122 45790
rect 19058 45726 19070 45778
rect 19122 45726 19134 45778
rect 26674 45726 26686 45778
rect 26738 45726 26750 45778
rect 29138 45726 29150 45778
rect 29202 45726 29214 45778
rect 10894 45714 10946 45726
rect 33070 45714 33122 45726
rect 33742 45778 33794 45790
rect 33742 45714 33794 45726
rect 34414 45778 34466 45790
rect 34414 45714 34466 45726
rect 37886 45778 37938 45790
rect 37886 45714 37938 45726
rect 41582 45778 41634 45790
rect 41582 45714 41634 45726
rect 41694 45778 41746 45790
rect 41694 45714 41746 45726
rect 41806 45778 41858 45790
rect 41806 45714 41858 45726
rect 45502 45778 45554 45790
rect 45502 45714 45554 45726
rect 45838 45778 45890 45790
rect 45838 45714 45890 45726
rect 47406 45778 47458 45790
rect 47406 45714 47458 45726
rect 11118 45666 11170 45678
rect 33406 45666 33458 45678
rect 19842 45614 19854 45666
rect 19906 45614 19918 45666
rect 20066 45614 20078 45666
rect 20130 45614 20142 45666
rect 31378 45614 31390 45666
rect 31442 45614 31454 45666
rect 11118 45602 11170 45614
rect 33406 45602 33458 45614
rect 33854 45666 33906 45678
rect 33854 45602 33906 45614
rect 33966 45666 34018 45678
rect 33966 45602 34018 45614
rect 34526 45666 34578 45678
rect 34526 45602 34578 45614
rect 34638 45666 34690 45678
rect 34638 45602 34690 45614
rect 37998 45666 38050 45678
rect 45950 45666 46002 45678
rect 46846 45666 46898 45678
rect 42242 45614 42254 45666
rect 42306 45614 42318 45666
rect 43586 45614 43598 45666
rect 43650 45614 43662 45666
rect 46498 45614 46510 45666
rect 46562 45614 46574 45666
rect 37998 45602 38050 45614
rect 45950 45602 46002 45614
rect 46846 45602 46898 45614
rect 47518 45666 47570 45678
rect 47518 45602 47570 45614
rect 47630 45666 47682 45678
rect 47630 45602 47682 45614
rect 48190 45666 48242 45678
rect 48190 45602 48242 45614
rect 1344 45498 48608 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 48608 45498
rect 1344 45412 48608 45446
rect 18846 45330 18898 45342
rect 17490 45278 17502 45330
rect 17554 45278 17566 45330
rect 18846 45266 18898 45278
rect 24670 45330 24722 45342
rect 31938 45278 31950 45330
rect 32002 45278 32014 45330
rect 24670 45266 24722 45278
rect 20514 45166 20526 45218
rect 20578 45166 20590 45218
rect 21970 45166 21982 45218
rect 22034 45166 22046 45218
rect 39106 45166 39118 45218
rect 39170 45166 39182 45218
rect 17838 45106 17890 45118
rect 18398 45106 18450 45118
rect 22430 45106 22482 45118
rect 25454 45106 25506 45118
rect 13458 45054 13470 45106
rect 13522 45054 13534 45106
rect 13794 45054 13806 45106
rect 13858 45054 13870 45106
rect 18162 45054 18174 45106
rect 18226 45054 18238 45106
rect 19730 45054 19742 45106
rect 19794 45054 19806 45106
rect 21410 45054 21422 45106
rect 21474 45054 21486 45106
rect 23202 45054 23214 45106
rect 23266 45054 23278 45106
rect 25218 45054 25230 45106
rect 25282 45054 25294 45106
rect 17838 45042 17890 45054
rect 18398 45042 18450 45054
rect 22430 45042 22482 45054
rect 25454 45042 25506 45054
rect 25678 45106 25730 45118
rect 25678 45042 25730 45054
rect 25790 45106 25842 45118
rect 25790 45042 25842 45054
rect 26350 45106 26402 45118
rect 31390 45106 31442 45118
rect 32286 45106 32338 45118
rect 41022 45106 41074 45118
rect 48190 45106 48242 45118
rect 27682 45054 27694 45106
rect 27746 45054 27758 45106
rect 31602 45054 31614 45106
rect 31666 45054 31678 45106
rect 36306 45054 36318 45106
rect 36370 45054 36382 45106
rect 39890 45054 39902 45106
rect 39954 45054 39966 45106
rect 42914 45054 42926 45106
rect 42978 45054 42990 45106
rect 26350 45042 26402 45054
rect 31390 45042 31442 45054
rect 32286 45042 32338 45054
rect 41022 45042 41074 45054
rect 48190 45042 48242 45054
rect 19406 44994 19458 45006
rect 10546 44942 10558 44994
rect 10610 44942 10622 44994
rect 12674 44942 12686 44994
rect 12738 44942 12750 44994
rect 14578 44942 14590 44994
rect 14642 44942 14654 44994
rect 16706 44942 16718 44994
rect 16770 44942 16782 44994
rect 19406 44930 19458 44942
rect 24558 44994 24610 45006
rect 24558 44930 24610 44942
rect 25566 44994 25618 45006
rect 31054 44994 31106 45006
rect 28466 44942 28478 44994
rect 28530 44942 28542 44994
rect 30594 44942 30606 44994
rect 30658 44942 30670 44994
rect 25566 44930 25618 44942
rect 31054 44930 31106 44942
rect 32510 44994 32562 45006
rect 41694 44994 41746 45006
rect 47630 44994 47682 45006
rect 33394 44942 33406 44994
rect 33458 44942 33470 44994
rect 35522 44942 35534 44994
rect 35586 44942 35598 44994
rect 36978 44942 36990 44994
rect 37042 44942 37054 44994
rect 44818 44942 44830 44994
rect 44882 44942 44894 44994
rect 32510 44930 32562 44942
rect 41694 44930 41746 44942
rect 47630 44930 47682 44942
rect 18510 44882 18562 44894
rect 18510 44818 18562 44830
rect 31166 44882 31218 44894
rect 31166 44818 31218 44830
rect 40910 44882 40962 44894
rect 40910 44818 40962 44830
rect 1344 44714 48608 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 48608 44714
rect 1344 44628 48608 44662
rect 16158 44546 16210 44558
rect 16158 44482 16210 44494
rect 20750 44546 20802 44558
rect 20750 44482 20802 44494
rect 32286 44546 32338 44558
rect 32286 44482 32338 44494
rect 32622 44546 32674 44558
rect 32622 44482 32674 44494
rect 33854 44546 33906 44558
rect 33854 44482 33906 44494
rect 34190 44546 34242 44558
rect 34190 44482 34242 44494
rect 12014 44434 12066 44446
rect 15150 44434 15202 44446
rect 30942 44434 30994 44446
rect 7634 44382 7646 44434
rect 7698 44382 7710 44434
rect 12674 44382 12686 44434
rect 12738 44382 12750 44434
rect 17378 44382 17390 44434
rect 17442 44382 17454 44434
rect 12014 44370 12066 44382
rect 15150 44370 15202 44382
rect 30942 44370 30994 44382
rect 33182 44434 33234 44446
rect 33182 44370 33234 44382
rect 34078 44434 34130 44446
rect 34078 44370 34130 44382
rect 37998 44434 38050 44446
rect 43810 44382 43822 44434
rect 43874 44382 43886 44434
rect 47730 44382 47742 44434
rect 47794 44382 47806 44434
rect 37998 44370 38050 44382
rect 11566 44322 11618 44334
rect 14366 44322 14418 44334
rect 15822 44322 15874 44334
rect 10434 44270 10446 44322
rect 10498 44270 10510 44322
rect 14130 44270 14142 44322
rect 14194 44270 14206 44322
rect 15586 44270 15598 44322
rect 15650 44270 15662 44322
rect 11566 44258 11618 44270
rect 14366 44258 14418 44270
rect 15822 44258 15874 44270
rect 16046 44322 16098 44334
rect 16718 44322 16770 44334
rect 16482 44270 16494 44322
rect 16546 44270 16558 44322
rect 16046 44258 16098 44270
rect 16718 44258 16770 44270
rect 16942 44322 16994 44334
rect 31950 44322 32002 44334
rect 20290 44270 20302 44322
rect 20354 44270 20366 44322
rect 26562 44270 26574 44322
rect 26626 44270 26638 44322
rect 31490 44270 31502 44322
rect 31554 44270 31566 44322
rect 16942 44258 16994 44270
rect 31950 44258 32002 44270
rect 32510 44322 32562 44334
rect 37102 44322 37154 44334
rect 40126 44322 40178 44334
rect 33618 44270 33630 44322
rect 33682 44270 33694 44322
rect 37426 44270 37438 44322
rect 37490 44270 37502 44322
rect 38546 44270 38558 44322
rect 38610 44270 38622 44322
rect 39778 44270 39790 44322
rect 39842 44270 39854 44322
rect 41010 44270 41022 44322
rect 41074 44270 41086 44322
rect 44818 44270 44830 44322
rect 44882 44270 44894 44322
rect 32510 44258 32562 44270
rect 37102 44258 37154 44270
rect 40126 44258 40178 44270
rect 11342 44210 11394 44222
rect 9762 44158 9774 44210
rect 9826 44158 9838 44210
rect 11342 44146 11394 44158
rect 11454 44210 11506 44222
rect 11454 44146 11506 44158
rect 12910 44210 12962 44222
rect 12910 44146 12962 44158
rect 13470 44210 13522 44222
rect 13470 44146 13522 44158
rect 15038 44210 15090 44222
rect 15038 44146 15090 44158
rect 15262 44210 15314 44222
rect 15262 44146 15314 44158
rect 17054 44210 17106 44222
rect 20638 44210 20690 44222
rect 30270 44210 30322 44222
rect 31278 44210 31330 44222
rect 19506 44158 19518 44210
rect 19570 44158 19582 44210
rect 24546 44158 24558 44210
rect 24610 44158 24622 44210
rect 31042 44158 31054 44210
rect 31106 44158 31118 44210
rect 17054 44146 17106 44158
rect 20638 44146 20690 44158
rect 30270 44146 30322 44158
rect 31278 44146 31330 44158
rect 39342 44210 39394 44222
rect 39342 44146 39394 44158
rect 40574 44210 40626 44222
rect 41682 44158 41694 44210
rect 41746 44158 41758 44210
rect 45602 44158 45614 44210
rect 45666 44158 45678 44210
rect 40574 44146 40626 44158
rect 12126 44098 12178 44110
rect 10882 44046 10894 44098
rect 10946 44046 10958 44098
rect 12126 44034 12178 44046
rect 12686 44098 12738 44110
rect 12686 44034 12738 44046
rect 27134 44098 27186 44110
rect 27134 44034 27186 44046
rect 30606 44098 30658 44110
rect 30606 44034 30658 44046
rect 32622 44098 32674 44110
rect 36206 44098 36258 44110
rect 40462 44098 40514 44110
rect 35858 44046 35870 44098
rect 35922 44046 35934 44098
rect 38322 44046 38334 44098
rect 38386 44046 38398 44098
rect 32622 44034 32674 44046
rect 36206 44034 36258 44046
rect 40462 44034 40514 44046
rect 48190 44098 48242 44110
rect 48190 44034 48242 44046
rect 1344 43930 48608 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 48608 43930
rect 1344 43844 48608 43878
rect 17278 43762 17330 43774
rect 16034 43710 16046 43762
rect 16098 43710 16110 43762
rect 17278 43698 17330 43710
rect 25790 43762 25842 43774
rect 25790 43698 25842 43710
rect 33182 43762 33234 43774
rect 33182 43698 33234 43710
rect 33742 43762 33794 43774
rect 33742 43698 33794 43710
rect 35422 43762 35474 43774
rect 38222 43762 38274 43774
rect 36978 43710 36990 43762
rect 37042 43710 37054 43762
rect 41122 43710 41134 43762
rect 41186 43710 41198 43762
rect 35422 43698 35474 43710
rect 38222 43698 38274 43710
rect 13582 43650 13634 43662
rect 13582 43586 13634 43598
rect 16606 43650 16658 43662
rect 18062 43650 18114 43662
rect 17826 43598 17838 43650
rect 17890 43598 17902 43650
rect 16606 43586 16658 43598
rect 18062 43586 18114 43598
rect 23886 43650 23938 43662
rect 23886 43586 23938 43598
rect 24334 43650 24386 43662
rect 24334 43586 24386 43598
rect 25230 43650 25282 43662
rect 25230 43586 25282 43598
rect 35646 43650 35698 43662
rect 35646 43586 35698 43598
rect 39006 43650 39058 43662
rect 39006 43586 39058 43598
rect 40350 43650 40402 43662
rect 44830 43650 44882 43662
rect 41010 43598 41022 43650
rect 41074 43598 41086 43650
rect 42466 43598 42478 43650
rect 42530 43598 42542 43650
rect 40350 43586 40402 43598
rect 44830 43586 44882 43598
rect 11902 43538 11954 43550
rect 16494 43538 16546 43550
rect 5954 43486 5966 43538
rect 6018 43486 6030 43538
rect 11330 43486 11342 43538
rect 11394 43486 11406 43538
rect 12562 43486 12574 43538
rect 12626 43486 12638 43538
rect 11902 43474 11954 43486
rect 16494 43474 16546 43486
rect 16718 43538 16770 43550
rect 18174 43538 18226 43550
rect 24110 43538 24162 43550
rect 17714 43486 17726 43538
rect 17778 43486 17790 43538
rect 20402 43486 20414 43538
rect 20466 43486 20478 43538
rect 21634 43486 21646 43538
rect 21698 43486 21710 43538
rect 21970 43486 21982 43538
rect 22034 43486 22046 43538
rect 22642 43486 22654 43538
rect 22706 43486 22718 43538
rect 16718 43474 16770 43486
rect 18174 43474 18226 43486
rect 24110 43474 24162 43486
rect 24446 43538 24498 43550
rect 24446 43474 24498 43486
rect 25454 43538 25506 43550
rect 25454 43474 25506 43486
rect 25678 43538 25730 43550
rect 25678 43474 25730 43486
rect 26350 43538 26402 43550
rect 34526 43538 34578 43550
rect 31938 43486 31950 43538
rect 32002 43486 32014 43538
rect 33394 43486 33406 43538
rect 33458 43486 33470 43538
rect 33954 43486 33966 43538
rect 34018 43486 34030 43538
rect 26350 43474 26402 43486
rect 34526 43474 34578 43486
rect 34750 43538 34802 43550
rect 36430 43538 36482 43550
rect 34962 43486 34974 43538
rect 35026 43486 35038 43538
rect 34750 43474 34802 43486
rect 36430 43474 36482 43486
rect 36654 43538 36706 43550
rect 36654 43474 36706 43486
rect 38110 43538 38162 43550
rect 38110 43474 38162 43486
rect 38446 43538 38498 43550
rect 38446 43474 38498 43486
rect 38558 43538 38610 43550
rect 38558 43474 38610 43486
rect 39230 43538 39282 43550
rect 39230 43474 39282 43486
rect 39678 43538 39730 43550
rect 39678 43474 39730 43486
rect 39790 43538 39842 43550
rect 40898 43486 40910 43538
rect 40962 43486 40974 43538
rect 42018 43486 42030 43538
rect 42082 43486 42094 43538
rect 43810 43486 43822 43538
rect 43874 43486 43886 43538
rect 48066 43486 48078 43538
rect 48130 43486 48142 43538
rect 39790 43474 39842 43486
rect 9550 43426 9602 43438
rect 6626 43374 6638 43426
rect 6690 43374 6702 43426
rect 8866 43374 8878 43426
rect 8930 43374 8942 43426
rect 9550 43362 9602 43374
rect 10446 43426 10498 43438
rect 10446 43362 10498 43374
rect 11566 43426 11618 43438
rect 11566 43362 11618 43374
rect 12238 43426 12290 43438
rect 12238 43362 12290 43374
rect 12350 43426 12402 43438
rect 18734 43426 18786 43438
rect 24222 43426 24274 43438
rect 13906 43374 13918 43426
rect 13970 43374 13982 43426
rect 20066 43374 20078 43426
rect 20130 43374 20142 43426
rect 23202 43374 23214 43426
rect 23266 43374 23278 43426
rect 12350 43362 12402 43374
rect 18734 43362 18786 43374
rect 24222 43362 24274 43374
rect 25566 43426 25618 43438
rect 38782 43426 38834 43438
rect 44270 43426 44322 43438
rect 27234 43374 27246 43426
rect 27298 43374 27310 43426
rect 35298 43374 35310 43426
rect 35362 43374 35374 43426
rect 43362 43374 43374 43426
rect 43426 43374 43438 43426
rect 25566 43362 25618 43374
rect 38782 43362 38834 43374
rect 44270 43362 44322 43374
rect 44606 43426 44658 43438
rect 44930 43374 44942 43426
rect 44994 43374 45006 43426
rect 45266 43374 45278 43426
rect 45330 43374 45342 43426
rect 47394 43374 47406 43426
rect 47458 43374 47470 43426
rect 44606 43362 44658 43374
rect 9774 43314 9826 43326
rect 10558 43314 10610 43326
rect 10098 43262 10110 43314
rect 10162 43262 10174 43314
rect 9774 43250 9826 43262
rect 10558 43250 10610 43262
rect 10782 43314 10834 43326
rect 10782 43250 10834 43262
rect 10894 43314 10946 43326
rect 10894 43250 10946 43262
rect 11790 43314 11842 43326
rect 11790 43250 11842 43262
rect 33070 43314 33122 43326
rect 33070 43250 33122 43262
rect 34414 43314 34466 43326
rect 34414 43250 34466 43262
rect 40014 43314 40066 43326
rect 40014 43250 40066 43262
rect 40238 43314 40290 43326
rect 40238 43250 40290 43262
rect 1344 43146 48608 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 48608 43146
rect 1344 43060 48608 43094
rect 24558 42978 24610 42990
rect 31390 42978 31442 42990
rect 39790 42978 39842 42990
rect 22642 42926 22654 42978
rect 22706 42926 22718 42978
rect 29698 42926 29710 42978
rect 29762 42926 29774 42978
rect 31714 42926 31726 42978
rect 31778 42926 31790 42978
rect 24558 42914 24610 42926
rect 31390 42914 31442 42926
rect 39790 42914 39842 42926
rect 47406 42978 47458 42990
rect 47406 42914 47458 42926
rect 47518 42978 47570 42990
rect 47518 42914 47570 42926
rect 16830 42866 16882 42878
rect 25118 42866 25170 42878
rect 30158 42866 30210 42878
rect 9986 42814 9998 42866
rect 10050 42814 10062 42866
rect 16370 42814 16382 42866
rect 16434 42814 16446 42866
rect 19394 42814 19406 42866
rect 19458 42814 19470 42866
rect 20402 42814 20414 42866
rect 20466 42814 20478 42866
rect 21298 42814 21310 42866
rect 21362 42814 21374 42866
rect 28578 42814 28590 42866
rect 28642 42814 28654 42866
rect 16830 42802 16882 42814
rect 25118 42802 25170 42814
rect 30158 42802 30210 42814
rect 31166 42866 31218 42878
rect 31166 42802 31218 42814
rect 33070 42866 33122 42878
rect 34290 42814 34302 42866
rect 34354 42814 34366 42866
rect 36418 42814 36430 42866
rect 36482 42814 36494 42866
rect 44258 42814 44270 42866
rect 44322 42814 44334 42866
rect 33070 42802 33122 42814
rect 16942 42754 16994 42766
rect 12898 42702 12910 42754
rect 12962 42702 12974 42754
rect 13570 42702 13582 42754
rect 13634 42702 13646 42754
rect 16942 42690 16994 42702
rect 17278 42754 17330 42766
rect 22318 42754 22370 42766
rect 23998 42754 24050 42766
rect 19170 42702 19182 42754
rect 19234 42702 19246 42754
rect 20178 42702 20190 42754
rect 20242 42702 20254 42754
rect 22754 42702 22766 42754
rect 22818 42702 22830 42754
rect 23538 42702 23550 42754
rect 23602 42702 23614 42754
rect 17278 42690 17330 42702
rect 22318 42690 22370 42702
rect 23998 42690 24050 42702
rect 24670 42754 24722 42766
rect 29150 42754 29202 42766
rect 25778 42702 25790 42754
rect 25842 42702 25854 42754
rect 24670 42690 24722 42702
rect 29150 42690 29202 42702
rect 29374 42754 29426 42766
rect 29374 42690 29426 42702
rect 30382 42754 30434 42766
rect 39566 42754 39618 42766
rect 40574 42754 40626 42766
rect 30594 42702 30606 42754
rect 30658 42702 30670 42754
rect 33618 42702 33630 42754
rect 33682 42702 33694 42754
rect 39330 42702 39342 42754
rect 39394 42702 39406 42754
rect 40226 42702 40238 42754
rect 40290 42702 40302 42754
rect 30382 42690 30434 42702
rect 39566 42690 39618 42702
rect 40574 42690 40626 42702
rect 40686 42754 40738 42766
rect 45614 42754 45666 42766
rect 41458 42702 41470 42754
rect 41522 42702 41534 42754
rect 40686 42690 40738 42702
rect 45614 42690 45666 42702
rect 45726 42754 45778 42766
rect 45726 42690 45778 42702
rect 46398 42754 46450 42766
rect 46398 42690 46450 42702
rect 46846 42754 46898 42766
rect 46846 42690 46898 42702
rect 47742 42754 47794 42766
rect 47742 42690 47794 42702
rect 47854 42754 47906 42766
rect 47854 42690 47906 42702
rect 16718 42642 16770 42654
rect 21646 42642 21698 42654
rect 14242 42590 14254 42642
rect 14306 42590 14318 42642
rect 17602 42590 17614 42642
rect 17666 42590 17678 42642
rect 19618 42590 19630 42642
rect 19682 42590 19694 42642
rect 16718 42578 16770 42590
rect 21646 42578 21698 42590
rect 24558 42642 24610 42654
rect 30046 42642 30098 42654
rect 39902 42642 39954 42654
rect 26450 42590 26462 42642
rect 26514 42590 26526 42642
rect 37874 42590 37886 42642
rect 37938 42590 37950 42642
rect 24558 42578 24610 42590
rect 30046 42578 30098 42590
rect 39902 42578 39954 42590
rect 41022 42642 41074 42654
rect 44942 42642 44994 42654
rect 42130 42590 42142 42642
rect 42194 42590 42206 42642
rect 41022 42578 41074 42590
rect 44942 42578 44994 42590
rect 45502 42642 45554 42654
rect 45502 42578 45554 42590
rect 47070 42642 47122 42654
rect 47070 42578 47122 42590
rect 17950 42530 18002 42542
rect 17950 42466 18002 42478
rect 25006 42530 25058 42542
rect 25006 42466 25058 42478
rect 32398 42530 32450 42542
rect 32398 42466 32450 42478
rect 33182 42530 33234 42542
rect 33182 42466 33234 42478
rect 37550 42530 37602 42542
rect 44830 42530 44882 42542
rect 46734 42530 46786 42542
rect 40786 42478 40798 42530
rect 40850 42478 40862 42530
rect 46162 42478 46174 42530
rect 46226 42478 46238 42530
rect 37550 42466 37602 42478
rect 44830 42466 44882 42478
rect 46734 42466 46786 42478
rect 1344 42362 48608 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 48608 42362
rect 1344 42276 48608 42310
rect 14030 42194 14082 42206
rect 14030 42130 14082 42142
rect 40238 42194 40290 42206
rect 40238 42130 40290 42142
rect 41582 42194 41634 42206
rect 41582 42130 41634 42142
rect 10782 42082 10834 42094
rect 10782 42018 10834 42030
rect 11902 42082 11954 42094
rect 11902 42018 11954 42030
rect 12574 42082 12626 42094
rect 12574 42018 12626 42030
rect 16830 42082 16882 42094
rect 16830 42018 16882 42030
rect 18622 42082 18674 42094
rect 18622 42018 18674 42030
rect 18734 42082 18786 42094
rect 18734 42018 18786 42030
rect 30830 42082 30882 42094
rect 41358 42082 41410 42094
rect 36978 42030 36990 42082
rect 37042 42030 37054 42082
rect 30830 42018 30882 42030
rect 41358 42018 41410 42030
rect 42030 42082 42082 42094
rect 47954 42030 47966 42082
rect 48018 42030 48030 42082
rect 42030 42018 42082 42030
rect 10110 41970 10162 41982
rect 6066 41918 6078 41970
rect 6130 41918 6142 41970
rect 6850 41918 6862 41970
rect 6914 41918 6926 41970
rect 10110 41906 10162 41918
rect 11678 41970 11730 41982
rect 11678 41906 11730 41918
rect 12462 41970 12514 41982
rect 14142 41970 14194 41982
rect 13794 41918 13806 41970
rect 13858 41918 13870 41970
rect 12462 41906 12514 41918
rect 14142 41906 14194 41918
rect 15374 41970 15426 41982
rect 16718 41970 16770 41982
rect 16034 41918 16046 41970
rect 16098 41918 16110 41970
rect 15374 41906 15426 41918
rect 16718 41906 16770 41918
rect 18958 41970 19010 41982
rect 24558 41970 24610 41982
rect 19170 41918 19182 41970
rect 19234 41918 19246 41970
rect 19618 41918 19630 41970
rect 19682 41918 19694 41970
rect 21074 41918 21086 41970
rect 21138 41918 21150 41970
rect 22194 41918 22206 41970
rect 22258 41918 22270 41970
rect 18958 41906 19010 41918
rect 24558 41906 24610 41918
rect 24670 41970 24722 41982
rect 24670 41906 24722 41918
rect 26126 41970 26178 41982
rect 26126 41906 26178 41918
rect 26462 41970 26514 41982
rect 30494 41970 30546 41982
rect 27234 41918 27246 41970
rect 27298 41918 27310 41970
rect 26462 41906 26514 41918
rect 30494 41906 30546 41918
rect 36654 41970 36706 41982
rect 36654 41906 36706 41918
rect 37886 41970 37938 41982
rect 41022 41970 41074 41982
rect 38434 41918 38446 41970
rect 38498 41918 38510 41970
rect 37886 41906 37938 41918
rect 41022 41906 41074 41918
rect 42142 41970 42194 41982
rect 42578 41918 42590 41970
rect 42642 41918 42654 41970
rect 43026 41918 43038 41970
rect 43090 41918 43102 41970
rect 42142 41906 42194 41918
rect 9886 41858 9938 41870
rect 11230 41858 11282 41870
rect 8978 41806 8990 41858
rect 9042 41806 9054 41858
rect 10434 41806 10446 41858
rect 10498 41806 10510 41858
rect 9886 41794 9938 41806
rect 11230 41794 11282 41806
rect 11790 41858 11842 41870
rect 11790 41794 11842 41806
rect 13134 41858 13186 41870
rect 17838 41858 17890 41870
rect 16258 41806 16270 41858
rect 16322 41806 16334 41858
rect 13134 41794 13186 41806
rect 17838 41794 17890 41806
rect 18398 41858 18450 41870
rect 24110 41858 24162 41870
rect 20738 41806 20750 41858
rect 20802 41806 20814 41858
rect 22642 41806 22654 41858
rect 22706 41806 22718 41858
rect 18398 41794 18450 41806
rect 24110 41794 24162 41806
rect 25454 41858 25506 41870
rect 31278 41858 31330 41870
rect 28018 41806 28030 41858
rect 28082 41806 28094 41858
rect 30146 41806 30158 41858
rect 30210 41806 30222 41858
rect 25454 41794 25506 41806
rect 31278 41794 31330 41806
rect 33070 41858 33122 41870
rect 33070 41794 33122 41806
rect 39902 41858 39954 41870
rect 39902 41794 39954 41806
rect 40350 41858 40402 41870
rect 40350 41794 40402 41806
rect 10894 41746 10946 41758
rect 10894 41682 10946 41694
rect 11118 41746 11170 41758
rect 11118 41682 11170 41694
rect 12574 41746 12626 41758
rect 12574 41682 12626 41694
rect 23998 41746 24050 41758
rect 23998 41682 24050 41694
rect 26350 41746 26402 41758
rect 26350 41682 26402 41694
rect 26686 41746 26738 41758
rect 26686 41682 26738 41694
rect 26798 41746 26850 41758
rect 26798 41682 26850 41694
rect 33182 41746 33234 41758
rect 33182 41682 33234 41694
rect 37326 41746 37378 41758
rect 37326 41682 37378 41694
rect 37662 41746 37714 41758
rect 37662 41682 37714 41694
rect 38446 41746 38498 41758
rect 38446 41682 38498 41694
rect 38782 41746 38834 41758
rect 38782 41682 38834 41694
rect 40910 41746 40962 41758
rect 40910 41682 40962 41694
rect 41694 41746 41746 41758
rect 41694 41682 41746 41694
rect 42366 41746 42418 41758
rect 42366 41682 42418 41694
rect 1344 41578 48608 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 48608 41578
rect 1344 41492 48608 41526
rect 19854 41410 19906 41422
rect 19854 41346 19906 41358
rect 30718 41410 30770 41422
rect 30718 41346 30770 41358
rect 34302 41410 34354 41422
rect 34302 41346 34354 41358
rect 40686 41410 40738 41422
rect 40686 41346 40738 41358
rect 29486 41298 29538 41310
rect 6066 41246 6078 41298
rect 6130 41246 6142 41298
rect 12002 41246 12014 41298
rect 12066 41246 12078 41298
rect 14466 41246 14478 41298
rect 14530 41246 14542 41298
rect 21746 41246 21758 41298
rect 21810 41246 21822 41298
rect 23874 41246 23886 41298
rect 23938 41246 23950 41298
rect 26450 41246 26462 41298
rect 26514 41246 26526 41298
rect 28578 41246 28590 41298
rect 28642 41246 28654 41298
rect 38098 41246 38110 41298
rect 38162 41246 38174 41298
rect 40226 41246 40238 41298
rect 40290 41246 40302 41298
rect 41346 41246 41358 41298
rect 41410 41246 41422 41298
rect 43474 41246 43486 41298
rect 43538 41246 43550 41298
rect 45266 41246 45278 41298
rect 45330 41246 45342 41298
rect 47394 41246 47406 41298
rect 47458 41246 47470 41298
rect 29486 41234 29538 41246
rect 13582 41186 13634 41198
rect 21422 41186 21474 41198
rect 30942 41186 30994 41198
rect 10882 41134 10894 41186
rect 10946 41134 10958 41186
rect 12338 41134 12350 41186
rect 12402 41134 12414 41186
rect 19506 41134 19518 41186
rect 19570 41134 19582 41186
rect 24546 41134 24558 41186
rect 24610 41134 24622 41186
rect 25778 41134 25790 41186
rect 25842 41134 25854 41186
rect 29698 41134 29710 41186
rect 29762 41134 29774 41186
rect 13582 41122 13634 41134
rect 21422 41122 21474 41134
rect 30942 41122 30994 41134
rect 31166 41186 31218 41198
rect 32286 41186 32338 41198
rect 32846 41186 32898 41198
rect 33742 41186 33794 41198
rect 31826 41134 31838 41186
rect 31890 41134 31902 41186
rect 32498 41134 32510 41186
rect 32562 41134 32574 41186
rect 33282 41134 33294 41186
rect 33346 41134 33358 41186
rect 34290 41134 34302 41186
rect 34354 41134 34366 41186
rect 37314 41134 37326 41186
rect 37378 41134 37390 41186
rect 44258 41134 44270 41186
rect 44322 41134 44334 41186
rect 48066 41134 48078 41186
rect 48130 41134 48142 41186
rect 31166 41122 31218 41134
rect 32286 41122 32338 41134
rect 32846 41122 32898 41134
rect 33742 41122 33794 41134
rect 12910 41074 12962 41086
rect 12910 41010 12962 41022
rect 13470 41074 13522 41086
rect 13470 41010 13522 41022
rect 13694 41074 13746 41086
rect 13694 41010 13746 41022
rect 19966 41074 20018 41086
rect 19966 41010 20018 41022
rect 20526 41074 20578 41086
rect 20526 41010 20578 41022
rect 20750 41074 20802 41086
rect 20750 41010 20802 41022
rect 29374 41074 29426 41086
rect 29374 41010 29426 41022
rect 32958 41074 33010 41086
rect 32958 41010 33010 41022
rect 33854 41074 33906 41086
rect 33854 41010 33906 41022
rect 34638 41074 34690 41086
rect 34638 41010 34690 41022
rect 35086 41074 35138 41086
rect 35086 41010 35138 41022
rect 36094 41074 36146 41086
rect 36094 41010 36146 41022
rect 40574 41074 40626 41086
rect 40574 41010 40626 41022
rect 11342 40962 11394 40974
rect 11342 40898 11394 40910
rect 20638 40962 20690 40974
rect 20638 40898 20690 40910
rect 25230 40962 25282 40974
rect 25230 40898 25282 40910
rect 31278 40962 31330 40974
rect 31278 40898 31330 40910
rect 31390 40962 31442 40974
rect 31390 40898 31442 40910
rect 32062 40962 32114 40974
rect 32062 40898 32114 40910
rect 32174 40962 32226 40974
rect 32174 40898 32226 40910
rect 33518 40962 33570 40974
rect 33518 40898 33570 40910
rect 33630 40962 33682 40974
rect 33630 40898 33682 40910
rect 34974 40962 35026 40974
rect 34974 40898 35026 40910
rect 35982 40962 36034 40974
rect 35982 40898 36034 40910
rect 40686 40962 40738 40974
rect 40686 40898 40738 40910
rect 1344 40794 48608 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 48608 40794
rect 1344 40708 48608 40742
rect 24446 40626 24498 40638
rect 18722 40574 18734 40626
rect 18786 40574 18798 40626
rect 18946 40574 18958 40626
rect 19010 40574 19022 40626
rect 24446 40562 24498 40574
rect 25902 40626 25954 40638
rect 25902 40562 25954 40574
rect 27694 40626 27746 40638
rect 27694 40562 27746 40574
rect 28926 40626 28978 40638
rect 28926 40562 28978 40574
rect 30494 40626 30546 40638
rect 30494 40562 30546 40574
rect 30606 40626 30658 40638
rect 30606 40562 30658 40574
rect 31614 40626 31666 40638
rect 31614 40562 31666 40574
rect 32398 40626 32450 40638
rect 32398 40562 32450 40574
rect 12798 40514 12850 40526
rect 14142 40514 14194 40526
rect 23998 40514 24050 40526
rect 31390 40514 31442 40526
rect 10322 40462 10334 40514
rect 10386 40462 10398 40514
rect 13122 40462 13134 40514
rect 13186 40462 13198 40514
rect 13794 40462 13806 40514
rect 13858 40462 13870 40514
rect 15922 40462 15934 40514
rect 15986 40462 15998 40514
rect 18050 40462 18062 40514
rect 18114 40462 18126 40514
rect 20178 40462 20190 40514
rect 20242 40462 20254 40514
rect 21746 40462 21758 40514
rect 21810 40462 21822 40514
rect 22642 40462 22654 40514
rect 22706 40462 22718 40514
rect 25554 40462 25566 40514
rect 25618 40462 25630 40514
rect 12798 40450 12850 40462
rect 14142 40450 14194 40462
rect 23998 40450 24050 40462
rect 31390 40450 31442 40462
rect 32286 40514 32338 40526
rect 34526 40514 34578 40526
rect 47070 40514 47122 40526
rect 33842 40462 33854 40514
rect 33906 40462 33918 40514
rect 36530 40462 36542 40514
rect 36594 40462 36606 40514
rect 32286 40450 32338 40462
rect 34526 40450 34578 40462
rect 47070 40450 47122 40462
rect 47966 40514 48018 40526
rect 47966 40450 48018 40462
rect 24222 40402 24274 40414
rect 25230 40402 25282 40414
rect 4610 40350 4622 40402
rect 4674 40350 4686 40402
rect 9650 40350 9662 40402
rect 9714 40350 9726 40402
rect 15698 40350 15710 40402
rect 15762 40350 15774 40402
rect 16258 40350 16270 40402
rect 16322 40350 16334 40402
rect 18162 40350 18174 40402
rect 18226 40350 18238 40402
rect 18498 40350 18510 40402
rect 18562 40350 18574 40402
rect 20066 40350 20078 40402
rect 20130 40350 20142 40402
rect 21186 40350 21198 40402
rect 21250 40350 21262 40402
rect 23202 40350 23214 40402
rect 23266 40350 23278 40402
rect 24658 40350 24670 40402
rect 24722 40350 24734 40402
rect 24222 40338 24274 40350
rect 25230 40338 25282 40350
rect 26014 40402 26066 40414
rect 27246 40402 27298 40414
rect 26674 40350 26686 40402
rect 26738 40350 26750 40402
rect 26014 40338 26066 40350
rect 27246 40338 27298 40350
rect 27470 40402 27522 40414
rect 27470 40338 27522 40350
rect 27806 40402 27858 40414
rect 27806 40338 27858 40350
rect 28030 40402 28082 40414
rect 28702 40402 28754 40414
rect 30382 40402 30434 40414
rect 28466 40350 28478 40402
rect 28530 40350 28542 40402
rect 29138 40350 29150 40402
rect 29202 40350 29214 40402
rect 30146 40350 30158 40402
rect 30210 40350 30222 40402
rect 28030 40338 28082 40350
rect 28702 40338 28754 40350
rect 30382 40338 30434 40350
rect 30718 40402 30770 40414
rect 30718 40338 30770 40350
rect 31502 40402 31554 40414
rect 31502 40338 31554 40350
rect 32062 40402 32114 40414
rect 34302 40402 34354 40414
rect 40910 40402 40962 40414
rect 33618 40350 33630 40402
rect 33682 40350 33694 40402
rect 38882 40350 38894 40402
rect 38946 40350 38958 40402
rect 32062 40338 32114 40350
rect 34302 40338 34354 40350
rect 40910 40338 40962 40350
rect 41470 40402 41522 40414
rect 41470 40338 41522 40350
rect 41918 40402 41970 40414
rect 41918 40338 41970 40350
rect 42590 40402 42642 40414
rect 42590 40338 42642 40350
rect 44606 40402 44658 40414
rect 45614 40402 45666 40414
rect 45042 40350 45054 40402
rect 45106 40350 45118 40402
rect 44606 40338 44658 40350
rect 45614 40338 45666 40350
rect 45726 40402 45778 40414
rect 47294 40402 47346 40414
rect 46610 40350 46622 40402
rect 46674 40350 46686 40402
rect 45726 40338 45778 40350
rect 47294 40338 47346 40350
rect 47742 40402 47794 40414
rect 47742 40338 47794 40350
rect 24334 40290 24386 40302
rect 34414 40290 34466 40302
rect 47518 40290 47570 40302
rect 1698 40238 1710 40290
rect 1762 40238 1774 40290
rect 3826 40238 3838 40290
rect 3890 40238 3902 40290
rect 26450 40238 26462 40290
rect 26514 40238 26526 40290
rect 28914 40238 28926 40290
rect 28978 40238 28990 40290
rect 46274 40238 46286 40290
rect 46338 40238 46350 40290
rect 12450 40182 12462 40234
rect 12514 40182 12526 40234
rect 24334 40226 24386 40238
rect 34414 40226 34466 40238
rect 47518 40226 47570 40238
rect 16494 40178 16546 40190
rect 16494 40114 16546 40126
rect 16718 40178 16770 40190
rect 16718 40114 16770 40126
rect 16830 40178 16882 40190
rect 16830 40114 16882 40126
rect 32398 40178 32450 40190
rect 32398 40114 32450 40126
rect 34078 40178 34130 40190
rect 34078 40114 34130 40126
rect 1344 40010 48608 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 48608 40010
rect 1344 39924 48608 39958
rect 19070 39842 19122 39854
rect 19070 39778 19122 39790
rect 29150 39842 29202 39854
rect 29150 39778 29202 39790
rect 30270 39842 30322 39854
rect 30270 39778 30322 39790
rect 32062 39842 32114 39854
rect 32062 39778 32114 39790
rect 44942 39842 44994 39854
rect 44942 39778 44994 39790
rect 26910 39730 26962 39742
rect 4162 39678 4174 39730
rect 4226 39678 4238 39730
rect 9650 39678 9662 39730
rect 9714 39678 9726 39730
rect 16706 39678 16718 39730
rect 16770 39678 16782 39730
rect 18834 39678 18846 39730
rect 18898 39678 18910 39730
rect 26002 39678 26014 39730
rect 26066 39678 26078 39730
rect 26910 39666 26962 39678
rect 31838 39730 31890 39742
rect 31838 39666 31890 39678
rect 35982 39730 36034 39742
rect 35982 39666 36034 39678
rect 36318 39730 36370 39742
rect 36318 39666 36370 39678
rect 37326 39730 37378 39742
rect 37326 39666 37378 39678
rect 38782 39730 38834 39742
rect 39666 39678 39678 39730
rect 39730 39678 39742 39730
rect 41682 39678 41694 39730
rect 41746 39678 41758 39730
rect 45266 39678 45278 39730
rect 45330 39678 45342 39730
rect 47394 39678 47406 39730
rect 47458 39678 47470 39730
rect 38782 39666 38834 39678
rect 2718 39618 2770 39630
rect 10222 39618 10274 39630
rect 6738 39566 6750 39618
rect 6802 39566 6814 39618
rect 2718 39554 2770 39566
rect 10222 39554 10274 39566
rect 14478 39618 14530 39630
rect 20078 39618 20130 39630
rect 27246 39618 27298 39630
rect 15922 39566 15934 39618
rect 15986 39566 15998 39618
rect 19506 39566 19518 39618
rect 19570 39566 19582 39618
rect 21298 39566 21310 39618
rect 21362 39566 21374 39618
rect 22194 39566 22206 39618
rect 22258 39566 22270 39618
rect 23090 39566 23102 39618
rect 23154 39566 23166 39618
rect 14478 39554 14530 39566
rect 20078 39554 20130 39566
rect 27246 39554 27298 39566
rect 27694 39618 27746 39630
rect 27694 39554 27746 39566
rect 28478 39618 28530 39630
rect 28478 39554 28530 39566
rect 29262 39618 29314 39630
rect 29262 39554 29314 39566
rect 29710 39618 29762 39630
rect 30494 39618 30546 39630
rect 30034 39566 30046 39618
rect 30098 39566 30110 39618
rect 29710 39554 29762 39566
rect 30494 39554 30546 39566
rect 30718 39618 30770 39630
rect 30718 39554 30770 39566
rect 32286 39618 32338 39630
rect 35646 39618 35698 39630
rect 35298 39566 35310 39618
rect 35362 39566 35374 39618
rect 32286 39554 32338 39566
rect 35646 39554 35698 39566
rect 37438 39618 37490 39630
rect 42030 39618 42082 39630
rect 37650 39566 37662 39618
rect 37714 39566 37726 39618
rect 39442 39566 39454 39618
rect 39506 39566 39518 39618
rect 40898 39566 40910 39618
rect 40962 39566 40974 39618
rect 41234 39566 41246 39618
rect 41298 39566 41310 39618
rect 37438 39554 37490 39566
rect 42030 39554 42082 39566
rect 42590 39618 42642 39630
rect 42590 39554 42642 39566
rect 44830 39618 44882 39630
rect 48066 39566 48078 39618
rect 48130 39566 48142 39618
rect 44830 39554 44882 39566
rect 3390 39506 3442 39518
rect 3390 39442 3442 39454
rect 3502 39506 3554 39518
rect 3502 39442 3554 39454
rect 3838 39506 3890 39518
rect 3838 39442 3890 39454
rect 4510 39506 4562 39518
rect 4510 39442 4562 39454
rect 4734 39506 4786 39518
rect 10110 39506 10162 39518
rect 7522 39454 7534 39506
rect 7586 39454 7598 39506
rect 4734 39442 4786 39454
rect 10110 39442 10162 39454
rect 15486 39506 15538 39518
rect 19854 39506 19906 39518
rect 32734 39506 32786 39518
rect 19618 39454 19630 39506
rect 19682 39454 19694 39506
rect 20738 39454 20750 39506
rect 20802 39454 20814 39506
rect 21410 39454 21422 39506
rect 21474 39454 21486 39506
rect 23874 39454 23886 39506
rect 23938 39454 23950 39506
rect 15486 39442 15538 39454
rect 19854 39442 19906 39454
rect 32734 39442 32786 39454
rect 32958 39506 33010 39518
rect 32958 39442 33010 39454
rect 34526 39506 34578 39518
rect 34526 39442 34578 39454
rect 34638 39506 34690 39518
rect 34638 39442 34690 39454
rect 34862 39506 34914 39518
rect 34862 39442 34914 39454
rect 35758 39506 35810 39518
rect 35758 39442 35810 39454
rect 36430 39506 36482 39518
rect 36430 39442 36482 39454
rect 36990 39506 37042 39518
rect 42478 39506 42530 39518
rect 41346 39454 41358 39506
rect 41410 39454 41422 39506
rect 36990 39442 37042 39454
rect 42478 39442 42530 39454
rect 44046 39506 44098 39518
rect 44046 39442 44098 39454
rect 2830 39394 2882 39406
rect 2830 39330 2882 39342
rect 3054 39394 3106 39406
rect 3054 39330 3106 39342
rect 3166 39394 3218 39406
rect 3166 39330 3218 39342
rect 4062 39394 4114 39406
rect 4062 39330 4114 39342
rect 4622 39394 4674 39406
rect 4622 39330 4674 39342
rect 9998 39394 10050 39406
rect 9998 39330 10050 39342
rect 10446 39394 10498 39406
rect 10446 39330 10498 39342
rect 12350 39394 12402 39406
rect 12350 39330 12402 39342
rect 14142 39394 14194 39406
rect 14142 39330 14194 39342
rect 15374 39394 15426 39406
rect 15374 39330 15426 39342
rect 20414 39394 20466 39406
rect 26686 39394 26738 39406
rect 22418 39342 22430 39394
rect 22482 39342 22494 39394
rect 22642 39342 22654 39394
rect 22706 39342 22718 39394
rect 20414 39330 20466 39342
rect 26686 39330 26738 39342
rect 28590 39394 28642 39406
rect 28590 39330 28642 39342
rect 30830 39394 30882 39406
rect 30830 39330 30882 39342
rect 33070 39394 33122 39406
rect 33070 39330 33122 39342
rect 34190 39394 34242 39406
rect 34190 39330 34242 39342
rect 34974 39394 35026 39406
rect 34974 39330 35026 39342
rect 37214 39394 37266 39406
rect 42366 39394 42418 39406
rect 40450 39342 40462 39394
rect 40514 39342 40526 39394
rect 37214 39330 37266 39342
rect 42366 39330 42418 39342
rect 43822 39394 43874 39406
rect 43822 39330 43874 39342
rect 44158 39394 44210 39406
rect 44158 39330 44210 39342
rect 44382 39394 44434 39406
rect 44382 39330 44434 39342
rect 1344 39226 48608 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 48608 39226
rect 1344 39140 48608 39174
rect 8542 39058 8594 39070
rect 8542 38994 8594 39006
rect 10110 39058 10162 39070
rect 10110 38994 10162 39006
rect 29374 39058 29426 39070
rect 29374 38994 29426 39006
rect 31278 39058 31330 39070
rect 31278 38994 31330 39006
rect 31950 39058 32002 39070
rect 31950 38994 32002 39006
rect 39790 39058 39842 39070
rect 39790 38994 39842 39006
rect 43150 39058 43202 39070
rect 43150 38994 43202 39006
rect 45838 39058 45890 39070
rect 45838 38994 45890 39006
rect 46734 39058 46786 39070
rect 46734 38994 46786 39006
rect 46846 39058 46898 39070
rect 46846 38994 46898 39006
rect 9662 38946 9714 38958
rect 6066 38894 6078 38946
rect 6130 38894 6142 38946
rect 9662 38882 9714 38894
rect 10334 38946 10386 38958
rect 10334 38882 10386 38894
rect 10446 38946 10498 38958
rect 12910 38946 12962 38958
rect 11666 38894 11678 38946
rect 11730 38894 11742 38946
rect 10446 38882 10498 38894
rect 12910 38882 12962 38894
rect 13134 38946 13186 38958
rect 13134 38882 13186 38894
rect 18174 38946 18226 38958
rect 18174 38882 18226 38894
rect 18286 38946 18338 38958
rect 27694 38946 27746 38958
rect 20066 38894 20078 38946
rect 20130 38894 20142 38946
rect 18286 38882 18338 38894
rect 27694 38882 27746 38894
rect 29710 38946 29762 38958
rect 29710 38882 29762 38894
rect 31726 38946 31778 38958
rect 31726 38882 31778 38894
rect 32174 38946 32226 38958
rect 32174 38882 32226 38894
rect 32398 38946 32450 38958
rect 35870 38946 35922 38958
rect 33282 38894 33294 38946
rect 33346 38894 33358 38946
rect 32398 38882 32450 38894
rect 35870 38882 35922 38894
rect 38446 38946 38498 38958
rect 45390 38946 45442 38958
rect 45042 38894 45054 38946
rect 45106 38894 45118 38946
rect 38446 38882 38498 38894
rect 45390 38882 45442 38894
rect 46398 38946 46450 38958
rect 46398 38882 46450 38894
rect 46622 38946 46674 38958
rect 47842 38894 47854 38946
rect 47906 38894 47918 38946
rect 46622 38882 46674 38894
rect 8878 38834 8930 38846
rect 4610 38782 4622 38834
rect 4674 38782 4686 38834
rect 5282 38782 5294 38834
rect 5346 38782 5358 38834
rect 8878 38770 8930 38782
rect 11006 38834 11058 38846
rect 11006 38770 11058 38782
rect 12014 38834 12066 38846
rect 12014 38770 12066 38782
rect 12462 38834 12514 38846
rect 16942 38834 16994 38846
rect 13570 38782 13582 38834
rect 13634 38782 13646 38834
rect 12462 38770 12514 38782
rect 16942 38770 16994 38782
rect 18398 38834 18450 38846
rect 23214 38834 23266 38846
rect 26238 38834 26290 38846
rect 35198 38834 35250 38846
rect 19842 38782 19854 38834
rect 19906 38782 19918 38834
rect 20514 38782 20526 38834
rect 20578 38782 20590 38834
rect 21298 38782 21310 38834
rect 21362 38782 21374 38834
rect 22530 38782 22542 38834
rect 22594 38782 22606 38834
rect 24434 38782 24446 38834
rect 24498 38782 24510 38834
rect 26002 38782 26014 38834
rect 26066 38782 26078 38834
rect 27122 38782 27134 38834
rect 27186 38782 27198 38834
rect 29138 38782 29150 38834
rect 29202 38782 29214 38834
rect 33170 38782 33182 38834
rect 33234 38782 33246 38834
rect 33730 38782 33742 38834
rect 33794 38782 33806 38834
rect 34066 38782 34078 38834
rect 34130 38782 34142 38834
rect 18398 38770 18450 38782
rect 23214 38770 23266 38782
rect 26238 38770 26290 38782
rect 35198 38770 35250 38782
rect 36094 38834 36146 38846
rect 36094 38770 36146 38782
rect 36990 38834 37042 38846
rect 36990 38770 37042 38782
rect 37214 38834 37266 38846
rect 37774 38834 37826 38846
rect 37538 38782 37550 38834
rect 37602 38782 37614 38834
rect 37214 38770 37266 38782
rect 37774 38770 37826 38782
rect 37998 38834 38050 38846
rect 37998 38770 38050 38782
rect 38110 38834 38162 38846
rect 38110 38770 38162 38782
rect 39678 38834 39730 38846
rect 39678 38770 39730 38782
rect 39902 38834 39954 38846
rect 43038 38834 43090 38846
rect 41122 38782 41134 38834
rect 41186 38782 41198 38834
rect 42130 38782 42142 38834
rect 42194 38782 42206 38834
rect 39902 38770 39954 38782
rect 43038 38770 43090 38782
rect 43374 38834 43426 38846
rect 45614 38834 45666 38846
rect 43698 38782 43710 38834
rect 43762 38782 43774 38834
rect 44146 38782 44158 38834
rect 44210 38782 44222 38834
rect 44930 38782 44942 38834
rect 44994 38782 45006 38834
rect 43374 38770 43426 38782
rect 45614 38770 45666 38782
rect 45726 38834 45778 38846
rect 45726 38770 45778 38782
rect 45950 38834 46002 38846
rect 45950 38770 46002 38782
rect 46958 38834 47010 38846
rect 46958 38770 47010 38782
rect 47406 38834 47458 38846
rect 47406 38770 47458 38782
rect 48190 38834 48242 38846
rect 48190 38770 48242 38782
rect 9886 38722 9938 38734
rect 1698 38670 1710 38722
rect 1762 38670 1774 38722
rect 3826 38670 3838 38722
rect 3890 38670 3902 38722
rect 8194 38670 8206 38722
rect 8258 38670 8270 38722
rect 9538 38670 9550 38722
rect 9602 38670 9614 38722
rect 9886 38658 9938 38670
rect 10782 38722 10834 38734
rect 12686 38722 12738 38734
rect 17838 38722 17890 38734
rect 25342 38722 25394 38734
rect 11330 38670 11342 38722
rect 11394 38670 11406 38722
rect 14242 38670 14254 38722
rect 14306 38670 14318 38722
rect 16370 38670 16382 38722
rect 16434 38670 16446 38722
rect 19954 38670 19966 38722
rect 20018 38670 20030 38722
rect 20850 38670 20862 38722
rect 20914 38670 20926 38722
rect 10782 38658 10834 38670
rect 12686 38658 12738 38670
rect 17838 38658 17890 38670
rect 25342 38658 25394 38670
rect 26798 38722 26850 38734
rect 26798 38658 26850 38670
rect 31390 38722 31442 38734
rect 31390 38658 31442 38670
rect 36430 38722 36482 38734
rect 36430 38658 36482 38670
rect 40126 38722 40178 38734
rect 40126 38658 40178 38670
rect 40350 38722 40402 38734
rect 47518 38722 47570 38734
rect 41346 38670 41358 38722
rect 41410 38670 41422 38722
rect 41906 38670 41918 38722
rect 41970 38670 41982 38722
rect 40350 38658 40402 38670
rect 47518 38658 47570 38670
rect 32286 38610 32338 38622
rect 18834 38558 18846 38610
rect 18898 38558 18910 38610
rect 21746 38558 21758 38610
rect 21810 38558 21822 38610
rect 32286 38546 32338 38558
rect 35086 38610 35138 38622
rect 42018 38558 42030 38610
rect 42082 38558 42094 38610
rect 44370 38558 44382 38610
rect 44434 38558 44446 38610
rect 35086 38546 35138 38558
rect 1344 38442 48608 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 48608 38442
rect 1344 38356 48608 38390
rect 19406 38274 19458 38286
rect 19406 38210 19458 38222
rect 19630 38274 19682 38286
rect 19630 38210 19682 38222
rect 20190 38274 20242 38286
rect 20190 38210 20242 38222
rect 21422 38274 21474 38286
rect 21422 38210 21474 38222
rect 22206 38274 22258 38286
rect 22206 38210 22258 38222
rect 29150 38274 29202 38286
rect 29150 38210 29202 38222
rect 30382 38274 30434 38286
rect 30382 38210 30434 38222
rect 30830 38274 30882 38286
rect 32498 38222 32510 38274
rect 32562 38271 32574 38274
rect 32946 38271 32958 38274
rect 32562 38225 32958 38271
rect 32562 38222 32574 38225
rect 32946 38222 32958 38225
rect 33010 38222 33022 38274
rect 30830 38210 30882 38222
rect 2718 38162 2770 38174
rect 10446 38162 10498 38174
rect 6066 38110 6078 38162
rect 6130 38110 6142 38162
rect 2718 38098 2770 38110
rect 10446 38098 10498 38110
rect 10894 38162 10946 38174
rect 10894 38098 10946 38110
rect 11566 38162 11618 38174
rect 11566 38098 11618 38110
rect 12462 38162 12514 38174
rect 20302 38162 20354 38174
rect 17266 38110 17278 38162
rect 17330 38110 17342 38162
rect 12462 38098 12514 38110
rect 20302 38098 20354 38110
rect 29374 38162 29426 38174
rect 29374 38098 29426 38110
rect 29710 38162 29762 38174
rect 29710 38098 29762 38110
rect 32734 38162 32786 38174
rect 32734 38098 32786 38110
rect 33182 38162 33234 38174
rect 43598 38162 43650 38174
rect 34290 38110 34302 38162
rect 34354 38110 34366 38162
rect 36418 38110 36430 38162
rect 36482 38110 36494 38162
rect 39666 38110 39678 38162
rect 39730 38110 39742 38162
rect 43138 38110 43150 38162
rect 43202 38110 43214 38162
rect 47394 38110 47406 38162
rect 47458 38110 47470 38162
rect 33182 38098 33234 38110
rect 43598 38098 43650 38110
rect 3278 38050 3330 38062
rect 7310 38050 7362 38062
rect 3826 37998 3838 38050
rect 3890 37998 3902 38050
rect 3278 37986 3330 37998
rect 7310 37986 7362 37998
rect 8094 38050 8146 38062
rect 13694 38050 13746 38062
rect 18622 38050 18674 38062
rect 8418 37998 8430 38050
rect 8482 37998 8494 38050
rect 8754 37998 8766 38050
rect 8818 37998 8830 38050
rect 9650 37998 9662 38050
rect 9714 37998 9726 38050
rect 12226 37998 12238 38050
rect 12290 37998 12302 38050
rect 14354 37998 14366 38050
rect 14418 37998 14430 38050
rect 8094 37986 8146 37998
rect 13694 37986 13746 37998
rect 18622 37986 18674 37998
rect 18846 38050 18898 38062
rect 18846 37986 18898 37998
rect 19070 38050 19122 38062
rect 19070 37986 19122 37998
rect 19742 38050 19794 38062
rect 19742 37986 19794 37998
rect 21534 38050 21586 38062
rect 29598 38050 29650 38062
rect 26562 37998 26574 38050
rect 26626 37998 26638 38050
rect 21534 37986 21586 37998
rect 29598 37986 29650 37998
rect 32062 38050 32114 38062
rect 32062 37986 32114 37998
rect 32398 38050 32450 38062
rect 43486 38050 43538 38062
rect 33618 37998 33630 38050
rect 33682 37998 33694 38050
rect 40114 37998 40126 38050
rect 40178 37998 40190 38050
rect 41234 37998 41246 38050
rect 41298 37998 41310 38050
rect 41906 37998 41918 38050
rect 41970 37998 41982 38050
rect 43026 37998 43038 38050
rect 43090 37998 43102 38050
rect 32398 37986 32450 37998
rect 43486 37986 43538 37998
rect 44158 38050 44210 38062
rect 44818 37998 44830 38050
rect 44882 37998 44894 38050
rect 45714 37998 45726 38050
rect 45778 37998 45790 38050
rect 46722 37998 46734 38050
rect 46786 37998 46798 38050
rect 47506 37998 47518 38050
rect 47570 37998 47582 38050
rect 44158 37986 44210 37998
rect 2830 37938 2882 37950
rect 2830 37874 2882 37886
rect 3166 37938 3218 37950
rect 3166 37874 3218 37886
rect 6190 37938 6242 37950
rect 6190 37874 6242 37886
rect 6414 37938 6466 37950
rect 6414 37874 6466 37886
rect 7870 37938 7922 37950
rect 10334 37938 10386 37950
rect 9202 37886 9214 37938
rect 9266 37886 9278 37938
rect 9874 37886 9886 37938
rect 9938 37886 9950 37938
rect 7870 37874 7922 37886
rect 10334 37874 10386 37886
rect 12574 37938 12626 37950
rect 17726 37938 17778 37950
rect 15138 37886 15150 37938
rect 15202 37886 15214 37938
rect 12574 37874 12626 37886
rect 17726 37874 17778 37886
rect 18398 37938 18450 37950
rect 18398 37874 18450 37886
rect 19294 37938 19346 37950
rect 19294 37874 19346 37886
rect 20414 37938 20466 37950
rect 20414 37874 20466 37886
rect 21422 37938 21474 37950
rect 21422 37874 21474 37886
rect 22094 37938 22146 37950
rect 22094 37874 22146 37886
rect 22206 37938 22258 37950
rect 30270 37938 30322 37950
rect 22978 37886 22990 37938
rect 23042 37886 23054 37938
rect 22206 37874 22258 37886
rect 30270 37874 30322 37886
rect 30382 37938 30434 37950
rect 30382 37874 30434 37886
rect 30942 37938 30994 37950
rect 30942 37874 30994 37886
rect 32174 37938 32226 37950
rect 45826 37886 45838 37938
rect 45890 37886 45902 37938
rect 47618 37886 47630 37938
rect 47682 37886 47694 37938
rect 32174 37874 32226 37886
rect 2606 37826 2658 37838
rect 7982 37826 8034 37838
rect 6962 37774 6974 37826
rect 7026 37774 7038 37826
rect 2606 37762 2658 37774
rect 7982 37762 8034 37774
rect 18062 37826 18114 37838
rect 18062 37762 18114 37774
rect 28590 37826 28642 37838
rect 28590 37762 28642 37774
rect 29822 37826 29874 37838
rect 29822 37762 29874 37774
rect 31502 37826 31554 37838
rect 31502 37762 31554 37774
rect 43710 37826 43762 37838
rect 43710 37762 43762 37774
rect 45054 37826 45106 37838
rect 46846 37826 46898 37838
rect 45154 37774 45166 37826
rect 45218 37774 45230 37826
rect 45054 37762 45106 37774
rect 46846 37762 46898 37774
rect 1344 37658 48608 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 48608 37658
rect 1344 37572 48608 37606
rect 17838 37490 17890 37502
rect 17838 37426 17890 37438
rect 19406 37490 19458 37502
rect 19406 37426 19458 37438
rect 19630 37490 19682 37502
rect 19630 37426 19682 37438
rect 23662 37490 23714 37502
rect 23662 37426 23714 37438
rect 25678 37490 25730 37502
rect 25678 37426 25730 37438
rect 27582 37490 27634 37502
rect 27582 37426 27634 37438
rect 33742 37490 33794 37502
rect 33742 37426 33794 37438
rect 34750 37490 34802 37502
rect 34750 37426 34802 37438
rect 34862 37490 34914 37502
rect 34862 37426 34914 37438
rect 35646 37490 35698 37502
rect 35646 37426 35698 37438
rect 36094 37490 36146 37502
rect 36094 37426 36146 37438
rect 41022 37490 41074 37502
rect 41022 37426 41074 37438
rect 42590 37490 42642 37502
rect 42590 37426 42642 37438
rect 46286 37490 46338 37502
rect 47058 37438 47070 37490
rect 47122 37438 47134 37490
rect 46286 37426 46338 37438
rect 8542 37378 8594 37390
rect 5730 37326 5742 37378
rect 5794 37326 5806 37378
rect 8542 37314 8594 37326
rect 15150 37378 15202 37390
rect 15150 37314 15202 37326
rect 23886 37378 23938 37390
rect 23886 37314 23938 37326
rect 23998 37378 24050 37390
rect 23998 37314 24050 37326
rect 26574 37378 26626 37390
rect 26574 37314 26626 37326
rect 34190 37378 34242 37390
rect 34190 37314 34242 37326
rect 35198 37378 35250 37390
rect 35198 37314 35250 37326
rect 43038 37378 43090 37390
rect 43038 37314 43090 37326
rect 44494 37378 44546 37390
rect 44494 37314 44546 37326
rect 46174 37378 46226 37390
rect 46174 37314 46226 37326
rect 46958 37378 47010 37390
rect 47730 37326 47742 37378
rect 47794 37326 47806 37378
rect 46958 37314 47010 37326
rect 3054 37266 3106 37278
rect 8094 37266 8146 37278
rect 3490 37214 3502 37266
rect 3554 37214 3566 37266
rect 5058 37214 5070 37266
rect 5122 37214 5134 37266
rect 3054 37202 3106 37214
rect 8094 37202 8146 37214
rect 8766 37266 8818 37278
rect 14142 37266 14194 37278
rect 9762 37214 9774 37266
rect 9826 37214 9838 37266
rect 8766 37202 8818 37214
rect 14142 37202 14194 37214
rect 14814 37266 14866 37278
rect 14814 37202 14866 37214
rect 16494 37266 16546 37278
rect 16494 37202 16546 37214
rect 16830 37266 16882 37278
rect 16830 37202 16882 37214
rect 17502 37266 17554 37278
rect 19070 37266 19122 37278
rect 18610 37214 18622 37266
rect 18674 37214 18686 37266
rect 17502 37202 17554 37214
rect 19070 37202 19122 37214
rect 19742 37266 19794 37278
rect 25566 37266 25618 37278
rect 27806 37266 27858 37278
rect 33630 37266 33682 37278
rect 22978 37214 22990 37266
rect 23042 37214 23054 37266
rect 27570 37214 27582 37266
rect 27634 37214 27646 37266
rect 28578 37214 28590 37266
rect 28642 37263 28654 37266
rect 28914 37263 28926 37266
rect 28642 37217 28926 37263
rect 28642 37214 28654 37217
rect 28914 37214 28926 37217
rect 28978 37214 28990 37266
rect 29138 37214 29150 37266
rect 29202 37214 29214 37266
rect 19742 37202 19794 37214
rect 25566 37202 25618 37214
rect 27806 37202 27858 37214
rect 33630 37202 33682 37214
rect 33966 37266 34018 37278
rect 33966 37202 34018 37214
rect 34638 37266 34690 37278
rect 34638 37202 34690 37214
rect 34974 37266 35026 37278
rect 41918 37266 41970 37278
rect 37090 37214 37102 37266
rect 37154 37214 37166 37266
rect 34974 37202 35026 37214
rect 41918 37202 41970 37214
rect 43934 37266 43986 37278
rect 47058 37214 47070 37266
rect 47122 37214 47134 37266
rect 47842 37214 47854 37266
rect 47906 37214 47918 37266
rect 43934 37202 43986 37214
rect 8654 37154 8706 37166
rect 13918 37154 13970 37166
rect 7858 37102 7870 37154
rect 7922 37102 7934 37154
rect 10546 37102 10558 37154
rect 10610 37102 10622 37154
rect 12674 37102 12686 37154
rect 12738 37102 12750 37154
rect 8654 37090 8706 37102
rect 13918 37090 13970 37102
rect 14478 37154 14530 37166
rect 14478 37090 14530 37102
rect 18174 37154 18226 37166
rect 23550 37154 23602 37166
rect 20066 37102 20078 37154
rect 20130 37102 20142 37154
rect 22194 37102 22206 37154
rect 22258 37102 22270 37154
rect 18174 37090 18226 37102
rect 23550 37090 23602 37102
rect 24670 37154 24722 37166
rect 33182 37154 33234 37166
rect 29922 37102 29934 37154
rect 29986 37102 29998 37154
rect 32050 37102 32062 37154
rect 32114 37102 32126 37154
rect 24670 37090 24722 37102
rect 33182 37090 33234 37102
rect 33854 37154 33906 37166
rect 40910 37154 40962 37166
rect 37874 37102 37886 37154
rect 37938 37102 37950 37154
rect 40002 37102 40014 37154
rect 40066 37102 40078 37154
rect 33854 37090 33906 37102
rect 40910 37090 40962 37102
rect 2942 37042 2994 37054
rect 2942 36978 2994 36990
rect 3278 37042 3330 37054
rect 3278 36978 3330 36990
rect 33070 37042 33122 37054
rect 33070 36978 33122 36990
rect 46286 37042 46338 37054
rect 46286 36978 46338 36990
rect 1344 36874 48608 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 48608 36874
rect 1344 36788 48608 36822
rect 19854 36706 19906 36718
rect 18498 36654 18510 36706
rect 18562 36654 18574 36706
rect 19854 36642 19906 36654
rect 38110 36706 38162 36718
rect 38110 36642 38162 36654
rect 40350 36706 40402 36718
rect 40350 36642 40402 36654
rect 43038 36706 43090 36718
rect 43038 36642 43090 36654
rect 44942 36594 44994 36606
rect 1698 36542 1710 36594
rect 1762 36542 1774 36594
rect 3826 36542 3838 36594
rect 3890 36542 3902 36594
rect 14914 36542 14926 36594
rect 14978 36542 14990 36594
rect 17042 36542 17054 36594
rect 17106 36542 17118 36594
rect 18162 36542 18174 36594
rect 18226 36542 18238 36594
rect 25330 36542 25342 36594
rect 25394 36542 25406 36594
rect 25666 36542 25678 36594
rect 25730 36542 25742 36594
rect 30594 36542 30606 36594
rect 30658 36542 30670 36594
rect 32610 36542 32622 36594
rect 32674 36542 32686 36594
rect 34738 36542 34750 36594
rect 34802 36542 34814 36594
rect 37874 36542 37886 36594
rect 37938 36542 37950 36594
rect 41346 36542 41358 36594
rect 41410 36542 41422 36594
rect 43810 36542 43822 36594
rect 43874 36542 43886 36594
rect 48178 36542 48190 36594
rect 48242 36542 48254 36594
rect 44942 36530 44994 36542
rect 20526 36482 20578 36494
rect 4610 36430 4622 36482
rect 4674 36430 4686 36482
rect 12002 36430 12014 36482
rect 12066 36430 12078 36482
rect 14130 36430 14142 36482
rect 14194 36430 14206 36482
rect 18050 36430 18062 36482
rect 18114 36430 18126 36482
rect 18834 36430 18846 36482
rect 18898 36430 18910 36482
rect 19282 36430 19294 36482
rect 19346 36430 19358 36482
rect 20526 36418 20578 36430
rect 20862 36482 20914 36494
rect 20862 36418 20914 36430
rect 21534 36482 21586 36494
rect 31054 36482 31106 36494
rect 37662 36482 37714 36494
rect 22530 36430 22542 36482
rect 22594 36430 22606 36482
rect 28578 36430 28590 36482
rect 28642 36430 28654 36482
rect 29250 36430 29262 36482
rect 29314 36430 29326 36482
rect 31938 36430 31950 36482
rect 32002 36430 32014 36482
rect 21534 36418 21586 36430
rect 31054 36418 31106 36430
rect 37662 36418 37714 36430
rect 38334 36482 38386 36494
rect 38334 36418 38386 36430
rect 40574 36482 40626 36494
rect 43250 36430 43262 36482
rect 43314 36430 43326 36482
rect 43922 36430 43934 36482
rect 43986 36430 43998 36482
rect 45378 36430 45390 36482
rect 45442 36430 45454 36482
rect 40574 36418 40626 36430
rect 5742 36370 5794 36382
rect 19966 36370 20018 36382
rect 29710 36370 29762 36382
rect 9762 36318 9774 36370
rect 9826 36318 9838 36370
rect 23202 36318 23214 36370
rect 23266 36318 23278 36370
rect 27794 36318 27806 36370
rect 27858 36318 27870 36370
rect 5742 36306 5794 36318
rect 19966 36306 20018 36318
rect 29710 36306 29762 36318
rect 36990 36370 37042 36382
rect 36990 36306 37042 36318
rect 37326 36370 37378 36382
rect 37326 36306 37378 36318
rect 37550 36370 37602 36382
rect 37550 36306 37602 36318
rect 39790 36370 39842 36382
rect 39790 36306 39842 36318
rect 40014 36370 40066 36382
rect 40014 36306 40066 36318
rect 40126 36370 40178 36382
rect 40126 36306 40178 36318
rect 41022 36370 41074 36382
rect 46050 36318 46062 36370
rect 46114 36318 46126 36370
rect 41022 36306 41074 36318
rect 5630 36258 5682 36270
rect 5630 36194 5682 36206
rect 12574 36258 12626 36270
rect 12574 36194 12626 36206
rect 20638 36258 20690 36270
rect 20638 36194 20690 36206
rect 21646 36258 21698 36270
rect 21646 36194 21698 36206
rect 21758 36258 21810 36270
rect 21758 36194 21810 36206
rect 21982 36258 22034 36270
rect 21982 36194 22034 36206
rect 29486 36258 29538 36270
rect 29486 36194 29538 36206
rect 29598 36258 29650 36270
rect 29598 36194 29650 36206
rect 29822 36258 29874 36270
rect 29822 36194 29874 36206
rect 30606 36258 30658 36270
rect 30606 36194 30658 36206
rect 30718 36258 30770 36270
rect 30718 36194 30770 36206
rect 30942 36258 30994 36270
rect 30942 36194 30994 36206
rect 36430 36258 36482 36270
rect 36430 36194 36482 36206
rect 37102 36258 37154 36270
rect 37102 36194 37154 36206
rect 42254 36258 42306 36270
rect 42254 36194 42306 36206
rect 42702 36258 42754 36270
rect 42702 36194 42754 36206
rect 44830 36258 44882 36270
rect 44830 36194 44882 36206
rect 1344 36090 48608 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 48608 36090
rect 1344 36004 48608 36038
rect 3278 35922 3330 35934
rect 3278 35858 3330 35870
rect 7086 35922 7138 35934
rect 7086 35858 7138 35870
rect 7198 35922 7250 35934
rect 7198 35858 7250 35870
rect 7310 35922 7362 35934
rect 7310 35858 7362 35870
rect 8206 35922 8258 35934
rect 8206 35858 8258 35870
rect 8878 35922 8930 35934
rect 8878 35858 8930 35870
rect 18174 35922 18226 35934
rect 18174 35858 18226 35870
rect 22654 35922 22706 35934
rect 22654 35858 22706 35870
rect 23998 35922 24050 35934
rect 23998 35858 24050 35870
rect 24558 35922 24610 35934
rect 28142 35922 28194 35934
rect 26898 35870 26910 35922
rect 26962 35870 26974 35922
rect 24558 35858 24610 35870
rect 28142 35858 28194 35870
rect 28814 35922 28866 35934
rect 28814 35858 28866 35870
rect 29150 35922 29202 35934
rect 29150 35858 29202 35870
rect 29598 35922 29650 35934
rect 29598 35858 29650 35870
rect 29934 35922 29986 35934
rect 29934 35858 29986 35870
rect 30830 35922 30882 35934
rect 30830 35858 30882 35870
rect 32062 35922 32114 35934
rect 36094 35922 36146 35934
rect 33394 35870 33406 35922
rect 33458 35870 33470 35922
rect 32062 35858 32114 35870
rect 36094 35858 36146 35870
rect 39902 35922 39954 35934
rect 39902 35858 39954 35870
rect 41694 35922 41746 35934
rect 41694 35858 41746 35870
rect 41918 35922 41970 35934
rect 41918 35858 41970 35870
rect 47518 35922 47570 35934
rect 47518 35858 47570 35870
rect 48190 35922 48242 35934
rect 48190 35858 48242 35870
rect 3726 35810 3778 35822
rect 4398 35810 4450 35822
rect 4162 35758 4174 35810
rect 4226 35758 4238 35810
rect 3726 35746 3778 35758
rect 4398 35746 4450 35758
rect 8654 35810 8706 35822
rect 8654 35746 8706 35758
rect 8990 35810 9042 35822
rect 25566 35810 25618 35822
rect 28254 35810 28306 35822
rect 21298 35758 21310 35810
rect 21362 35758 21374 35810
rect 27346 35758 27358 35810
rect 27410 35758 27422 35810
rect 8990 35746 9042 35758
rect 25566 35746 25618 35758
rect 28254 35746 28306 35758
rect 30046 35810 30098 35822
rect 46286 35810 46338 35822
rect 31378 35758 31390 35810
rect 31442 35758 31454 35810
rect 30046 35746 30098 35758
rect 46286 35746 46338 35758
rect 47070 35810 47122 35822
rect 47070 35746 47122 35758
rect 47406 35810 47458 35822
rect 47842 35758 47854 35810
rect 47906 35758 47918 35810
rect 47406 35746 47458 35758
rect 3166 35698 3218 35710
rect 3166 35634 3218 35646
rect 3502 35698 3554 35710
rect 3502 35634 3554 35646
rect 4062 35698 4114 35710
rect 4062 35634 4114 35646
rect 4846 35698 4898 35710
rect 4846 35634 4898 35646
rect 6862 35698 6914 35710
rect 6862 35634 6914 35646
rect 7982 35698 8034 35710
rect 7982 35634 8034 35646
rect 8094 35698 8146 35710
rect 8094 35634 8146 35646
rect 8430 35698 8482 35710
rect 22542 35698 22594 35710
rect 13794 35646 13806 35698
rect 13858 35646 13870 35698
rect 22082 35646 22094 35698
rect 22146 35646 22158 35698
rect 8430 35634 8482 35646
rect 22542 35634 22594 35646
rect 22766 35698 22818 35710
rect 22766 35634 22818 35646
rect 23214 35698 23266 35710
rect 23214 35634 23266 35646
rect 23774 35698 23826 35710
rect 23774 35634 23826 35646
rect 24110 35698 24162 35710
rect 24110 35634 24162 35646
rect 24446 35698 24498 35710
rect 24446 35634 24498 35646
rect 24782 35698 24834 35710
rect 24782 35634 24834 35646
rect 25230 35698 25282 35710
rect 25230 35634 25282 35646
rect 25342 35698 25394 35710
rect 25342 35634 25394 35646
rect 25790 35698 25842 35710
rect 30606 35698 30658 35710
rect 26674 35646 26686 35698
rect 26738 35646 26750 35698
rect 27682 35646 27694 35698
rect 27746 35646 27758 35698
rect 30370 35646 30382 35698
rect 30434 35646 30446 35698
rect 25790 35634 25842 35646
rect 30606 35634 30658 35646
rect 30718 35698 30770 35710
rect 31726 35698 31778 35710
rect 31042 35646 31054 35698
rect 31106 35646 31118 35698
rect 30718 35634 30770 35646
rect 31726 35634 31778 35646
rect 32174 35698 32226 35710
rect 32174 35634 32226 35646
rect 33070 35698 33122 35710
rect 33070 35634 33122 35646
rect 35982 35698 36034 35710
rect 35982 35634 36034 35646
rect 36318 35698 36370 35710
rect 39790 35698 39842 35710
rect 36530 35646 36542 35698
rect 36594 35646 36606 35698
rect 36318 35634 36370 35646
rect 39790 35634 39842 35646
rect 42030 35698 42082 35710
rect 46062 35698 46114 35710
rect 42466 35646 42478 35698
rect 42530 35646 42542 35698
rect 42030 35634 42082 35646
rect 46062 35634 46114 35646
rect 46398 35698 46450 35710
rect 46398 35634 46450 35646
rect 17726 35586 17778 35598
rect 10882 35534 10894 35586
rect 10946 35534 10958 35586
rect 13010 35534 13022 35586
rect 13074 35534 13086 35586
rect 17726 35522 17778 35534
rect 18062 35586 18114 35598
rect 18062 35522 18114 35534
rect 18734 35586 18786 35598
rect 18734 35522 18786 35534
rect 19182 35586 19234 35598
rect 19182 35522 19234 35534
rect 23662 35586 23714 35598
rect 23662 35522 23714 35534
rect 26014 35586 26066 35598
rect 26014 35522 26066 35534
rect 34078 35586 34130 35598
rect 34078 35522 34130 35534
rect 34526 35586 34578 35598
rect 46958 35586 47010 35598
rect 37314 35534 37326 35586
rect 37378 35534 37390 35586
rect 39442 35534 39454 35586
rect 39506 35534 39518 35586
rect 43138 35534 43150 35586
rect 43202 35534 43214 35586
rect 45266 35534 45278 35586
rect 45330 35534 45342 35586
rect 34526 35522 34578 35534
rect 46958 35522 47010 35534
rect 5070 35474 5122 35486
rect 5070 35410 5122 35422
rect 6638 35474 6690 35486
rect 6638 35410 6690 35422
rect 33966 35474 34018 35486
rect 33966 35410 34018 35422
rect 45838 35474 45890 35486
rect 45838 35410 45890 35422
rect 46622 35474 46674 35486
rect 46622 35410 46674 35422
rect 1344 35306 48608 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 48608 35306
rect 1344 35220 48608 35254
rect 11902 35138 11954 35150
rect 3938 35086 3950 35138
rect 4002 35086 4014 35138
rect 11902 35074 11954 35086
rect 12238 35138 12290 35150
rect 12238 35074 12290 35086
rect 12910 35138 12962 35150
rect 12910 35074 12962 35086
rect 23774 35138 23826 35150
rect 23774 35074 23826 35086
rect 25006 35138 25058 35150
rect 25006 35074 25058 35086
rect 36990 35138 37042 35150
rect 36990 35074 37042 35086
rect 37550 35138 37602 35150
rect 37550 35074 37602 35086
rect 37774 35138 37826 35150
rect 37774 35074 37826 35086
rect 43262 35138 43314 35150
rect 43262 35074 43314 35086
rect 3054 35026 3106 35038
rect 3054 34962 3106 34974
rect 8094 35026 8146 35038
rect 19966 35026 20018 35038
rect 8866 34974 8878 35026
rect 8930 34974 8942 35026
rect 9538 34974 9550 35026
rect 9602 34974 9614 35026
rect 17938 34974 17950 35026
rect 18002 34974 18014 35026
rect 8094 34962 8146 34974
rect 19966 34962 20018 34974
rect 20302 35026 20354 35038
rect 26350 35026 26402 35038
rect 23538 34974 23550 35026
rect 23602 34974 23614 35026
rect 20302 34962 20354 34974
rect 26350 34962 26402 34974
rect 29262 35026 29314 35038
rect 29262 34962 29314 34974
rect 35422 35026 35474 35038
rect 44942 35026 44994 35038
rect 37314 34974 37326 35026
rect 37378 34974 37390 35026
rect 40450 34974 40462 35026
rect 40514 34974 40526 35026
rect 42578 34974 42590 35026
rect 42642 34974 42654 35026
rect 43474 34974 43486 35026
rect 43538 34974 43550 35026
rect 48178 34974 48190 35026
rect 48242 34974 48254 35026
rect 35422 34962 35474 34974
rect 44942 34962 44994 34974
rect 2158 34914 2210 34926
rect 2158 34850 2210 34862
rect 3614 34914 3666 34926
rect 3614 34850 3666 34862
rect 4398 34914 4450 34926
rect 4398 34850 4450 34862
rect 4622 34914 4674 34926
rect 4622 34850 4674 34862
rect 6750 34914 6802 34926
rect 6750 34850 6802 34862
rect 7086 34914 7138 34926
rect 7086 34850 7138 34862
rect 7310 34914 7362 34926
rect 9214 34914 9266 34926
rect 11454 34914 11506 34926
rect 14030 34914 14082 34926
rect 22094 34914 22146 34926
rect 8754 34862 8766 34914
rect 8818 34862 8830 34914
rect 9986 34862 9998 34914
rect 10050 34862 10062 34914
rect 13458 34862 13470 34914
rect 13522 34862 13534 34914
rect 15138 34862 15150 34914
rect 15202 34862 15214 34914
rect 18274 34862 18286 34914
rect 18338 34862 18350 34914
rect 7310 34850 7362 34862
rect 9214 34850 9266 34862
rect 11454 34850 11506 34862
rect 14030 34850 14082 34862
rect 22094 34850 22146 34862
rect 22430 34914 22482 34926
rect 37102 34914 37154 34926
rect 23426 34862 23438 34914
rect 23490 34862 23502 34914
rect 34178 34862 34190 34914
rect 34242 34862 34254 34914
rect 22430 34850 22482 34862
rect 37102 34850 37154 34862
rect 38558 34914 38610 34926
rect 43038 34914 43090 34926
rect 39778 34862 39790 34914
rect 39842 34862 39854 34914
rect 45378 34862 45390 34914
rect 45442 34862 45454 34914
rect 38558 34850 38610 34862
rect 43038 34850 43090 34862
rect 2270 34802 2322 34814
rect 2270 34738 2322 34750
rect 2606 34802 2658 34814
rect 2606 34738 2658 34750
rect 2942 34802 2994 34814
rect 2942 34738 2994 34750
rect 3166 34802 3218 34814
rect 3166 34738 3218 34750
rect 4510 34802 4562 34814
rect 4510 34738 4562 34750
rect 5630 34802 5682 34814
rect 5630 34738 5682 34750
rect 5966 34802 6018 34814
rect 5966 34738 6018 34750
rect 7758 34802 7810 34814
rect 7758 34738 7810 34750
rect 7982 34802 8034 34814
rect 7982 34738 8034 34750
rect 8206 34802 8258 34814
rect 8206 34738 8258 34750
rect 11230 34802 11282 34814
rect 11230 34738 11282 34750
rect 11566 34802 11618 34814
rect 11566 34738 11618 34750
rect 12462 34802 12514 34814
rect 12462 34738 12514 34750
rect 12798 34802 12850 34814
rect 12798 34738 12850 34750
rect 13806 34802 13858 34814
rect 19406 34802 19458 34814
rect 15810 34750 15822 34802
rect 15874 34750 15886 34802
rect 13806 34738 13858 34750
rect 19406 34738 19458 34750
rect 22206 34802 22258 34814
rect 22206 34738 22258 34750
rect 24222 34802 24274 34814
rect 24222 34738 24274 34750
rect 24558 34802 24610 34814
rect 24558 34738 24610 34750
rect 24894 34802 24946 34814
rect 24894 34738 24946 34750
rect 25790 34802 25842 34814
rect 25790 34738 25842 34750
rect 27022 34802 27074 34814
rect 38222 34802 38274 34814
rect 29922 34750 29934 34802
rect 29986 34750 29998 34802
rect 27022 34738 27074 34750
rect 38222 34738 38274 34750
rect 38334 34802 38386 34814
rect 38334 34738 38386 34750
rect 43598 34802 43650 34814
rect 43598 34738 43650 34750
rect 43822 34802 43874 34814
rect 46050 34750 46062 34802
rect 46114 34750 46126 34802
rect 43822 34738 43874 34750
rect 2494 34690 2546 34702
rect 2494 34626 2546 34638
rect 6862 34690 6914 34702
rect 6862 34626 6914 34638
rect 13694 34690 13746 34702
rect 13694 34626 13746 34638
rect 13918 34690 13970 34702
rect 13918 34626 13970 34638
rect 14702 34690 14754 34702
rect 14702 34626 14754 34638
rect 18510 34690 18562 34702
rect 18510 34626 18562 34638
rect 18622 34690 18674 34702
rect 18622 34626 18674 34638
rect 18734 34690 18786 34702
rect 18734 34626 18786 34638
rect 18846 34690 18898 34702
rect 18846 34626 18898 34638
rect 19294 34690 19346 34702
rect 19294 34626 19346 34638
rect 20862 34690 20914 34702
rect 20862 34626 20914 34638
rect 21870 34690 21922 34702
rect 21870 34626 21922 34638
rect 23214 34690 23266 34702
rect 23214 34626 23266 34638
rect 25006 34690 25058 34702
rect 25006 34626 25058 34638
rect 25454 34690 25506 34702
rect 25454 34626 25506 34638
rect 25678 34690 25730 34702
rect 25678 34626 25730 34638
rect 26910 34690 26962 34702
rect 26910 34626 26962 34638
rect 27470 34690 27522 34702
rect 27470 34626 27522 34638
rect 27918 34690 27970 34702
rect 27918 34626 27970 34638
rect 29374 34690 29426 34702
rect 36430 34690 36482 34702
rect 36082 34638 36094 34690
rect 36146 34638 36158 34690
rect 29374 34626 29426 34638
rect 36430 34626 36482 34638
rect 38894 34690 38946 34702
rect 38894 34626 38946 34638
rect 39342 34690 39394 34702
rect 39342 34626 39394 34638
rect 44270 34690 44322 34702
rect 44270 34626 44322 34638
rect 1344 34522 48608 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 48608 34522
rect 1344 34436 48608 34470
rect 13246 34354 13298 34366
rect 13246 34290 13298 34302
rect 13582 34354 13634 34366
rect 13582 34290 13634 34302
rect 16382 34354 16434 34366
rect 16382 34290 16434 34302
rect 18398 34354 18450 34366
rect 18398 34290 18450 34302
rect 19294 34354 19346 34366
rect 19294 34290 19346 34302
rect 23998 34354 24050 34366
rect 36654 34354 36706 34366
rect 32162 34302 32174 34354
rect 32226 34302 32238 34354
rect 41234 34302 41246 34354
rect 41298 34302 41310 34354
rect 23998 34290 24050 34302
rect 36654 34290 36706 34302
rect 13470 34242 13522 34254
rect 2482 34190 2494 34242
rect 2546 34190 2558 34242
rect 5954 34190 5966 34242
rect 6018 34190 6030 34242
rect 13470 34178 13522 34190
rect 14142 34242 14194 34254
rect 14142 34178 14194 34190
rect 16494 34242 16546 34254
rect 16494 34178 16546 34190
rect 17950 34242 18002 34254
rect 17950 34178 18002 34190
rect 18958 34242 19010 34254
rect 18958 34178 19010 34190
rect 23774 34242 23826 34254
rect 23774 34178 23826 34190
rect 24110 34242 24162 34254
rect 39678 34242 39730 34254
rect 26450 34190 26462 34242
rect 26514 34190 26526 34242
rect 29698 34190 29710 34242
rect 29762 34190 29774 34242
rect 33842 34190 33854 34242
rect 33906 34190 33918 34242
rect 24110 34178 24162 34190
rect 39678 34178 39730 34190
rect 40014 34242 40066 34254
rect 40910 34242 40962 34254
rect 40338 34190 40350 34242
rect 40402 34190 40414 34242
rect 40014 34178 40066 34190
rect 40910 34178 40962 34190
rect 18174 34130 18226 34142
rect 19182 34130 19234 34142
rect 1810 34078 1822 34130
rect 1874 34078 1886 34130
rect 5170 34078 5182 34130
rect 5234 34078 5246 34130
rect 9762 34078 9774 34130
rect 9826 34078 9838 34130
rect 13010 34078 13022 34130
rect 13074 34078 13086 34130
rect 18610 34078 18622 34130
rect 18674 34078 18686 34130
rect 18174 34066 18226 34078
rect 19182 34066 19234 34078
rect 19406 34130 19458 34142
rect 24334 34130 24386 34142
rect 36542 34130 36594 34142
rect 19618 34078 19630 34130
rect 19682 34078 19694 34130
rect 20514 34078 20526 34130
rect 20578 34078 20590 34130
rect 25778 34078 25790 34130
rect 25842 34078 25854 34130
rect 29026 34078 29038 34130
rect 29090 34078 29102 34130
rect 32386 34078 32398 34130
rect 32450 34078 32462 34130
rect 33058 34078 33070 34130
rect 33122 34078 33134 34130
rect 36306 34078 36318 34130
rect 36370 34078 36382 34130
rect 19406 34066 19458 34078
rect 24334 34066 24386 34078
rect 36542 34066 36594 34078
rect 36766 34130 36818 34142
rect 36978 34078 36990 34130
rect 37042 34078 37054 34130
rect 42130 34078 42142 34130
rect 42194 34078 42206 34130
rect 43138 34078 43150 34130
rect 43202 34078 43214 34130
rect 36766 34066 36818 34078
rect 13358 34018 13410 34030
rect 4610 33966 4622 34018
rect 4674 33966 4686 34018
rect 8082 33966 8094 34018
rect 8146 33966 8158 34018
rect 10546 33966 10558 34018
rect 10610 33966 10622 34018
rect 12674 33966 12686 34018
rect 12738 33966 12750 34018
rect 13358 33954 13410 33966
rect 14478 34018 14530 34030
rect 14478 33954 14530 33966
rect 15038 34018 15090 34030
rect 15038 33954 15090 33966
rect 15822 34018 15874 34030
rect 15822 33954 15874 33966
rect 18286 34018 18338 34030
rect 18286 33954 18338 33966
rect 20078 34018 20130 34030
rect 25454 34018 25506 34030
rect 37438 34018 37490 34030
rect 21298 33966 21310 34018
rect 21362 33966 21374 34018
rect 23426 33966 23438 34018
rect 23490 33966 23502 34018
rect 28578 33966 28590 34018
rect 28642 33966 28654 34018
rect 31826 33966 31838 34018
rect 31890 33966 31902 34018
rect 35970 33966 35982 34018
rect 36034 33966 36046 34018
rect 20078 33954 20130 33966
rect 25454 33954 25506 33966
rect 37438 33954 37490 33966
rect 38670 34018 38722 34030
rect 38670 33954 38722 33966
rect 39342 34018 39394 34030
rect 39342 33954 39394 33966
rect 41694 34018 41746 34030
rect 42466 33966 42478 34018
rect 42530 33966 42542 34018
rect 46946 33966 46958 34018
rect 47010 33966 47022 34018
rect 41694 33954 41746 33966
rect 14590 33906 14642 33918
rect 14590 33842 14642 33854
rect 1344 33738 48608 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 48608 33738
rect 1344 33652 48608 33686
rect 11118 33570 11170 33582
rect 44158 33570 44210 33582
rect 30258 33518 30270 33570
rect 30322 33567 30334 33570
rect 30706 33567 30718 33570
rect 30322 33521 30718 33567
rect 30322 33518 30334 33521
rect 30706 33518 30718 33521
rect 30770 33567 30782 33570
rect 31602 33567 31614 33570
rect 30770 33521 31614 33567
rect 30770 33518 30782 33521
rect 31602 33518 31614 33521
rect 31666 33518 31678 33570
rect 11118 33506 11170 33518
rect 44158 33506 44210 33518
rect 46398 33570 46450 33582
rect 46398 33506 46450 33518
rect 46622 33570 46674 33582
rect 46622 33506 46674 33518
rect 48078 33570 48130 33582
rect 48078 33506 48130 33518
rect 9438 33458 9490 33470
rect 11230 33458 11282 33470
rect 22430 33458 22482 33470
rect 29486 33458 29538 33470
rect 7970 33406 7982 33458
rect 8034 33406 8046 33458
rect 10322 33406 10334 33458
rect 10386 33406 10398 33458
rect 13570 33406 13582 33458
rect 13634 33406 13646 33458
rect 15698 33406 15710 33458
rect 15762 33406 15774 33458
rect 20402 33406 20414 33458
rect 20466 33406 20478 33458
rect 26898 33406 26910 33458
rect 26962 33406 26974 33458
rect 9438 33394 9490 33406
rect 11230 33394 11282 33406
rect 22430 33394 22482 33406
rect 29486 33394 29538 33406
rect 30718 33458 30770 33470
rect 30718 33394 30770 33406
rect 31166 33458 31218 33470
rect 44942 33458 44994 33470
rect 32050 33406 32062 33458
rect 32114 33406 32126 33458
rect 33058 33406 33070 33458
rect 33122 33406 33134 33458
rect 43698 33406 43710 33458
rect 43762 33406 43774 33458
rect 46050 33406 46062 33458
rect 46114 33406 46126 33458
rect 31166 33394 31218 33406
rect 44942 33394 44994 33406
rect 22318 33346 22370 33358
rect 7746 33294 7758 33346
rect 7810 33294 7822 33346
rect 9874 33294 9886 33346
rect 9938 33294 9950 33346
rect 16370 33294 16382 33346
rect 16434 33294 16446 33346
rect 17490 33294 17502 33346
rect 17554 33294 17566 33346
rect 21522 33294 21534 33346
rect 21586 33294 21598 33346
rect 22318 33282 22370 33294
rect 22542 33346 22594 33358
rect 22542 33282 22594 33294
rect 22878 33346 22930 33358
rect 22878 33282 22930 33294
rect 23550 33346 23602 33358
rect 23550 33282 23602 33294
rect 23886 33346 23938 33358
rect 27582 33346 27634 33358
rect 24322 33294 24334 33346
rect 24386 33294 24398 33346
rect 26002 33294 26014 33346
rect 26066 33294 26078 33346
rect 23886 33282 23938 33294
rect 27582 33282 27634 33294
rect 28254 33346 28306 33358
rect 28254 33282 28306 33294
rect 29262 33346 29314 33358
rect 29262 33282 29314 33294
rect 29374 33346 29426 33358
rect 37326 33346 37378 33358
rect 29810 33294 29822 33346
rect 29874 33294 29886 33346
rect 35970 33294 35982 33346
rect 36034 33294 36046 33346
rect 29374 33282 29426 33294
rect 37326 33282 37378 33294
rect 37550 33346 37602 33358
rect 37550 33282 37602 33294
rect 38222 33346 38274 33358
rect 38222 33282 38274 33294
rect 38782 33346 38834 33358
rect 38782 33282 38834 33294
rect 39790 33346 39842 33358
rect 39790 33282 39842 33294
rect 40014 33346 40066 33358
rect 44046 33346 44098 33358
rect 40898 33294 40910 33346
rect 40962 33294 40974 33346
rect 41570 33294 41582 33346
rect 41634 33294 41646 33346
rect 40014 33282 40066 33294
rect 44046 33282 44098 33294
rect 45502 33346 45554 33358
rect 45502 33282 45554 33294
rect 47070 33346 47122 33358
rect 47070 33282 47122 33294
rect 47630 33346 47682 33358
rect 47630 33282 47682 33294
rect 7086 33234 7138 33246
rect 23214 33234 23266 33246
rect 32286 33234 32338 33246
rect 37886 33234 37938 33246
rect 39230 33234 39282 33246
rect 18274 33182 18286 33234
rect 18338 33182 18350 33234
rect 21298 33182 21310 33234
rect 21362 33182 21374 33234
rect 24546 33182 24558 33234
rect 24610 33182 24622 33234
rect 25218 33182 25230 33234
rect 25282 33182 25294 33234
rect 35186 33182 35198 33234
rect 35250 33182 35262 33234
rect 38546 33182 38558 33234
rect 38610 33182 38622 33234
rect 7086 33170 7138 33182
rect 23214 33170 23266 33182
rect 32286 33170 32338 33182
rect 37886 33170 37938 33182
rect 39230 33170 39282 33182
rect 39454 33234 39506 33246
rect 39454 33170 39506 33182
rect 39902 33234 39954 33246
rect 39902 33170 39954 33182
rect 40350 33234 40402 33246
rect 40350 33170 40402 33182
rect 45838 33234 45890 33246
rect 45838 33170 45890 33182
rect 46062 33234 46114 33246
rect 48078 33234 48130 33246
rect 46062 33170 46114 33182
rect 47966 33178 48018 33190
rect 6750 33122 6802 33134
rect 6750 33058 6802 33070
rect 6974 33122 7026 33134
rect 6974 33058 7026 33070
rect 8990 33122 9042 33134
rect 8990 33058 9042 33070
rect 23550 33122 23602 33134
rect 23550 33058 23602 33070
rect 24894 33122 24946 33134
rect 27358 33122 27410 33134
rect 26226 33070 26238 33122
rect 26290 33070 26302 33122
rect 24894 33058 24946 33070
rect 27358 33058 27410 33070
rect 27694 33122 27746 33134
rect 27694 33058 27746 33070
rect 27918 33122 27970 33134
rect 27918 33058 27970 33070
rect 28590 33122 28642 33134
rect 28590 33058 28642 33070
rect 29598 33122 29650 33134
rect 29598 33058 29650 33070
rect 30382 33122 30434 33134
rect 30382 33058 30434 33070
rect 31614 33122 31666 33134
rect 31614 33058 31666 33070
rect 32062 33122 32114 33134
rect 32062 33058 32114 33070
rect 36430 33122 36482 33134
rect 36430 33058 36482 33070
rect 37438 33122 37490 33134
rect 37438 33058 37490 33070
rect 39118 33122 39170 33134
rect 39118 33058 39170 33070
rect 44158 33122 44210 33134
rect 48078 33170 48130 33182
rect 47966 33114 48018 33126
rect 44158 33058 44210 33070
rect 1344 32954 48608 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 48608 32954
rect 1344 32868 48608 32902
rect 14478 32786 14530 32798
rect 14478 32722 14530 32734
rect 14590 32786 14642 32798
rect 18174 32786 18226 32798
rect 15138 32734 15150 32786
rect 15202 32734 15214 32786
rect 14590 32722 14642 32734
rect 18174 32722 18226 32734
rect 30270 32786 30322 32798
rect 30270 32722 30322 32734
rect 33966 32786 34018 32798
rect 33966 32722 34018 32734
rect 34078 32786 34130 32798
rect 34078 32722 34130 32734
rect 34862 32786 34914 32798
rect 34862 32722 34914 32734
rect 39790 32786 39842 32798
rect 44482 32734 44494 32786
rect 44546 32734 44558 32786
rect 39790 32722 39842 32734
rect 8766 32674 8818 32686
rect 4946 32622 4958 32674
rect 5010 32622 5022 32674
rect 8766 32610 8818 32622
rect 14142 32674 14194 32686
rect 24558 32674 24610 32686
rect 29822 32674 29874 32686
rect 33742 32674 33794 32686
rect 20178 32622 20190 32674
rect 20242 32622 20254 32674
rect 26674 32622 26686 32674
rect 26738 32622 26750 32674
rect 27906 32622 27918 32674
rect 27970 32622 27982 32674
rect 33394 32622 33406 32674
rect 33458 32622 33470 32674
rect 14142 32610 14194 32622
rect 24558 32610 24610 32622
rect 29822 32610 29874 32622
rect 33742 32610 33794 32622
rect 34750 32674 34802 32686
rect 40238 32674 40290 32686
rect 37202 32622 37214 32674
rect 37266 32622 37278 32674
rect 34750 32610 34802 32622
rect 40238 32610 40290 32622
rect 44942 32674 44994 32686
rect 48066 32622 48078 32674
rect 48130 32622 48142 32674
rect 44942 32610 44994 32622
rect 8878 32562 8930 32574
rect 13918 32562 13970 32574
rect 8306 32510 8318 32562
rect 8370 32510 8382 32562
rect 10434 32510 10446 32562
rect 10498 32510 10510 32562
rect 8878 32498 8930 32510
rect 13918 32498 13970 32510
rect 14366 32562 14418 32574
rect 16830 32562 16882 32574
rect 18398 32562 18450 32574
rect 24670 32562 24722 32574
rect 28814 32562 28866 32574
rect 14802 32510 14814 32562
rect 14866 32510 14878 32562
rect 15362 32510 15374 32562
rect 15426 32510 15438 32562
rect 17938 32510 17950 32562
rect 18002 32510 18014 32562
rect 18610 32510 18622 32562
rect 18674 32510 18686 32562
rect 23538 32510 23550 32562
rect 23602 32510 23614 32562
rect 25218 32510 25230 32562
rect 25282 32510 25294 32562
rect 28466 32510 28478 32562
rect 28530 32510 28542 32562
rect 14366 32498 14418 32510
rect 16830 32498 16882 32510
rect 18398 32498 18450 32510
rect 24670 32498 24722 32510
rect 28814 32498 28866 32510
rect 29038 32562 29090 32574
rect 29038 32498 29090 32510
rect 29374 32562 29426 32574
rect 29374 32498 29426 32510
rect 33070 32562 33122 32574
rect 33070 32498 33122 32510
rect 34190 32562 34242 32574
rect 34190 32498 34242 32510
rect 34302 32562 34354 32574
rect 34302 32498 34354 32510
rect 35422 32562 35474 32574
rect 39678 32562 39730 32574
rect 36530 32510 36542 32562
rect 36594 32510 36606 32562
rect 35422 32498 35474 32510
rect 39678 32498 39730 32510
rect 39902 32562 39954 32574
rect 41122 32510 41134 32562
rect 41186 32510 41198 32562
rect 45938 32510 45950 32562
rect 46002 32510 46014 32562
rect 48178 32510 48190 32562
rect 48242 32510 48254 32562
rect 39902 32498 39954 32510
rect 9662 32450 9714 32462
rect 16046 32450 16098 32462
rect 11106 32398 11118 32450
rect 11170 32398 11182 32450
rect 13234 32398 13246 32450
rect 13298 32398 13310 32450
rect 9662 32386 9714 32398
rect 16046 32386 16098 32398
rect 16382 32450 16434 32462
rect 16382 32386 16434 32398
rect 17502 32450 17554 32462
rect 17502 32386 17554 32398
rect 18286 32450 18338 32462
rect 29262 32450 29314 32462
rect 28018 32398 28030 32450
rect 28082 32398 28094 32450
rect 18286 32386 18338 32398
rect 29262 32386 29314 32398
rect 35982 32450 36034 32462
rect 39330 32398 39342 32450
rect 39394 32398 39406 32450
rect 41906 32398 41918 32450
rect 41970 32398 41982 32450
rect 44034 32398 44046 32450
rect 44098 32398 44110 32450
rect 35982 32386 36034 32398
rect 8766 32338 8818 32350
rect 8766 32274 8818 32286
rect 17390 32338 17442 32350
rect 17390 32274 17442 32286
rect 1344 32170 48608 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 48608 32170
rect 1344 32084 48608 32118
rect 43362 31950 43374 32002
rect 43426 31999 43438 32002
rect 44034 31999 44046 32002
rect 43426 31953 44046 31999
rect 43426 31950 43438 31953
rect 44034 31950 44046 31953
rect 44098 31950 44110 32002
rect 26014 31890 26066 31902
rect 38334 31890 38386 31902
rect 43038 31890 43090 31902
rect 4610 31838 4622 31890
rect 4674 31838 4686 31890
rect 7746 31838 7758 31890
rect 7810 31838 7822 31890
rect 15362 31838 15374 31890
rect 15426 31838 15438 31890
rect 17490 31838 17502 31890
rect 17554 31838 17566 31890
rect 17826 31838 17838 31890
rect 17890 31838 17902 31890
rect 22866 31838 22878 31890
rect 22930 31838 22942 31890
rect 24994 31838 25006 31890
rect 25058 31838 25070 31890
rect 29922 31838 29934 31890
rect 29986 31838 29998 31890
rect 32050 31838 32062 31890
rect 32114 31838 32126 31890
rect 33954 31838 33966 31890
rect 34018 31838 34030 31890
rect 42354 31838 42366 31890
rect 42418 31838 42430 31890
rect 26014 31826 26066 31838
rect 38334 31826 38386 31838
rect 43038 31826 43090 31838
rect 44270 31890 44322 31902
rect 44270 31826 44322 31838
rect 5966 31778 6018 31790
rect 1810 31726 1822 31778
rect 1874 31726 1886 31778
rect 5966 31714 6018 31726
rect 6414 31778 6466 31790
rect 13918 31778 13970 31790
rect 25902 31778 25954 31790
rect 10546 31726 10558 31778
rect 10610 31726 10622 31778
rect 13458 31726 13470 31778
rect 13522 31726 13534 31778
rect 14130 31726 14142 31778
rect 14194 31726 14206 31778
rect 14578 31726 14590 31778
rect 14642 31726 14654 31778
rect 20626 31726 20638 31778
rect 20690 31726 20702 31778
rect 22082 31726 22094 31778
rect 22146 31726 22158 31778
rect 6414 31714 6466 31726
rect 13918 31714 13970 31726
rect 25902 31714 25954 31726
rect 26126 31778 26178 31790
rect 26126 31714 26178 31726
rect 26798 31778 26850 31790
rect 26798 31714 26850 31726
rect 26910 31778 26962 31790
rect 26910 31714 26962 31726
rect 27358 31778 27410 31790
rect 27358 31714 27410 31726
rect 27694 31778 27746 31790
rect 27694 31714 27746 31726
rect 27918 31778 27970 31790
rect 45054 31778 45106 31790
rect 29138 31726 29150 31778
rect 29202 31726 29214 31778
rect 39554 31726 39566 31778
rect 39618 31726 39630 31778
rect 44818 31726 44830 31778
rect 44882 31726 44894 31778
rect 27918 31714 27970 31726
rect 45054 31714 45106 31726
rect 45390 31778 45442 31790
rect 45390 31714 45442 31726
rect 45726 31778 45778 31790
rect 45726 31714 45778 31726
rect 46062 31778 46114 31790
rect 46062 31714 46114 31726
rect 47406 31778 47458 31790
rect 47406 31714 47458 31726
rect 5630 31666 5682 31678
rect 2482 31614 2494 31666
rect 2546 31614 2558 31666
rect 5630 31602 5682 31614
rect 5742 31666 5794 31678
rect 5742 31602 5794 31614
rect 6190 31666 6242 31678
rect 6190 31602 6242 31614
rect 6862 31666 6914 31678
rect 6862 31602 6914 31614
rect 7086 31666 7138 31678
rect 11790 31666 11842 31678
rect 9874 31614 9886 31666
rect 9938 31614 9950 31666
rect 7086 31602 7138 31614
rect 11790 31602 11842 31614
rect 11902 31666 11954 31678
rect 11902 31602 11954 31614
rect 13806 31666 13858 31678
rect 21646 31666 21698 31678
rect 19954 31614 19966 31666
rect 20018 31614 20030 31666
rect 21298 31614 21310 31666
rect 21362 31614 21374 31666
rect 13806 31602 13858 31614
rect 21646 31602 21698 31614
rect 38670 31666 38722 31678
rect 43150 31666 43202 31678
rect 40226 31614 40238 31666
rect 40290 31614 40302 31666
rect 38670 31602 38722 31614
rect 43150 31602 43202 31614
rect 43710 31666 43762 31678
rect 43710 31602 43762 31614
rect 45166 31666 45218 31678
rect 45166 31602 45218 31614
rect 45950 31666 46002 31678
rect 45950 31602 46002 31614
rect 46398 31666 46450 31678
rect 46398 31602 46450 31614
rect 46846 31666 46898 31678
rect 46846 31602 46898 31614
rect 6638 31554 6690 31566
rect 6638 31490 6690 31502
rect 13694 31554 13746 31566
rect 13694 31490 13746 31502
rect 25678 31554 25730 31566
rect 25678 31490 25730 31502
rect 26574 31554 26626 31566
rect 26574 31490 26626 31502
rect 27022 31554 27074 31566
rect 27022 31490 27074 31502
rect 27806 31554 27858 31566
rect 27806 31490 27858 31502
rect 28366 31554 28418 31566
rect 28366 31490 28418 31502
rect 33182 31554 33234 31566
rect 33182 31490 33234 31502
rect 33518 31554 33570 31566
rect 33518 31490 33570 31502
rect 34638 31554 34690 31566
rect 34638 31490 34690 31502
rect 35198 31554 35250 31566
rect 35198 31490 35250 31502
rect 35982 31554 36034 31566
rect 35982 31490 36034 31502
rect 36542 31554 36594 31566
rect 36542 31490 36594 31502
rect 37102 31554 37154 31566
rect 37774 31554 37826 31566
rect 37426 31502 37438 31554
rect 37490 31502 37502 31554
rect 37102 31490 37154 31502
rect 37774 31490 37826 31502
rect 38782 31554 38834 31566
rect 38782 31490 38834 31502
rect 45278 31554 45330 31566
rect 45278 31490 45330 31502
rect 46510 31554 46562 31566
rect 46510 31490 46562 31502
rect 46958 31554 47010 31566
rect 46958 31490 47010 31502
rect 47966 31554 48018 31566
rect 47966 31490 48018 31502
rect 1344 31386 48608 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 48608 31386
rect 1344 31300 48608 31334
rect 6974 31218 7026 31230
rect 6974 31154 7026 31166
rect 7198 31218 7250 31230
rect 7198 31154 7250 31166
rect 8094 31218 8146 31230
rect 8094 31154 8146 31166
rect 8654 31218 8706 31230
rect 8654 31154 8706 31166
rect 16270 31218 16322 31230
rect 16270 31154 16322 31166
rect 20638 31218 20690 31230
rect 20638 31154 20690 31166
rect 21422 31218 21474 31230
rect 21422 31154 21474 31166
rect 22654 31218 22706 31230
rect 25902 31218 25954 31230
rect 25554 31166 25566 31218
rect 25618 31166 25630 31218
rect 22654 31154 22706 31166
rect 25902 31154 25954 31166
rect 26574 31218 26626 31230
rect 26574 31154 26626 31166
rect 26798 31218 26850 31230
rect 26798 31154 26850 31166
rect 27134 31218 27186 31230
rect 27134 31154 27186 31166
rect 27358 31218 27410 31230
rect 41358 31218 41410 31230
rect 32274 31166 32286 31218
rect 32338 31166 32350 31218
rect 27358 31154 27410 31166
rect 41358 31154 41410 31166
rect 41918 31218 41970 31230
rect 41918 31154 41970 31166
rect 43038 31218 43090 31230
rect 43038 31154 43090 31166
rect 43150 31218 43202 31230
rect 43150 31154 43202 31166
rect 43262 31218 43314 31230
rect 43262 31154 43314 31166
rect 44046 31218 44098 31230
rect 44046 31154 44098 31166
rect 44158 31218 44210 31230
rect 44158 31154 44210 31166
rect 7310 31106 7362 31118
rect 4386 31054 4398 31106
rect 4450 31054 4462 31106
rect 7310 31042 7362 31054
rect 7758 31106 7810 31118
rect 7758 31042 7810 31054
rect 7870 31106 7922 31118
rect 7870 31042 7922 31054
rect 8542 31106 8594 31118
rect 8542 31042 8594 31054
rect 8878 31106 8930 31118
rect 8878 31042 8930 31054
rect 10782 31106 10834 31118
rect 10782 31042 10834 31054
rect 14926 31106 14978 31118
rect 14926 31042 14978 31054
rect 20750 31106 20802 31118
rect 20750 31042 20802 31054
rect 27582 31106 27634 31118
rect 31614 31106 31666 31118
rect 29026 31054 29038 31106
rect 29090 31054 29102 31106
rect 27582 31042 27634 31054
rect 31614 31042 31666 31054
rect 44270 31106 44322 31118
rect 47170 31054 47182 31106
rect 47234 31054 47246 31106
rect 44270 31042 44322 31054
rect 8318 30994 8370 31006
rect 3714 30942 3726 30994
rect 3778 30942 3790 30994
rect 8318 30930 8370 30942
rect 11118 30994 11170 31006
rect 11118 30930 11170 30942
rect 11566 30994 11618 31006
rect 11566 30930 11618 30942
rect 12126 30994 12178 31006
rect 26126 30994 26178 31006
rect 31726 30994 31778 31006
rect 15474 30942 15486 30994
rect 15538 30942 15550 30994
rect 17378 30942 17390 30994
rect 17442 30942 17454 30994
rect 21858 30942 21870 30994
rect 21922 30942 21934 30994
rect 23650 30942 23662 30994
rect 23714 30942 23726 30994
rect 28018 30991 28030 30994
rect 12126 30930 12178 30942
rect 26126 30930 26178 30942
rect 27921 30945 28030 30991
rect 12574 30882 12626 30894
rect 6514 30830 6526 30882
rect 6578 30830 6590 30882
rect 12574 30818 12626 30830
rect 14142 30882 14194 30894
rect 14142 30818 14194 30830
rect 14590 30882 14642 30894
rect 14590 30818 14642 30830
rect 15150 30882 15202 30894
rect 22318 30882 22370 30894
rect 24222 30882 24274 30894
rect 16706 30830 16718 30882
rect 16770 30830 16782 30882
rect 18162 30830 18174 30882
rect 18226 30830 18238 30882
rect 20290 30830 20302 30882
rect 20354 30830 20366 30882
rect 23090 30830 23102 30882
rect 23154 30830 23166 30882
rect 15150 30818 15202 30830
rect 22318 30818 22370 30830
rect 24222 30818 24274 30830
rect 24670 30882 24722 30894
rect 24670 30818 24722 30830
rect 26686 30882 26738 30894
rect 26686 30818 26738 30830
rect 27246 30882 27298 30894
rect 27682 30830 27694 30882
rect 27746 30879 27758 30882
rect 27921 30879 27967 30945
rect 28018 30942 28030 30945
rect 28082 30942 28094 30994
rect 28242 30942 28254 30994
rect 28306 30942 28318 30994
rect 31726 30930 31778 30942
rect 31838 30994 31890 31006
rect 31838 30930 31890 30942
rect 34862 30994 34914 31006
rect 41134 30994 41186 31006
rect 43374 30994 43426 31006
rect 35298 30942 35310 30994
rect 35362 30942 35374 30994
rect 36530 30942 36542 30994
rect 36594 30942 36606 30994
rect 37426 30942 37438 30994
rect 37490 30942 37502 30994
rect 40898 30942 40910 30994
rect 40962 30942 40974 30994
rect 41570 30942 41582 30994
rect 41634 30942 41646 30994
rect 42802 30942 42814 30994
rect 42866 30942 42878 30994
rect 34862 30930 34914 30942
rect 41134 30930 41186 30942
rect 43374 30930 43426 30942
rect 43934 30994 43986 31006
rect 44482 30942 44494 30994
rect 44546 30942 44558 30994
rect 47954 30942 47966 30994
rect 48018 30942 48030 30994
rect 43934 30930 43986 30942
rect 33406 30882 33458 30894
rect 27746 30833 27967 30879
rect 27746 30830 27758 30833
rect 31154 30830 31166 30882
rect 31218 30830 31230 30882
rect 27246 30818 27298 30830
rect 33406 30818 33458 30830
rect 34302 30882 34354 30894
rect 34302 30818 34354 30830
rect 35758 30882 35810 30894
rect 41246 30882 41298 30894
rect 36194 30830 36206 30882
rect 36258 30830 36270 30882
rect 38098 30830 38110 30882
rect 38162 30830 38174 30882
rect 40226 30830 40238 30882
rect 40290 30830 40302 30882
rect 35758 30818 35810 30830
rect 41246 30818 41298 30830
rect 42030 30882 42082 30894
rect 42030 30818 42082 30830
rect 42478 30882 42530 30894
rect 45042 30830 45054 30882
rect 45106 30830 45118 30882
rect 42478 30818 42530 30830
rect 23998 30770 24050 30782
rect 23998 30706 24050 30718
rect 1344 30602 48608 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 48608 30602
rect 1344 30516 48608 30550
rect 25454 30434 25506 30446
rect 25454 30370 25506 30382
rect 27918 30434 27970 30446
rect 27918 30370 27970 30382
rect 31390 30434 31442 30446
rect 31390 30370 31442 30382
rect 34078 30434 34130 30446
rect 34078 30370 34130 30382
rect 13806 30322 13858 30334
rect 4610 30270 4622 30322
rect 4674 30270 4686 30322
rect 13806 30258 13858 30270
rect 22542 30322 22594 30334
rect 22542 30258 22594 30270
rect 30270 30322 30322 30334
rect 30270 30258 30322 30270
rect 32062 30322 32114 30334
rect 45266 30270 45278 30322
rect 45330 30270 45342 30322
rect 32062 30258 32114 30270
rect 5630 30210 5682 30222
rect 1810 30158 1822 30210
rect 1874 30158 1886 30210
rect 5630 30146 5682 30158
rect 6190 30210 6242 30222
rect 6190 30146 6242 30158
rect 6414 30210 6466 30222
rect 6414 30146 6466 30158
rect 7310 30210 7362 30222
rect 7310 30146 7362 30158
rect 8542 30210 8594 30222
rect 8542 30146 8594 30158
rect 9214 30210 9266 30222
rect 22990 30210 23042 30222
rect 20738 30158 20750 30210
rect 20802 30158 20814 30210
rect 9214 30146 9266 30158
rect 22990 30146 23042 30158
rect 25566 30210 25618 30222
rect 25566 30146 25618 30158
rect 26462 30210 26514 30222
rect 26462 30146 26514 30158
rect 26798 30210 26850 30222
rect 26798 30146 26850 30158
rect 27134 30210 27186 30222
rect 27134 30146 27186 30158
rect 27470 30210 27522 30222
rect 27470 30146 27522 30158
rect 30718 30210 30770 30222
rect 34750 30210 34802 30222
rect 31042 30158 31054 30210
rect 31106 30158 31118 30210
rect 34066 30158 34078 30210
rect 34130 30158 34142 30210
rect 30718 30146 30770 30158
rect 34750 30146 34802 30158
rect 36430 30210 36482 30222
rect 43486 30210 43538 30222
rect 36978 30158 36990 30210
rect 37042 30158 37054 30210
rect 47394 30158 47406 30210
rect 47458 30158 47470 30210
rect 48066 30158 48078 30210
rect 48130 30158 48142 30210
rect 36430 30146 36482 30158
rect 43486 30146 43538 30158
rect 5742 30098 5794 30110
rect 2482 30046 2494 30098
rect 2546 30046 2558 30098
rect 5742 30034 5794 30046
rect 5966 30098 6018 30110
rect 5966 30034 6018 30046
rect 6638 30098 6690 30110
rect 6638 30034 6690 30046
rect 6750 30098 6802 30110
rect 6750 30034 6802 30046
rect 6974 30098 7026 30110
rect 6974 30034 7026 30046
rect 7534 30098 7586 30110
rect 7534 30034 7586 30046
rect 7870 30098 7922 30110
rect 7870 30034 7922 30046
rect 8430 30098 8482 30110
rect 8430 30034 8482 30046
rect 14926 30098 14978 30110
rect 25902 30098 25954 30110
rect 18722 30046 18734 30098
rect 18786 30046 18798 30098
rect 14926 30034 14978 30046
rect 25902 30034 25954 30046
rect 26238 30098 26290 30110
rect 26238 30034 26290 30046
rect 27694 30098 27746 30110
rect 27694 30034 27746 30046
rect 30382 30098 30434 30110
rect 30382 30034 30434 30046
rect 31502 30098 31554 30110
rect 31502 30034 31554 30046
rect 31726 30098 31778 30110
rect 31726 30034 31778 30046
rect 33406 30098 33458 30110
rect 33406 30034 33458 30046
rect 33742 30098 33794 30110
rect 33742 30034 33794 30046
rect 35086 30098 35138 30110
rect 35410 30046 35422 30098
rect 35474 30046 35486 30098
rect 41794 30046 41806 30098
rect 41858 30046 41870 30098
rect 35086 30034 35138 30046
rect 7198 29986 7250 29998
rect 7198 29922 7250 29934
rect 7758 29986 7810 29998
rect 7758 29922 7810 29934
rect 8206 29986 8258 29998
rect 8206 29922 8258 29934
rect 11342 29986 11394 29998
rect 11342 29922 11394 29934
rect 12910 29986 12962 29998
rect 12910 29922 12962 29934
rect 13694 29986 13746 29998
rect 13694 29922 13746 29934
rect 13918 29986 13970 29998
rect 13918 29922 13970 29934
rect 14142 29986 14194 29998
rect 14142 29922 14194 29934
rect 14590 29986 14642 29998
rect 14590 29922 14642 29934
rect 21422 29986 21474 29998
rect 21422 29922 21474 29934
rect 24110 29986 24162 29998
rect 24110 29922 24162 29934
rect 24558 29986 24610 29998
rect 24558 29922 24610 29934
rect 25006 29986 25058 29998
rect 25006 29922 25058 29934
rect 25454 29986 25506 29998
rect 25454 29922 25506 29934
rect 26014 29986 26066 29998
rect 26014 29922 26066 29934
rect 27246 29986 27298 29998
rect 30830 29986 30882 29998
rect 28242 29934 28254 29986
rect 28306 29934 28318 29986
rect 27246 29922 27298 29934
rect 30830 29922 30882 29934
rect 32174 29986 32226 29998
rect 35870 29986 35922 29998
rect 33058 29934 33070 29986
rect 33122 29934 33134 29986
rect 34402 29934 34414 29986
rect 34466 29934 34478 29986
rect 32174 29922 32226 29934
rect 35870 29922 35922 29934
rect 1344 29818 48608 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 48608 29818
rect 1344 29732 48608 29766
rect 5070 29650 5122 29662
rect 5070 29586 5122 29598
rect 5966 29650 6018 29662
rect 5966 29586 6018 29598
rect 6190 29650 6242 29662
rect 6190 29586 6242 29598
rect 6974 29650 7026 29662
rect 6974 29586 7026 29598
rect 16830 29650 16882 29662
rect 18958 29650 19010 29662
rect 33630 29650 33682 29662
rect 17714 29598 17726 29650
rect 17778 29598 17790 29650
rect 32274 29598 32286 29650
rect 32338 29598 32350 29650
rect 16830 29586 16882 29598
rect 18958 29586 19010 29598
rect 33630 29586 33682 29598
rect 33854 29650 33906 29662
rect 33854 29586 33906 29598
rect 5630 29538 5682 29550
rect 5630 29474 5682 29486
rect 5742 29538 5794 29550
rect 5742 29474 5794 29486
rect 6302 29538 6354 29550
rect 6302 29474 6354 29486
rect 8990 29538 9042 29550
rect 33742 29538 33794 29550
rect 12786 29486 12798 29538
rect 12850 29486 12862 29538
rect 27346 29486 27358 29538
rect 27410 29486 27422 29538
rect 8990 29474 9042 29486
rect 33742 29474 33794 29486
rect 39790 29538 39842 29550
rect 39790 29474 39842 29486
rect 40350 29538 40402 29550
rect 40350 29474 40402 29486
rect 40910 29538 40962 29550
rect 40910 29474 40962 29486
rect 41246 29538 41298 29550
rect 41246 29474 41298 29486
rect 42702 29538 42754 29550
rect 42702 29474 42754 29486
rect 4846 29426 4898 29438
rect 1810 29374 1822 29426
rect 1874 29374 1886 29426
rect 4846 29362 4898 29374
rect 5182 29426 5234 29438
rect 7534 29426 7586 29438
rect 6738 29374 6750 29426
rect 6802 29374 6814 29426
rect 7298 29374 7310 29426
rect 7362 29374 7374 29426
rect 5182 29362 5234 29374
rect 7534 29362 7586 29374
rect 7758 29426 7810 29438
rect 7758 29362 7810 29374
rect 7982 29426 8034 29438
rect 7982 29362 8034 29374
rect 8318 29426 8370 29438
rect 8318 29362 8370 29374
rect 8654 29426 8706 29438
rect 13134 29426 13186 29438
rect 24222 29426 24274 29438
rect 42590 29426 42642 29438
rect 12450 29374 12462 29426
rect 12514 29374 12526 29426
rect 13570 29374 13582 29426
rect 13634 29374 13646 29426
rect 17714 29374 17726 29426
rect 17778 29374 17790 29426
rect 17938 29374 17950 29426
rect 18002 29374 18014 29426
rect 23202 29374 23214 29426
rect 23266 29374 23278 29426
rect 25330 29374 25342 29426
rect 25394 29374 25406 29426
rect 33394 29374 33406 29426
rect 33458 29374 33470 29426
rect 34066 29374 34078 29426
rect 34130 29374 34142 29426
rect 34514 29374 34526 29426
rect 34578 29374 34590 29426
rect 38770 29374 38782 29426
rect 38834 29374 38846 29426
rect 8654 29362 8706 29374
rect 13134 29362 13186 29374
rect 24222 29362 24274 29374
rect 42590 29362 42642 29374
rect 42926 29426 42978 29438
rect 42926 29362 42978 29374
rect 43262 29426 43314 29438
rect 43698 29374 43710 29426
rect 43762 29374 43774 29426
rect 45378 29374 45390 29426
rect 45442 29374 45454 29426
rect 43262 29362 43314 29374
rect 8542 29314 8594 29326
rect 19070 29314 19122 29326
rect 24446 29314 24498 29326
rect 2482 29262 2494 29314
rect 2546 29262 2558 29314
rect 4610 29262 4622 29314
rect 4674 29262 4686 29314
rect 9538 29262 9550 29314
rect 9602 29262 9614 29314
rect 11666 29262 11678 29314
rect 11730 29262 11742 29314
rect 14242 29262 14254 29314
rect 14306 29262 14318 29314
rect 16370 29262 16382 29314
rect 16434 29262 16446 29314
rect 17490 29262 17502 29314
rect 17554 29262 17566 29314
rect 20290 29262 20302 29314
rect 20354 29262 20366 29314
rect 22418 29262 22430 29314
rect 22482 29262 22494 29314
rect 8542 29250 8594 29262
rect 19070 29250 19122 29262
rect 24446 29250 24498 29262
rect 31726 29314 31778 29326
rect 37886 29314 37938 29326
rect 39230 29314 39282 29326
rect 35186 29262 35198 29314
rect 35250 29262 35262 29314
rect 37314 29262 37326 29314
rect 37378 29262 37390 29314
rect 38322 29262 38334 29314
rect 38386 29262 38398 29314
rect 31726 29250 31778 29262
rect 37886 29250 37938 29262
rect 39230 29250 39282 29262
rect 39566 29314 39618 29326
rect 40238 29314 40290 29326
rect 39890 29262 39902 29314
rect 39954 29262 39966 29314
rect 39566 29250 39618 29262
rect 40238 29250 40290 29262
rect 41694 29314 41746 29326
rect 41694 29250 41746 29262
rect 44158 29314 44210 29326
rect 46050 29262 46062 29314
rect 46114 29262 46126 29314
rect 48178 29262 48190 29314
rect 48242 29262 48254 29314
rect 44158 29250 44210 29262
rect 5630 29202 5682 29214
rect 5630 29138 5682 29150
rect 8094 29202 8146 29214
rect 31950 29202 32002 29214
rect 23874 29150 23886 29202
rect 23938 29150 23950 29202
rect 8094 29138 8146 29150
rect 31950 29138 32002 29150
rect 41582 29202 41634 29214
rect 41582 29138 41634 29150
rect 1344 29034 48608 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 48608 29034
rect 1344 28948 48608 28982
rect 33518 28866 33570 28878
rect 35198 28866 35250 28878
rect 45726 28866 45778 28878
rect 19058 28814 19070 28866
rect 19122 28863 19134 28866
rect 19282 28863 19294 28866
rect 19122 28817 19294 28863
rect 19122 28814 19134 28817
rect 19282 28814 19294 28817
rect 19346 28814 19358 28866
rect 33842 28814 33854 28866
rect 33906 28814 33918 28866
rect 43698 28814 43710 28866
rect 43762 28863 43774 28866
rect 44034 28863 44046 28866
rect 43762 28817 44046 28863
rect 43762 28814 43774 28817
rect 44034 28814 44046 28817
rect 44098 28814 44110 28866
rect 33518 28802 33570 28814
rect 35198 28802 35250 28814
rect 45726 28802 45778 28814
rect 46062 28866 46114 28878
rect 46062 28802 46114 28814
rect 3726 28754 3778 28766
rect 3726 28690 3778 28702
rect 11678 28754 11730 28766
rect 11678 28690 11730 28702
rect 12798 28754 12850 28766
rect 19182 28754 19234 28766
rect 20638 28754 20690 28766
rect 17378 28702 17390 28754
rect 17442 28702 17454 28754
rect 19618 28702 19630 28754
rect 19682 28702 19694 28754
rect 12798 28690 12850 28702
rect 19182 28690 19234 28702
rect 20638 28690 20690 28702
rect 21534 28754 21586 28766
rect 21534 28690 21586 28702
rect 22430 28754 22482 28766
rect 43710 28754 43762 28766
rect 23986 28702 23998 28754
rect 24050 28702 24062 28754
rect 26114 28702 26126 28754
rect 26178 28702 26190 28754
rect 27458 28702 27470 28754
rect 27522 28702 27534 28754
rect 35970 28702 35982 28754
rect 36034 28702 36046 28754
rect 22430 28690 22482 28702
rect 43710 28690 43762 28702
rect 44158 28754 44210 28766
rect 44158 28690 44210 28702
rect 47630 28754 47682 28766
rect 47630 28690 47682 28702
rect 3614 28642 3666 28654
rect 3614 28578 3666 28590
rect 4062 28642 4114 28654
rect 4062 28578 4114 28590
rect 4622 28642 4674 28654
rect 4622 28578 4674 28590
rect 4734 28642 4786 28654
rect 4734 28578 4786 28590
rect 5070 28642 5122 28654
rect 8654 28642 8706 28654
rect 6178 28590 6190 28642
rect 6242 28590 6254 28642
rect 7298 28590 7310 28642
rect 7362 28590 7374 28642
rect 5070 28578 5122 28590
rect 8654 28578 8706 28590
rect 11790 28642 11842 28654
rect 12350 28642 12402 28654
rect 12002 28590 12014 28642
rect 12066 28590 12078 28642
rect 11790 28578 11842 28590
rect 12350 28578 12402 28590
rect 12686 28642 12738 28654
rect 12686 28578 12738 28590
rect 13022 28642 13074 28654
rect 22094 28642 22146 28654
rect 14914 28590 14926 28642
rect 14978 28590 14990 28642
rect 19506 28590 19518 28642
rect 19570 28590 19582 28642
rect 20178 28590 20190 28642
rect 20242 28590 20254 28642
rect 13022 28578 13074 28590
rect 22094 28578 22146 28590
rect 22542 28642 22594 28654
rect 23202 28602 23214 28654
rect 23266 28602 23278 28654
rect 27582 28642 27634 28654
rect 27122 28590 27134 28642
rect 27186 28590 27198 28642
rect 22542 28578 22594 28590
rect 27582 28578 27634 28590
rect 28478 28642 28530 28654
rect 33294 28642 33346 28654
rect 29138 28590 29150 28642
rect 29202 28590 29214 28642
rect 31154 28590 31166 28642
rect 31218 28590 31230 28642
rect 28478 28578 28530 28590
rect 33294 28578 33346 28590
rect 34190 28642 34242 28654
rect 34190 28578 34242 28590
rect 34750 28642 34802 28654
rect 34750 28578 34802 28590
rect 35086 28642 35138 28654
rect 35086 28578 35138 28590
rect 36430 28642 36482 28654
rect 43374 28642 43426 28654
rect 41794 28590 41806 28642
rect 41858 28590 41870 28642
rect 36430 28578 36482 28590
rect 43374 28578 43426 28590
rect 44830 28642 44882 28654
rect 44830 28578 44882 28590
rect 45054 28642 45106 28654
rect 47406 28642 47458 28654
rect 46050 28590 46062 28642
rect 46114 28590 46126 28642
rect 45054 28578 45106 28590
rect 47406 28578 47458 28590
rect 48190 28642 48242 28654
rect 48190 28578 48242 28590
rect 3054 28530 3106 28542
rect 3054 28466 3106 28478
rect 3166 28530 3218 28542
rect 3166 28466 3218 28478
rect 3390 28530 3442 28542
rect 3390 28466 3442 28478
rect 3950 28530 4002 28542
rect 3950 28466 4002 28478
rect 4510 28530 4562 28542
rect 8318 28530 8370 28542
rect 5618 28478 5630 28530
rect 5682 28478 5694 28530
rect 7186 28478 7198 28530
rect 7250 28478 7262 28530
rect 7970 28478 7982 28530
rect 8034 28478 8046 28530
rect 4510 28466 4562 28478
rect 8318 28466 8370 28478
rect 8430 28530 8482 28542
rect 8430 28466 8482 28478
rect 9102 28530 9154 28542
rect 9102 28466 9154 28478
rect 19742 28530 19794 28542
rect 19742 28466 19794 28478
rect 19966 28530 20018 28542
rect 19966 28466 20018 28478
rect 21422 28530 21474 28542
rect 21422 28466 21474 28478
rect 21646 28530 21698 28542
rect 21646 28466 21698 28478
rect 22318 28530 22370 28542
rect 22318 28466 22370 28478
rect 22878 28530 22930 28542
rect 22878 28466 22930 28478
rect 28590 28530 28642 28542
rect 32286 28530 32338 28542
rect 42814 28530 42866 28542
rect 29250 28478 29262 28530
rect 29314 28478 29326 28530
rect 38658 28478 38670 28530
rect 38722 28478 38734 28530
rect 28590 28466 28642 28478
rect 32286 28466 32338 28478
rect 42814 28466 42866 28478
rect 7646 28418 7698 28430
rect 6626 28366 6638 28418
rect 6690 28366 6702 28418
rect 7646 28354 7698 28366
rect 8766 28418 8818 28430
rect 8766 28354 8818 28366
rect 8990 28418 9042 28430
rect 8990 28354 9042 28366
rect 10782 28418 10834 28430
rect 10782 28354 10834 28366
rect 27918 28418 27970 28430
rect 43038 28418 43090 28430
rect 30594 28366 30606 28418
rect 30658 28366 30670 28418
rect 27918 28354 27970 28366
rect 43038 28354 43090 28366
rect 43262 28418 43314 28430
rect 45378 28366 45390 28418
rect 45442 28366 45454 28418
rect 43262 28354 43314 28366
rect 1344 28250 48608 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 48608 28250
rect 1344 28164 48608 28198
rect 9662 28082 9714 28094
rect 9662 28018 9714 28030
rect 10558 28082 10610 28094
rect 10558 28018 10610 28030
rect 15822 28082 15874 28094
rect 15822 28018 15874 28030
rect 18846 28082 18898 28094
rect 18846 28018 18898 28030
rect 22878 28082 22930 28094
rect 22878 28018 22930 28030
rect 23438 28082 23490 28094
rect 23438 28018 23490 28030
rect 26238 28082 26290 28094
rect 26238 28018 26290 28030
rect 26574 28082 26626 28094
rect 29374 28082 29426 28094
rect 28018 28030 28030 28082
rect 28082 28030 28094 28082
rect 26574 28018 26626 28030
rect 29374 28018 29426 28030
rect 30046 28082 30098 28094
rect 30046 28018 30098 28030
rect 31278 28082 31330 28094
rect 31278 28018 31330 28030
rect 40350 28082 40402 28094
rect 40350 28018 40402 28030
rect 41246 28082 41298 28094
rect 41246 28018 41298 28030
rect 41470 28082 41522 28094
rect 41470 28018 41522 28030
rect 41582 28082 41634 28094
rect 41582 28018 41634 28030
rect 42142 28082 42194 28094
rect 42466 28030 42478 28082
rect 42530 28030 42542 28082
rect 42142 28018 42194 28030
rect 14814 27970 14866 27982
rect 11666 27918 11678 27970
rect 11730 27918 11742 27970
rect 14814 27906 14866 27918
rect 14926 27970 14978 27982
rect 14926 27906 14978 27918
rect 26686 27970 26738 27982
rect 26686 27906 26738 27918
rect 29486 27970 29538 27982
rect 29486 27906 29538 27918
rect 29822 27970 29874 27982
rect 29822 27906 29874 27918
rect 40238 27970 40290 27982
rect 40238 27906 40290 27918
rect 19070 27858 19122 27870
rect 8642 27806 8654 27858
rect 8706 27806 8718 27858
rect 10322 27806 10334 27858
rect 10386 27806 10398 27858
rect 10994 27806 11006 27858
rect 11058 27806 11070 27858
rect 14578 27806 14590 27858
rect 14642 27806 14654 27858
rect 15698 27806 15710 27858
rect 15762 27806 15774 27858
rect 18610 27806 18622 27858
rect 18674 27806 18686 27858
rect 19070 27794 19122 27806
rect 19182 27858 19234 27870
rect 21758 27858 21810 27870
rect 20066 27806 20078 27858
rect 20130 27806 20142 27858
rect 20290 27806 20302 27858
rect 20354 27806 20366 27858
rect 21074 27806 21086 27858
rect 21138 27806 21150 27858
rect 19182 27794 19234 27806
rect 21758 27794 21810 27806
rect 22654 27858 22706 27870
rect 22654 27794 22706 27806
rect 22990 27858 23042 27870
rect 22990 27794 23042 27806
rect 27582 27858 27634 27870
rect 31726 27858 31778 27870
rect 27794 27806 27806 27858
rect 27858 27806 27870 27858
rect 29138 27806 29150 27858
rect 29202 27806 29214 27858
rect 30706 27806 30718 27858
rect 30770 27806 30782 27858
rect 31154 27806 31166 27858
rect 31218 27806 31230 27858
rect 27582 27794 27634 27806
rect 31726 27794 31778 27806
rect 31950 27858 32002 27870
rect 41134 27858 41186 27870
rect 33730 27806 33742 27858
rect 33794 27806 33806 27858
rect 36978 27806 36990 27858
rect 37042 27806 37054 27858
rect 43586 27806 43598 27858
rect 43650 27806 43662 27858
rect 31950 27794 32002 27806
rect 41134 27794 41186 27806
rect 16158 27746 16210 27758
rect 6066 27694 6078 27746
rect 6130 27694 6142 27746
rect 13794 27694 13806 27746
rect 13858 27694 13870 27746
rect 16158 27682 16210 27694
rect 16830 27746 16882 27758
rect 16830 27682 16882 27694
rect 17502 27746 17554 27758
rect 17502 27682 17554 27694
rect 18958 27746 19010 27758
rect 22430 27746 22482 27758
rect 20626 27694 20638 27746
rect 20690 27694 20702 27746
rect 18958 27682 19010 27694
rect 22430 27682 22482 27694
rect 24334 27746 24386 27758
rect 24334 27682 24386 27694
rect 25342 27746 25394 27758
rect 33182 27746 33234 27758
rect 27682 27694 27694 27746
rect 27746 27694 27758 27746
rect 30146 27694 30158 27746
rect 30210 27694 30222 27746
rect 25342 27682 25394 27694
rect 33182 27682 33234 27694
rect 33294 27746 33346 27758
rect 34402 27694 34414 27746
rect 34466 27694 34478 27746
rect 36530 27694 36542 27746
rect 36594 27694 36606 27746
rect 37650 27694 37662 27746
rect 37714 27694 37726 27746
rect 39778 27694 39790 27746
rect 39842 27694 39854 27746
rect 41570 27694 41582 27746
rect 41634 27694 41646 27746
rect 45378 27694 45390 27746
rect 45442 27694 45454 27746
rect 33294 27682 33346 27694
rect 15934 27634 15986 27646
rect 15362 27582 15374 27634
rect 15426 27582 15438 27634
rect 15934 27570 15986 27582
rect 17390 27634 17442 27646
rect 21870 27634 21922 27646
rect 20738 27582 20750 27634
rect 20802 27582 20814 27634
rect 17390 27570 17442 27582
rect 21870 27570 21922 27582
rect 25230 27634 25282 27646
rect 32274 27582 32286 27634
rect 32338 27582 32350 27634
rect 25230 27570 25282 27582
rect 1344 27466 48608 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 48608 27466
rect 1344 27380 48608 27414
rect 30158 27298 30210 27310
rect 30158 27234 30210 27246
rect 37438 27298 37490 27310
rect 37438 27234 37490 27246
rect 37774 27298 37826 27310
rect 37774 27234 37826 27246
rect 14366 27186 14418 27198
rect 19630 27186 19682 27198
rect 2482 27134 2494 27186
rect 2546 27134 2558 27186
rect 4610 27134 4622 27186
rect 4674 27134 4686 27186
rect 8978 27134 8990 27186
rect 9042 27134 9054 27186
rect 9314 27134 9326 27186
rect 9378 27134 9390 27186
rect 16706 27134 16718 27186
rect 16770 27134 16782 27186
rect 18834 27134 18846 27186
rect 18898 27134 18910 27186
rect 14366 27122 14418 27134
rect 19630 27122 19682 27134
rect 20414 27186 20466 27198
rect 27358 27186 27410 27198
rect 21298 27134 21310 27186
rect 21362 27134 21374 27186
rect 25666 27134 25678 27186
rect 25730 27134 25742 27186
rect 20414 27122 20466 27134
rect 27358 27122 27410 27134
rect 30382 27186 30434 27198
rect 30382 27122 30434 27134
rect 31502 27186 31554 27198
rect 31502 27122 31554 27134
rect 32286 27186 32338 27198
rect 34974 27186 35026 27198
rect 32722 27134 32734 27186
rect 32786 27134 32798 27186
rect 33954 27134 33966 27186
rect 34018 27134 34030 27186
rect 32286 27122 32338 27134
rect 34974 27122 35026 27134
rect 35422 27186 35474 27198
rect 35422 27122 35474 27134
rect 38446 27186 38498 27198
rect 38446 27122 38498 27134
rect 40686 27186 40738 27198
rect 42466 27134 42478 27186
rect 42530 27134 42542 27186
rect 48066 27134 48078 27186
rect 48130 27134 48142 27186
rect 40686 27122 40738 27134
rect 14814 27074 14866 27086
rect 26014 27074 26066 27086
rect 32846 27074 32898 27086
rect 1810 27022 1822 27074
rect 1874 27022 1886 27074
rect 6066 27022 6078 27074
rect 6130 27022 6142 27074
rect 12226 27022 12238 27074
rect 12290 27022 12302 27074
rect 16034 27022 16046 27074
rect 16098 27022 16110 27074
rect 24210 27022 24222 27074
rect 24274 27022 24286 27074
rect 32610 27022 32622 27074
rect 32674 27022 32686 27074
rect 14814 27010 14866 27022
rect 26014 27010 26066 27022
rect 32846 27010 32898 27022
rect 33182 27074 33234 27086
rect 34078 27074 34130 27086
rect 33842 27022 33854 27074
rect 33906 27022 33918 27074
rect 33182 27010 33234 27022
rect 34078 27010 34130 27022
rect 34302 27074 34354 27086
rect 37550 27074 37602 27086
rect 39230 27074 39282 27086
rect 34514 27022 34526 27074
rect 34578 27022 34590 27074
rect 37986 27022 37998 27074
rect 38050 27022 38062 27074
rect 38658 27022 38670 27074
rect 38722 27022 38734 27074
rect 34302 27010 34354 27022
rect 37550 27010 37602 27022
rect 39230 27010 39282 27022
rect 39342 27074 39394 27086
rect 39342 27010 39394 27022
rect 39566 27074 39618 27086
rect 39566 27010 39618 27022
rect 40350 27074 40402 27086
rect 40350 27010 40402 27022
rect 41358 27074 41410 27086
rect 41358 27010 41410 27022
rect 42254 27074 42306 27086
rect 43150 27074 43202 27086
rect 42690 27022 42702 27074
rect 42754 27022 42766 27074
rect 42254 27010 42306 27022
rect 43150 27010 43202 27022
rect 43598 27074 43650 27086
rect 43598 27010 43650 27022
rect 43934 27074 43986 27086
rect 45266 27022 45278 27074
rect 45330 27022 45342 27074
rect 43934 27010 43986 27022
rect 14254 26962 14306 26974
rect 6850 26910 6862 26962
rect 6914 26910 6926 26962
rect 11442 26910 11454 26962
rect 11506 26910 11518 26962
rect 14254 26898 14306 26910
rect 14590 26962 14642 26974
rect 14590 26898 14642 26910
rect 19854 26962 19906 26974
rect 24894 26962 24946 26974
rect 23426 26910 23438 26962
rect 23490 26910 23502 26962
rect 24546 26910 24558 26962
rect 24610 26910 24622 26962
rect 19854 26898 19906 26910
rect 24894 26898 24946 26910
rect 25678 26962 25730 26974
rect 25678 26898 25730 26910
rect 26238 26962 26290 26974
rect 38334 26962 38386 26974
rect 26562 26910 26574 26962
rect 26626 26910 26638 26962
rect 29810 26910 29822 26962
rect 29874 26910 29886 26962
rect 26238 26898 26290 26910
rect 38334 26898 38386 26910
rect 40126 26962 40178 26974
rect 42030 26962 42082 26974
rect 41010 26910 41022 26962
rect 41074 26910 41086 26962
rect 40126 26898 40178 26910
rect 42030 26898 42082 26910
rect 42926 26962 42978 26974
rect 43810 26910 43822 26962
rect 43874 26910 43886 26962
rect 45938 26910 45950 26962
rect 46002 26910 46014 26962
rect 42926 26898 42978 26910
rect 19966 26850 20018 26862
rect 19966 26786 20018 26798
rect 25790 26850 25842 26862
rect 25790 26786 25842 26798
rect 26910 26850 26962 26862
rect 26910 26786 26962 26798
rect 31390 26850 31442 26862
rect 31390 26786 31442 26798
rect 33070 26850 33122 26862
rect 33070 26786 33122 26798
rect 39454 26850 39506 26862
rect 39454 26786 39506 26798
rect 39678 26850 39730 26862
rect 39678 26786 39730 26798
rect 42478 26850 42530 26862
rect 42478 26786 42530 26798
rect 1344 26682 48608 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 48608 26682
rect 1344 26596 48608 26630
rect 6302 26514 6354 26526
rect 5954 26462 5966 26514
rect 6018 26462 6030 26514
rect 6302 26450 6354 26462
rect 7758 26514 7810 26526
rect 7758 26450 7810 26462
rect 7870 26514 7922 26526
rect 7870 26450 7922 26462
rect 8430 26514 8482 26526
rect 8430 26450 8482 26462
rect 10558 26514 10610 26526
rect 10558 26450 10610 26462
rect 16270 26514 16322 26526
rect 16270 26450 16322 26462
rect 16606 26514 16658 26526
rect 16606 26450 16658 26462
rect 18062 26514 18114 26526
rect 18062 26450 18114 26462
rect 25790 26514 25842 26526
rect 33854 26514 33906 26526
rect 29586 26462 29598 26514
rect 29650 26462 29662 26514
rect 25790 26450 25842 26462
rect 33854 26450 33906 26462
rect 34638 26514 34690 26526
rect 34638 26450 34690 26462
rect 37550 26514 37602 26526
rect 37550 26450 37602 26462
rect 38446 26514 38498 26526
rect 38446 26450 38498 26462
rect 39790 26514 39842 26526
rect 39790 26450 39842 26462
rect 43934 26514 43986 26526
rect 43934 26450 43986 26462
rect 44382 26514 44434 26526
rect 44382 26450 44434 26462
rect 44942 26514 44994 26526
rect 44942 26450 44994 26462
rect 8318 26402 8370 26414
rect 8318 26338 8370 26350
rect 8542 26402 8594 26414
rect 8542 26338 8594 26350
rect 9886 26402 9938 26414
rect 9886 26338 9938 26350
rect 10110 26402 10162 26414
rect 16382 26402 16434 26414
rect 13682 26350 13694 26402
rect 13746 26350 13758 26402
rect 10110 26338 10162 26350
rect 16382 26338 16434 26350
rect 17614 26402 17666 26414
rect 40910 26402 40962 26414
rect 42030 26402 42082 26414
rect 21410 26350 21422 26402
rect 21474 26350 21486 26402
rect 22306 26350 22318 26402
rect 22370 26350 22382 26402
rect 24546 26350 24558 26402
rect 24610 26350 24622 26402
rect 27346 26350 27358 26402
rect 27410 26350 27422 26402
rect 39218 26350 39230 26402
rect 39282 26350 39294 26402
rect 41794 26350 41806 26402
rect 41858 26350 41870 26402
rect 17614 26338 17666 26350
rect 40910 26338 40962 26350
rect 42030 26338 42082 26350
rect 42814 26402 42866 26414
rect 42814 26338 42866 26350
rect 43038 26402 43090 26414
rect 43038 26338 43090 26350
rect 43486 26402 43538 26414
rect 43486 26338 43538 26350
rect 44046 26402 44098 26414
rect 44046 26338 44098 26350
rect 44494 26402 44546 26414
rect 44494 26338 44546 26350
rect 47630 26402 47682 26414
rect 47630 26338 47682 26350
rect 48078 26402 48130 26414
rect 48078 26338 48130 26350
rect 4846 26290 4898 26302
rect 4610 26238 4622 26290
rect 4674 26238 4686 26290
rect 4846 26226 4898 26238
rect 5182 26290 5234 26302
rect 5182 26226 5234 26238
rect 5406 26290 5458 26302
rect 5406 26226 5458 26238
rect 7086 26290 7138 26302
rect 7086 26226 7138 26238
rect 7310 26290 7362 26302
rect 7310 26226 7362 26238
rect 7982 26290 8034 26302
rect 7982 26226 8034 26238
rect 9774 26290 9826 26302
rect 9774 26226 9826 26238
rect 10222 26290 10274 26302
rect 10222 26226 10274 26238
rect 10670 26290 10722 26302
rect 10670 26226 10722 26238
rect 10782 26290 10834 26302
rect 25230 26290 25282 26302
rect 12898 26238 12910 26290
rect 12962 26238 12974 26290
rect 16818 26238 16830 26290
rect 16882 26238 16894 26290
rect 18610 26238 18622 26290
rect 18674 26238 18686 26290
rect 19058 26238 19070 26290
rect 19122 26238 19134 26290
rect 19618 26238 19630 26290
rect 19682 26238 19694 26290
rect 20626 26238 20638 26290
rect 20690 26238 20702 26290
rect 22194 26238 22206 26290
rect 22258 26238 22270 26290
rect 23986 26238 23998 26290
rect 24050 26238 24062 26290
rect 10782 26226 10834 26238
rect 25230 26226 25282 26238
rect 25678 26290 25730 26302
rect 25678 26226 25730 26238
rect 25902 26290 25954 26302
rect 33630 26290 33682 26302
rect 38334 26290 38386 26302
rect 26674 26238 26686 26290
rect 26738 26238 26750 26290
rect 33394 26238 33406 26290
rect 33458 26238 33470 26290
rect 34066 26238 34078 26290
rect 34130 26238 34142 26290
rect 25902 26226 25954 26238
rect 33630 26226 33682 26238
rect 38334 26226 38386 26238
rect 38782 26290 38834 26302
rect 38782 26226 38834 26238
rect 39006 26290 39058 26302
rect 41022 26290 41074 26302
rect 42142 26290 42194 26302
rect 39330 26238 39342 26290
rect 39394 26238 39406 26290
rect 41682 26238 41694 26290
rect 41746 26238 41758 26290
rect 39006 26226 39058 26238
rect 41022 26226 41074 26238
rect 42142 26226 42194 26238
rect 42590 26290 42642 26302
rect 42590 26226 42642 26238
rect 43598 26290 43650 26302
rect 45054 26290 45106 26302
rect 44818 26238 44830 26290
rect 44882 26238 44894 26290
rect 43598 26226 43650 26238
rect 45054 26226 45106 26238
rect 46510 26290 46562 26302
rect 46510 26226 46562 26238
rect 46622 26290 46674 26302
rect 47182 26290 47234 26302
rect 46946 26238 46958 26290
rect 47010 26238 47022 26290
rect 46622 26226 46674 26238
rect 47182 26226 47234 26238
rect 47406 26290 47458 26302
rect 47406 26226 47458 26238
rect 5070 26178 5122 26190
rect 16494 26178 16546 26190
rect 25454 26178 25506 26190
rect 37886 26178 37938 26190
rect 1698 26126 1710 26178
rect 1762 26126 1774 26178
rect 3826 26126 3838 26178
rect 3890 26126 3902 26178
rect 15810 26126 15822 26178
rect 15874 26126 15886 26178
rect 19394 26126 19406 26178
rect 19458 26126 19470 26178
rect 33506 26126 33518 26178
rect 33570 26126 33582 26178
rect 5070 26114 5122 26126
rect 16494 26114 16546 26126
rect 25454 26114 25506 26126
rect 37886 26114 37938 26126
rect 42702 26178 42754 26190
rect 47966 26178 48018 26190
rect 47058 26126 47070 26178
rect 47122 26126 47134 26178
rect 42702 26114 42754 26126
rect 47966 26114 48018 26126
rect 37998 26066 38050 26078
rect 19506 26014 19518 26066
rect 19570 26014 19582 26066
rect 37998 26002 38050 26014
rect 41246 26066 41298 26078
rect 41246 26002 41298 26014
rect 45278 26066 45330 26078
rect 45278 26002 45330 26014
rect 1344 25898 48608 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 48608 25898
rect 1344 25812 48608 25846
rect 3502 25730 3554 25742
rect 3502 25666 3554 25678
rect 28030 25730 28082 25742
rect 28030 25666 28082 25678
rect 38782 25730 38834 25742
rect 38782 25666 38834 25678
rect 7310 25618 7362 25630
rect 7310 25554 7362 25566
rect 16382 25618 16434 25630
rect 20638 25618 20690 25630
rect 33294 25618 33346 25630
rect 20290 25566 20302 25618
rect 20354 25566 20366 25618
rect 30818 25566 30830 25618
rect 30882 25566 30894 25618
rect 32946 25566 32958 25618
rect 33010 25566 33022 25618
rect 16382 25554 16434 25566
rect 20638 25554 20690 25566
rect 33294 25554 33346 25566
rect 33742 25618 33794 25630
rect 39106 25566 39118 25618
rect 39170 25566 39182 25618
rect 48178 25566 48190 25618
rect 48242 25566 48254 25618
rect 33742 25554 33794 25566
rect 3054 25506 3106 25518
rect 3054 25442 3106 25454
rect 3950 25506 4002 25518
rect 3950 25442 4002 25454
rect 4286 25506 4338 25518
rect 4286 25442 4338 25454
rect 4398 25506 4450 25518
rect 4398 25442 4450 25454
rect 4734 25506 4786 25518
rect 10670 25506 10722 25518
rect 36430 25506 36482 25518
rect 37214 25506 37266 25518
rect 7074 25454 7086 25506
rect 7138 25454 7150 25506
rect 13458 25454 13470 25506
rect 13522 25454 13534 25506
rect 17490 25454 17502 25506
rect 17554 25454 17566 25506
rect 25106 25454 25118 25506
rect 25170 25454 25182 25506
rect 27234 25454 27246 25506
rect 27298 25454 27310 25506
rect 30146 25454 30158 25506
rect 30210 25454 30222 25506
rect 36978 25454 36990 25506
rect 37042 25454 37054 25506
rect 4734 25442 4786 25454
rect 10670 25442 10722 25454
rect 36430 25442 36482 25454
rect 37214 25442 37266 25454
rect 37326 25506 37378 25518
rect 37326 25442 37378 25454
rect 39790 25506 39842 25518
rect 39790 25442 39842 25454
rect 40238 25506 40290 25518
rect 40238 25442 40290 25454
rect 40686 25506 40738 25518
rect 40686 25442 40738 25454
rect 41022 25506 41074 25518
rect 41022 25442 41074 25454
rect 41358 25506 41410 25518
rect 41358 25442 41410 25454
rect 42030 25506 42082 25518
rect 42030 25442 42082 25454
rect 43150 25506 43202 25518
rect 44046 25506 44098 25518
rect 43586 25454 43598 25506
rect 43650 25454 43662 25506
rect 45378 25454 45390 25506
rect 45442 25454 45454 25506
rect 43150 25442 43202 25454
rect 44046 25442 44098 25454
rect 3614 25394 3666 25406
rect 3614 25330 3666 25342
rect 4622 25394 4674 25406
rect 6750 25394 6802 25406
rect 5618 25342 5630 25394
rect 5682 25342 5694 25394
rect 4622 25330 4674 25342
rect 6750 25330 6802 25342
rect 7422 25394 7474 25406
rect 7422 25330 7474 25342
rect 8430 25394 8482 25406
rect 8430 25330 8482 25342
rect 8654 25394 8706 25406
rect 8654 25330 8706 25342
rect 8878 25394 8930 25406
rect 8878 25330 8930 25342
rect 8990 25394 9042 25406
rect 8990 25330 9042 25342
rect 9774 25394 9826 25406
rect 9774 25330 9826 25342
rect 10334 25394 10386 25406
rect 10334 25330 10386 25342
rect 10446 25394 10498 25406
rect 10446 25330 10498 25342
rect 11118 25394 11170 25406
rect 27806 25394 27858 25406
rect 14242 25342 14254 25394
rect 14306 25342 14318 25394
rect 18162 25342 18174 25394
rect 18226 25342 18238 25394
rect 21970 25342 21982 25394
rect 22034 25342 22046 25394
rect 27010 25342 27022 25394
rect 27074 25342 27086 25394
rect 11118 25330 11170 25342
rect 27806 25330 27858 25342
rect 28478 25394 28530 25406
rect 28478 25330 28530 25342
rect 38110 25394 38162 25406
rect 38110 25330 38162 25342
rect 38446 25394 38498 25406
rect 38446 25330 38498 25342
rect 39006 25394 39058 25406
rect 39006 25330 39058 25342
rect 39678 25394 39730 25406
rect 39678 25330 39730 25342
rect 42366 25394 42418 25406
rect 42366 25330 42418 25342
rect 42590 25394 42642 25406
rect 42590 25330 42642 25342
rect 44270 25394 44322 25406
rect 44270 25330 44322 25342
rect 44830 25394 44882 25406
rect 44830 25330 44882 25342
rect 44942 25394 44994 25406
rect 46050 25342 46062 25394
rect 46114 25342 46126 25394
rect 44942 25330 44994 25342
rect 2718 25282 2770 25294
rect 2718 25218 2770 25230
rect 2942 25282 2994 25294
rect 2942 25218 2994 25230
rect 3502 25282 3554 25294
rect 3502 25218 3554 25230
rect 4062 25282 4114 25294
rect 4062 25218 4114 25230
rect 5966 25282 6018 25294
rect 5966 25218 6018 25230
rect 6414 25282 6466 25294
rect 6414 25218 6466 25230
rect 7758 25282 7810 25294
rect 9886 25282 9938 25294
rect 8082 25230 8094 25282
rect 8146 25230 8158 25282
rect 7758 25218 7810 25230
rect 9886 25218 9938 25230
rect 10110 25282 10162 25294
rect 10110 25218 10162 25230
rect 11230 25282 11282 25294
rect 11230 25218 11282 25230
rect 11454 25282 11506 25294
rect 11454 25218 11506 25230
rect 20750 25282 20802 25294
rect 20750 25218 20802 25230
rect 27918 25282 27970 25294
rect 27918 25218 27970 25230
rect 29710 25282 29762 25294
rect 29710 25218 29762 25230
rect 33406 25282 33458 25294
rect 33406 25218 33458 25230
rect 33854 25282 33906 25294
rect 39566 25282 39618 25294
rect 37762 25230 37774 25282
rect 37826 25230 37838 25282
rect 33854 25218 33906 25230
rect 39566 25218 39618 25230
rect 41022 25282 41074 25294
rect 41022 25218 41074 25230
rect 42254 25282 42306 25294
rect 42254 25218 42306 25230
rect 42814 25282 42866 25294
rect 42814 25218 42866 25230
rect 43038 25282 43090 25294
rect 43038 25218 43090 25230
rect 43822 25282 43874 25294
rect 43822 25218 43874 25230
rect 43934 25282 43986 25294
rect 43934 25218 43986 25230
rect 1344 25114 48608 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 48608 25114
rect 1344 25028 48608 25062
rect 5966 24946 6018 24958
rect 5966 24882 6018 24894
rect 8206 24946 8258 24958
rect 8206 24882 8258 24894
rect 10222 24946 10274 24958
rect 10222 24882 10274 24894
rect 11790 24946 11842 24958
rect 11790 24882 11842 24894
rect 16382 24946 16434 24958
rect 16382 24882 16434 24894
rect 24446 24946 24498 24958
rect 24446 24882 24498 24894
rect 32510 24946 32562 24958
rect 32510 24882 32562 24894
rect 39790 24946 39842 24958
rect 39790 24882 39842 24894
rect 42590 24946 42642 24958
rect 42590 24882 42642 24894
rect 44046 24946 44098 24958
rect 44046 24882 44098 24894
rect 45950 24946 46002 24958
rect 45950 24882 46002 24894
rect 9886 24834 9938 24846
rect 9886 24770 9938 24782
rect 9998 24834 10050 24846
rect 9998 24770 10050 24782
rect 11342 24834 11394 24846
rect 11342 24770 11394 24782
rect 11566 24834 11618 24846
rect 11566 24770 11618 24782
rect 12238 24834 12290 24846
rect 12238 24770 12290 24782
rect 12350 24834 12402 24846
rect 12350 24770 12402 24782
rect 16718 24834 16770 24846
rect 16718 24770 16770 24782
rect 24334 24834 24386 24846
rect 39902 24834 39954 24846
rect 28578 24782 28590 24834
rect 28642 24782 28654 24834
rect 33842 24782 33854 24834
rect 33906 24782 33918 24834
rect 24334 24770 24386 24782
rect 39902 24770 39954 24782
rect 42478 24834 42530 24846
rect 42478 24770 42530 24782
rect 43150 24834 43202 24846
rect 43150 24770 43202 24782
rect 46062 24834 46114 24846
rect 46062 24770 46114 24782
rect 4846 24722 4898 24734
rect 1810 24670 1822 24722
rect 1874 24670 1886 24722
rect 4846 24658 4898 24670
rect 5182 24722 5234 24734
rect 5182 24658 5234 24670
rect 5406 24722 5458 24734
rect 5406 24658 5458 24670
rect 6302 24722 6354 24734
rect 6302 24658 6354 24670
rect 8318 24722 8370 24734
rect 8318 24658 8370 24670
rect 8542 24722 8594 24734
rect 10334 24722 10386 24734
rect 8754 24670 8766 24722
rect 8818 24670 8830 24722
rect 8542 24658 8594 24670
rect 10334 24658 10386 24670
rect 10670 24722 10722 24734
rect 10670 24658 10722 24670
rect 10894 24722 10946 24734
rect 10894 24658 10946 24670
rect 12014 24722 12066 24734
rect 25342 24722 25394 24734
rect 31278 24722 31330 24734
rect 20178 24670 20190 24722
rect 20242 24670 20254 24722
rect 23538 24670 23550 24722
rect 23602 24670 23614 24722
rect 25778 24670 25790 24722
rect 25842 24670 25854 24722
rect 12014 24658 12066 24670
rect 25342 24658 25394 24670
rect 31278 24658 31330 24670
rect 31502 24722 31554 24734
rect 39454 24722 39506 24734
rect 33058 24670 33070 24722
rect 33122 24670 33134 24722
rect 36306 24670 36318 24722
rect 36370 24670 36382 24722
rect 31502 24658 31554 24670
rect 39454 24658 39506 24670
rect 40014 24722 40066 24734
rect 44818 24670 44830 24722
rect 44882 24670 44894 24722
rect 40014 24658 40066 24670
rect 5070 24610 5122 24622
rect 2482 24558 2494 24610
rect 2546 24558 2558 24610
rect 4610 24558 4622 24610
rect 4674 24558 4686 24610
rect 5070 24546 5122 24558
rect 6750 24610 6802 24622
rect 6750 24546 6802 24558
rect 10558 24610 10610 24622
rect 10558 24546 10610 24558
rect 16830 24610 16882 24622
rect 44158 24610 44210 24622
rect 45502 24610 45554 24622
rect 17378 24558 17390 24610
rect 17442 24558 17454 24610
rect 19506 24558 19518 24610
rect 19570 24558 19582 24610
rect 20738 24558 20750 24610
rect 20802 24558 20814 24610
rect 22866 24558 22878 24610
rect 22930 24558 22942 24610
rect 35970 24558 35982 24610
rect 36034 24558 36046 24610
rect 37090 24558 37102 24610
rect 37154 24558 37166 24610
rect 39218 24558 39230 24610
rect 39282 24558 39294 24610
rect 45042 24558 45054 24610
rect 45106 24558 45118 24610
rect 16830 24546 16882 24558
rect 44158 24546 44210 24558
rect 45502 24546 45554 24558
rect 45838 24610 45890 24622
rect 45838 24546 45890 24558
rect 8094 24498 8146 24510
rect 8094 24434 8146 24446
rect 12350 24498 12402 24510
rect 12350 24434 12402 24446
rect 24446 24498 24498 24510
rect 43038 24498 43090 24510
rect 31826 24446 31838 24498
rect 31890 24446 31902 24498
rect 24446 24434 24498 24446
rect 43038 24434 43090 24446
rect 1344 24330 48608 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 48608 24330
rect 1344 24244 48608 24278
rect 21310 24162 21362 24174
rect 21310 24098 21362 24110
rect 30494 24162 30546 24174
rect 30494 24098 30546 24110
rect 21534 24050 21586 24062
rect 30270 24050 30322 24062
rect 38334 24050 38386 24062
rect 9986 23998 9998 24050
rect 10050 23998 10062 24050
rect 12114 23998 12126 24050
rect 12178 23998 12190 24050
rect 16370 23998 16382 24050
rect 16434 23998 16446 24050
rect 19730 23998 19742 24050
rect 19794 23998 19806 24050
rect 24546 23998 24558 24050
rect 24610 23998 24622 24050
rect 26674 23998 26686 24050
rect 26738 23998 26750 24050
rect 37986 23998 37998 24050
rect 38050 23998 38062 24050
rect 42578 23998 42590 24050
rect 42642 23998 42654 24050
rect 45266 23998 45278 24050
rect 45330 23998 45342 24050
rect 21534 23986 21586 23998
rect 30270 23986 30322 23998
rect 38334 23986 38386 23998
rect 4510 23938 4562 23950
rect 4510 23874 4562 23886
rect 5966 23938 6018 23950
rect 5966 23874 6018 23886
rect 8206 23938 8258 23950
rect 8206 23874 8258 23886
rect 8654 23938 8706 23950
rect 21870 23938 21922 23950
rect 8978 23886 8990 23938
rect 9042 23886 9054 23938
rect 12786 23886 12798 23938
rect 12850 23886 12862 23938
rect 13570 23886 13582 23938
rect 13634 23886 13646 23938
rect 16818 23886 16830 23938
rect 16882 23886 16894 23938
rect 20738 23886 20750 23938
rect 20802 23886 20814 23938
rect 8654 23874 8706 23886
rect 21870 23874 21922 23886
rect 21982 23938 22034 23950
rect 21982 23874 22034 23886
rect 22542 23938 22594 23950
rect 22542 23874 22594 23886
rect 22766 23938 22818 23950
rect 22766 23874 22818 23886
rect 22990 23938 23042 23950
rect 27246 23938 27298 23950
rect 28142 23938 28194 23950
rect 29374 23938 29426 23950
rect 23874 23886 23886 23938
rect 23938 23886 23950 23938
rect 27682 23886 27694 23938
rect 27746 23886 27758 23938
rect 29138 23886 29150 23938
rect 29202 23886 29214 23938
rect 22990 23874 23042 23886
rect 27246 23874 27298 23886
rect 28142 23874 28194 23886
rect 29374 23874 29426 23886
rect 29598 23938 29650 23950
rect 39342 23938 39394 23950
rect 29810 23886 29822 23938
rect 29874 23886 29886 23938
rect 36418 23886 36430 23938
rect 36482 23886 36494 23938
rect 37874 23886 37886 23938
rect 37938 23886 37950 23938
rect 29598 23874 29650 23886
rect 39342 23874 39394 23886
rect 40014 23938 40066 23950
rect 40014 23874 40066 23886
rect 41246 23938 41298 23950
rect 41246 23874 41298 23886
rect 41806 23938 41858 23950
rect 41806 23874 41858 23886
rect 42030 23938 42082 23950
rect 43598 23938 43650 23950
rect 43138 23886 43150 23938
rect 43202 23886 43214 23938
rect 48066 23886 48078 23938
rect 48130 23886 48142 23938
rect 42030 23874 42082 23886
rect 43598 23874 43650 23886
rect 4174 23826 4226 23838
rect 4174 23762 4226 23774
rect 6750 23826 6802 23838
rect 6750 23762 6802 23774
rect 7086 23826 7138 23838
rect 23102 23826 23154 23838
rect 7746 23774 7758 23826
rect 7810 23774 7822 23826
rect 8418 23774 8430 23826
rect 8482 23774 8494 23826
rect 14242 23774 14254 23826
rect 14306 23774 14318 23826
rect 17602 23774 17614 23826
rect 17666 23774 17678 23826
rect 20402 23774 20414 23826
rect 20466 23774 20478 23826
rect 7086 23762 7138 23774
rect 23102 23762 23154 23774
rect 27022 23826 27074 23838
rect 27022 23762 27074 23774
rect 28478 23826 28530 23838
rect 28478 23762 28530 23774
rect 29486 23826 29538 23838
rect 41694 23826 41746 23838
rect 31938 23774 31950 23826
rect 32002 23774 32014 23826
rect 29486 23762 29538 23774
rect 41694 23762 41746 23774
rect 42926 23826 42978 23838
rect 42926 23762 42978 23774
rect 43710 23826 43762 23838
rect 43710 23762 43762 23774
rect 43822 23826 43874 23838
rect 47394 23774 47406 23826
rect 47458 23774 47470 23826
rect 43822 23762 43874 23774
rect 4286 23714 4338 23726
rect 7422 23714 7474 23726
rect 21758 23714 21810 23726
rect 5618 23662 5630 23714
rect 5682 23662 5694 23714
rect 8530 23662 8542 23714
rect 8594 23662 8606 23714
rect 20178 23662 20190 23714
rect 20242 23662 20254 23714
rect 4286 23650 4338 23662
rect 7422 23650 7474 23662
rect 21758 23650 21810 23662
rect 23214 23714 23266 23726
rect 23214 23650 23266 23662
rect 27358 23714 27410 23726
rect 27358 23650 27410 23662
rect 27470 23714 27522 23726
rect 27470 23650 27522 23662
rect 28030 23714 28082 23726
rect 28030 23650 28082 23662
rect 28590 23714 28642 23726
rect 38782 23714 38834 23726
rect 30818 23662 30830 23714
rect 30882 23662 30894 23714
rect 28590 23650 28642 23662
rect 38782 23650 38834 23662
rect 39454 23714 39506 23726
rect 39454 23650 39506 23662
rect 39566 23714 39618 23726
rect 39566 23650 39618 23662
rect 41022 23714 41074 23726
rect 41022 23650 41074 23662
rect 42590 23714 42642 23726
rect 42590 23650 42642 23662
rect 42702 23714 42754 23726
rect 44258 23662 44270 23714
rect 44322 23662 44334 23714
rect 42702 23650 42754 23662
rect 1344 23546 48608 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 48608 23546
rect 1344 23460 48608 23494
rect 3950 23378 4002 23390
rect 13582 23378 13634 23390
rect 5842 23326 5854 23378
rect 5906 23326 5918 23378
rect 3950 23314 4002 23326
rect 13582 23314 13634 23326
rect 14366 23378 14418 23390
rect 14366 23314 14418 23326
rect 14590 23378 14642 23390
rect 14590 23314 14642 23326
rect 17950 23378 18002 23390
rect 17950 23314 18002 23326
rect 24558 23378 24610 23390
rect 24558 23314 24610 23326
rect 36990 23378 37042 23390
rect 41806 23378 41858 23390
rect 38434 23326 38446 23378
rect 38498 23326 38510 23378
rect 36990 23314 37042 23326
rect 41806 23314 41858 23326
rect 42254 23378 42306 23390
rect 42254 23314 42306 23326
rect 42702 23378 42754 23390
rect 42702 23314 42754 23326
rect 44494 23378 44546 23390
rect 47842 23326 47854 23378
rect 47906 23326 47918 23378
rect 44494 23314 44546 23326
rect 3278 23266 3330 23278
rect 3278 23202 3330 23214
rect 3390 23266 3442 23278
rect 6526 23266 6578 23278
rect 4498 23214 4510 23266
rect 4562 23214 4574 23266
rect 5954 23214 5966 23266
rect 6018 23214 6030 23266
rect 3390 23202 3442 23214
rect 6526 23202 6578 23214
rect 6862 23266 6914 23278
rect 6862 23202 6914 23214
rect 8654 23266 8706 23278
rect 8654 23202 8706 23214
rect 8766 23266 8818 23278
rect 8766 23202 8818 23214
rect 13470 23266 13522 23278
rect 13470 23202 13522 23214
rect 14142 23266 14194 23278
rect 23102 23266 23154 23278
rect 14914 23214 14926 23266
rect 14978 23214 14990 23266
rect 16146 23214 16158 23266
rect 16210 23214 16222 23266
rect 18610 23214 18622 23266
rect 18674 23214 18686 23266
rect 20514 23214 20526 23266
rect 20578 23214 20590 23266
rect 14142 23202 14194 23214
rect 23102 23202 23154 23214
rect 23998 23266 24050 23278
rect 23998 23202 24050 23214
rect 24110 23266 24162 23278
rect 24110 23202 24162 23214
rect 24670 23266 24722 23278
rect 24670 23202 24722 23214
rect 25230 23266 25282 23278
rect 25230 23202 25282 23214
rect 25790 23266 25842 23278
rect 25790 23202 25842 23214
rect 26238 23266 26290 23278
rect 26238 23202 26290 23214
rect 26462 23266 26514 23278
rect 36542 23266 36594 23278
rect 44942 23266 44994 23278
rect 29586 23214 29598 23266
rect 29650 23214 29662 23266
rect 39442 23214 39454 23266
rect 39506 23214 39518 23266
rect 26462 23202 26514 23214
rect 36542 23202 36594 23214
rect 44942 23202 44994 23214
rect 46398 23266 46450 23278
rect 46398 23202 46450 23214
rect 3614 23154 3666 23166
rect 3614 23090 3666 23102
rect 4062 23154 4114 23166
rect 15262 23154 15314 23166
rect 21310 23154 21362 23166
rect 27134 23154 27186 23166
rect 30718 23154 30770 23166
rect 4386 23102 4398 23154
rect 4450 23102 4462 23154
rect 5394 23102 5406 23154
rect 5458 23102 5470 23154
rect 15922 23102 15934 23154
rect 15986 23102 15998 23154
rect 18946 23102 18958 23154
rect 19010 23102 19022 23154
rect 20290 23102 20302 23154
rect 20354 23102 20366 23154
rect 22754 23102 22766 23154
rect 22818 23102 22830 23154
rect 30258 23102 30270 23154
rect 30322 23102 30334 23154
rect 4062 23090 4114 23102
rect 15262 23090 15314 23102
rect 21310 23090 21362 23102
rect 27134 23090 27186 23102
rect 30718 23090 30770 23102
rect 31278 23154 31330 23166
rect 31278 23090 31330 23102
rect 31614 23154 31666 23166
rect 31614 23090 31666 23102
rect 31838 23154 31890 23166
rect 31838 23090 31890 23102
rect 33070 23154 33122 23166
rect 34974 23154 35026 23166
rect 33282 23102 33294 23154
rect 33346 23102 33358 23154
rect 34290 23102 34302 23154
rect 34354 23102 34366 23154
rect 33070 23090 33122 23102
rect 34974 23090 35026 23102
rect 35422 23154 35474 23166
rect 35422 23090 35474 23102
rect 35534 23154 35586 23166
rect 35534 23090 35586 23102
rect 35646 23154 35698 23166
rect 35646 23090 35698 23102
rect 35982 23154 36034 23166
rect 35982 23090 36034 23102
rect 36318 23154 36370 23166
rect 37326 23154 37378 23166
rect 36866 23102 36878 23154
rect 36930 23102 36942 23154
rect 36318 23090 36370 23102
rect 37326 23090 37378 23102
rect 38782 23154 38834 23166
rect 38782 23090 38834 23102
rect 39118 23154 39170 23166
rect 39118 23090 39170 23102
rect 41470 23154 41522 23166
rect 41470 23090 41522 23102
rect 41694 23154 41746 23166
rect 42478 23154 42530 23166
rect 41906 23102 41918 23154
rect 41970 23102 41982 23154
rect 41694 23090 41746 23102
rect 42478 23090 42530 23102
rect 45166 23154 45218 23166
rect 45166 23090 45218 23102
rect 45390 23154 45442 23166
rect 48190 23154 48242 23166
rect 45826 23102 45838 23154
rect 45890 23102 45902 23154
rect 45390 23090 45442 23102
rect 48190 23090 48242 23102
rect 14478 23042 14530 23054
rect 14478 22978 14530 22990
rect 15486 23042 15538 23054
rect 15486 22978 15538 22990
rect 16830 23042 16882 23054
rect 26350 23042 26402 23054
rect 33854 23042 33906 23054
rect 17490 22990 17502 23042
rect 17554 22990 17566 23042
rect 27458 22990 27470 23042
rect 27522 22990 27534 23042
rect 16830 22978 16882 22990
rect 26350 22978 26402 22990
rect 33854 22978 33906 22990
rect 34750 23042 34802 23054
rect 34750 22978 34802 22990
rect 36094 23042 36146 23054
rect 36094 22978 36146 22990
rect 37102 23042 37154 23054
rect 37102 22978 37154 22990
rect 37886 23042 37938 23054
rect 37886 22978 37938 22990
rect 42366 23042 42418 23054
rect 42366 22978 42418 22990
rect 45054 23042 45106 23054
rect 45054 22978 45106 22990
rect 47630 23042 47682 23054
rect 47630 22978 47682 22990
rect 3950 22930 4002 22942
rect 3950 22866 4002 22878
rect 8654 22930 8706 22942
rect 8654 22866 8706 22878
rect 13694 22930 13746 22942
rect 13694 22866 13746 22878
rect 23214 22930 23266 22942
rect 23214 22866 23266 22878
rect 23998 22930 24050 22942
rect 23998 22866 24050 22878
rect 24558 22930 24610 22942
rect 24558 22866 24610 22878
rect 25342 22930 25394 22942
rect 25342 22866 25394 22878
rect 25678 22930 25730 22942
rect 44270 22930 44322 22942
rect 32162 22878 32174 22930
rect 32226 22878 32238 22930
rect 25678 22866 25730 22878
rect 44270 22866 44322 22878
rect 44606 22930 44658 22942
rect 44606 22866 44658 22878
rect 46062 22930 46114 22942
rect 46062 22866 46114 22878
rect 46286 22930 46338 22942
rect 46286 22866 46338 22878
rect 1344 22762 48608 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 48608 22762
rect 1344 22676 48608 22710
rect 17390 22594 17442 22606
rect 17390 22530 17442 22542
rect 43934 22594 43986 22606
rect 43934 22530 43986 22542
rect 15710 22482 15762 22494
rect 4610 22430 4622 22482
rect 4674 22430 4686 22482
rect 10882 22430 10894 22482
rect 10946 22430 10958 22482
rect 15710 22418 15762 22430
rect 16270 22482 16322 22494
rect 21646 22482 21698 22494
rect 17826 22430 17838 22482
rect 17890 22430 17902 22482
rect 16270 22418 16322 22430
rect 21646 22418 21698 22430
rect 21982 22482 22034 22494
rect 43710 22482 43762 22494
rect 24546 22430 24558 22482
rect 24610 22430 24622 22482
rect 26674 22430 26686 22482
rect 26738 22430 26750 22482
rect 29138 22430 29150 22482
rect 29202 22430 29214 22482
rect 36082 22430 36094 22482
rect 36146 22430 36158 22482
rect 39890 22430 39902 22482
rect 39954 22430 39966 22482
rect 45266 22430 45278 22482
rect 45330 22430 45342 22482
rect 21982 22418 22034 22430
rect 43710 22418 43762 22430
rect 5630 22370 5682 22382
rect 1698 22318 1710 22370
rect 1762 22318 1774 22370
rect 5630 22306 5682 22318
rect 6414 22370 6466 22382
rect 6414 22306 6466 22318
rect 7422 22370 7474 22382
rect 14478 22370 14530 22382
rect 17166 22370 17218 22382
rect 21422 22370 21474 22382
rect 8082 22318 8094 22370
rect 8146 22318 8158 22370
rect 16930 22318 16942 22370
rect 16994 22318 17006 22370
rect 20738 22318 20750 22370
rect 20802 22318 20814 22370
rect 7422 22306 7474 22318
rect 14478 22306 14530 22318
rect 17166 22306 17218 22318
rect 21422 22306 21474 22318
rect 22990 22370 23042 22382
rect 23438 22370 23490 22382
rect 42814 22370 42866 22382
rect 23090 22318 23102 22370
rect 23154 22318 23166 22370
rect 23762 22318 23774 22370
rect 23826 22318 23838 22370
rect 31938 22318 31950 22370
rect 32002 22318 32014 22370
rect 33170 22318 33182 22370
rect 33234 22318 33246 22370
rect 36978 22318 36990 22370
rect 37042 22318 37054 22370
rect 40450 22318 40462 22370
rect 40514 22318 40526 22370
rect 41346 22318 41358 22370
rect 41410 22318 41422 22370
rect 42018 22318 42030 22370
rect 42082 22318 42094 22370
rect 22990 22306 23042 22318
rect 23438 22306 23490 22318
rect 42814 22306 42866 22318
rect 43262 22370 43314 22382
rect 48066 22318 48078 22370
rect 48130 22318 48142 22370
rect 43262 22306 43314 22318
rect 6302 22258 6354 22270
rect 2482 22206 2494 22258
rect 2546 22206 2558 22258
rect 6302 22194 6354 22206
rect 7534 22258 7586 22270
rect 17502 22258 17554 22270
rect 22878 22258 22930 22270
rect 32286 22258 32338 22270
rect 8754 22206 8766 22258
rect 8818 22206 8830 22258
rect 19954 22206 19966 22258
rect 20018 22206 20030 22258
rect 31266 22206 31278 22258
rect 31330 22206 31342 22258
rect 7534 22194 7586 22206
rect 17502 22194 17554 22206
rect 22878 22194 22930 22206
rect 32286 22194 32338 22206
rect 32846 22258 32898 22270
rect 42926 22258 42978 22270
rect 33954 22206 33966 22258
rect 34018 22206 34030 22258
rect 37762 22206 37774 22258
rect 37826 22206 37838 22258
rect 40226 22206 40238 22258
rect 40290 22206 40302 22258
rect 42354 22206 42366 22258
rect 42418 22206 42430 22258
rect 32846 22194 32898 22206
rect 42926 22194 42978 22206
rect 43374 22258 43426 22270
rect 47394 22206 47406 22258
rect 47458 22206 47470 22258
rect 43374 22194 43426 22206
rect 5742 22146 5794 22158
rect 5742 22082 5794 22094
rect 5966 22146 6018 22158
rect 5966 22082 6018 22094
rect 6078 22146 6130 22158
rect 6078 22082 6130 22094
rect 7758 22146 7810 22158
rect 7758 22082 7810 22094
rect 14590 22146 14642 22158
rect 14590 22082 14642 22094
rect 14702 22146 14754 22158
rect 14702 22082 14754 22094
rect 14926 22146 14978 22158
rect 14926 22082 14978 22094
rect 16718 22146 16770 22158
rect 16718 22082 16770 22094
rect 21870 22146 21922 22158
rect 21870 22082 21922 22094
rect 22094 22146 22146 22158
rect 22094 22082 22146 22094
rect 22766 22146 22818 22158
rect 22766 22082 22818 22094
rect 27358 22146 27410 22158
rect 27358 22082 27410 22094
rect 27470 22146 27522 22158
rect 27470 22082 27522 22094
rect 27582 22146 27634 22158
rect 27582 22082 27634 22094
rect 27806 22146 27858 22158
rect 27806 22082 27858 22094
rect 28478 22146 28530 22158
rect 28478 22082 28530 22094
rect 32398 22146 32450 22158
rect 32398 22082 32450 22094
rect 32622 22146 32674 22158
rect 41458 22094 41470 22146
rect 41522 22094 41534 22146
rect 44258 22094 44270 22146
rect 44322 22094 44334 22146
rect 32622 22082 32674 22094
rect 1344 21978 48608 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 48608 21978
rect 1344 21892 48608 21926
rect 3838 21810 3890 21822
rect 3838 21746 3890 21758
rect 6862 21810 6914 21822
rect 6862 21746 6914 21758
rect 8654 21810 8706 21822
rect 8654 21746 8706 21758
rect 16718 21810 16770 21822
rect 16718 21746 16770 21758
rect 23102 21810 23154 21822
rect 23102 21746 23154 21758
rect 23326 21810 23378 21822
rect 23326 21746 23378 21758
rect 24334 21810 24386 21822
rect 24334 21746 24386 21758
rect 24446 21810 24498 21822
rect 24446 21746 24498 21758
rect 28814 21810 28866 21822
rect 28814 21746 28866 21758
rect 29486 21810 29538 21822
rect 29486 21746 29538 21758
rect 30158 21810 30210 21822
rect 30158 21746 30210 21758
rect 31726 21810 31778 21822
rect 31726 21746 31778 21758
rect 32398 21810 32450 21822
rect 32398 21746 32450 21758
rect 33070 21810 33122 21822
rect 33070 21746 33122 21758
rect 35534 21810 35586 21822
rect 35534 21746 35586 21758
rect 38110 21810 38162 21822
rect 38110 21746 38162 21758
rect 38782 21810 38834 21822
rect 38782 21746 38834 21758
rect 41806 21810 41858 21822
rect 41806 21746 41858 21758
rect 41918 21810 41970 21822
rect 41918 21746 41970 21758
rect 47966 21810 48018 21822
rect 47966 21746 48018 21758
rect 3166 21698 3218 21710
rect 3166 21634 3218 21646
rect 3278 21698 3330 21710
rect 3278 21634 3330 21646
rect 3502 21698 3554 21710
rect 3502 21634 3554 21646
rect 4958 21698 5010 21710
rect 4958 21634 5010 21646
rect 6078 21698 6130 21710
rect 6078 21634 6130 21646
rect 6750 21698 6802 21710
rect 6750 21634 6802 21646
rect 7534 21698 7586 21710
rect 7534 21634 7586 21646
rect 8430 21698 8482 21710
rect 8430 21634 8482 21646
rect 14030 21698 14082 21710
rect 14030 21634 14082 21646
rect 14254 21698 14306 21710
rect 23438 21698 23490 21710
rect 34190 21698 34242 21710
rect 18050 21646 18062 21698
rect 18114 21646 18126 21698
rect 27346 21646 27358 21698
rect 27410 21646 27422 21698
rect 30482 21646 30494 21698
rect 30546 21646 30558 21698
rect 33394 21646 33406 21698
rect 33458 21646 33470 21698
rect 14254 21634 14306 21646
rect 23438 21634 23490 21646
rect 34190 21634 34242 21646
rect 34638 21698 34690 21710
rect 34638 21634 34690 21646
rect 39118 21698 39170 21710
rect 39118 21634 39170 21646
rect 44494 21698 44546 21710
rect 44494 21634 44546 21646
rect 44606 21698 44658 21710
rect 44606 21634 44658 21646
rect 45614 21698 45666 21710
rect 45614 21634 45666 21646
rect 3614 21586 3666 21598
rect 3614 21522 3666 21534
rect 3950 21586 4002 21598
rect 3950 21522 4002 21534
rect 4286 21586 4338 21598
rect 4286 21522 4338 21534
rect 4510 21586 4562 21598
rect 4510 21522 4562 21534
rect 5182 21586 5234 21598
rect 5182 21522 5234 21534
rect 5854 21586 5906 21598
rect 5854 21522 5906 21534
rect 6526 21586 6578 21598
rect 6526 21522 6578 21534
rect 7870 21586 7922 21598
rect 7870 21522 7922 21534
rect 8206 21586 8258 21598
rect 8206 21522 8258 21534
rect 8878 21586 8930 21598
rect 14814 21586 14866 21598
rect 16382 21586 16434 21598
rect 10770 21534 10782 21586
rect 10834 21534 10846 21586
rect 15810 21534 15822 21586
rect 15874 21534 15886 21586
rect 8878 21522 8930 21534
rect 14814 21522 14866 21534
rect 16382 21522 16434 21534
rect 16606 21586 16658 21598
rect 16606 21522 16658 21534
rect 16942 21586 16994 21598
rect 23998 21586 24050 21598
rect 22418 21534 22430 21586
rect 22482 21534 22494 21586
rect 16942 21522 16994 21534
rect 23998 21522 24050 21534
rect 24222 21586 24274 21598
rect 28478 21586 28530 21598
rect 28018 21534 28030 21586
rect 28082 21534 28094 21586
rect 24222 21522 24274 21534
rect 28478 21522 28530 21534
rect 28814 21586 28866 21598
rect 28814 21522 28866 21534
rect 29038 21586 29090 21598
rect 29038 21522 29090 21534
rect 30830 21586 30882 21598
rect 30830 21522 30882 21534
rect 31278 21586 31330 21598
rect 31278 21522 31330 21534
rect 31838 21586 31890 21598
rect 31838 21522 31890 21534
rect 32286 21586 32338 21598
rect 32286 21522 32338 21534
rect 32510 21586 32562 21598
rect 34414 21586 34466 21598
rect 33954 21534 33966 21586
rect 34018 21534 34030 21586
rect 32510 21522 32562 21534
rect 34414 21522 34466 21534
rect 35086 21586 35138 21598
rect 37438 21586 37490 21598
rect 41694 21586 41746 21598
rect 43038 21586 43090 21598
rect 36306 21534 36318 21586
rect 36370 21534 36382 21586
rect 38322 21534 38334 21586
rect 38386 21534 38398 21586
rect 41458 21534 41470 21586
rect 41522 21534 41534 21586
rect 42130 21534 42142 21586
rect 42194 21534 42206 21586
rect 35086 21522 35138 21534
rect 37438 21522 37490 21534
rect 41694 21522 41746 21534
rect 43038 21522 43090 21534
rect 44830 21586 44882 21598
rect 45502 21586 45554 21598
rect 45042 21534 45054 21586
rect 45106 21534 45118 21586
rect 44830 21522 44882 21534
rect 45502 21522 45554 21534
rect 46062 21586 46114 21598
rect 46062 21522 46114 21534
rect 46398 21586 46450 21598
rect 46398 21522 46450 21534
rect 46734 21586 46786 21598
rect 46734 21522 46786 21534
rect 47182 21586 47234 21598
rect 47182 21522 47234 21534
rect 47294 21586 47346 21598
rect 47294 21522 47346 21534
rect 4734 21474 4786 21486
rect 4734 21410 4786 21422
rect 6302 21474 6354 21486
rect 6302 21410 6354 21422
rect 9662 21474 9714 21486
rect 14590 21474 14642 21486
rect 11442 21422 11454 21474
rect 11506 21422 11518 21474
rect 13570 21422 13582 21474
rect 13634 21422 13646 21474
rect 13906 21422 13918 21474
rect 13970 21422 13982 21474
rect 9662 21410 9714 21422
rect 14590 21410 14642 21422
rect 15598 21474 15650 21486
rect 31054 21474 31106 21486
rect 25218 21422 25230 21474
rect 25282 21422 25294 21474
rect 15598 21410 15650 21422
rect 31054 21410 31106 21422
rect 34302 21474 34354 21486
rect 36878 21474 36930 21486
rect 35970 21422 35982 21474
rect 36034 21422 36046 21474
rect 34302 21410 34354 21422
rect 36878 21410 36930 21422
rect 37214 21474 37266 21486
rect 37214 21410 37266 21422
rect 37774 21474 37826 21486
rect 37774 21410 37826 21422
rect 42478 21474 42530 21486
rect 42478 21410 42530 21422
rect 42590 21474 42642 21486
rect 42590 21410 42642 21422
rect 45278 21474 45330 21486
rect 45278 21410 45330 21422
rect 46958 21474 47010 21486
rect 46958 21410 47010 21422
rect 47742 21474 47794 21486
rect 47742 21410 47794 21422
rect 47854 21474 47906 21486
rect 47854 21410 47906 21422
rect 6862 21362 6914 21374
rect 15486 21362 15538 21374
rect 15138 21310 15150 21362
rect 15202 21310 15214 21362
rect 6862 21298 6914 21310
rect 15486 21298 15538 21310
rect 23774 21362 23826 21374
rect 23774 21298 23826 21310
rect 34974 21362 35026 21374
rect 34974 21298 35026 21310
rect 42926 21362 42978 21374
rect 42926 21298 42978 21310
rect 45950 21362 46002 21374
rect 45950 21298 46002 21310
rect 46286 21362 46338 21374
rect 46286 21298 46338 21310
rect 1344 21194 48608 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 48608 21194
rect 1344 21108 48608 21142
rect 10782 21026 10834 21038
rect 29486 21026 29538 21038
rect 19282 20974 19294 21026
rect 19346 20974 19358 21026
rect 27122 20974 27134 21026
rect 27186 20974 27198 21026
rect 10782 20962 10834 20974
rect 29486 20962 29538 20974
rect 43934 21026 43986 21038
rect 44258 20974 44270 21026
rect 44322 20974 44334 21026
rect 43934 20962 43986 20974
rect 11454 20914 11506 20926
rect 2482 20862 2494 20914
rect 2546 20862 2558 20914
rect 4610 20862 4622 20914
rect 4674 20862 4686 20914
rect 6402 20862 6414 20914
rect 6466 20862 6478 20914
rect 8530 20862 8542 20914
rect 8594 20862 8606 20914
rect 9650 20862 9662 20914
rect 9714 20862 9726 20914
rect 11454 20850 11506 20862
rect 14702 20914 14754 20926
rect 20638 20914 20690 20926
rect 18386 20862 18398 20914
rect 18450 20862 18462 20914
rect 14702 20850 14754 20862
rect 20638 20850 20690 20862
rect 32062 20914 32114 20926
rect 42926 20914 42978 20926
rect 41794 20862 41806 20914
rect 41858 20862 41870 20914
rect 32062 20850 32114 20862
rect 42926 20850 42978 20862
rect 43710 20914 43762 20926
rect 46050 20862 46062 20914
rect 46114 20862 46126 20914
rect 48178 20862 48190 20914
rect 48242 20862 48254 20914
rect 43710 20850 43762 20862
rect 11006 20802 11058 20814
rect 1698 20750 1710 20802
rect 1762 20750 1774 20802
rect 5730 20750 5742 20802
rect 5794 20750 5806 20802
rect 11006 20738 11058 20750
rect 14142 20802 14194 20814
rect 14142 20738 14194 20750
rect 14814 20802 14866 20814
rect 19966 20802 20018 20814
rect 15138 20750 15150 20802
rect 15202 20750 15214 20802
rect 17154 20750 17166 20802
rect 17218 20750 17230 20802
rect 14814 20738 14866 20750
rect 19966 20738 20018 20750
rect 21646 20802 21698 20814
rect 21646 20738 21698 20750
rect 21982 20802 22034 20814
rect 27806 20802 27858 20814
rect 23202 20750 23214 20802
rect 23266 20750 23278 20802
rect 25106 20750 25118 20802
rect 25170 20750 25182 20802
rect 26450 20750 26462 20802
rect 26514 20750 26526 20802
rect 21982 20738 22034 20750
rect 27806 20738 27858 20750
rect 33966 20802 34018 20814
rect 41682 20750 41694 20802
rect 41746 20750 41758 20802
rect 45378 20750 45390 20802
rect 45442 20750 45454 20802
rect 33966 20738 34018 20750
rect 9998 20690 10050 20702
rect 18286 20690 18338 20702
rect 9202 20638 9214 20690
rect 9266 20687 9278 20690
rect 9538 20687 9550 20690
rect 9266 20641 9550 20687
rect 9266 20638 9278 20641
rect 9538 20638 9550 20641
rect 9602 20638 9614 20690
rect 15250 20638 15262 20690
rect 15314 20638 15326 20690
rect 9998 20626 10050 20638
rect 18286 20626 18338 20638
rect 19742 20690 19794 20702
rect 19742 20626 19794 20638
rect 19854 20690 19906 20702
rect 19854 20626 19906 20638
rect 21310 20690 21362 20702
rect 21310 20626 21362 20638
rect 21422 20690 21474 20702
rect 21422 20626 21474 20638
rect 21870 20690 21922 20702
rect 27582 20690 27634 20702
rect 23538 20638 23550 20690
rect 23602 20638 23614 20690
rect 25890 20638 25902 20690
rect 25954 20638 25966 20690
rect 21870 20626 21922 20638
rect 27582 20626 27634 20638
rect 27694 20690 27746 20702
rect 27694 20626 27746 20638
rect 29598 20690 29650 20702
rect 41246 20690 41298 20702
rect 29922 20638 29934 20690
rect 29986 20638 29998 20690
rect 29598 20626 29650 20638
rect 41246 20626 41298 20638
rect 41358 20690 41410 20702
rect 41358 20626 41410 20638
rect 42142 20690 42194 20702
rect 42142 20626 42194 20638
rect 42814 20690 42866 20702
rect 42814 20626 42866 20638
rect 8990 20578 9042 20590
rect 8990 20514 9042 20526
rect 9774 20578 9826 20590
rect 14590 20578 14642 20590
rect 10434 20526 10446 20578
rect 10498 20526 10510 20578
rect 9774 20514 9826 20526
rect 14590 20514 14642 20526
rect 20750 20578 20802 20590
rect 28366 20578 28418 20590
rect 22866 20526 22878 20578
rect 22930 20526 22942 20578
rect 20750 20514 20802 20526
rect 28366 20514 28418 20526
rect 30270 20578 30322 20590
rect 30270 20514 30322 20526
rect 30718 20578 30770 20590
rect 30718 20514 30770 20526
rect 31166 20578 31218 20590
rect 31166 20514 31218 20526
rect 35534 20578 35586 20590
rect 35534 20514 35586 20526
rect 36094 20578 36146 20590
rect 36094 20514 36146 20526
rect 37214 20578 37266 20590
rect 37214 20514 37266 20526
rect 41022 20578 41074 20590
rect 41022 20514 41074 20526
rect 42254 20578 42306 20590
rect 42254 20514 42306 20526
rect 42366 20578 42418 20590
rect 42366 20514 42418 20526
rect 43374 20578 43426 20590
rect 43374 20514 43426 20526
rect 1344 20410 48608 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 48608 20410
rect 1344 20324 48608 20358
rect 9886 20242 9938 20254
rect 33294 20242 33346 20254
rect 16258 20190 16270 20242
rect 16322 20190 16334 20242
rect 9886 20178 9938 20190
rect 33294 20178 33346 20190
rect 33630 20242 33682 20254
rect 33630 20178 33682 20190
rect 41246 20242 41298 20254
rect 41246 20178 41298 20190
rect 9774 20130 9826 20142
rect 23102 20130 23154 20142
rect 25902 20130 25954 20142
rect 12786 20078 12798 20130
rect 12850 20078 12862 20130
rect 23874 20078 23886 20130
rect 23938 20078 23950 20130
rect 9774 20066 9826 20078
rect 23102 20066 23154 20078
rect 25902 20066 25954 20078
rect 30382 20130 30434 20142
rect 30382 20066 30434 20078
rect 31838 20130 31890 20142
rect 31838 20066 31890 20078
rect 33854 20130 33906 20142
rect 33854 20066 33906 20078
rect 35310 20130 35362 20142
rect 35310 20066 35362 20078
rect 41918 20130 41970 20142
rect 41918 20066 41970 20078
rect 9998 20018 10050 20030
rect 8194 19966 8206 20018
rect 8258 19966 8270 20018
rect 9998 19954 10050 19966
rect 10446 20018 10498 20030
rect 16606 20018 16658 20030
rect 15922 19966 15934 20018
rect 15986 19966 15998 20018
rect 10446 19954 10498 19966
rect 16606 19954 16658 19966
rect 16830 20018 16882 20030
rect 23550 20018 23602 20030
rect 18834 19966 18846 20018
rect 18898 19966 18910 20018
rect 16830 19954 16882 19966
rect 23550 19954 23602 19966
rect 25566 20018 25618 20030
rect 25566 19954 25618 19966
rect 26798 20018 26850 20030
rect 26798 19954 26850 19966
rect 28366 20018 28418 20030
rect 28366 19954 28418 19966
rect 33406 20018 33458 20030
rect 33406 19954 33458 19966
rect 34302 20018 34354 20030
rect 40014 20018 40066 20030
rect 41134 20018 41186 20030
rect 36530 19966 36542 20018
rect 36594 19966 36606 20018
rect 40338 19966 40350 20018
rect 40402 19966 40414 20018
rect 40898 19966 40910 20018
rect 40962 19966 40974 20018
rect 34302 19954 34354 19966
rect 40014 19954 40066 19966
rect 41134 19954 41186 19966
rect 41358 20018 41410 20030
rect 42142 20018 42194 20030
rect 41570 19966 41582 20018
rect 41634 19966 41646 20018
rect 43362 19966 43374 20018
rect 43426 19966 43438 20018
rect 41358 19954 41410 19966
rect 42142 19954 42194 19966
rect 8878 19906 8930 19918
rect 24334 19906 24386 19918
rect 3378 19854 3390 19906
rect 3442 19854 3454 19906
rect 22418 19854 22430 19906
rect 22482 19854 22494 19906
rect 8878 19842 8930 19854
rect 24334 19842 24386 19854
rect 26350 19906 26402 19918
rect 26350 19842 26402 19854
rect 29486 19906 29538 19918
rect 29486 19842 29538 19854
rect 31502 19906 31554 19918
rect 31502 19842 31554 19854
rect 32398 19906 32450 19918
rect 32398 19842 32450 19854
rect 33518 19906 33570 19918
rect 33518 19842 33570 19854
rect 34974 19906 35026 19918
rect 34974 19842 35026 19854
rect 35982 19906 36034 19918
rect 35982 19842 36034 19854
rect 36094 19906 36146 19918
rect 42478 19906 42530 19918
rect 37202 19854 37214 19906
rect 37266 19854 37278 19906
rect 39330 19854 39342 19906
rect 39394 19854 39406 19906
rect 40226 19854 40238 19906
rect 40290 19854 40302 19906
rect 46834 19854 46846 19906
rect 46898 19854 46910 19906
rect 36094 19842 36146 19854
rect 42478 19842 42530 19854
rect 8766 19794 8818 19806
rect 8766 19730 8818 19742
rect 31950 19794 32002 19806
rect 31950 19730 32002 19742
rect 32510 19794 32562 19806
rect 34626 19742 34638 19794
rect 34690 19791 34702 19794
rect 35298 19791 35310 19794
rect 34690 19745 35310 19791
rect 34690 19742 34702 19745
rect 35298 19742 35310 19745
rect 35362 19742 35374 19794
rect 32510 19730 32562 19742
rect 1344 19626 48608 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 48608 19626
rect 1344 19540 48608 19574
rect 7422 19458 7474 19470
rect 7074 19406 7086 19458
rect 7138 19406 7150 19458
rect 7422 19394 7474 19406
rect 20750 19458 20802 19470
rect 20750 19394 20802 19406
rect 31054 19458 31106 19470
rect 31054 19394 31106 19406
rect 42590 19458 42642 19470
rect 42590 19394 42642 19406
rect 16382 19346 16434 19358
rect 20638 19346 20690 19358
rect 44942 19346 44994 19358
rect 4610 19294 4622 19346
rect 4674 19294 4686 19346
rect 8978 19294 8990 19346
rect 9042 19294 9054 19346
rect 11106 19294 11118 19346
rect 11170 19294 11182 19346
rect 13458 19294 13470 19346
rect 13522 19294 13534 19346
rect 15698 19294 15710 19346
rect 15762 19294 15774 19346
rect 18162 19294 18174 19346
rect 18226 19294 18238 19346
rect 20290 19294 20302 19346
rect 20354 19294 20366 19346
rect 21410 19294 21422 19346
rect 21474 19294 21486 19346
rect 23538 19294 23550 19346
rect 23602 19294 23614 19346
rect 25666 19294 25678 19346
rect 25730 19294 25742 19346
rect 27794 19294 27806 19346
rect 27858 19294 27870 19346
rect 32610 19294 32622 19346
rect 32674 19294 32686 19346
rect 34738 19294 34750 19346
rect 34802 19294 34814 19346
rect 42018 19294 42030 19346
rect 42082 19294 42094 19346
rect 44146 19294 44158 19346
rect 44210 19294 44222 19346
rect 46050 19294 46062 19346
rect 46114 19294 46126 19346
rect 48178 19294 48190 19346
rect 48242 19294 48254 19346
rect 16382 19282 16434 19294
rect 20638 19282 20690 19294
rect 44942 19282 44994 19294
rect 6526 19234 6578 19246
rect 1810 19182 1822 19234
rect 1874 19182 1886 19234
rect 6526 19170 6578 19182
rect 6862 19234 6914 19246
rect 6862 19170 6914 19182
rect 7646 19234 7698 19246
rect 30046 19234 30098 19246
rect 35422 19234 35474 19246
rect 44830 19234 44882 19246
rect 8306 19182 8318 19234
rect 8370 19182 8382 19234
rect 15250 19182 15262 19234
rect 15314 19182 15326 19234
rect 17490 19182 17502 19234
rect 17554 19182 17566 19234
rect 7646 19170 7698 19182
rect 24322 19170 24334 19222
rect 24386 19170 24398 19222
rect 24882 19182 24894 19234
rect 24946 19182 24958 19234
rect 30370 19182 30382 19234
rect 30434 19182 30446 19234
rect 30706 19182 30718 19234
rect 30770 19182 30782 19234
rect 31938 19182 31950 19234
rect 32002 19182 32014 19234
rect 37314 19182 37326 19234
rect 37378 19182 37390 19234
rect 43922 19182 43934 19234
rect 43986 19182 43998 19234
rect 45378 19182 45390 19234
rect 45442 19182 45454 19234
rect 30046 19170 30098 19182
rect 35422 19170 35474 19182
rect 44830 19170 44882 19182
rect 5630 19122 5682 19134
rect 2482 19070 2494 19122
rect 2546 19070 2558 19122
rect 5630 19058 5682 19070
rect 13806 19122 13858 19134
rect 13806 19058 13858 19070
rect 14814 19122 14866 19134
rect 14814 19058 14866 19070
rect 29150 19122 29202 19134
rect 29150 19058 29202 19070
rect 29710 19122 29762 19134
rect 29710 19058 29762 19070
rect 30158 19122 30210 19134
rect 30158 19058 30210 19070
rect 35534 19122 35586 19134
rect 35534 19058 35586 19070
rect 35758 19122 35810 19134
rect 35758 19058 35810 19070
rect 36206 19122 36258 19134
rect 36206 19058 36258 19070
rect 42814 19122 42866 19134
rect 42814 19058 42866 19070
rect 43262 19122 43314 19134
rect 43262 19058 43314 19070
rect 5742 19010 5794 19022
rect 5742 18946 5794 18958
rect 5854 19010 5906 19022
rect 5854 18946 5906 18958
rect 6638 19010 6690 19022
rect 6638 18946 6690 18958
rect 13582 19010 13634 19022
rect 13582 18946 13634 18958
rect 14366 19010 14418 19022
rect 14366 18946 14418 18958
rect 29262 19010 29314 19022
rect 29262 18946 29314 18958
rect 29934 19010 29986 19022
rect 29934 18946 29986 18958
rect 30942 19010 30994 19022
rect 30942 18946 30994 18958
rect 31502 19010 31554 19022
rect 31502 18946 31554 18958
rect 35198 19010 35250 19022
rect 35198 18946 35250 18958
rect 35310 19010 35362 19022
rect 35310 18946 35362 18958
rect 36318 19010 36370 19022
rect 36318 18946 36370 18958
rect 42702 19010 42754 19022
rect 42702 18946 42754 18958
rect 1344 18842 48608 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 48608 18842
rect 1344 18756 48608 18790
rect 4398 18674 4450 18686
rect 4398 18610 4450 18622
rect 4622 18674 4674 18686
rect 24670 18674 24722 18686
rect 21858 18622 21870 18674
rect 21922 18622 21934 18674
rect 4622 18610 4674 18622
rect 24670 18610 24722 18622
rect 35646 18674 35698 18686
rect 35646 18610 35698 18622
rect 36542 18674 36594 18686
rect 36542 18610 36594 18622
rect 47518 18674 47570 18686
rect 47518 18610 47570 18622
rect 33630 18562 33682 18574
rect 17490 18510 17502 18562
rect 17554 18510 17566 18562
rect 20962 18510 20974 18562
rect 21026 18510 21038 18562
rect 28018 18510 28030 18562
rect 28082 18510 28094 18562
rect 31154 18510 31166 18562
rect 31218 18510 31230 18562
rect 31490 18510 31502 18562
rect 31554 18510 31566 18562
rect 33630 18498 33682 18510
rect 33854 18562 33906 18574
rect 33854 18498 33906 18510
rect 35422 18562 35474 18574
rect 35422 18498 35474 18510
rect 35870 18562 35922 18574
rect 35870 18498 35922 18510
rect 36430 18562 36482 18574
rect 36430 18498 36482 18510
rect 47630 18562 47682 18574
rect 47630 18498 47682 18510
rect 3502 18450 3554 18462
rect 3154 18398 3166 18450
rect 3218 18398 3230 18450
rect 3502 18386 3554 18398
rect 3726 18450 3778 18462
rect 4510 18450 4562 18462
rect 17838 18450 17890 18462
rect 21310 18450 21362 18462
rect 4050 18398 4062 18450
rect 4114 18398 4126 18450
rect 5282 18398 5294 18450
rect 5346 18398 5358 18450
rect 10658 18398 10670 18450
rect 10722 18398 10734 18450
rect 11442 18398 11454 18450
rect 11506 18398 11518 18450
rect 12114 18398 12126 18450
rect 12178 18398 12190 18450
rect 18610 18398 18622 18450
rect 18674 18398 18686 18450
rect 20066 18398 20078 18450
rect 20130 18398 20142 18450
rect 3726 18386 3778 18398
rect 4510 18386 4562 18398
rect 17838 18386 17890 18398
rect 21310 18386 21362 18398
rect 22206 18450 22258 18462
rect 22206 18386 22258 18398
rect 22654 18450 22706 18462
rect 22654 18386 22706 18398
rect 23214 18450 23266 18462
rect 23214 18386 23266 18398
rect 23550 18450 23602 18462
rect 32286 18450 32338 18462
rect 25218 18398 25230 18450
rect 25282 18398 25294 18450
rect 30930 18398 30942 18450
rect 30994 18398 31006 18450
rect 31714 18398 31726 18450
rect 31778 18398 31790 18450
rect 23550 18386 23602 18398
rect 32286 18386 32338 18398
rect 34862 18450 34914 18462
rect 35534 18450 35586 18462
rect 35186 18398 35198 18450
rect 35250 18398 35262 18450
rect 34862 18386 34914 18398
rect 35534 18386 35586 18398
rect 36766 18450 36818 18462
rect 37090 18398 37102 18450
rect 37154 18398 37166 18450
rect 40898 18398 40910 18450
rect 40962 18398 40974 18450
rect 44258 18398 44270 18450
rect 44322 18398 44334 18450
rect 36766 18386 36818 18398
rect 8654 18338 8706 18350
rect 15710 18338 15762 18350
rect 6066 18286 6078 18338
rect 6130 18286 6142 18338
rect 8194 18286 8206 18338
rect 8258 18286 8270 18338
rect 14242 18286 14254 18338
rect 14306 18286 14318 18338
rect 8654 18274 8706 18286
rect 15710 18274 15762 18286
rect 16942 18338 16994 18350
rect 24110 18338 24162 18350
rect 19954 18286 19966 18338
rect 20018 18286 20030 18338
rect 16942 18274 16994 18286
rect 24110 18274 24162 18286
rect 33182 18338 33234 18350
rect 33182 18274 33234 18286
rect 34302 18338 34354 18350
rect 40238 18338 40290 18350
rect 48190 18338 48242 18350
rect 37762 18286 37774 18338
rect 37826 18286 37838 18338
rect 39890 18286 39902 18338
rect 39954 18286 39966 18338
rect 41682 18286 41694 18338
rect 41746 18286 41758 18338
rect 43810 18286 43822 18338
rect 43874 18286 43886 18338
rect 44930 18286 44942 18338
rect 44994 18286 45006 18338
rect 47058 18286 47070 18338
rect 47122 18286 47134 18338
rect 34302 18274 34354 18286
rect 40238 18274 40290 18286
rect 48190 18274 48242 18286
rect 10670 18226 10722 18238
rect 10670 18162 10722 18174
rect 11006 18226 11058 18238
rect 11006 18162 11058 18174
rect 15934 18226 15986 18238
rect 33966 18226 34018 18238
rect 16258 18174 16270 18226
rect 16322 18174 16334 18226
rect 18274 18174 18286 18226
rect 18338 18174 18350 18226
rect 15934 18162 15986 18174
rect 33966 18162 34018 18174
rect 40350 18226 40402 18238
rect 40350 18162 40402 18174
rect 1344 18058 48608 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 48608 18058
rect 1344 17972 48608 18006
rect 23326 17890 23378 17902
rect 43710 17890 43762 17902
rect 23650 17838 23662 17890
rect 23714 17887 23726 17890
rect 24210 17887 24222 17890
rect 23714 17841 24222 17887
rect 23714 17838 23726 17841
rect 24210 17838 24222 17841
rect 24274 17887 24286 17890
rect 25330 17887 25342 17890
rect 24274 17841 25342 17887
rect 24274 17838 24286 17841
rect 25330 17838 25342 17841
rect 25394 17838 25406 17890
rect 23326 17826 23378 17838
rect 43710 17826 43762 17838
rect 20862 17778 20914 17790
rect 4610 17726 4622 17778
rect 4674 17726 4686 17778
rect 10546 17726 10558 17778
rect 10610 17726 10622 17778
rect 12674 17726 12686 17778
rect 12738 17726 12750 17778
rect 14130 17726 14142 17778
rect 14194 17726 14206 17778
rect 20862 17714 20914 17726
rect 23438 17778 23490 17790
rect 23438 17714 23490 17726
rect 23886 17778 23938 17790
rect 23886 17714 23938 17726
rect 24334 17778 24386 17790
rect 24334 17714 24386 17726
rect 25342 17778 25394 17790
rect 25342 17714 25394 17726
rect 28030 17778 28082 17790
rect 34526 17778 34578 17790
rect 29138 17726 29150 17778
rect 29202 17726 29214 17778
rect 33506 17726 33518 17778
rect 33570 17726 33582 17778
rect 28030 17714 28082 17726
rect 34526 17714 34578 17726
rect 37214 17778 37266 17790
rect 43598 17778 43650 17790
rect 46174 17778 46226 17790
rect 40898 17726 40910 17778
rect 40962 17726 40974 17778
rect 45714 17726 45726 17778
rect 45778 17726 45790 17778
rect 37214 17714 37266 17726
rect 43598 17714 43650 17726
rect 46174 17714 46226 17726
rect 47182 17778 47234 17790
rect 47182 17714 47234 17726
rect 25790 17666 25842 17678
rect 27134 17666 27186 17678
rect 1810 17614 1822 17666
rect 1874 17614 1886 17666
rect 8866 17614 8878 17666
rect 8930 17614 8942 17666
rect 9874 17614 9886 17666
rect 9938 17614 9950 17666
rect 17042 17614 17054 17666
rect 17106 17614 17118 17666
rect 19058 17614 19070 17666
rect 19122 17614 19134 17666
rect 19618 17614 19630 17666
rect 19682 17614 19694 17666
rect 26338 17614 26350 17666
rect 26402 17614 26414 17666
rect 25790 17602 25842 17614
rect 27134 17602 27186 17614
rect 27694 17666 27746 17678
rect 32398 17666 32450 17678
rect 34862 17666 34914 17678
rect 32050 17614 32062 17666
rect 32114 17614 32126 17666
rect 33170 17614 33182 17666
rect 33234 17614 33246 17666
rect 27694 17602 27746 17614
rect 32398 17602 32450 17614
rect 34862 17602 34914 17614
rect 35422 17666 35474 17678
rect 45278 17666 45330 17678
rect 37874 17614 37886 17666
rect 37938 17614 37950 17666
rect 43362 17614 43374 17666
rect 43426 17614 43438 17666
rect 35422 17602 35474 17614
rect 45278 17602 45330 17614
rect 45614 17666 45666 17678
rect 45614 17602 45666 17614
rect 9214 17554 9266 17566
rect 17390 17554 17442 17566
rect 2482 17502 2494 17554
rect 2546 17502 2558 17554
rect 16258 17502 16270 17554
rect 16322 17502 16334 17554
rect 9214 17490 9266 17502
rect 17390 17490 17442 17502
rect 17502 17554 17554 17566
rect 17502 17490 17554 17502
rect 17614 17554 17666 17566
rect 21870 17554 21922 17566
rect 19954 17502 19966 17554
rect 20018 17502 20030 17554
rect 17614 17490 17666 17502
rect 21870 17490 21922 17502
rect 22430 17554 22482 17566
rect 22430 17490 22482 17502
rect 22766 17554 22818 17566
rect 22766 17490 22818 17502
rect 22990 17554 23042 17566
rect 22990 17490 23042 17502
rect 25678 17554 25730 17566
rect 25678 17490 25730 17502
rect 27246 17554 27298 17566
rect 27246 17490 27298 17502
rect 28590 17554 28642 17566
rect 44158 17554 44210 17566
rect 31266 17502 31278 17554
rect 31330 17502 31342 17554
rect 36418 17502 36430 17554
rect 36482 17502 36494 17554
rect 28590 17490 28642 17502
rect 44158 17490 44210 17502
rect 46622 17554 46674 17566
rect 48190 17554 48242 17566
rect 47842 17502 47854 17554
rect 47906 17502 47918 17554
rect 46622 17490 46674 17502
rect 48190 17490 48242 17502
rect 5966 17442 6018 17454
rect 5618 17390 5630 17442
rect 5682 17390 5694 17442
rect 5966 17378 6018 17390
rect 6974 17442 7026 17454
rect 6974 17378 7026 17390
rect 9102 17442 9154 17454
rect 9102 17378 9154 17390
rect 18174 17442 18226 17454
rect 21310 17442 21362 17454
rect 18610 17390 18622 17442
rect 18674 17390 18686 17442
rect 19618 17390 19630 17442
rect 19682 17390 19694 17442
rect 18174 17378 18226 17390
rect 21310 17378 21362 17390
rect 22654 17442 22706 17454
rect 22654 17378 22706 17390
rect 24894 17442 24946 17454
rect 24894 17378 24946 17390
rect 27358 17442 27410 17454
rect 27358 17378 27410 17390
rect 28254 17442 28306 17454
rect 28254 17378 28306 17390
rect 28478 17442 28530 17454
rect 28478 17378 28530 17390
rect 32734 17442 32786 17454
rect 32734 17378 32786 17390
rect 33966 17442 34018 17454
rect 33966 17378 34018 17390
rect 36094 17442 36146 17454
rect 36094 17378 36146 17390
rect 44046 17442 44098 17454
rect 44046 17378 44098 17390
rect 45390 17442 45442 17454
rect 45390 17378 45442 17390
rect 45726 17442 45778 17454
rect 45726 17378 45778 17390
rect 46286 17442 46338 17454
rect 46286 17378 46338 17390
rect 46734 17442 46786 17454
rect 46734 17378 46786 17390
rect 1344 17274 48608 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 48608 17274
rect 1344 17188 48608 17222
rect 9662 17106 9714 17118
rect 9662 17042 9714 17054
rect 12014 17106 12066 17118
rect 12014 17042 12066 17054
rect 16046 17106 16098 17118
rect 16046 17042 16098 17054
rect 16270 17106 16322 17118
rect 16270 17042 16322 17054
rect 20638 17106 20690 17118
rect 20638 17042 20690 17054
rect 26910 17106 26962 17118
rect 26910 17042 26962 17054
rect 31054 17106 31106 17118
rect 31054 17042 31106 17054
rect 31838 17106 31890 17118
rect 31838 17042 31890 17054
rect 40350 17106 40402 17118
rect 40350 17042 40402 17054
rect 41134 17106 41186 17118
rect 41134 17042 41186 17054
rect 42142 17106 42194 17118
rect 42142 17042 42194 17054
rect 42590 17106 42642 17118
rect 42590 17042 42642 17054
rect 3390 16994 3442 17006
rect 3390 16930 3442 16942
rect 4062 16994 4114 17006
rect 30830 16994 30882 17006
rect 4834 16942 4846 16994
rect 4898 16942 4910 16994
rect 6850 16942 6862 16994
rect 6914 16942 6926 16994
rect 13122 16942 13134 16994
rect 13186 16942 13198 16994
rect 23650 16942 23662 16994
rect 23714 16942 23726 16994
rect 29474 16942 29486 16994
rect 29538 16942 29550 16994
rect 4062 16930 4114 16942
rect 30830 16930 30882 16942
rect 31166 16994 31218 17006
rect 31166 16930 31218 16942
rect 31950 16994 32002 17006
rect 31950 16930 32002 16942
rect 32286 16994 32338 17006
rect 41582 16994 41634 17006
rect 38658 16942 38670 16994
rect 38722 16942 38734 16994
rect 39890 16942 39902 16994
rect 39954 16942 39966 16994
rect 32286 16930 32338 16942
rect 41582 16930 41634 16942
rect 4286 16882 4338 16894
rect 4286 16818 4338 16830
rect 4510 16882 4562 16894
rect 4510 16818 4562 16830
rect 5406 16882 5458 16894
rect 9550 16882 9602 16894
rect 6066 16830 6078 16882
rect 6130 16830 6142 16882
rect 5406 16818 5458 16830
rect 9550 16818 9602 16830
rect 9774 16882 9826 16894
rect 9774 16818 9826 16830
rect 10222 16882 10274 16894
rect 10222 16818 10274 16830
rect 11342 16882 11394 16894
rect 11342 16818 11394 16830
rect 11790 16882 11842 16894
rect 15598 16882 15650 16894
rect 12338 16830 12350 16882
rect 12402 16830 12414 16882
rect 11790 16818 11842 16830
rect 15598 16818 15650 16830
rect 18062 16882 18114 16894
rect 18062 16818 18114 16830
rect 18398 16882 18450 16894
rect 19966 16882 20018 16894
rect 25342 16882 25394 16894
rect 18610 16830 18622 16882
rect 18674 16830 18686 16882
rect 24434 16830 24446 16882
rect 24498 16830 24510 16882
rect 18398 16818 18450 16830
rect 19966 16818 20018 16830
rect 25342 16818 25394 16830
rect 26014 16882 26066 16894
rect 31278 16882 31330 16894
rect 39566 16882 39618 16894
rect 41358 16882 41410 16894
rect 30258 16830 30270 16882
rect 30322 16830 30334 16882
rect 31490 16830 31502 16882
rect 31554 16830 31566 16882
rect 37874 16830 37886 16882
rect 37938 16830 37950 16882
rect 38882 16830 38894 16882
rect 38946 16830 38958 16882
rect 40898 16830 40910 16882
rect 40962 16830 40974 16882
rect 42914 16830 42926 16882
rect 42978 16830 42990 16882
rect 26014 16818 26066 16830
rect 31278 16818 31330 16830
rect 39566 16818 39618 16830
rect 41358 16818 41410 16830
rect 4398 16770 4450 16782
rect 11902 16770 11954 16782
rect 16158 16770 16210 16782
rect 3266 16718 3278 16770
rect 3330 16718 3342 16770
rect 8978 16718 8990 16770
rect 9042 16718 9054 16770
rect 15250 16718 15262 16770
rect 15314 16718 15326 16770
rect 4398 16706 4450 16718
rect 11902 16706 11954 16718
rect 16158 16706 16210 16718
rect 19518 16770 19570 16782
rect 26238 16770 26290 16782
rect 21074 16718 21086 16770
rect 21138 16718 21150 16770
rect 21522 16718 21534 16770
rect 21586 16718 21598 16770
rect 27346 16718 27358 16770
rect 27410 16718 27422 16770
rect 35074 16718 35086 16770
rect 35138 16718 35150 16770
rect 41010 16718 41022 16770
rect 41074 16718 41086 16770
rect 44930 16718 44942 16770
rect 44994 16718 45006 16770
rect 19518 16706 19570 16718
rect 26238 16706 26290 16718
rect 3614 16658 3666 16670
rect 3614 16594 3666 16606
rect 5182 16658 5234 16670
rect 19742 16658 19794 16670
rect 19058 16606 19070 16658
rect 19122 16606 19134 16658
rect 5182 16594 5234 16606
rect 19742 16594 19794 16606
rect 20414 16658 20466 16670
rect 20414 16594 20466 16606
rect 25678 16658 25730 16670
rect 25678 16594 25730 16606
rect 32398 16658 32450 16670
rect 32398 16594 32450 16606
rect 1344 16490 48608 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 48608 16490
rect 1344 16404 48608 16438
rect 10110 16322 10162 16334
rect 9538 16270 9550 16322
rect 9602 16270 9614 16322
rect 34962 16270 34974 16322
rect 35026 16319 35038 16322
rect 35298 16319 35310 16322
rect 35026 16273 35310 16319
rect 35026 16270 35038 16273
rect 35298 16270 35310 16273
rect 35362 16270 35374 16322
rect 10110 16258 10162 16270
rect 4846 16210 4898 16222
rect 3042 16158 3054 16210
rect 3106 16158 3118 16210
rect 4846 16146 4898 16158
rect 5854 16210 5906 16222
rect 5854 16146 5906 16158
rect 8990 16210 9042 16222
rect 8990 16146 9042 16158
rect 9214 16210 9266 16222
rect 9214 16146 9266 16158
rect 11118 16210 11170 16222
rect 12910 16210 12962 16222
rect 23214 16210 23266 16222
rect 29150 16210 29202 16222
rect 12338 16158 12350 16210
rect 12402 16158 12414 16210
rect 19618 16158 19630 16210
rect 19682 16158 19694 16210
rect 21970 16158 21982 16210
rect 22034 16158 22046 16210
rect 28130 16158 28142 16210
rect 28194 16158 28206 16210
rect 11118 16146 11170 16158
rect 12910 16146 12962 16158
rect 23214 16146 23266 16158
rect 29150 16146 29202 16158
rect 29374 16210 29426 16222
rect 29374 16146 29426 16158
rect 29710 16210 29762 16222
rect 29710 16146 29762 16158
rect 30382 16210 30434 16222
rect 34974 16210 35026 16222
rect 30706 16158 30718 16210
rect 30770 16158 30782 16210
rect 32834 16158 32846 16210
rect 32898 16158 32910 16210
rect 30382 16146 30434 16158
rect 34974 16146 35026 16158
rect 35870 16210 35922 16222
rect 35870 16146 35922 16158
rect 36430 16210 36482 16222
rect 37762 16158 37774 16210
rect 37826 16158 37838 16210
rect 39890 16184 39902 16236
rect 39954 16184 39966 16236
rect 41134 16210 41186 16222
rect 44942 16210 44994 16222
rect 41346 16158 41358 16210
rect 41410 16158 41422 16210
rect 43474 16158 43486 16210
rect 43538 16158 43550 16210
rect 45266 16158 45278 16210
rect 45330 16158 45342 16210
rect 47394 16158 47406 16210
rect 47458 16158 47470 16210
rect 36430 16146 36482 16158
rect 41134 16146 41186 16158
rect 44942 16146 44994 16158
rect 3390 16098 3442 16110
rect 3390 16034 3442 16046
rect 3838 16098 3890 16110
rect 3838 16034 3890 16046
rect 4398 16098 4450 16110
rect 9886 16098 9938 16110
rect 12686 16098 12738 16110
rect 6402 16046 6414 16098
rect 6466 16046 6478 16098
rect 11778 16046 11790 16098
rect 11842 16046 11854 16098
rect 4398 16034 4450 16046
rect 9886 16034 9938 16046
rect 12686 16034 12738 16046
rect 13582 16098 13634 16110
rect 13582 16034 13634 16046
rect 14478 16098 14530 16110
rect 14478 16034 14530 16046
rect 15150 16098 15202 16110
rect 15150 16034 15202 16046
rect 18174 16098 18226 16110
rect 18174 16034 18226 16046
rect 18398 16098 18450 16110
rect 21198 16098 21250 16110
rect 19058 16046 19070 16098
rect 19122 16046 19134 16098
rect 19394 16046 19406 16098
rect 19458 16046 19470 16098
rect 18398 16034 18450 16046
rect 21198 16034 21250 16046
rect 21534 16098 21586 16110
rect 23102 16098 23154 16110
rect 22306 16046 22318 16098
rect 22370 16046 22382 16098
rect 21534 16034 21586 16046
rect 23102 16034 23154 16046
rect 23326 16098 23378 16110
rect 23326 16034 23378 16046
rect 23774 16098 23826 16110
rect 23774 16034 23826 16046
rect 24558 16098 24610 16110
rect 28590 16098 28642 16110
rect 35422 16098 35474 16110
rect 25218 16046 25230 16098
rect 25282 16046 25294 16098
rect 33618 16046 33630 16098
rect 33682 16046 33694 16098
rect 24558 16034 24610 16046
rect 28590 16034 28642 16046
rect 35422 16034 35474 16046
rect 35646 16098 35698 16110
rect 37090 16046 37102 16098
rect 37154 16046 37166 16098
rect 44258 16046 44270 16098
rect 44322 16046 44334 16098
rect 48066 16046 48078 16098
rect 48130 16046 48142 16098
rect 35646 16034 35698 16046
rect 3726 15986 3778 15998
rect 12014 15986 12066 15998
rect 14254 15986 14306 15998
rect 6178 15934 6190 15986
rect 6242 15934 6254 15986
rect 13906 15934 13918 15986
rect 13970 15934 13982 15986
rect 3726 15922 3778 15934
rect 12014 15922 12066 15934
rect 14254 15922 14306 15934
rect 14814 15986 14866 15998
rect 14814 15922 14866 15934
rect 20302 15986 20354 15998
rect 20302 15922 20354 15934
rect 20526 15986 20578 15998
rect 20526 15922 20578 15934
rect 21422 15986 21474 15998
rect 28478 15986 28530 15998
rect 26002 15934 26014 15986
rect 26066 15934 26078 15986
rect 21422 15922 21474 15934
rect 28478 15922 28530 15934
rect 34526 15986 34578 15998
rect 34526 15922 34578 15934
rect 35982 15986 36034 15998
rect 40562 15934 40574 15986
rect 40626 15934 40638 15986
rect 35982 15922 36034 15934
rect 3166 15874 3218 15886
rect 3166 15810 3218 15822
rect 3950 15874 4002 15886
rect 14478 15874 14530 15886
rect 17950 15874 18002 15886
rect 10434 15822 10446 15874
rect 10498 15822 10510 15874
rect 15474 15822 15486 15874
rect 15538 15822 15550 15874
rect 3950 15810 4002 15822
rect 14478 15810 14530 15822
rect 17950 15810 18002 15822
rect 18286 15874 18338 15886
rect 20414 15874 20466 15886
rect 19058 15822 19070 15874
rect 19122 15822 19134 15874
rect 18286 15810 18338 15822
rect 20414 15810 20466 15822
rect 23998 15874 24050 15886
rect 23998 15810 24050 15822
rect 29598 15874 29650 15886
rect 29598 15810 29650 15822
rect 29822 15874 29874 15886
rect 29822 15810 29874 15822
rect 30270 15874 30322 15886
rect 30270 15810 30322 15822
rect 33966 15874 34018 15886
rect 33966 15810 34018 15822
rect 40238 15874 40290 15886
rect 40238 15810 40290 15822
rect 44830 15874 44882 15886
rect 44830 15810 44882 15822
rect 1344 15706 48608 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 48608 15706
rect 1344 15620 48608 15654
rect 5742 15538 5794 15550
rect 5742 15474 5794 15486
rect 9550 15538 9602 15550
rect 9550 15474 9602 15486
rect 9774 15538 9826 15550
rect 9774 15474 9826 15486
rect 10670 15538 10722 15550
rect 10670 15474 10722 15486
rect 11342 15538 11394 15550
rect 11342 15474 11394 15486
rect 11790 15538 11842 15550
rect 11790 15474 11842 15486
rect 18398 15538 18450 15550
rect 18398 15474 18450 15486
rect 18846 15538 18898 15550
rect 18846 15474 18898 15486
rect 20974 15538 21026 15550
rect 20974 15474 21026 15486
rect 21870 15538 21922 15550
rect 21870 15474 21922 15486
rect 22878 15538 22930 15550
rect 22878 15474 22930 15486
rect 23438 15538 23490 15550
rect 23438 15474 23490 15486
rect 24110 15538 24162 15550
rect 24110 15474 24162 15486
rect 24446 15538 24498 15550
rect 24446 15474 24498 15486
rect 29038 15538 29090 15550
rect 29038 15474 29090 15486
rect 29262 15538 29314 15550
rect 29262 15474 29314 15486
rect 31614 15538 31666 15550
rect 31614 15474 31666 15486
rect 31838 15538 31890 15550
rect 31838 15474 31890 15486
rect 33854 15538 33906 15550
rect 33854 15474 33906 15486
rect 35422 15538 35474 15550
rect 35422 15474 35474 15486
rect 36542 15538 36594 15550
rect 36542 15474 36594 15486
rect 39118 15538 39170 15550
rect 39118 15474 39170 15486
rect 40014 15538 40066 15550
rect 40014 15474 40066 15486
rect 19966 15426 20018 15438
rect 2482 15374 2494 15426
rect 2546 15374 2558 15426
rect 15698 15374 15710 15426
rect 15762 15374 15774 15426
rect 19730 15374 19742 15426
rect 19794 15374 19806 15426
rect 19966 15362 20018 15374
rect 20750 15426 20802 15438
rect 20750 15362 20802 15374
rect 26126 15426 26178 15438
rect 26126 15362 26178 15374
rect 26910 15426 26962 15438
rect 26910 15362 26962 15374
rect 27022 15426 27074 15438
rect 27022 15362 27074 15374
rect 27134 15426 27186 15438
rect 27134 15362 27186 15374
rect 28702 15426 28754 15438
rect 28702 15362 28754 15374
rect 29374 15426 29426 15438
rect 29374 15362 29426 15374
rect 31278 15426 31330 15438
rect 31278 15362 31330 15374
rect 31726 15426 31778 15438
rect 36094 15426 36146 15438
rect 33506 15374 33518 15426
rect 33570 15374 33582 15426
rect 35074 15374 35086 15426
rect 35138 15374 35150 15426
rect 31726 15362 31778 15374
rect 36094 15362 36146 15374
rect 36990 15426 37042 15438
rect 36990 15362 37042 15374
rect 38334 15426 38386 15438
rect 47394 15374 47406 15426
rect 47458 15374 47470 15426
rect 38334 15362 38386 15374
rect 10222 15314 10274 15326
rect 1810 15262 1822 15314
rect 1874 15262 1886 15314
rect 5506 15262 5518 15314
rect 5570 15262 5582 15314
rect 6066 15262 6078 15314
rect 6130 15262 6142 15314
rect 6850 15262 6862 15314
rect 6914 15262 6926 15314
rect 10222 15250 10274 15262
rect 10558 15314 10610 15326
rect 10558 15250 10610 15262
rect 11566 15314 11618 15326
rect 20190 15314 20242 15326
rect 16370 15262 16382 15314
rect 16434 15262 16446 15314
rect 19506 15262 19518 15314
rect 19570 15262 19582 15314
rect 11566 15250 11618 15262
rect 20190 15250 20242 15262
rect 20638 15314 20690 15326
rect 22430 15314 22482 15326
rect 21186 15262 21198 15314
rect 21250 15262 21262 15314
rect 20638 15250 20690 15262
rect 22430 15250 22482 15262
rect 23550 15314 23602 15326
rect 26014 15314 26066 15326
rect 25554 15262 25566 15314
rect 25618 15262 25630 15314
rect 23550 15250 23602 15262
rect 26014 15250 26066 15262
rect 27694 15314 27746 15326
rect 27694 15250 27746 15262
rect 27918 15314 27970 15326
rect 28590 15314 28642 15326
rect 28130 15262 28142 15314
rect 28194 15262 28206 15314
rect 27918 15250 27970 15262
rect 28590 15250 28642 15262
rect 30046 15314 30098 15326
rect 30046 15250 30098 15262
rect 30606 15314 30658 15326
rect 30606 15250 30658 15262
rect 31502 15314 31554 15326
rect 31502 15250 31554 15262
rect 34190 15314 34242 15326
rect 34190 15250 34242 15262
rect 34750 15314 34802 15326
rect 35858 15262 35870 15314
rect 35922 15262 35934 15314
rect 37426 15262 37438 15314
rect 37490 15262 37502 15314
rect 38546 15262 38558 15314
rect 38610 15262 38622 15314
rect 43810 15262 43822 15314
rect 43874 15262 43886 15314
rect 48066 15262 48078 15314
rect 48130 15262 48142 15314
rect 34750 15250 34802 15262
rect 9662 15202 9714 15214
rect 4610 15150 4622 15202
rect 4674 15150 4686 15202
rect 8978 15150 8990 15202
rect 9042 15150 9054 15202
rect 9662 15138 9714 15150
rect 10446 15202 10498 15214
rect 10446 15138 10498 15150
rect 11678 15202 11730 15214
rect 18734 15202 18786 15214
rect 13570 15150 13582 15202
rect 13634 15150 13646 15202
rect 11678 15138 11730 15150
rect 18734 15138 18786 15150
rect 20862 15202 20914 15214
rect 20862 15138 20914 15150
rect 25790 15202 25842 15214
rect 28478 15202 28530 15214
rect 39566 15202 39618 15214
rect 44718 15202 44770 15214
rect 26450 15150 26462 15202
rect 26514 15150 26526 15202
rect 37762 15150 37774 15202
rect 37826 15150 37838 15202
rect 40898 15150 40910 15202
rect 40962 15150 40974 15202
rect 43026 15150 43038 15202
rect 43090 15150 43102 15202
rect 45266 15150 45278 15202
rect 45330 15150 45342 15202
rect 25790 15138 25842 15150
rect 28478 15138 28530 15150
rect 39566 15138 39618 15150
rect 44718 15138 44770 15150
rect 19182 15090 19234 15102
rect 19182 15026 19234 15038
rect 23438 15090 23490 15102
rect 23438 15026 23490 15038
rect 27582 15090 27634 15102
rect 27582 15026 27634 15038
rect 39454 15090 39506 15102
rect 39454 15026 39506 15038
rect 44606 15090 44658 15102
rect 44606 15026 44658 15038
rect 1344 14922 48608 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 48608 14922
rect 1344 14836 48608 14870
rect 3838 14754 3890 14766
rect 3490 14702 3502 14754
rect 3554 14702 3566 14754
rect 3838 14690 3890 14702
rect 11790 14754 11842 14766
rect 11790 14690 11842 14702
rect 19630 14754 19682 14766
rect 19630 14690 19682 14702
rect 28254 14754 28306 14766
rect 28254 14690 28306 14702
rect 4062 14642 4114 14654
rect 14926 14642 14978 14654
rect 24670 14642 24722 14654
rect 34750 14642 34802 14654
rect 6066 14590 6078 14642
rect 6130 14590 6142 14642
rect 18722 14590 18734 14642
rect 18786 14590 18798 14642
rect 21298 14590 21310 14642
rect 21362 14590 21374 14642
rect 23426 14590 23438 14642
rect 23490 14590 23502 14642
rect 24994 14590 25006 14642
rect 25058 14590 25070 14642
rect 27122 14590 27134 14642
rect 27186 14590 27198 14642
rect 29698 14590 29710 14642
rect 29762 14590 29774 14642
rect 4062 14578 4114 14590
rect 14926 14578 14978 14590
rect 24670 14578 24722 14590
rect 34750 14578 34802 14590
rect 38222 14642 38274 14654
rect 38222 14578 38274 14590
rect 42590 14642 42642 14654
rect 43362 14590 43374 14642
rect 43426 14590 43438 14642
rect 45714 14590 45726 14642
rect 45778 14590 45790 14642
rect 42590 14578 42642 14590
rect 4398 14530 4450 14542
rect 11566 14530 11618 14542
rect 10882 14478 10894 14530
rect 10946 14478 10958 14530
rect 4398 14466 4450 14478
rect 11566 14466 11618 14478
rect 15038 14530 15090 14542
rect 15038 14466 15090 14478
rect 15486 14530 15538 14542
rect 19854 14530 19906 14542
rect 35870 14530 35922 14542
rect 15922 14478 15934 14530
rect 15986 14478 15998 14530
rect 19394 14478 19406 14530
rect 19458 14478 19470 14530
rect 24098 14478 24110 14530
rect 24162 14478 24174 14530
rect 27794 14478 27806 14530
rect 27858 14478 27870 14530
rect 29362 14478 29374 14530
rect 29426 14478 29438 14530
rect 30594 14478 30606 14530
rect 30658 14478 30670 14530
rect 35298 14478 35310 14530
rect 35362 14478 35374 14530
rect 15486 14466 15538 14478
rect 19854 14466 19906 14478
rect 35870 14466 35922 14478
rect 36542 14530 36594 14542
rect 36542 14466 36594 14478
rect 37214 14530 37266 14542
rect 37214 14466 37266 14478
rect 37998 14530 38050 14542
rect 39006 14530 39058 14542
rect 39902 14530 39954 14542
rect 38322 14478 38334 14530
rect 38386 14478 38398 14530
rect 39330 14478 39342 14530
rect 39394 14478 39406 14530
rect 37998 14466 38050 14478
rect 39006 14466 39058 14478
rect 39902 14466 39954 14478
rect 40238 14530 40290 14542
rect 40238 14466 40290 14478
rect 40462 14530 40514 14542
rect 43150 14530 43202 14542
rect 42914 14478 42926 14530
rect 42978 14478 42990 14530
rect 40462 14466 40514 14478
rect 43150 14466 43202 14478
rect 43486 14530 43538 14542
rect 43486 14466 43538 14478
rect 45278 14530 45330 14542
rect 45278 14466 45330 14478
rect 45390 14530 45442 14542
rect 45390 14466 45442 14478
rect 45614 14530 45666 14542
rect 45614 14466 45666 14478
rect 46958 14530 47010 14542
rect 46958 14466 47010 14478
rect 4846 14418 4898 14430
rect 12574 14418 12626 14430
rect 12114 14366 12126 14418
rect 12178 14366 12190 14418
rect 4846 14354 4898 14366
rect 12574 14354 12626 14366
rect 13470 14418 13522 14430
rect 13470 14354 13522 14366
rect 13582 14418 13634 14430
rect 13582 14354 13634 14366
rect 14814 14418 14866 14430
rect 20302 14418 20354 14430
rect 30158 14418 30210 14430
rect 16594 14366 16606 14418
rect 16658 14366 16670 14418
rect 19170 14415 19182 14418
rect 18961 14369 19182 14415
rect 14814 14354 14866 14366
rect 4510 14306 4562 14318
rect 4510 14242 4562 14254
rect 4622 14306 4674 14318
rect 12910 14306 12962 14318
rect 10882 14254 10894 14306
rect 10946 14303 10958 14306
rect 11330 14303 11342 14306
rect 10946 14257 11342 14303
rect 10946 14254 10958 14257
rect 11330 14254 11342 14257
rect 11394 14254 11406 14306
rect 4622 14242 4674 14254
rect 12910 14242 12962 14254
rect 13806 14306 13858 14318
rect 18961 14306 19007 14369
rect 19170 14366 19182 14369
rect 19234 14415 19246 14418
rect 19394 14415 19406 14418
rect 19234 14369 19406 14415
rect 19234 14366 19246 14369
rect 19394 14366 19406 14369
rect 19458 14366 19470 14418
rect 29474 14366 29486 14418
rect 29538 14366 29550 14418
rect 20302 14354 20354 14366
rect 30158 14354 30210 14366
rect 35982 14418 36034 14430
rect 35982 14354 36034 14366
rect 37102 14418 37154 14430
rect 37102 14354 37154 14366
rect 37326 14418 37378 14430
rect 41134 14418 41186 14430
rect 40786 14366 40798 14418
rect 40850 14366 40862 14418
rect 37326 14354 37378 14366
rect 41134 14354 41186 14366
rect 41470 14418 41522 14430
rect 41470 14354 41522 14366
rect 43934 14418 43986 14430
rect 43934 14354 43986 14366
rect 46174 14418 46226 14430
rect 46174 14354 46226 14366
rect 19518 14306 19570 14318
rect 18946 14254 18958 14306
rect 19010 14254 19022 14306
rect 13806 14242 13858 14254
rect 19518 14242 19570 14254
rect 20414 14306 20466 14318
rect 20414 14242 20466 14254
rect 20526 14306 20578 14318
rect 20526 14242 20578 14254
rect 28366 14306 28418 14318
rect 28366 14242 28418 14254
rect 28478 14306 28530 14318
rect 36094 14306 36146 14318
rect 38558 14306 38610 14318
rect 35074 14254 35086 14306
rect 35138 14254 35150 14306
rect 37762 14254 37774 14306
rect 37826 14254 37838 14306
rect 28478 14242 28530 14254
rect 36094 14242 36146 14254
rect 38558 14242 38610 14254
rect 42030 14306 42082 14318
rect 42030 14242 42082 14254
rect 43374 14306 43426 14318
rect 43374 14242 43426 14254
rect 44046 14306 44098 14318
rect 44046 14242 44098 14254
rect 44270 14306 44322 14318
rect 44270 14242 44322 14254
rect 45726 14306 45778 14318
rect 45726 14242 45778 14254
rect 46510 14306 46562 14318
rect 46510 14242 46562 14254
rect 1344 14138 48608 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 48608 14138
rect 1344 14052 48608 14086
rect 15710 13970 15762 13982
rect 27470 13970 27522 13982
rect 6514 13918 6526 13970
rect 6578 13918 6590 13970
rect 10882 13918 10894 13970
rect 10946 13918 10958 13970
rect 18386 13918 18398 13970
rect 18450 13918 18462 13970
rect 25890 13918 25902 13970
rect 25954 13918 25966 13970
rect 15710 13906 15762 13918
rect 27470 13906 27522 13918
rect 28030 13970 28082 13982
rect 28030 13906 28082 13918
rect 28366 13970 28418 13982
rect 28366 13906 28418 13918
rect 28702 13970 28754 13982
rect 28702 13906 28754 13918
rect 31950 13970 32002 13982
rect 31950 13906 32002 13918
rect 41022 13970 41074 13982
rect 41022 13906 41074 13918
rect 42590 13970 42642 13982
rect 44482 13918 44494 13970
rect 44546 13918 44558 13970
rect 42590 13906 42642 13918
rect 11902 13858 11954 13870
rect 11902 13794 11954 13806
rect 14030 13858 14082 13870
rect 14030 13794 14082 13806
rect 17950 13858 18002 13870
rect 17950 13794 18002 13806
rect 18958 13858 19010 13870
rect 27806 13858 27858 13870
rect 21746 13806 21758 13858
rect 21810 13806 21822 13858
rect 18958 13794 19010 13806
rect 27806 13794 27858 13806
rect 28254 13858 28306 13870
rect 39454 13858 39506 13870
rect 29922 13806 29934 13858
rect 29986 13806 29998 13858
rect 30594 13806 30606 13858
rect 30658 13806 30670 13858
rect 36306 13806 36318 13858
rect 36370 13806 36382 13858
rect 39218 13806 39230 13858
rect 39282 13806 39294 13858
rect 47394 13806 47406 13858
rect 47458 13806 47470 13858
rect 28254 13794 28306 13806
rect 39454 13794 39506 13806
rect 4958 13746 5010 13758
rect 1810 13694 1822 13746
rect 1874 13694 1886 13746
rect 4958 13682 5010 13694
rect 5182 13746 5234 13758
rect 5182 13682 5234 13694
rect 7086 13746 7138 13758
rect 7086 13682 7138 13694
rect 7534 13746 7586 13758
rect 7534 13682 7586 13694
rect 10222 13746 10274 13758
rect 10222 13682 10274 13694
rect 11230 13746 11282 13758
rect 14142 13746 14194 13758
rect 12226 13694 12238 13746
rect 12290 13694 12302 13746
rect 11230 13682 11282 13694
rect 14142 13682 14194 13694
rect 14590 13746 14642 13758
rect 14590 13682 14642 13694
rect 17838 13746 17890 13758
rect 26238 13746 26290 13758
rect 23874 13694 23886 13746
rect 23938 13694 23950 13746
rect 17838 13682 17890 13694
rect 26238 13682 26290 13694
rect 26462 13746 26514 13758
rect 26462 13682 26514 13694
rect 27694 13746 27746 13758
rect 27694 13682 27746 13694
rect 28590 13746 28642 13758
rect 31614 13746 31666 13758
rect 28802 13694 28814 13746
rect 28866 13694 28878 13746
rect 30146 13694 30158 13746
rect 30210 13694 30222 13746
rect 30706 13694 30718 13746
rect 30770 13694 30782 13746
rect 31378 13694 31390 13746
rect 31442 13694 31454 13746
rect 28590 13682 28642 13694
rect 31614 13682 31666 13694
rect 31838 13746 31890 13758
rect 31838 13682 31890 13694
rect 33182 13746 33234 13758
rect 39118 13746 39170 13758
rect 42814 13746 42866 13758
rect 35522 13694 35534 13746
rect 35586 13694 35598 13746
rect 39666 13694 39678 13746
rect 39730 13694 39742 13746
rect 33182 13682 33234 13694
rect 39118 13682 39170 13694
rect 42814 13682 42866 13694
rect 43822 13746 43874 13758
rect 43822 13682 43874 13694
rect 43934 13746 43986 13758
rect 43934 13682 43986 13694
rect 44046 13746 44098 13758
rect 48066 13694 48078 13746
rect 48130 13694 48142 13746
rect 44046 13682 44098 13694
rect 12014 13634 12066 13646
rect 2482 13582 2494 13634
rect 2546 13582 2558 13634
rect 4610 13582 4622 13634
rect 4674 13582 4686 13634
rect 12014 13570 12066 13582
rect 13806 13634 13858 13646
rect 13806 13570 13858 13582
rect 25342 13634 25394 13646
rect 25342 13570 25394 13582
rect 31726 13634 31778 13646
rect 31726 13570 31778 13582
rect 32398 13634 32450 13646
rect 32398 13570 32450 13582
rect 34302 13634 34354 13646
rect 40126 13634 40178 13646
rect 38434 13582 38446 13634
rect 38498 13582 38510 13634
rect 34302 13570 34354 13582
rect 40126 13570 40178 13582
rect 41694 13634 41746 13646
rect 41694 13570 41746 13582
rect 43038 13634 43090 13646
rect 43038 13570 43090 13582
rect 43374 13634 43426 13646
rect 45266 13582 45278 13634
rect 45330 13582 45342 13634
rect 43374 13570 43426 13582
rect 6862 13522 6914 13534
rect 5506 13470 5518 13522
rect 5570 13470 5582 13522
rect 6862 13458 6914 13470
rect 10334 13522 10386 13534
rect 10334 13458 10386 13470
rect 14814 13522 14866 13534
rect 14814 13458 14866 13470
rect 17950 13522 18002 13534
rect 17950 13458 18002 13470
rect 18734 13522 18786 13534
rect 18734 13458 18786 13470
rect 32510 13522 32562 13534
rect 32510 13458 32562 13470
rect 34190 13522 34242 13534
rect 34190 13458 34242 13470
rect 1344 13354 48608 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 48608 13354
rect 1344 13268 48608 13302
rect 3726 13186 3778 13198
rect 3726 13122 3778 13134
rect 4062 13186 4114 13198
rect 4062 13122 4114 13134
rect 38110 13186 38162 13198
rect 38110 13122 38162 13134
rect 7086 13074 7138 13086
rect 7086 13010 7138 13022
rect 7758 13074 7810 13086
rect 12126 13074 12178 13086
rect 16270 13074 16322 13086
rect 21310 13074 21362 13086
rect 9090 13022 9102 13074
rect 9154 13022 9166 13074
rect 11218 13022 11230 13074
rect 11282 13022 11294 13074
rect 13682 13022 13694 13074
rect 13746 13022 13758 13074
rect 15138 13022 15150 13074
rect 15202 13022 15214 13074
rect 18722 13022 18734 13074
rect 18786 13022 18798 13074
rect 7758 13010 7810 13022
rect 12126 13010 12178 13022
rect 16270 13010 16322 13022
rect 21310 13010 21362 13022
rect 22430 13074 22482 13086
rect 23774 13074 23826 13086
rect 23314 13022 23326 13074
rect 23378 13022 23390 13074
rect 22430 13010 22482 13022
rect 23774 13010 23826 13022
rect 29374 13074 29426 13086
rect 29374 13010 29426 13022
rect 29710 13074 29762 13086
rect 38894 13074 38946 13086
rect 31042 13022 31054 13074
rect 31106 13022 31118 13074
rect 33170 13022 33182 13074
rect 33234 13022 33246 13074
rect 34402 13022 34414 13074
rect 34466 13022 34478 13074
rect 29710 13010 29762 13022
rect 38894 13010 38946 13022
rect 40462 13074 40514 13086
rect 40462 13010 40514 13022
rect 6302 12962 6354 12974
rect 6302 12898 6354 12910
rect 6750 12962 6802 12974
rect 6750 12898 6802 12910
rect 6862 12962 6914 12974
rect 17726 12962 17778 12974
rect 8306 12910 8318 12962
rect 8370 12910 8382 12962
rect 11666 12910 11678 12962
rect 11730 12910 11742 12962
rect 12674 12910 12686 12962
rect 12738 12910 12750 12962
rect 14018 12910 14030 12962
rect 14082 12910 14094 12962
rect 6862 12898 6914 12910
rect 17726 12898 17778 12910
rect 17950 12962 18002 12974
rect 17950 12898 18002 12910
rect 18286 12962 18338 12974
rect 20302 12962 20354 12974
rect 26014 12962 26066 12974
rect 18946 12910 18958 12962
rect 19010 12910 19022 12962
rect 19842 12910 19854 12962
rect 19906 12910 19918 12962
rect 23090 12910 23102 12962
rect 23154 12910 23166 12962
rect 24322 12910 24334 12962
rect 24386 12910 24398 12962
rect 18286 12898 18338 12910
rect 20302 12898 20354 12910
rect 26014 12898 26066 12910
rect 26238 12962 26290 12974
rect 26238 12898 26290 12910
rect 26574 12962 26626 12974
rect 26574 12898 26626 12910
rect 29150 12962 29202 12974
rect 34750 12962 34802 12974
rect 33842 12910 33854 12962
rect 33906 12910 33918 12962
rect 29150 12898 29202 12910
rect 34750 12898 34802 12910
rect 38222 12962 38274 12974
rect 38222 12898 38274 12910
rect 40574 12962 40626 12974
rect 44270 12962 44322 12974
rect 41906 12910 41918 12962
rect 41970 12910 41982 12962
rect 42466 12910 42478 12962
rect 42530 12910 42542 12962
rect 42690 12910 42702 12962
rect 42754 12910 42766 12962
rect 43586 12910 43598 12962
rect 43650 12910 43662 12962
rect 44034 12910 44046 12962
rect 44098 12910 44110 12962
rect 40574 12898 40626 12910
rect 44270 12898 44322 12910
rect 45166 12962 45218 12974
rect 45166 12898 45218 12910
rect 45390 12962 45442 12974
rect 45390 12898 45442 12910
rect 3838 12850 3890 12862
rect 3838 12786 3890 12798
rect 4734 12850 4786 12862
rect 4734 12786 4786 12798
rect 5070 12850 5122 12862
rect 5070 12786 5122 12798
rect 5630 12850 5682 12862
rect 5630 12786 5682 12798
rect 7198 12850 7250 12862
rect 7198 12786 7250 12798
rect 14478 12850 14530 12862
rect 14478 12786 14530 12798
rect 14814 12850 14866 12862
rect 14814 12786 14866 12798
rect 15038 12850 15090 12862
rect 15038 12786 15090 12798
rect 18174 12850 18226 12862
rect 26910 12850 26962 12862
rect 19058 12798 19070 12850
rect 19122 12798 19134 12850
rect 18174 12786 18226 12798
rect 26910 12786 26962 12798
rect 27022 12850 27074 12862
rect 27022 12786 27074 12798
rect 34974 12850 35026 12862
rect 34974 12786 35026 12798
rect 40014 12850 40066 12862
rect 46062 12850 46114 12862
rect 45714 12798 45726 12850
rect 45778 12798 45790 12850
rect 47842 12798 47854 12850
rect 47906 12798 47918 12850
rect 40014 12786 40066 12798
rect 46062 12786 46114 12798
rect 5742 12738 5794 12750
rect 5742 12674 5794 12686
rect 5854 12738 5906 12750
rect 15598 12738 15650 12750
rect 12450 12686 12462 12738
rect 12514 12686 12526 12738
rect 5854 12674 5906 12686
rect 15598 12674 15650 12686
rect 17614 12738 17666 12750
rect 17614 12674 17666 12686
rect 20862 12738 20914 12750
rect 20862 12674 20914 12686
rect 21870 12738 21922 12750
rect 21870 12674 21922 12686
rect 24110 12738 24162 12750
rect 24110 12674 24162 12686
rect 25454 12738 25506 12750
rect 25454 12674 25506 12686
rect 25678 12738 25730 12750
rect 25678 12674 25730 12686
rect 25902 12738 25954 12750
rect 25902 12674 25954 12686
rect 26462 12738 26514 12750
rect 26462 12674 26514 12686
rect 29598 12738 29650 12750
rect 29598 12674 29650 12686
rect 29822 12738 29874 12750
rect 29822 12674 29874 12686
rect 34414 12738 34466 12750
rect 34414 12674 34466 12686
rect 34526 12738 34578 12750
rect 34526 12674 34578 12686
rect 40126 12738 40178 12750
rect 40126 12674 40178 12686
rect 42142 12738 42194 12750
rect 42142 12674 42194 12686
rect 42926 12738 42978 12750
rect 42926 12674 42978 12686
rect 43038 12738 43090 12750
rect 43038 12674 43090 12686
rect 46398 12738 46450 12750
rect 46398 12674 46450 12686
rect 47630 12738 47682 12750
rect 47630 12674 47682 12686
rect 48190 12738 48242 12750
rect 48190 12674 48242 12686
rect 1344 12570 48608 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 48608 12570
rect 1344 12484 48608 12518
rect 5294 12402 5346 12414
rect 5294 12338 5346 12350
rect 9886 12402 9938 12414
rect 9886 12338 9938 12350
rect 11342 12402 11394 12414
rect 11342 12338 11394 12350
rect 16718 12402 16770 12414
rect 16718 12338 16770 12350
rect 31166 12402 31218 12414
rect 31166 12338 31218 12350
rect 31390 12402 31442 12414
rect 31390 12338 31442 12350
rect 32062 12402 32114 12414
rect 32062 12338 32114 12350
rect 41134 12402 41186 12414
rect 41134 12338 41186 12350
rect 41358 12402 41410 12414
rect 42242 12350 42254 12402
rect 42306 12350 42318 12402
rect 42466 12350 42478 12402
rect 42530 12350 42542 12402
rect 41358 12338 41410 12350
rect 5406 12290 5458 12302
rect 11678 12290 11730 12302
rect 8082 12238 8094 12290
rect 8146 12238 8158 12290
rect 9538 12238 9550 12290
rect 9602 12238 9614 12290
rect 5406 12226 5458 12238
rect 11678 12226 11730 12238
rect 12014 12290 12066 12302
rect 17614 12290 17666 12302
rect 15474 12238 15486 12290
rect 15538 12238 15550 12290
rect 12014 12226 12066 12238
rect 17614 12226 17666 12238
rect 17950 12290 18002 12302
rect 25790 12290 25842 12302
rect 22530 12238 22542 12290
rect 22594 12238 22606 12290
rect 17950 12226 18002 12238
rect 25790 12226 25842 12238
rect 26686 12290 26738 12302
rect 26686 12226 26738 12238
rect 29038 12290 29090 12302
rect 29038 12226 29090 12238
rect 31278 12290 31330 12302
rect 31278 12226 31330 12238
rect 40126 12290 40178 12302
rect 43586 12238 43598 12290
rect 43650 12238 43662 12290
rect 47394 12238 47406 12290
rect 47458 12238 47470 12290
rect 40126 12226 40178 12238
rect 4958 12178 5010 12190
rect 1810 12126 1822 12178
rect 1874 12126 1886 12178
rect 4958 12114 5010 12126
rect 5630 12178 5682 12190
rect 10782 12178 10834 12190
rect 8754 12126 8766 12178
rect 8818 12126 8830 12178
rect 10322 12126 10334 12178
rect 10386 12126 10398 12178
rect 5630 12114 5682 12126
rect 10782 12114 10834 12126
rect 12350 12178 12402 12190
rect 16606 12178 16658 12190
rect 16258 12126 16270 12178
rect 16322 12126 16334 12178
rect 12350 12114 12402 12126
rect 16606 12114 16658 12126
rect 16942 12178 16994 12190
rect 16942 12114 16994 12126
rect 17390 12178 17442 12190
rect 25566 12178 25618 12190
rect 21410 12126 21422 12178
rect 21474 12126 21486 12178
rect 21746 12126 21758 12178
rect 21810 12126 21822 12178
rect 17390 12114 17442 12126
rect 25566 12114 25618 12126
rect 26238 12178 26290 12190
rect 26238 12114 26290 12126
rect 26798 12178 26850 12190
rect 26798 12114 26850 12126
rect 30382 12178 30434 12190
rect 37326 12178 37378 12190
rect 30930 12126 30942 12178
rect 30994 12126 31006 12178
rect 31602 12126 31614 12178
rect 31666 12126 31678 12178
rect 33282 12126 33294 12178
rect 33346 12126 33358 12178
rect 34066 12126 34078 12178
rect 34130 12126 34142 12178
rect 30382 12114 30434 12126
rect 37326 12114 37378 12126
rect 37774 12178 37826 12190
rect 37774 12114 37826 12126
rect 37998 12178 38050 12190
rect 39230 12178 39282 12190
rect 38994 12126 39006 12178
rect 39058 12126 39070 12178
rect 37998 12114 38050 12126
rect 39230 12114 39282 12126
rect 39454 12178 39506 12190
rect 40014 12178 40066 12190
rect 43934 12178 43986 12190
rect 39666 12126 39678 12178
rect 39730 12126 39742 12178
rect 40898 12126 40910 12178
rect 40962 12126 40974 12178
rect 41570 12126 41582 12178
rect 41634 12126 41646 12178
rect 42690 12126 42702 12178
rect 42754 12126 42766 12178
rect 43474 12126 43486 12178
rect 43538 12126 43550 12178
rect 39454 12114 39506 12126
rect 40014 12114 40066 12126
rect 43934 12114 43986 12126
rect 44158 12178 44210 12190
rect 48066 12126 48078 12178
rect 48130 12126 48142 12178
rect 44158 12114 44210 12126
rect 12798 12066 12850 12078
rect 17838 12066 17890 12078
rect 26462 12066 26514 12078
rect 2482 12014 2494 12066
rect 2546 12014 2558 12066
rect 4610 12014 4622 12066
rect 4674 12014 4686 12066
rect 5954 12014 5966 12066
rect 6018 12014 6030 12066
rect 13346 12014 13358 12066
rect 13410 12014 13422 12066
rect 18498 12014 18510 12066
rect 18562 12014 18574 12066
rect 20626 12014 20638 12066
rect 20690 12014 20702 12066
rect 24658 12014 24670 12066
rect 24722 12014 24734 12066
rect 12798 12002 12850 12014
rect 17838 12002 17890 12014
rect 26462 12002 26514 12014
rect 28926 12066 28978 12078
rect 36654 12066 36706 12078
rect 36194 12014 36206 12066
rect 36258 12014 36270 12066
rect 28926 12002 28978 12014
rect 36654 12002 36706 12014
rect 37550 12066 37602 12078
rect 37550 12002 37602 12014
rect 37886 12066 37938 12078
rect 37886 12002 37938 12014
rect 39342 12066 39394 12078
rect 44942 12066 44994 12078
rect 41010 12014 41022 12066
rect 41074 12014 41086 12066
rect 45266 12014 45278 12066
rect 45330 12014 45342 12066
rect 39342 12002 39394 12014
rect 44942 12002 44994 12014
rect 25230 11954 25282 11966
rect 25230 11890 25282 11902
rect 30494 11954 30546 11966
rect 30494 11890 30546 11902
rect 36542 11954 36594 11966
rect 44482 11902 44494 11954
rect 44546 11902 44558 11954
rect 36542 11890 36594 11902
rect 1344 11786 48608 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 48608 11786
rect 1344 11700 48608 11734
rect 3614 11618 3666 11630
rect 24110 11618 24162 11630
rect 6402 11566 6414 11618
rect 6466 11566 6478 11618
rect 3614 11554 3666 11566
rect 24110 11554 24162 11566
rect 42254 11618 42306 11630
rect 42254 11554 42306 11566
rect 43822 11618 43874 11630
rect 43822 11554 43874 11566
rect 45054 11618 45106 11630
rect 45054 11554 45106 11566
rect 4398 11506 4450 11518
rect 29598 11506 29650 11518
rect 10210 11454 10222 11506
rect 10274 11454 10286 11506
rect 16706 11454 16718 11506
rect 16770 11454 16782 11506
rect 18834 11454 18846 11506
rect 18898 11454 18910 11506
rect 22194 11454 22206 11506
rect 22258 11454 22270 11506
rect 26450 11454 26462 11506
rect 26514 11454 26526 11506
rect 28578 11454 28590 11506
rect 28642 11454 28654 11506
rect 4398 11442 4450 11454
rect 29598 11442 29650 11454
rect 30270 11506 30322 11518
rect 30270 11442 30322 11454
rect 42142 11506 42194 11518
rect 42142 11442 42194 11454
rect 3390 11394 3442 11406
rect 3390 11330 3442 11342
rect 4286 11394 4338 11406
rect 4286 11330 4338 11342
rect 4622 11394 4674 11406
rect 4622 11330 4674 11342
rect 4846 11394 4898 11406
rect 5854 11394 5906 11406
rect 5618 11342 5630 11394
rect 5682 11342 5694 11394
rect 4846 11330 4898 11342
rect 5854 11330 5906 11342
rect 5966 11394 6018 11406
rect 10894 11394 10946 11406
rect 7298 11342 7310 11394
rect 7362 11342 7374 11394
rect 5966 11330 6018 11342
rect 10894 11330 10946 11342
rect 11118 11394 11170 11406
rect 11118 11330 11170 11342
rect 12126 11394 12178 11406
rect 23214 11394 23266 11406
rect 15362 11342 15374 11394
rect 15426 11342 15438 11394
rect 16034 11342 16046 11394
rect 16098 11342 16110 11394
rect 21858 11342 21870 11394
rect 21922 11342 21934 11394
rect 12126 11330 12178 11342
rect 23214 11330 23266 11342
rect 23326 11394 23378 11406
rect 23326 11330 23378 11342
rect 23438 11394 23490 11406
rect 30494 11394 30546 11406
rect 36990 11394 37042 11406
rect 40798 11394 40850 11406
rect 23762 11342 23774 11394
rect 23826 11342 23838 11394
rect 25778 11342 25790 11394
rect 25842 11342 25854 11394
rect 36418 11342 36430 11394
rect 36482 11342 36494 11394
rect 37762 11342 37774 11394
rect 37826 11342 37838 11394
rect 38434 11342 38446 11394
rect 38498 11342 38510 11394
rect 39330 11342 39342 11394
rect 39394 11342 39406 11394
rect 23438 11330 23490 11342
rect 30494 11330 30546 11342
rect 36990 11330 37042 11342
rect 40798 11330 40850 11342
rect 42702 11394 42754 11406
rect 42702 11330 42754 11342
rect 42814 11394 42866 11406
rect 45278 11394 45330 11406
rect 43138 11342 43150 11394
rect 43202 11342 43214 11394
rect 44818 11342 44830 11394
rect 44882 11342 44894 11394
rect 42814 11330 42866 11342
rect 45278 11330 45330 11342
rect 45502 11394 45554 11406
rect 45502 11330 45554 11342
rect 46734 11394 46786 11406
rect 46734 11330 46786 11342
rect 11566 11282 11618 11294
rect 8082 11230 8094 11282
rect 8146 11230 8158 11282
rect 11566 11218 11618 11230
rect 11678 11282 11730 11294
rect 11678 11218 11730 11230
rect 12238 11282 12290 11294
rect 29934 11282 29986 11294
rect 37102 11282 37154 11294
rect 40238 11282 40290 11294
rect 43934 11282 43986 11294
rect 15586 11230 15598 11282
rect 15650 11230 15662 11282
rect 31938 11230 31950 11282
rect 32002 11230 32014 11282
rect 37650 11230 37662 11282
rect 37714 11230 37726 11282
rect 38658 11230 38670 11282
rect 38722 11230 38734 11282
rect 43026 11230 43038 11282
rect 43090 11230 43102 11282
rect 12238 11218 12290 11230
rect 29934 11218 29986 11230
rect 37102 11218 37154 11230
rect 40238 11218 40290 11230
rect 43934 11218 43986 11230
rect 45614 11282 45666 11294
rect 45614 11218 45666 11230
rect 45950 11282 46002 11294
rect 45950 11218 46002 11230
rect 10670 11170 10722 11182
rect 3938 11118 3950 11170
rect 4002 11118 4014 11170
rect 10670 11106 10722 11118
rect 11006 11170 11058 11182
rect 11006 11106 11058 11118
rect 11902 11170 11954 11182
rect 11902 11106 11954 11118
rect 12350 11170 12402 11182
rect 12350 11106 12402 11118
rect 12574 11170 12626 11182
rect 12574 11106 12626 11118
rect 22766 11170 22818 11182
rect 37326 11170 37378 11182
rect 40126 11170 40178 11182
rect 30818 11118 30830 11170
rect 30882 11118 30894 11170
rect 38210 11118 38222 11170
rect 38274 11118 38286 11170
rect 22766 11106 22818 11118
rect 37326 11106 37378 11118
rect 40126 11106 40178 11118
rect 40350 11170 40402 11182
rect 40350 11106 40402 11118
rect 41806 11170 41858 11182
rect 41806 11106 41858 11118
rect 43598 11170 43650 11182
rect 43598 11106 43650 11118
rect 46286 11170 46338 11182
rect 46286 11106 46338 11118
rect 1344 11002 48608 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 48608 11002
rect 1344 10916 48608 10950
rect 6526 10834 6578 10846
rect 6526 10770 6578 10782
rect 9662 10834 9714 10846
rect 9662 10770 9714 10782
rect 12574 10834 12626 10846
rect 12574 10770 12626 10782
rect 21534 10834 21586 10846
rect 21534 10770 21586 10782
rect 33406 10834 33458 10846
rect 33406 10770 33458 10782
rect 33630 10834 33682 10846
rect 33630 10770 33682 10782
rect 33742 10834 33794 10846
rect 33742 10770 33794 10782
rect 37662 10834 37714 10846
rect 37662 10770 37714 10782
rect 38334 10834 38386 10846
rect 38334 10770 38386 10782
rect 39230 10834 39282 10846
rect 39230 10770 39282 10782
rect 39790 10834 39842 10846
rect 39790 10770 39842 10782
rect 42030 10834 42082 10846
rect 42030 10770 42082 10782
rect 5182 10722 5234 10734
rect 5182 10658 5234 10670
rect 9550 10722 9602 10734
rect 9550 10658 9602 10670
rect 9886 10722 9938 10734
rect 9886 10658 9938 10670
rect 10110 10722 10162 10734
rect 10110 10658 10162 10670
rect 15038 10722 15090 10734
rect 32510 10722 32562 10734
rect 31266 10670 31278 10722
rect 31330 10670 31342 10722
rect 15038 10658 15090 10670
rect 32510 10658 32562 10670
rect 33966 10722 34018 10734
rect 33966 10658 34018 10670
rect 39902 10722 39954 10734
rect 39902 10658 39954 10670
rect 40238 10722 40290 10734
rect 40238 10658 40290 10670
rect 40910 10722 40962 10734
rect 40910 10658 40962 10670
rect 41470 10722 41522 10734
rect 41470 10658 41522 10670
rect 42478 10722 42530 10734
rect 47954 10670 47966 10722
rect 48018 10670 48030 10722
rect 42478 10658 42530 10670
rect 6750 10610 6802 10622
rect 4610 10558 4622 10610
rect 4674 10558 4686 10610
rect 6750 10546 6802 10558
rect 7198 10610 7250 10622
rect 7198 10546 7250 10558
rect 12238 10610 12290 10622
rect 21310 10610 21362 10622
rect 12674 10558 12686 10610
rect 12738 10558 12750 10610
rect 15250 10558 15262 10610
rect 15314 10558 15326 10610
rect 18162 10558 18174 10610
rect 18226 10558 18238 10610
rect 12238 10546 12290 10558
rect 21310 10546 21362 10558
rect 25342 10610 25394 10622
rect 25342 10546 25394 10558
rect 25566 10610 25618 10622
rect 25566 10546 25618 10558
rect 25790 10610 25842 10622
rect 33518 10610 33570 10622
rect 37998 10610 38050 10622
rect 31938 10558 31950 10610
rect 32002 10558 32014 10610
rect 36418 10558 36430 10610
rect 36482 10558 36494 10610
rect 37090 10558 37102 10610
rect 37154 10558 37166 10610
rect 25790 10546 25842 10558
rect 33518 10546 33570 10558
rect 37998 10546 38050 10558
rect 38334 10610 38386 10622
rect 38334 10546 38386 10558
rect 38670 10610 38722 10622
rect 38670 10546 38722 10558
rect 39566 10610 39618 10622
rect 39566 10546 39618 10558
rect 41246 10610 41298 10622
rect 43474 10558 43486 10610
rect 43538 10558 43550 10610
rect 41246 10546 41298 10558
rect 5070 10498 5122 10510
rect 1698 10446 1710 10498
rect 1762 10446 1774 10498
rect 3826 10446 3838 10498
rect 3890 10446 3902 10498
rect 5070 10434 5122 10446
rect 6638 10498 6690 10510
rect 21422 10498 21474 10510
rect 18834 10446 18846 10498
rect 18898 10446 18910 10498
rect 20962 10446 20974 10498
rect 21026 10446 21038 10498
rect 6638 10434 6690 10446
rect 21422 10434 21474 10446
rect 25678 10498 25730 10510
rect 39006 10498 39058 10510
rect 29138 10446 29150 10498
rect 29202 10446 29214 10498
rect 34290 10446 34302 10498
rect 34354 10446 34366 10498
rect 37426 10446 37438 10498
rect 37490 10446 37502 10498
rect 25678 10434 25730 10446
rect 4958 10386 5010 10398
rect 4958 10322 5010 10334
rect 12462 10386 12514 10398
rect 12462 10322 12514 10334
rect 32398 10386 32450 10398
rect 37441 10383 37487 10446
rect 39006 10434 39058 10446
rect 39118 10498 39170 10510
rect 39118 10434 39170 10446
rect 40350 10498 40402 10510
rect 40350 10434 40402 10446
rect 41022 10498 41074 10510
rect 41022 10434 41074 10446
rect 42142 10498 42194 10510
rect 42142 10434 42194 10446
rect 42590 10386 42642 10398
rect 37874 10383 37886 10386
rect 37441 10337 37886 10383
rect 37874 10334 37886 10337
rect 37938 10334 37950 10386
rect 41570 10334 41582 10386
rect 41634 10383 41646 10386
rect 41794 10383 41806 10386
rect 41634 10337 41806 10383
rect 41634 10334 41646 10337
rect 41794 10334 41806 10337
rect 41858 10334 41870 10386
rect 32398 10322 32450 10334
rect 42590 10322 42642 10334
rect 1344 10218 48608 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 48608 10218
rect 1344 10132 48608 10166
rect 12238 10050 12290 10062
rect 12238 9986 12290 9998
rect 13582 10050 13634 10062
rect 13582 9986 13634 9998
rect 18846 10050 18898 10062
rect 18846 9986 18898 9998
rect 27918 10050 27970 10062
rect 39342 10050 39394 10062
rect 37202 9998 37214 10050
rect 37266 10047 37278 10050
rect 37538 10047 37550 10050
rect 37266 10001 37550 10047
rect 37266 9998 37278 10001
rect 37538 9998 37550 10001
rect 37602 9998 37614 10050
rect 41570 9998 41582 10050
rect 41634 9998 41646 10050
rect 27918 9986 27970 9998
rect 39342 9986 39394 9998
rect 3502 9938 3554 9950
rect 3502 9874 3554 9886
rect 4398 9938 4450 9950
rect 11342 9938 11394 9950
rect 8530 9886 8542 9938
rect 8594 9886 8606 9938
rect 4398 9874 4450 9886
rect 11342 9874 11394 9886
rect 13694 9938 13746 9950
rect 23438 9938 23490 9950
rect 14802 9886 14814 9938
rect 14866 9886 14878 9938
rect 16930 9886 16942 9938
rect 16994 9886 17006 9938
rect 13694 9874 13746 9886
rect 23438 9874 23490 9886
rect 23886 9938 23938 9950
rect 35086 9938 35138 9950
rect 24994 9886 25006 9938
rect 25058 9886 25070 9938
rect 27122 9886 27134 9938
rect 27186 9886 27198 9938
rect 31490 9886 31502 9938
rect 31554 9886 31566 9938
rect 33618 9886 33630 9938
rect 33682 9886 33694 9938
rect 23886 9874 23938 9886
rect 35086 9874 35138 9886
rect 37550 9938 37602 9950
rect 37550 9874 37602 9886
rect 38894 9938 38946 9950
rect 38894 9874 38946 9886
rect 45054 9938 45106 9950
rect 45266 9886 45278 9938
rect 45330 9886 45342 9938
rect 47394 9886 47406 9938
rect 47458 9886 47470 9938
rect 45054 9874 45106 9886
rect 3390 9826 3442 9838
rect 3390 9762 3442 9774
rect 3614 9826 3666 9838
rect 3614 9762 3666 9774
rect 4062 9826 4114 9838
rect 10446 9826 10498 9838
rect 5618 9774 5630 9826
rect 5682 9774 5694 9826
rect 4062 9762 4114 9774
rect 10446 9762 10498 9774
rect 10670 9826 10722 9838
rect 10670 9762 10722 9774
rect 11006 9826 11058 9838
rect 18062 9826 18114 9838
rect 21870 9826 21922 9838
rect 27582 9826 27634 9838
rect 12562 9774 12574 9826
rect 12626 9774 12638 9826
rect 14130 9774 14142 9826
rect 14194 9774 14206 9826
rect 17490 9774 17502 9826
rect 17554 9774 17566 9826
rect 18834 9774 18846 9826
rect 18898 9774 18910 9826
rect 21298 9774 21310 9826
rect 21362 9774 21374 9826
rect 24210 9774 24222 9826
rect 24274 9774 24286 9826
rect 11006 9762 11058 9774
rect 18062 9762 18114 9774
rect 21870 9762 21922 9774
rect 27582 9762 27634 9774
rect 27806 9826 27858 9838
rect 34862 9826 34914 9838
rect 30706 9774 30718 9826
rect 30770 9774 30782 9826
rect 27806 9762 27858 9774
rect 34862 9762 34914 9774
rect 34974 9826 35026 9838
rect 35982 9826 36034 9838
rect 35410 9774 35422 9826
rect 35474 9774 35486 9826
rect 35746 9774 35758 9826
rect 35810 9774 35822 9826
rect 34974 9762 35026 9774
rect 35982 9762 36034 9774
rect 36206 9826 36258 9838
rect 39118 9826 39170 9838
rect 36418 9774 36430 9826
rect 36482 9774 36494 9826
rect 36206 9762 36258 9774
rect 39118 9762 39170 9774
rect 40798 9826 40850 9838
rect 41458 9774 41470 9826
rect 41522 9774 41534 9826
rect 42018 9774 42030 9826
rect 42082 9774 42094 9826
rect 43362 9774 43374 9826
rect 43426 9774 43438 9826
rect 44258 9774 44270 9826
rect 44322 9774 44334 9826
rect 48066 9774 48078 9826
rect 48130 9774 48142 9826
rect 40798 9762 40850 9774
rect 19182 9714 19234 9726
rect 6402 9662 6414 9714
rect 6466 9662 6478 9714
rect 19182 9650 19234 9662
rect 22654 9714 22706 9726
rect 22654 9650 22706 9662
rect 27470 9714 27522 9726
rect 41010 9662 41022 9714
rect 41074 9662 41086 9714
rect 43810 9662 43822 9714
rect 43874 9662 43886 9714
rect 27470 9650 27522 9662
rect 10782 9602 10834 9614
rect 10782 9538 10834 9550
rect 12350 9602 12402 9614
rect 12350 9538 12402 9550
rect 17278 9602 17330 9614
rect 17278 9538 17330 9550
rect 21534 9602 21586 9614
rect 21534 9538 21586 9550
rect 21646 9602 21698 9614
rect 21646 9538 21698 9550
rect 21758 9602 21810 9614
rect 21758 9538 21810 9550
rect 22766 9602 22818 9614
rect 22766 9538 22818 9550
rect 34414 9602 34466 9614
rect 34414 9538 34466 9550
rect 35198 9602 35250 9614
rect 35198 9538 35250 9550
rect 36094 9602 36146 9614
rect 36094 9538 36146 9550
rect 37102 9602 37154 9614
rect 37102 9538 37154 9550
rect 39790 9602 39842 9614
rect 42914 9550 42926 9602
rect 42978 9550 42990 9602
rect 43138 9550 43150 9602
rect 43202 9550 43214 9602
rect 39790 9538 39842 9550
rect 1344 9434 48608 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 48608 9434
rect 1344 9348 48608 9382
rect 6302 9266 6354 9278
rect 6302 9202 6354 9214
rect 9662 9266 9714 9278
rect 9662 9202 9714 9214
rect 10782 9266 10834 9278
rect 10782 9202 10834 9214
rect 10894 9266 10946 9278
rect 10894 9202 10946 9214
rect 16270 9266 16322 9278
rect 16270 9202 16322 9214
rect 16830 9266 16882 9278
rect 16830 9202 16882 9214
rect 24782 9266 24834 9278
rect 24782 9202 24834 9214
rect 25790 9266 25842 9278
rect 25790 9202 25842 9214
rect 26014 9266 26066 9278
rect 26014 9202 26066 9214
rect 32510 9266 32562 9278
rect 32510 9202 32562 9214
rect 39566 9266 39618 9278
rect 39566 9202 39618 9214
rect 40238 9266 40290 9278
rect 40238 9202 40290 9214
rect 40910 9266 40962 9278
rect 40910 9202 40962 9214
rect 42926 9266 42978 9278
rect 42926 9202 42978 9214
rect 6078 9154 6130 9166
rect 6078 9090 6130 9102
rect 6414 9154 6466 9166
rect 6414 9090 6466 9102
rect 6638 9154 6690 9166
rect 6638 9090 6690 9102
rect 7198 9154 7250 9166
rect 7198 9090 7250 9102
rect 7310 9154 7362 9166
rect 25902 9154 25954 9166
rect 35198 9154 35250 9166
rect 12338 9102 12350 9154
rect 12402 9102 12414 9154
rect 15922 9102 15934 9154
rect 15986 9102 15998 9154
rect 7310 9090 7362 9102
rect 25678 9098 25730 9110
rect 10670 9042 10722 9054
rect 28690 9102 28702 9154
rect 28754 9102 28766 9154
rect 25902 9090 25954 9102
rect 35198 9090 35250 9102
rect 35310 9154 35362 9166
rect 40350 9154 40402 9166
rect 36418 9102 36430 9154
rect 36482 9102 36494 9154
rect 35310 9090 35362 9102
rect 40350 9090 40402 9102
rect 41134 9154 41186 9166
rect 41134 9090 41186 9102
rect 41358 9154 41410 9166
rect 41358 9090 41410 9102
rect 43038 9154 43090 9166
rect 43038 9090 43090 9102
rect 6962 8990 6974 9042
rect 7026 8990 7038 9042
rect 10322 8990 10334 9042
rect 10386 8990 10398 9042
rect 11554 8990 11566 9042
rect 11618 8990 11630 9042
rect 17378 8990 17390 9042
rect 17442 8990 17454 9042
rect 24098 8990 24110 9042
rect 24162 8990 24174 9042
rect 25218 8990 25230 9042
rect 25282 8990 25294 9042
rect 25678 9034 25730 9046
rect 27022 9042 27074 9054
rect 26786 8990 26798 9042
rect 26850 8990 26862 9042
rect 10670 8978 10722 8990
rect 27022 8978 27074 8990
rect 27134 9042 27186 9054
rect 33294 9042 33346 9054
rect 39678 9042 39730 9054
rect 41918 9042 41970 9054
rect 27906 8990 27918 9042
rect 27970 8990 27982 9042
rect 33506 8990 33518 9042
rect 33570 8990 33582 9042
rect 35634 8990 35646 9042
rect 35698 8990 35710 9042
rect 40002 8990 40014 9042
rect 40066 8990 40078 9042
rect 27134 8978 27186 8990
rect 33294 8978 33346 8990
rect 39678 8978 39730 8990
rect 41918 8978 41970 8990
rect 42030 9042 42082 9054
rect 42030 8978 42082 8990
rect 42142 9042 42194 9054
rect 42142 8978 42194 8990
rect 42254 9042 42306 9054
rect 43150 9042 43202 9054
rect 42466 8990 42478 9042
rect 42530 8990 42542 9042
rect 42254 8978 42306 8990
rect 43150 8978 43202 8990
rect 43374 9042 43426 9054
rect 44258 8990 44270 9042
rect 44322 8990 44334 9042
rect 48066 8990 48078 9042
rect 48130 8990 48142 9042
rect 43374 8978 43426 8990
rect 4062 8930 4114 8942
rect 20862 8930 20914 8942
rect 34078 8930 34130 8942
rect 14466 8878 14478 8930
rect 14530 8878 14542 8930
rect 18162 8878 18174 8930
rect 18226 8878 18238 8930
rect 20290 8878 20302 8930
rect 20354 8878 20366 8930
rect 21186 8878 21198 8930
rect 21250 8878 21262 8930
rect 23314 8878 23326 8930
rect 23378 8878 23390 8930
rect 30818 8878 30830 8930
rect 30882 8878 30894 8930
rect 4062 8866 4114 8878
rect 20862 8866 20914 8878
rect 34078 8866 34130 8878
rect 34750 8930 34802 8942
rect 41022 8930 41074 8942
rect 44942 8930 44994 8942
rect 38546 8878 38558 8930
rect 38610 8878 38622 8930
rect 44146 8878 44158 8930
rect 44210 8878 44222 8930
rect 45266 8878 45278 8930
rect 45330 8878 45342 8930
rect 47394 8878 47406 8930
rect 47458 8878 47470 8930
rect 34750 8866 34802 8878
rect 41022 8866 41074 8878
rect 44942 8866 44994 8878
rect 3838 8818 3890 8830
rect 34862 8818 34914 8830
rect 3490 8766 3502 8818
rect 3554 8766 3566 8818
rect 7746 8766 7758 8818
rect 7810 8766 7822 8818
rect 27570 8766 27582 8818
rect 27634 8766 27646 8818
rect 3838 8754 3890 8766
rect 34862 8754 34914 8766
rect 43598 8818 43650 8830
rect 43598 8754 43650 8766
rect 1344 8650 48608 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 48608 8650
rect 1344 8564 48608 8598
rect 13582 8482 13634 8494
rect 13582 8418 13634 8430
rect 18398 8482 18450 8494
rect 47182 8482 47234 8494
rect 40338 8430 40350 8482
rect 40402 8430 40414 8482
rect 44146 8430 44158 8482
rect 44210 8430 44222 8482
rect 18398 8418 18450 8430
rect 47182 8418 47234 8430
rect 18734 8370 18786 8382
rect 24110 8370 24162 8382
rect 4610 8318 4622 8370
rect 4674 8318 4686 8370
rect 5842 8318 5854 8370
rect 5906 8318 5918 8370
rect 12114 8318 12126 8370
rect 12178 8318 12190 8370
rect 16706 8318 16718 8370
rect 16770 8318 16782 8370
rect 20178 8318 20190 8370
rect 20242 8318 20254 8370
rect 21410 8318 21422 8370
rect 21474 8318 21486 8370
rect 23762 8318 23774 8370
rect 23826 8318 23838 8370
rect 18734 8306 18786 8318
rect 24110 8306 24162 8318
rect 24558 8370 24610 8382
rect 29262 8370 29314 8382
rect 35646 8370 35698 8382
rect 27458 8318 27470 8370
rect 27522 8318 27534 8370
rect 30370 8318 30382 8370
rect 30434 8318 30446 8370
rect 34290 8318 34302 8370
rect 34354 8318 34366 8370
rect 24558 8306 24610 8318
rect 29262 8306 29314 8318
rect 35646 8306 35698 8318
rect 37214 8370 37266 8382
rect 37214 8306 37266 8318
rect 37438 8370 37490 8382
rect 37438 8306 37490 8318
rect 38334 8370 38386 8382
rect 43822 8370 43874 8382
rect 40226 8318 40238 8370
rect 40290 8318 40302 8370
rect 41570 8318 41582 8370
rect 41634 8318 41646 8370
rect 45502 8370 45554 8382
rect 38334 8306 38386 8318
rect 43822 8306 43874 8318
rect 45278 8314 45330 8326
rect 12910 8258 12962 8270
rect 1810 8206 1822 8258
rect 1874 8206 1886 8258
rect 10882 8206 10894 8258
rect 10946 8206 10958 8258
rect 11890 8206 11902 8258
rect 11954 8206 11966 8258
rect 12910 8194 12962 8206
rect 13694 8258 13746 8270
rect 13694 8194 13746 8206
rect 16270 8258 16322 8270
rect 16270 8194 16322 8206
rect 18062 8258 18114 8270
rect 20638 8258 20690 8270
rect 18386 8206 18398 8258
rect 18450 8206 18462 8258
rect 19618 8206 19630 8258
rect 19682 8206 19694 8258
rect 18062 8194 18114 8206
rect 20638 8194 20690 8206
rect 21534 8258 21586 8270
rect 22990 8258 23042 8270
rect 25902 8258 25954 8270
rect 29150 8258 29202 8270
rect 21970 8206 21982 8258
rect 22034 8206 22046 8258
rect 22754 8206 22766 8258
rect 22818 8206 22830 8258
rect 23202 8206 23214 8258
rect 23266 8206 23278 8258
rect 26226 8206 26238 8258
rect 26290 8206 26302 8258
rect 27682 8206 27694 8258
rect 27746 8206 27758 8258
rect 21534 8194 21586 8206
rect 22990 8194 23042 8206
rect 25902 8194 25954 8206
rect 29150 8194 29202 8206
rect 29598 8258 29650 8270
rect 35086 8258 35138 8270
rect 31490 8206 31502 8258
rect 31554 8206 31566 8258
rect 29598 8194 29650 8206
rect 35086 8194 35138 8206
rect 35198 8258 35250 8270
rect 35198 8194 35250 8206
rect 36430 8258 36482 8270
rect 36430 8194 36482 8206
rect 36990 8258 37042 8270
rect 36990 8194 37042 8206
rect 38782 8258 38834 8270
rect 42142 8258 42194 8270
rect 40114 8206 40126 8258
rect 40178 8206 40190 8258
rect 40898 8206 40910 8258
rect 40962 8206 40974 8258
rect 41234 8206 41246 8258
rect 41298 8206 41310 8258
rect 38782 8194 38834 8206
rect 42142 8194 42194 8206
rect 43598 8258 43650 8270
rect 45502 8306 45554 8318
rect 46846 8370 46898 8382
rect 46846 8306 46898 8318
rect 45278 8250 45330 8262
rect 43598 8194 43650 8206
rect 11230 8146 11282 8158
rect 2482 8094 2494 8146
rect 2546 8094 2558 8146
rect 11230 8082 11282 8094
rect 17278 8146 17330 8158
rect 17278 8082 17330 8094
rect 20302 8146 20354 8158
rect 20302 8082 20354 8094
rect 21422 8146 21474 8158
rect 21422 8082 21474 8094
rect 22542 8146 22594 8158
rect 22542 8082 22594 8094
rect 23886 8146 23938 8158
rect 23886 8082 23938 8094
rect 25230 8146 25282 8158
rect 25230 8082 25282 8094
rect 25566 8146 25618 8158
rect 25566 8082 25618 8094
rect 25678 8146 25730 8158
rect 25678 8082 25730 8094
rect 26798 8146 26850 8158
rect 26798 8082 26850 8094
rect 28478 8146 28530 8158
rect 28478 8082 28530 8094
rect 28590 8146 28642 8158
rect 28590 8082 28642 8094
rect 29486 8146 29538 8158
rect 29486 8082 29538 8094
rect 30046 8146 30098 8158
rect 37886 8146 37938 8158
rect 32162 8094 32174 8146
rect 32226 8094 32238 8146
rect 37650 8094 37662 8146
rect 37714 8094 37726 8146
rect 30046 8082 30098 8094
rect 37886 8082 37938 8094
rect 42366 8146 42418 8158
rect 42366 8082 42418 8094
rect 42590 8146 42642 8158
rect 42590 8082 42642 8094
rect 42814 8146 42866 8158
rect 42814 8082 42866 8094
rect 43150 8146 43202 8158
rect 43150 8082 43202 8094
rect 43262 8146 43314 8158
rect 46174 8146 46226 8158
rect 45826 8094 45838 8146
rect 45890 8094 45902 8146
rect 43262 8082 43314 8094
rect 46174 8082 46226 8094
rect 46510 8146 46562 8158
rect 46510 8082 46562 8094
rect 47854 8146 47906 8158
rect 47854 8082 47906 8094
rect 5070 8034 5122 8046
rect 5070 7970 5122 7982
rect 12574 8034 12626 8046
rect 12574 7970 12626 7982
rect 13582 8034 13634 8046
rect 13582 7970 13634 7982
rect 16046 8034 16098 8046
rect 16046 7970 16098 7982
rect 16158 8034 16210 8046
rect 16158 7970 16210 7982
rect 16718 8034 16770 8046
rect 16718 7970 16770 7982
rect 16830 8034 16882 8046
rect 16830 7970 16882 7982
rect 17054 8034 17106 8046
rect 17054 7970 17106 7982
rect 17838 8034 17890 8046
rect 17838 7970 17890 7982
rect 17950 8034 18002 8046
rect 20190 8034 20242 8046
rect 19394 7982 19406 8034
rect 19458 7982 19470 8034
rect 17950 7970 18002 7982
rect 20190 7970 20242 7982
rect 20526 8034 20578 8046
rect 20526 7970 20578 7982
rect 21758 8034 21810 8046
rect 21758 7970 21810 7982
rect 23326 8034 23378 8046
rect 28254 8034 28306 8046
rect 26450 7982 26462 8034
rect 26514 7982 26526 8034
rect 23326 7970 23378 7982
rect 28254 7970 28306 7982
rect 30270 8034 30322 8046
rect 30270 7970 30322 7982
rect 34750 8034 34802 8046
rect 34750 7970 34802 7982
rect 34862 8034 34914 8046
rect 34862 7970 34914 7982
rect 34974 8034 35026 8046
rect 34974 7970 35026 7982
rect 35758 8034 35810 8046
rect 44942 8034 44994 8046
rect 36082 7982 36094 8034
rect 36146 7982 36158 8034
rect 37538 7982 37550 8034
rect 37602 7982 37614 8034
rect 35758 7970 35810 7982
rect 44942 7970 44994 7982
rect 47070 8034 47122 8046
rect 47070 7970 47122 7982
rect 47518 8034 47570 8046
rect 47518 7970 47570 7982
rect 1344 7866 48608 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 48608 7866
rect 1344 7780 48608 7814
rect 3502 7698 3554 7710
rect 3502 7634 3554 7646
rect 3726 7698 3778 7710
rect 3726 7634 3778 7646
rect 4622 7698 4674 7710
rect 32398 7698 32450 7710
rect 22978 7646 22990 7698
rect 23042 7646 23054 7698
rect 4622 7634 4674 7646
rect 32398 7634 32450 7646
rect 39454 7698 39506 7710
rect 39454 7634 39506 7646
rect 41470 7698 41522 7710
rect 41470 7634 41522 7646
rect 42478 7698 42530 7710
rect 44718 7698 44770 7710
rect 42802 7646 42814 7698
rect 42866 7646 42878 7698
rect 42478 7634 42530 7646
rect 44718 7634 44770 7646
rect 2942 7586 2994 7598
rect 2942 7522 2994 7534
rect 8990 7586 9042 7598
rect 8990 7522 9042 7534
rect 12798 7586 12850 7598
rect 23774 7586 23826 7598
rect 14578 7534 14590 7586
rect 14642 7534 14654 7586
rect 17602 7534 17614 7586
rect 17666 7534 17678 7586
rect 12798 7522 12850 7534
rect 23774 7522 23826 7534
rect 24110 7586 24162 7598
rect 32510 7586 32562 7598
rect 43374 7586 43426 7598
rect 31154 7534 31166 7586
rect 31218 7534 31230 7586
rect 33506 7534 33518 7586
rect 33570 7534 33582 7586
rect 35522 7534 35534 7586
rect 35586 7534 35598 7586
rect 47394 7534 47406 7586
rect 47458 7534 47470 7586
rect 24110 7522 24162 7534
rect 32510 7522 32562 7534
rect 43374 7522 43426 7534
rect 4174 7474 4226 7486
rect 4174 7410 4226 7422
rect 4398 7474 4450 7486
rect 4398 7410 4450 7422
rect 5070 7474 5122 7486
rect 23326 7474 23378 7486
rect 5506 7422 5518 7474
rect 5570 7422 5582 7474
rect 8642 7422 8654 7474
rect 8706 7422 8718 7474
rect 9650 7422 9662 7474
rect 9714 7422 9726 7474
rect 13010 7422 13022 7474
rect 13074 7422 13086 7474
rect 13794 7422 13806 7474
rect 13858 7422 13870 7474
rect 22642 7422 22654 7474
rect 22706 7422 22718 7474
rect 5070 7410 5122 7422
rect 23326 7410 23378 7422
rect 23998 7474 24050 7486
rect 41358 7474 41410 7486
rect 25554 7422 25566 7474
rect 25618 7422 25630 7474
rect 31938 7422 31950 7474
rect 32002 7422 32014 7474
rect 33282 7422 33294 7474
rect 33346 7422 33358 7474
rect 37650 7422 37662 7474
rect 37714 7422 37726 7474
rect 23998 7410 24050 7422
rect 41358 7410 41410 7422
rect 41582 7474 41634 7486
rect 43262 7474 43314 7486
rect 41682 7422 41694 7474
rect 41746 7422 41758 7474
rect 41582 7410 41634 7422
rect 43262 7410 43314 7422
rect 43598 7474 43650 7486
rect 43598 7410 43650 7422
rect 43822 7474 43874 7486
rect 43822 7410 43874 7422
rect 44382 7474 44434 7486
rect 44818 7422 44830 7474
rect 44882 7422 44894 7474
rect 48066 7422 48078 7474
rect 48130 7422 48142 7474
rect 44382 7410 44434 7422
rect 3614 7362 3666 7374
rect 2818 7310 2830 7362
rect 2882 7310 2894 7362
rect 3614 7298 3666 7310
rect 4510 7362 4562 7374
rect 8878 7362 8930 7374
rect 39566 7362 39618 7374
rect 6178 7310 6190 7362
rect 6242 7310 6254 7362
rect 8306 7310 8318 7362
rect 8370 7310 8382 7362
rect 10322 7310 10334 7362
rect 10386 7310 10398 7362
rect 12450 7310 12462 7362
rect 12514 7310 12526 7362
rect 16706 7310 16718 7362
rect 16770 7310 16782 7362
rect 26226 7310 26238 7362
rect 26290 7310 26302 7362
rect 28354 7310 28366 7362
rect 28418 7310 28430 7362
rect 29026 7310 29038 7362
rect 29090 7310 29102 7362
rect 4510 7298 4562 7310
rect 8878 7298 8930 7310
rect 39566 7298 39618 7310
rect 40014 7362 40066 7374
rect 40014 7298 40066 7310
rect 44606 7362 44658 7374
rect 45266 7310 45278 7362
rect 45330 7310 45342 7362
rect 44606 7298 44658 7310
rect 3166 7250 3218 7262
rect 3166 7186 3218 7198
rect 24334 7250 24386 7262
rect 24334 7186 24386 7198
rect 24558 7250 24610 7262
rect 24558 7186 24610 7198
rect 42030 7250 42082 7262
rect 42030 7186 42082 7198
rect 44158 7250 44210 7262
rect 44158 7186 44210 7198
rect 1344 7082 48608 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 48608 7082
rect 1344 6996 48608 7030
rect 13022 6914 13074 6926
rect 13022 6850 13074 6862
rect 30270 6914 30322 6926
rect 30270 6850 30322 6862
rect 40238 6914 40290 6926
rect 40238 6850 40290 6862
rect 41022 6914 41074 6926
rect 41022 6850 41074 6862
rect 42254 6914 42306 6926
rect 42254 6850 42306 6862
rect 45054 6914 45106 6926
rect 45054 6850 45106 6862
rect 45278 6914 45330 6926
rect 45278 6850 45330 6862
rect 45502 6914 45554 6926
rect 45502 6850 45554 6862
rect 5182 6802 5234 6814
rect 4610 6750 4622 6802
rect 4674 6750 4686 6802
rect 5182 6738 5234 6750
rect 6414 6802 6466 6814
rect 12014 6802 12066 6814
rect 17054 6802 17106 6814
rect 29262 6802 29314 6814
rect 11106 6750 11118 6802
rect 11170 6750 11182 6802
rect 16370 6750 16382 6802
rect 16434 6750 16446 6802
rect 17826 6750 17838 6802
rect 17890 6750 17902 6802
rect 6414 6738 6466 6750
rect 12014 6738 12066 6750
rect 17054 6738 17106 6750
rect 29262 6738 29314 6750
rect 33854 6802 33906 6814
rect 46734 6802 46786 6814
rect 37762 6750 37774 6802
rect 37826 6750 37838 6802
rect 39890 6750 39902 6802
rect 39954 6750 39966 6802
rect 33854 6738 33906 6750
rect 46734 6738 46786 6750
rect 6862 6690 6914 6702
rect 1810 6638 1822 6690
rect 1874 6638 1886 6690
rect 6862 6626 6914 6638
rect 7310 6690 7362 6702
rect 7310 6626 7362 6638
rect 7870 6690 7922 6702
rect 29374 6690 29426 6702
rect 8194 6638 8206 6690
rect 8258 6638 8270 6690
rect 8978 6638 8990 6690
rect 9042 6638 9054 6690
rect 12562 6638 12574 6690
rect 12626 6638 12638 6690
rect 13570 6638 13582 6690
rect 13634 6638 13646 6690
rect 16706 6638 16718 6690
rect 16770 6638 16782 6690
rect 17378 6638 17390 6690
rect 17442 6638 17454 6690
rect 20738 6638 20750 6690
rect 20802 6638 20814 6690
rect 26002 6638 26014 6690
rect 26066 6638 26078 6690
rect 7870 6626 7922 6638
rect 29374 6626 29426 6638
rect 29598 6690 29650 6702
rect 29598 6626 29650 6638
rect 30046 6690 30098 6702
rect 30046 6626 30098 6638
rect 30942 6690 30994 6702
rect 30942 6626 30994 6638
rect 32174 6690 32226 6702
rect 32174 6626 32226 6638
rect 33294 6690 33346 6702
rect 43710 6690 43762 6702
rect 35746 6638 35758 6690
rect 35810 6638 35822 6690
rect 36978 6638 36990 6690
rect 37042 6638 37054 6690
rect 40226 6638 40238 6690
rect 40290 6638 40302 6690
rect 33294 6626 33346 6638
rect 43710 6626 43762 6638
rect 43822 6690 43874 6702
rect 47630 6690 47682 6702
rect 44034 6638 44046 6690
rect 44098 6638 44110 6690
rect 44818 6638 44830 6690
rect 44882 6638 44894 6690
rect 43822 6626 43874 6638
rect 47630 6626 47682 6638
rect 48190 6690 48242 6702
rect 48190 6626 48242 6638
rect 5630 6578 5682 6590
rect 2482 6526 2494 6578
rect 2546 6526 2558 6578
rect 5630 6514 5682 6526
rect 6302 6578 6354 6590
rect 6302 6514 6354 6526
rect 6638 6578 6690 6590
rect 21310 6578 21362 6590
rect 29150 6578 29202 6590
rect 40574 6578 40626 6590
rect 12114 6526 12126 6578
rect 12178 6526 12190 6578
rect 12450 6526 12462 6578
rect 12514 6526 12526 6578
rect 14242 6526 14254 6578
rect 14306 6526 14318 6578
rect 19954 6526 19966 6578
rect 20018 6526 20030 6578
rect 24210 6526 24222 6578
rect 24274 6526 24286 6578
rect 28242 6526 28254 6578
rect 28306 6526 28318 6578
rect 32946 6526 32958 6578
rect 33010 6526 33022 6578
rect 6638 6514 6690 6526
rect 21310 6514 21362 6526
rect 29150 6514 29202 6526
rect 40574 6514 40626 6526
rect 41134 6578 41186 6590
rect 41134 6514 41186 6526
rect 42366 6578 42418 6590
rect 42366 6514 42418 6526
rect 42926 6578 42978 6590
rect 45614 6578 45666 6590
rect 43250 6526 43262 6578
rect 43314 6526 43326 6578
rect 44146 6526 44158 6578
rect 44210 6575 44222 6578
rect 44370 6575 44382 6578
rect 44210 6529 44382 6575
rect 44210 6526 44222 6529
rect 44370 6526 44382 6529
rect 44434 6526 44446 6578
rect 42926 6514 42978 6526
rect 45614 6514 45666 6526
rect 45950 6578 46002 6590
rect 47842 6526 47854 6578
rect 47906 6526 47918 6578
rect 45950 6514 46002 6526
rect 5966 6466 6018 6478
rect 5966 6402 6018 6414
rect 7198 6466 7250 6478
rect 7198 6402 7250 6414
rect 7422 6466 7474 6478
rect 7422 6402 7474 6414
rect 16942 6466 16994 6478
rect 16942 6402 16994 6414
rect 17166 6466 17218 6478
rect 17166 6402 17218 6414
rect 21422 6466 21474 6478
rect 21422 6402 21474 6414
rect 21534 6466 21586 6478
rect 21534 6402 21586 6414
rect 28590 6466 28642 6478
rect 31054 6466 31106 6478
rect 30594 6414 30606 6466
rect 30658 6414 30670 6466
rect 28590 6402 28642 6414
rect 31054 6402 31106 6414
rect 31278 6466 31330 6478
rect 31278 6402 31330 6414
rect 31614 6466 31666 6478
rect 31614 6402 31666 6414
rect 32510 6466 32562 6478
rect 32510 6402 32562 6414
rect 41022 6466 41074 6478
rect 41022 6402 41074 6414
rect 41582 6466 41634 6478
rect 41582 6402 41634 6414
rect 41918 6466 41970 6478
rect 41918 6402 41970 6414
rect 42142 6466 42194 6478
rect 42142 6402 42194 6414
rect 42590 6466 42642 6478
rect 42590 6402 42642 6414
rect 42814 6466 42866 6478
rect 42814 6402 42866 6414
rect 46286 6466 46338 6478
rect 46286 6402 46338 6414
rect 1344 6298 48608 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 48608 6298
rect 1344 6212 48608 6246
rect 5182 6130 5234 6142
rect 4722 6078 4734 6130
rect 4786 6078 4798 6130
rect 5182 6066 5234 6078
rect 8766 6130 8818 6142
rect 8766 6066 8818 6078
rect 15598 6130 15650 6142
rect 15598 6066 15650 6078
rect 16270 6130 16322 6142
rect 26574 6130 26626 6142
rect 20850 6078 20862 6130
rect 20914 6078 20926 6130
rect 16270 6066 16322 6078
rect 26574 6066 26626 6078
rect 33742 6130 33794 6142
rect 33742 6066 33794 6078
rect 33966 6130 34018 6142
rect 33966 6066 34018 6078
rect 38670 6130 38722 6142
rect 38670 6066 38722 6078
rect 39342 6130 39394 6142
rect 39342 6066 39394 6078
rect 39454 6130 39506 6142
rect 44606 6130 44658 6142
rect 41234 6078 41246 6130
rect 41298 6078 41310 6130
rect 39454 6066 39506 6078
rect 44606 6066 44658 6078
rect 45054 6130 45106 6142
rect 45054 6066 45106 6078
rect 5070 6018 5122 6030
rect 5070 5954 5122 5966
rect 7982 6018 8034 6030
rect 7982 5954 8034 5966
rect 16158 6018 16210 6030
rect 16158 5954 16210 5966
rect 16382 6018 16434 6030
rect 26462 6018 26514 6030
rect 25218 5966 25230 6018
rect 25282 5966 25294 6018
rect 16382 5954 16434 5966
rect 26462 5954 26514 5966
rect 26686 6018 26738 6030
rect 26686 5954 26738 5966
rect 34974 6018 35026 6030
rect 36082 5966 36094 6018
rect 36146 5966 36158 6018
rect 41122 5966 41134 6018
rect 41186 5966 41198 6018
rect 47394 5966 47406 6018
rect 47458 5966 47470 6018
rect 34974 5954 35026 5966
rect 4174 5906 4226 5918
rect 7422 5906 7474 5918
rect 5394 5854 5406 5906
rect 5458 5854 5470 5906
rect 6514 5854 6526 5906
rect 6578 5854 6590 5906
rect 4174 5842 4226 5854
rect 7422 5842 7474 5854
rect 7870 5906 7922 5918
rect 7870 5842 7922 5854
rect 8094 5906 8146 5918
rect 21198 5906 21250 5918
rect 33630 5906 33682 5918
rect 34862 5906 34914 5918
rect 39230 5906 39282 5918
rect 15138 5854 15150 5906
rect 15202 5854 15214 5906
rect 17938 5854 17950 5906
rect 18002 5854 18014 5906
rect 21746 5854 21758 5906
rect 21810 5854 21822 5906
rect 25442 5854 25454 5906
rect 25506 5854 25518 5906
rect 32274 5854 32286 5906
rect 32338 5854 32350 5906
rect 34178 5854 34190 5906
rect 34242 5854 34254 5906
rect 35410 5854 35422 5906
rect 35474 5854 35486 5906
rect 8094 5842 8146 5854
rect 21198 5842 21250 5854
rect 33630 5842 33682 5854
rect 34862 5842 34914 5854
rect 39230 5842 39282 5854
rect 39566 5906 39618 5918
rect 40798 5906 40850 5918
rect 39778 5854 39790 5906
rect 39842 5854 39854 5906
rect 39566 5842 39618 5854
rect 40798 5842 40850 5854
rect 41806 5906 41858 5918
rect 41806 5842 41858 5854
rect 42702 5906 42754 5918
rect 42702 5842 42754 5854
rect 42814 5906 42866 5918
rect 43486 5906 43538 5918
rect 43026 5854 43038 5906
rect 43090 5854 43102 5906
rect 48066 5854 48078 5906
rect 48130 5854 48142 5906
rect 42814 5842 42866 5854
rect 43486 5842 43538 5854
rect 6974 5794 7026 5806
rect 17614 5794 17666 5806
rect 26014 5794 26066 5806
rect 33182 5794 33234 5806
rect 6178 5742 6190 5794
rect 6242 5742 6254 5794
rect 10098 5742 10110 5794
rect 10162 5742 10174 5794
rect 22418 5742 22430 5794
rect 22482 5742 22494 5794
rect 24546 5742 24558 5794
rect 24610 5742 24622 5794
rect 29250 5742 29262 5794
rect 29314 5742 29326 5794
rect 6974 5730 7026 5742
rect 17614 5730 17666 5742
rect 26014 5730 26066 5742
rect 33182 5730 33234 5742
rect 33854 5794 33906 5806
rect 40126 5794 40178 5806
rect 38210 5742 38222 5794
rect 38274 5742 38286 5794
rect 33854 5730 33906 5742
rect 40126 5730 40178 5742
rect 40238 5794 40290 5806
rect 40238 5730 40290 5742
rect 41582 5794 41634 5806
rect 45266 5742 45278 5794
rect 45330 5742 45342 5794
rect 41582 5730 41634 5742
rect 4398 5682 4450 5694
rect 4398 5618 4450 5630
rect 7198 5682 7250 5694
rect 7198 5618 7250 5630
rect 18958 5682 19010 5694
rect 18958 5618 19010 5630
rect 25902 5682 25954 5694
rect 25902 5618 25954 5630
rect 33070 5682 33122 5694
rect 33070 5618 33122 5630
rect 41358 5682 41410 5694
rect 43710 5682 43762 5694
rect 42242 5630 42254 5682
rect 42306 5630 42318 5682
rect 44034 5630 44046 5682
rect 44098 5630 44110 5682
rect 44370 5630 44382 5682
rect 44434 5679 44446 5682
rect 45042 5679 45054 5682
rect 44434 5633 45054 5679
rect 44434 5630 44446 5633
rect 45042 5630 45054 5633
rect 45106 5630 45118 5682
rect 41358 5618 41410 5630
rect 43710 5618 43762 5630
rect 1344 5514 48608 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 48608 5514
rect 1344 5428 48608 5462
rect 30270 5346 30322 5358
rect 22530 5294 22542 5346
rect 22594 5294 22606 5346
rect 30270 5282 30322 5294
rect 39902 5346 39954 5358
rect 39902 5282 39954 5294
rect 40238 5346 40290 5358
rect 40238 5282 40290 5294
rect 41582 5346 41634 5358
rect 41582 5282 41634 5294
rect 41918 5346 41970 5358
rect 41918 5282 41970 5294
rect 15262 5234 15314 5246
rect 21534 5234 21586 5246
rect 25118 5234 25170 5246
rect 9650 5182 9662 5234
rect 9714 5182 9726 5234
rect 10770 5182 10782 5234
rect 10834 5182 10846 5234
rect 12898 5182 12910 5234
rect 12962 5182 12974 5234
rect 14914 5182 14926 5234
rect 14978 5182 14990 5234
rect 15698 5182 15710 5234
rect 15762 5182 15774 5234
rect 19506 5182 19518 5234
rect 19570 5182 19582 5234
rect 20402 5182 20414 5234
rect 20466 5182 20478 5234
rect 23538 5182 23550 5234
rect 23602 5182 23614 5234
rect 24658 5182 24670 5234
rect 24722 5182 24734 5234
rect 15262 5170 15314 5182
rect 21534 5170 21586 5182
rect 25118 5170 25170 5182
rect 26462 5234 26514 5246
rect 26462 5170 26514 5182
rect 26910 5234 26962 5246
rect 26910 5170 26962 5182
rect 29150 5234 29202 5246
rect 31054 5234 31106 5246
rect 43486 5234 43538 5246
rect 29586 5182 29598 5234
rect 29650 5182 29662 5234
rect 32162 5182 32174 5234
rect 32226 5182 32238 5234
rect 34290 5182 34302 5234
rect 34354 5182 34366 5234
rect 34738 5182 34750 5234
rect 34802 5182 34814 5234
rect 35858 5182 35870 5234
rect 35922 5182 35934 5234
rect 42690 5182 42702 5234
rect 42754 5182 42766 5234
rect 29150 5170 29202 5182
rect 31054 5170 31106 5182
rect 43486 5170 43538 5182
rect 44382 5234 44434 5246
rect 44818 5182 44830 5234
rect 44882 5182 44894 5234
rect 44382 5170 44434 5182
rect 5854 5122 5906 5134
rect 5854 5058 5906 5070
rect 6190 5122 6242 5134
rect 16158 5122 16210 5134
rect 21646 5122 21698 5134
rect 6738 5070 6750 5122
rect 6802 5070 6814 5122
rect 10098 5070 10110 5122
rect 10162 5070 10174 5122
rect 16594 5070 16606 5122
rect 16658 5070 16670 5122
rect 19842 5070 19854 5122
rect 19906 5070 19918 5122
rect 20514 5070 20526 5122
rect 20578 5070 20590 5122
rect 21298 5070 21310 5122
rect 21362 5070 21374 5122
rect 6190 5058 6242 5070
rect 16158 5058 16210 5070
rect 21646 5058 21698 5070
rect 22318 5122 22370 5134
rect 23438 5122 23490 5134
rect 24782 5122 24834 5134
rect 22754 5070 22766 5122
rect 22818 5070 22830 5122
rect 23986 5070 23998 5122
rect 24050 5070 24062 5122
rect 22318 5058 22370 5070
rect 23438 5058 23490 5070
rect 24782 5058 24834 5070
rect 29486 5122 29538 5134
rect 35086 5122 35138 5134
rect 40686 5122 40738 5134
rect 31490 5070 31502 5122
rect 31554 5070 31566 5122
rect 34626 5070 34638 5122
rect 34690 5070 34702 5122
rect 35634 5070 35646 5122
rect 35698 5070 35710 5122
rect 36306 5070 36318 5122
rect 36370 5070 36382 5122
rect 36978 5070 36990 5122
rect 37042 5070 37054 5122
rect 40226 5070 40238 5122
rect 40290 5070 40302 5122
rect 29486 5058 29538 5070
rect 35086 5058 35138 5070
rect 40686 5058 40738 5070
rect 41358 5122 41410 5134
rect 42802 5070 42814 5122
rect 42866 5070 42878 5122
rect 46946 5070 46958 5122
rect 47010 5070 47022 5122
rect 47618 5070 47630 5122
rect 47682 5070 47694 5122
rect 41358 5058 41410 5070
rect 5966 5010 6018 5022
rect 15038 5010 15090 5022
rect 7522 4958 7534 5010
rect 7586 4958 7598 5010
rect 5966 4946 6018 4958
rect 15038 4946 15090 4958
rect 15710 5010 15762 5022
rect 15710 4946 15762 4958
rect 15822 5010 15874 5022
rect 20078 5010 20130 5022
rect 17378 4958 17390 5010
rect 17442 4958 17454 5010
rect 15822 4946 15874 4958
rect 20078 4946 20130 4958
rect 21982 5010 22034 5022
rect 21982 4946 22034 4958
rect 23774 5010 23826 5022
rect 30494 5010 30546 5022
rect 27794 4958 27806 5010
rect 27858 4958 27870 5010
rect 23774 4946 23826 4958
rect 30494 4946 30546 4958
rect 35310 5010 35362 5022
rect 35310 4946 35362 4958
rect 35870 5010 35922 5022
rect 35870 4946 35922 4958
rect 41022 5010 41074 5022
rect 41022 4946 41074 4958
rect 16046 4898 16098 4910
rect 16046 4834 16098 4846
rect 20302 4898 20354 4910
rect 23550 4898 23602 4910
rect 26014 4898 26066 4910
rect 22418 4846 22430 4898
rect 22482 4846 22494 4898
rect 25666 4846 25678 4898
rect 25730 4846 25742 4898
rect 20302 4834 20354 4846
rect 23550 4834 23602 4846
rect 26014 4834 26066 4846
rect 28142 4898 28194 4910
rect 28142 4834 28194 4846
rect 28590 4898 28642 4910
rect 28590 4834 28642 4846
rect 30382 4898 30434 4910
rect 30382 4834 30434 4846
rect 34862 4898 34914 4910
rect 34862 4834 34914 4846
rect 36094 4898 36146 4910
rect 36094 4834 36146 4846
rect 37998 4898 38050 4910
rect 37998 4834 38050 4846
rect 1344 4730 48608 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 48608 4730
rect 1344 4644 48608 4678
rect 7758 4562 7810 4574
rect 7758 4498 7810 4510
rect 17614 4562 17666 4574
rect 17614 4498 17666 4510
rect 17838 4562 17890 4574
rect 17838 4498 17890 4510
rect 17950 4562 18002 4574
rect 17950 4498 18002 4510
rect 33294 4562 33346 4574
rect 33294 4498 33346 4510
rect 7422 4450 7474 4462
rect 7422 4386 7474 4398
rect 8654 4450 8706 4462
rect 8654 4386 8706 4398
rect 8990 4450 9042 4462
rect 17390 4450 17442 4462
rect 25230 4450 25282 4462
rect 33518 4450 33570 4462
rect 40910 4450 40962 4462
rect 10994 4398 11006 4450
rect 11058 4398 11070 4450
rect 14242 4398 14254 4450
rect 14306 4398 14318 4450
rect 19282 4398 19294 4450
rect 19346 4398 19358 4450
rect 22530 4398 22542 4450
rect 22594 4398 22606 4450
rect 30034 4398 30046 4450
rect 30098 4398 30110 4450
rect 39554 4398 39566 4450
rect 39618 4398 39630 4450
rect 8990 4386 9042 4398
rect 17390 4386 17442 4398
rect 25230 4386 25282 4398
rect 33518 4386 33570 4398
rect 40910 4386 40962 4398
rect 41246 4450 41298 4462
rect 41246 4386 41298 4398
rect 41582 4450 41634 4462
rect 41582 4386 41634 4398
rect 42142 4450 42194 4462
rect 45378 4398 45390 4450
rect 45442 4398 45454 4450
rect 42142 4386 42194 4398
rect 4162 4286 4174 4338
rect 4226 4286 4238 4338
rect 10210 4286 10222 4338
rect 10274 4286 10286 4338
rect 13570 4286 13582 4338
rect 13634 4286 13646 4338
rect 18498 4286 18510 4338
rect 18562 4286 18574 4338
rect 21858 4286 21870 4338
rect 21922 4286 21934 4338
rect 25778 4286 25790 4338
rect 25842 4286 25854 4338
rect 29250 4286 29262 4338
rect 29314 4286 29326 4338
rect 34066 4286 34078 4338
rect 34130 4286 34142 4338
rect 40338 4286 40350 4338
rect 40402 4286 40414 4338
rect 43586 4286 43598 4338
rect 43650 4286 43662 4338
rect 17726 4226 17778 4238
rect 42030 4226 42082 4238
rect 4946 4174 4958 4226
rect 5010 4174 5022 4226
rect 7074 4174 7086 4226
rect 7138 4174 7150 4226
rect 13122 4174 13134 4226
rect 13186 4174 13198 4226
rect 16370 4174 16382 4226
rect 16434 4174 16446 4226
rect 21410 4174 21422 4226
rect 21474 4174 21486 4226
rect 24658 4174 24670 4226
rect 24722 4174 24734 4226
rect 26562 4174 26574 4226
rect 26626 4174 26638 4226
rect 28690 4174 28702 4226
rect 28754 4174 28766 4226
rect 32162 4174 32174 4226
rect 32226 4174 32238 4226
rect 34738 4174 34750 4226
rect 34802 4174 34814 4226
rect 36866 4174 36878 4226
rect 36930 4174 36942 4226
rect 37426 4174 37438 4226
rect 37490 4174 37502 4226
rect 17726 4162 17778 4174
rect 42030 4162 42082 4174
rect 33630 4114 33682 4126
rect 33630 4050 33682 4062
rect 1344 3946 48608 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 48608 3946
rect 1344 3860 48608 3894
rect 7422 3778 7474 3790
rect 7422 3714 7474 3726
rect 17278 3778 17330 3790
rect 17278 3714 17330 3726
rect 24558 3778 24610 3790
rect 24558 3714 24610 3726
rect 24894 3778 24946 3790
rect 24894 3714 24946 3726
rect 26574 3778 26626 3790
rect 26574 3714 26626 3726
rect 26910 3778 26962 3790
rect 26910 3714 26962 3726
rect 28702 3778 28754 3790
rect 28702 3714 28754 3726
rect 40014 3778 40066 3790
rect 40014 3714 40066 3726
rect 7534 3666 7586 3678
rect 7534 3602 7586 3614
rect 17166 3666 17218 3678
rect 17166 3602 17218 3614
rect 22094 3666 22146 3678
rect 22094 3602 22146 3614
rect 28590 3666 28642 3678
rect 36990 3666 37042 3678
rect 30258 3614 30270 3666
rect 30322 3614 30334 3666
rect 32946 3614 32958 3666
rect 33010 3614 33022 3666
rect 35074 3614 35086 3666
rect 35138 3614 35150 3666
rect 28590 3602 28642 3614
rect 36990 3602 37042 3614
rect 45502 3666 45554 3678
rect 45502 3602 45554 3614
rect 47630 3554 47682 3566
rect 7746 3502 7758 3554
rect 7810 3502 7822 3554
rect 16370 3502 16382 3554
rect 16434 3502 16446 3554
rect 17602 3502 17614 3554
rect 17666 3502 17678 3554
rect 21074 3502 21086 3554
rect 21138 3502 21150 3554
rect 26562 3502 26574 3554
rect 26626 3502 26638 3554
rect 29026 3502 29038 3554
rect 29090 3502 29102 3554
rect 32274 3502 32286 3554
rect 32338 3502 32350 3554
rect 35970 3502 35982 3554
rect 36034 3502 36046 3554
rect 42354 3502 42366 3554
rect 42418 3502 42430 3554
rect 43922 3502 43934 3554
rect 43986 3502 43998 3554
rect 47630 3490 47682 3502
rect 8206 3442 8258 3454
rect 8206 3378 8258 3390
rect 17054 3442 17106 3454
rect 24670 3442 24722 3454
rect 19282 3390 19294 3442
rect 19346 3390 19358 3442
rect 17054 3378 17106 3390
rect 24670 3378 24722 3390
rect 44158 3442 44210 3454
rect 48190 3442 48242 3454
rect 47842 3390 47854 3442
rect 47906 3390 47918 3442
rect 44158 3378 44210 3390
rect 48190 3378 48242 3390
rect 3838 3330 3890 3342
rect 3838 3266 3890 3278
rect 5518 3330 5570 3342
rect 5518 3266 5570 3278
rect 6974 3330 7026 3342
rect 6974 3266 7026 3278
rect 8542 3330 8594 3342
rect 8542 3266 8594 3278
rect 10110 3330 10162 3342
rect 10110 3266 10162 3278
rect 11678 3330 11730 3342
rect 11678 3266 11730 3278
rect 12574 3330 12626 3342
rect 12574 3266 12626 3278
rect 13470 3330 13522 3342
rect 13470 3266 13522 3278
rect 15374 3330 15426 3342
rect 15374 3266 15426 3278
rect 25230 3330 25282 3342
rect 25230 3266 25282 3278
rect 25790 3330 25842 3342
rect 25790 3266 25842 3278
rect 27358 3330 27410 3342
rect 27358 3266 27410 3278
rect 38894 3330 38946 3342
rect 38894 3266 38946 3278
rect 42702 3330 42754 3342
rect 42702 3266 42754 3278
rect 44494 3330 44546 3342
rect 44494 3266 44546 3278
rect 44942 3330 44994 3342
rect 44942 3266 44994 3278
rect 46174 3330 46226 3342
rect 46174 3266 46226 3278
rect 1344 3162 48608 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 48608 3162
rect 1344 3076 48608 3110
rect 13458 1710 13470 1762
rect 13522 1759 13534 1762
rect 14578 1759 14590 1762
rect 13522 1713 14590 1759
rect 13522 1710 13534 1713
rect 14578 1710 14590 1713
rect 14642 1710 14654 1762
<< via1 >>
rect 30942 46398 30994 46450
rect 32622 46398 32674 46450
rect 33182 46398 33234 46450
rect 40350 46398 40402 46450
rect 41806 46398 41858 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 18510 45950 18562 46002
rect 21534 45950 21586 46002
rect 23662 45950 23714 46002
rect 24558 45950 24610 46002
rect 43150 45950 43202 46002
rect 44942 45950 44994 46002
rect 11342 45838 11394 45890
rect 18734 45838 18786 45890
rect 19630 45838 19682 45890
rect 20862 45838 20914 45890
rect 27470 45838 27522 45890
rect 28366 45838 28418 45890
rect 32174 45838 32226 45890
rect 32622 45838 32674 45890
rect 38222 45838 38274 45890
rect 43822 45838 43874 45890
rect 45278 45838 45330 45890
rect 10670 45726 10722 45778
rect 10894 45726 10946 45778
rect 19070 45726 19122 45778
rect 26686 45726 26738 45778
rect 29150 45726 29202 45778
rect 33070 45726 33122 45778
rect 33742 45726 33794 45778
rect 34414 45726 34466 45778
rect 37886 45726 37938 45778
rect 41582 45726 41634 45778
rect 41694 45726 41746 45778
rect 41806 45726 41858 45778
rect 45502 45726 45554 45778
rect 45838 45726 45890 45778
rect 47406 45726 47458 45778
rect 11118 45614 11170 45666
rect 19854 45614 19906 45666
rect 20078 45614 20130 45666
rect 31390 45614 31442 45666
rect 33406 45614 33458 45666
rect 33854 45614 33906 45666
rect 33966 45614 34018 45666
rect 34526 45614 34578 45666
rect 34638 45614 34690 45666
rect 37998 45614 38050 45666
rect 42254 45614 42306 45666
rect 43598 45614 43650 45666
rect 45950 45614 46002 45666
rect 46510 45614 46562 45666
rect 46846 45614 46898 45666
rect 47518 45614 47570 45666
rect 47630 45614 47682 45666
rect 48190 45614 48242 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 17502 45278 17554 45330
rect 18846 45278 18898 45330
rect 24670 45278 24722 45330
rect 31950 45278 32002 45330
rect 20526 45166 20578 45218
rect 21982 45166 22034 45218
rect 39118 45166 39170 45218
rect 13470 45054 13522 45106
rect 13806 45054 13858 45106
rect 17838 45054 17890 45106
rect 18174 45054 18226 45106
rect 18398 45054 18450 45106
rect 19742 45054 19794 45106
rect 21422 45054 21474 45106
rect 22430 45054 22482 45106
rect 23214 45054 23266 45106
rect 25230 45054 25282 45106
rect 25454 45054 25506 45106
rect 25678 45054 25730 45106
rect 25790 45054 25842 45106
rect 26350 45054 26402 45106
rect 27694 45054 27746 45106
rect 31390 45054 31442 45106
rect 31614 45054 31666 45106
rect 32286 45054 32338 45106
rect 36318 45054 36370 45106
rect 39902 45054 39954 45106
rect 41022 45054 41074 45106
rect 42926 45054 42978 45106
rect 48190 45054 48242 45106
rect 10558 44942 10610 44994
rect 12686 44942 12738 44994
rect 14590 44942 14642 44994
rect 16718 44942 16770 44994
rect 19406 44942 19458 44994
rect 24558 44942 24610 44994
rect 25566 44942 25618 44994
rect 28478 44942 28530 44994
rect 30606 44942 30658 44994
rect 31054 44942 31106 44994
rect 32510 44942 32562 44994
rect 33406 44942 33458 44994
rect 35534 44942 35586 44994
rect 36990 44942 37042 44994
rect 41694 44942 41746 44994
rect 44830 44942 44882 44994
rect 47630 44942 47682 44994
rect 18510 44830 18562 44882
rect 31166 44830 31218 44882
rect 40910 44830 40962 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 16158 44494 16210 44546
rect 20750 44494 20802 44546
rect 32286 44494 32338 44546
rect 32622 44494 32674 44546
rect 33854 44494 33906 44546
rect 34190 44494 34242 44546
rect 7646 44382 7698 44434
rect 12014 44382 12066 44434
rect 12686 44382 12738 44434
rect 15150 44382 15202 44434
rect 17390 44382 17442 44434
rect 30942 44382 30994 44434
rect 33182 44382 33234 44434
rect 34078 44382 34130 44434
rect 37998 44382 38050 44434
rect 43822 44382 43874 44434
rect 47742 44382 47794 44434
rect 10446 44270 10498 44322
rect 11566 44270 11618 44322
rect 14142 44270 14194 44322
rect 14366 44270 14418 44322
rect 15598 44270 15650 44322
rect 15822 44270 15874 44322
rect 16046 44270 16098 44322
rect 16494 44270 16546 44322
rect 16718 44270 16770 44322
rect 16942 44270 16994 44322
rect 20302 44270 20354 44322
rect 26574 44270 26626 44322
rect 31502 44270 31554 44322
rect 31950 44270 32002 44322
rect 32510 44270 32562 44322
rect 33630 44270 33682 44322
rect 37102 44270 37154 44322
rect 37438 44270 37490 44322
rect 38558 44270 38610 44322
rect 39790 44270 39842 44322
rect 40126 44270 40178 44322
rect 41022 44270 41074 44322
rect 44830 44270 44882 44322
rect 9774 44158 9826 44210
rect 11342 44158 11394 44210
rect 11454 44158 11506 44210
rect 12910 44158 12962 44210
rect 13470 44158 13522 44210
rect 15038 44158 15090 44210
rect 15262 44158 15314 44210
rect 17054 44158 17106 44210
rect 19518 44158 19570 44210
rect 20638 44158 20690 44210
rect 24558 44158 24610 44210
rect 30270 44158 30322 44210
rect 31054 44158 31106 44210
rect 31278 44158 31330 44210
rect 39342 44158 39394 44210
rect 40574 44158 40626 44210
rect 41694 44158 41746 44210
rect 45614 44158 45666 44210
rect 10894 44046 10946 44098
rect 12126 44046 12178 44098
rect 12686 44046 12738 44098
rect 27134 44046 27186 44098
rect 30606 44046 30658 44098
rect 32622 44046 32674 44098
rect 35870 44046 35922 44098
rect 36206 44046 36258 44098
rect 38334 44046 38386 44098
rect 40462 44046 40514 44098
rect 48190 44046 48242 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 16046 43710 16098 43762
rect 17278 43710 17330 43762
rect 25790 43710 25842 43762
rect 33182 43710 33234 43762
rect 33742 43710 33794 43762
rect 35422 43710 35474 43762
rect 36990 43710 37042 43762
rect 38222 43710 38274 43762
rect 41134 43710 41186 43762
rect 13582 43598 13634 43650
rect 16606 43598 16658 43650
rect 17838 43598 17890 43650
rect 18062 43598 18114 43650
rect 23886 43598 23938 43650
rect 24334 43598 24386 43650
rect 25230 43598 25282 43650
rect 35646 43598 35698 43650
rect 39006 43598 39058 43650
rect 40350 43598 40402 43650
rect 41022 43598 41074 43650
rect 42478 43598 42530 43650
rect 44830 43598 44882 43650
rect 5966 43486 6018 43538
rect 11342 43486 11394 43538
rect 11902 43486 11954 43538
rect 12574 43486 12626 43538
rect 16494 43486 16546 43538
rect 16718 43486 16770 43538
rect 17726 43486 17778 43538
rect 18174 43486 18226 43538
rect 20414 43486 20466 43538
rect 21646 43486 21698 43538
rect 21982 43486 22034 43538
rect 22654 43486 22706 43538
rect 24110 43486 24162 43538
rect 24446 43486 24498 43538
rect 25454 43486 25506 43538
rect 25678 43486 25730 43538
rect 26350 43486 26402 43538
rect 31950 43486 32002 43538
rect 33406 43486 33458 43538
rect 33966 43486 34018 43538
rect 34526 43486 34578 43538
rect 34750 43486 34802 43538
rect 34974 43486 35026 43538
rect 36430 43486 36482 43538
rect 36654 43486 36706 43538
rect 38110 43486 38162 43538
rect 38446 43486 38498 43538
rect 38558 43486 38610 43538
rect 39230 43486 39282 43538
rect 39678 43486 39730 43538
rect 39790 43486 39842 43538
rect 40910 43486 40962 43538
rect 42030 43486 42082 43538
rect 43822 43486 43874 43538
rect 48078 43486 48130 43538
rect 6638 43374 6690 43426
rect 8878 43374 8930 43426
rect 9550 43374 9602 43426
rect 10446 43374 10498 43426
rect 11566 43374 11618 43426
rect 12238 43374 12290 43426
rect 12350 43374 12402 43426
rect 13918 43374 13970 43426
rect 18734 43374 18786 43426
rect 20078 43374 20130 43426
rect 23214 43374 23266 43426
rect 24222 43374 24274 43426
rect 25566 43374 25618 43426
rect 27246 43374 27298 43426
rect 35310 43374 35362 43426
rect 38782 43374 38834 43426
rect 43374 43374 43426 43426
rect 44270 43374 44322 43426
rect 44606 43374 44658 43426
rect 44942 43374 44994 43426
rect 45278 43374 45330 43426
rect 47406 43374 47458 43426
rect 9774 43262 9826 43314
rect 10110 43262 10162 43314
rect 10558 43262 10610 43314
rect 10782 43262 10834 43314
rect 10894 43262 10946 43314
rect 11790 43262 11842 43314
rect 33070 43262 33122 43314
rect 34414 43262 34466 43314
rect 40014 43262 40066 43314
rect 40238 43262 40290 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 22654 42926 22706 42978
rect 24558 42926 24610 42978
rect 29710 42926 29762 42978
rect 31390 42926 31442 42978
rect 31726 42926 31778 42978
rect 39790 42926 39842 42978
rect 47406 42926 47458 42978
rect 47518 42926 47570 42978
rect 9998 42814 10050 42866
rect 16382 42814 16434 42866
rect 16830 42814 16882 42866
rect 19406 42814 19458 42866
rect 20414 42814 20466 42866
rect 21310 42814 21362 42866
rect 25118 42814 25170 42866
rect 28590 42814 28642 42866
rect 30158 42814 30210 42866
rect 31166 42814 31218 42866
rect 33070 42814 33122 42866
rect 34302 42814 34354 42866
rect 36430 42814 36482 42866
rect 44270 42814 44322 42866
rect 12910 42702 12962 42754
rect 13582 42702 13634 42754
rect 16942 42702 16994 42754
rect 17278 42702 17330 42754
rect 19182 42702 19234 42754
rect 20190 42702 20242 42754
rect 22318 42702 22370 42754
rect 22766 42702 22818 42754
rect 23550 42702 23602 42754
rect 23998 42702 24050 42754
rect 24670 42702 24722 42754
rect 25790 42702 25842 42754
rect 29150 42702 29202 42754
rect 29374 42702 29426 42754
rect 30382 42702 30434 42754
rect 30606 42702 30658 42754
rect 33630 42702 33682 42754
rect 39342 42702 39394 42754
rect 39566 42702 39618 42754
rect 40238 42702 40290 42754
rect 40574 42702 40626 42754
rect 40686 42702 40738 42754
rect 41470 42702 41522 42754
rect 45614 42702 45666 42754
rect 45726 42702 45778 42754
rect 46398 42702 46450 42754
rect 46846 42702 46898 42754
rect 47742 42702 47794 42754
rect 47854 42702 47906 42754
rect 14254 42590 14306 42642
rect 16718 42590 16770 42642
rect 17614 42590 17666 42642
rect 19630 42590 19682 42642
rect 21646 42590 21698 42642
rect 24558 42590 24610 42642
rect 26462 42590 26514 42642
rect 30046 42590 30098 42642
rect 37886 42590 37938 42642
rect 39902 42590 39954 42642
rect 41022 42590 41074 42642
rect 42142 42590 42194 42642
rect 44942 42590 44994 42642
rect 45502 42590 45554 42642
rect 47070 42590 47122 42642
rect 17950 42478 18002 42530
rect 25006 42478 25058 42530
rect 32398 42478 32450 42530
rect 33182 42478 33234 42530
rect 37550 42478 37602 42530
rect 40798 42478 40850 42530
rect 44830 42478 44882 42530
rect 46174 42478 46226 42530
rect 46734 42478 46786 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 14030 42142 14082 42194
rect 40238 42142 40290 42194
rect 41582 42142 41634 42194
rect 10782 42030 10834 42082
rect 11902 42030 11954 42082
rect 12574 42030 12626 42082
rect 16830 42030 16882 42082
rect 18622 42030 18674 42082
rect 18734 42030 18786 42082
rect 30830 42030 30882 42082
rect 36990 42030 37042 42082
rect 41358 42030 41410 42082
rect 42030 42030 42082 42082
rect 47966 42030 48018 42082
rect 6078 41918 6130 41970
rect 6862 41918 6914 41970
rect 10110 41918 10162 41970
rect 11678 41918 11730 41970
rect 12462 41918 12514 41970
rect 13806 41918 13858 41970
rect 14142 41918 14194 41970
rect 15374 41918 15426 41970
rect 16046 41918 16098 41970
rect 16718 41918 16770 41970
rect 18958 41918 19010 41970
rect 19182 41918 19234 41970
rect 19630 41918 19682 41970
rect 21086 41918 21138 41970
rect 22206 41918 22258 41970
rect 24558 41918 24610 41970
rect 24670 41918 24722 41970
rect 26126 41918 26178 41970
rect 26462 41918 26514 41970
rect 27246 41918 27298 41970
rect 30494 41918 30546 41970
rect 36654 41918 36706 41970
rect 37886 41918 37938 41970
rect 38446 41918 38498 41970
rect 41022 41918 41074 41970
rect 42142 41918 42194 41970
rect 42590 41918 42642 41970
rect 43038 41918 43090 41970
rect 8990 41806 9042 41858
rect 9886 41806 9938 41858
rect 10446 41806 10498 41858
rect 11230 41806 11282 41858
rect 11790 41806 11842 41858
rect 13134 41806 13186 41858
rect 16270 41806 16322 41858
rect 17838 41806 17890 41858
rect 18398 41806 18450 41858
rect 20750 41806 20802 41858
rect 22654 41806 22706 41858
rect 24110 41806 24162 41858
rect 25454 41806 25506 41858
rect 28030 41806 28082 41858
rect 30158 41806 30210 41858
rect 31278 41806 31330 41858
rect 33070 41806 33122 41858
rect 39902 41806 39954 41858
rect 40350 41806 40402 41858
rect 10894 41694 10946 41746
rect 11118 41694 11170 41746
rect 12574 41694 12626 41746
rect 23998 41694 24050 41746
rect 26350 41694 26402 41746
rect 26686 41694 26738 41746
rect 26798 41694 26850 41746
rect 33182 41694 33234 41746
rect 37326 41694 37378 41746
rect 37662 41694 37714 41746
rect 38446 41694 38498 41746
rect 38782 41694 38834 41746
rect 40910 41694 40962 41746
rect 41694 41694 41746 41746
rect 42366 41694 42418 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 19854 41358 19906 41410
rect 30718 41358 30770 41410
rect 34302 41358 34354 41410
rect 40686 41358 40738 41410
rect 6078 41246 6130 41298
rect 12014 41246 12066 41298
rect 14478 41246 14530 41298
rect 21758 41246 21810 41298
rect 23886 41246 23938 41298
rect 26462 41246 26514 41298
rect 28590 41246 28642 41298
rect 29486 41246 29538 41298
rect 38110 41246 38162 41298
rect 40238 41246 40290 41298
rect 41358 41246 41410 41298
rect 43486 41246 43538 41298
rect 45278 41246 45330 41298
rect 47406 41246 47458 41298
rect 10894 41134 10946 41186
rect 12350 41134 12402 41186
rect 13582 41134 13634 41186
rect 19518 41134 19570 41186
rect 21422 41134 21474 41186
rect 24558 41134 24610 41186
rect 25790 41134 25842 41186
rect 29710 41134 29762 41186
rect 30942 41134 30994 41186
rect 31166 41134 31218 41186
rect 31838 41134 31890 41186
rect 32286 41134 32338 41186
rect 32510 41134 32562 41186
rect 32846 41134 32898 41186
rect 33294 41134 33346 41186
rect 33742 41134 33794 41186
rect 34302 41134 34354 41186
rect 37326 41134 37378 41186
rect 44270 41134 44322 41186
rect 48078 41134 48130 41186
rect 12910 41022 12962 41074
rect 13470 41022 13522 41074
rect 13694 41022 13746 41074
rect 19966 41022 20018 41074
rect 20526 41022 20578 41074
rect 20750 41022 20802 41074
rect 29374 41022 29426 41074
rect 32958 41022 33010 41074
rect 33854 41022 33906 41074
rect 34638 41022 34690 41074
rect 35086 41022 35138 41074
rect 36094 41022 36146 41074
rect 40574 41022 40626 41074
rect 11342 40910 11394 40962
rect 20638 40910 20690 40962
rect 25230 40910 25282 40962
rect 31278 40910 31330 40962
rect 31390 40910 31442 40962
rect 32062 40910 32114 40962
rect 32174 40910 32226 40962
rect 33518 40910 33570 40962
rect 33630 40910 33682 40962
rect 34974 40910 35026 40962
rect 35982 40910 36034 40962
rect 40686 40910 40738 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 18734 40574 18786 40626
rect 18958 40574 19010 40626
rect 24446 40574 24498 40626
rect 25902 40574 25954 40626
rect 27694 40574 27746 40626
rect 28926 40574 28978 40626
rect 30494 40574 30546 40626
rect 30606 40574 30658 40626
rect 31614 40574 31666 40626
rect 32398 40574 32450 40626
rect 10334 40462 10386 40514
rect 12798 40462 12850 40514
rect 13134 40462 13186 40514
rect 13806 40462 13858 40514
rect 14142 40462 14194 40514
rect 15934 40462 15986 40514
rect 18062 40462 18114 40514
rect 20190 40462 20242 40514
rect 21758 40462 21810 40514
rect 22654 40462 22706 40514
rect 23998 40462 24050 40514
rect 25566 40462 25618 40514
rect 31390 40462 31442 40514
rect 32286 40462 32338 40514
rect 33854 40462 33906 40514
rect 34526 40462 34578 40514
rect 36542 40462 36594 40514
rect 47070 40462 47122 40514
rect 47966 40462 48018 40514
rect 4622 40350 4674 40402
rect 9662 40350 9714 40402
rect 15710 40350 15762 40402
rect 16270 40350 16322 40402
rect 18174 40350 18226 40402
rect 18510 40350 18562 40402
rect 20078 40350 20130 40402
rect 21198 40350 21250 40402
rect 23214 40350 23266 40402
rect 24222 40350 24274 40402
rect 24670 40350 24722 40402
rect 25230 40350 25282 40402
rect 26014 40350 26066 40402
rect 26686 40350 26738 40402
rect 27246 40350 27298 40402
rect 27470 40350 27522 40402
rect 27806 40350 27858 40402
rect 28030 40350 28082 40402
rect 28478 40350 28530 40402
rect 28702 40350 28754 40402
rect 29150 40350 29202 40402
rect 30158 40350 30210 40402
rect 30382 40350 30434 40402
rect 30718 40350 30770 40402
rect 31502 40350 31554 40402
rect 32062 40350 32114 40402
rect 33630 40350 33682 40402
rect 34302 40350 34354 40402
rect 38894 40350 38946 40402
rect 40910 40350 40962 40402
rect 41470 40350 41522 40402
rect 41918 40350 41970 40402
rect 42590 40350 42642 40402
rect 44606 40350 44658 40402
rect 45054 40350 45106 40402
rect 45614 40350 45666 40402
rect 45726 40350 45778 40402
rect 46622 40350 46674 40402
rect 47294 40350 47346 40402
rect 47742 40350 47794 40402
rect 1710 40238 1762 40290
rect 3838 40238 3890 40290
rect 24334 40238 24386 40290
rect 26462 40238 26514 40290
rect 28926 40238 28978 40290
rect 34414 40238 34466 40290
rect 46286 40238 46338 40290
rect 47518 40238 47570 40290
rect 12462 40182 12514 40234
rect 16494 40126 16546 40178
rect 16718 40126 16770 40178
rect 16830 40126 16882 40178
rect 32398 40126 32450 40178
rect 34078 40126 34130 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 19070 39790 19122 39842
rect 29150 39790 29202 39842
rect 30270 39790 30322 39842
rect 32062 39790 32114 39842
rect 44942 39790 44994 39842
rect 4174 39678 4226 39730
rect 9662 39678 9714 39730
rect 16718 39678 16770 39730
rect 18846 39678 18898 39730
rect 26014 39678 26066 39730
rect 26910 39678 26962 39730
rect 31838 39678 31890 39730
rect 35982 39678 36034 39730
rect 36318 39678 36370 39730
rect 37326 39678 37378 39730
rect 38782 39678 38834 39730
rect 39678 39678 39730 39730
rect 41694 39678 41746 39730
rect 45278 39678 45330 39730
rect 47406 39678 47458 39730
rect 2718 39566 2770 39618
rect 6750 39566 6802 39618
rect 10222 39566 10274 39618
rect 14478 39566 14530 39618
rect 15934 39566 15986 39618
rect 19518 39566 19570 39618
rect 20078 39566 20130 39618
rect 21310 39566 21362 39618
rect 22206 39566 22258 39618
rect 23102 39566 23154 39618
rect 27246 39566 27298 39618
rect 27694 39566 27746 39618
rect 28478 39566 28530 39618
rect 29262 39566 29314 39618
rect 29710 39566 29762 39618
rect 30046 39566 30098 39618
rect 30494 39566 30546 39618
rect 30718 39566 30770 39618
rect 32286 39566 32338 39618
rect 35310 39566 35362 39618
rect 35646 39566 35698 39618
rect 37438 39566 37490 39618
rect 37662 39566 37714 39618
rect 39454 39566 39506 39618
rect 40910 39566 40962 39618
rect 41246 39566 41298 39618
rect 42030 39566 42082 39618
rect 42590 39566 42642 39618
rect 44830 39566 44882 39618
rect 48078 39566 48130 39618
rect 3390 39454 3442 39506
rect 3502 39454 3554 39506
rect 3838 39454 3890 39506
rect 4510 39454 4562 39506
rect 4734 39454 4786 39506
rect 7534 39454 7586 39506
rect 10110 39454 10162 39506
rect 15486 39454 15538 39506
rect 19630 39454 19682 39506
rect 19854 39454 19906 39506
rect 20750 39454 20802 39506
rect 21422 39454 21474 39506
rect 23886 39454 23938 39506
rect 32734 39454 32786 39506
rect 32958 39454 33010 39506
rect 34526 39454 34578 39506
rect 34638 39454 34690 39506
rect 34862 39454 34914 39506
rect 35758 39454 35810 39506
rect 36430 39454 36482 39506
rect 36990 39454 37042 39506
rect 41358 39454 41410 39506
rect 42478 39454 42530 39506
rect 44046 39454 44098 39506
rect 2830 39342 2882 39394
rect 3054 39342 3106 39394
rect 3166 39342 3218 39394
rect 4062 39342 4114 39394
rect 4622 39342 4674 39394
rect 9998 39342 10050 39394
rect 10446 39342 10498 39394
rect 12350 39342 12402 39394
rect 14142 39342 14194 39394
rect 15374 39342 15426 39394
rect 20414 39342 20466 39394
rect 22430 39342 22482 39394
rect 22654 39342 22706 39394
rect 26686 39342 26738 39394
rect 28590 39342 28642 39394
rect 30830 39342 30882 39394
rect 33070 39342 33122 39394
rect 34190 39342 34242 39394
rect 34974 39342 35026 39394
rect 37214 39342 37266 39394
rect 40462 39342 40514 39394
rect 42366 39342 42418 39394
rect 43822 39342 43874 39394
rect 44158 39342 44210 39394
rect 44382 39342 44434 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 8542 39006 8594 39058
rect 10110 39006 10162 39058
rect 29374 39006 29426 39058
rect 31278 39006 31330 39058
rect 31950 39006 32002 39058
rect 39790 39006 39842 39058
rect 43150 39006 43202 39058
rect 45838 39006 45890 39058
rect 46734 39006 46786 39058
rect 46846 39006 46898 39058
rect 6078 38894 6130 38946
rect 9662 38894 9714 38946
rect 10334 38894 10386 38946
rect 10446 38894 10498 38946
rect 11678 38894 11730 38946
rect 12910 38894 12962 38946
rect 13134 38894 13186 38946
rect 18174 38894 18226 38946
rect 18286 38894 18338 38946
rect 20078 38894 20130 38946
rect 27694 38894 27746 38946
rect 29710 38894 29762 38946
rect 31726 38894 31778 38946
rect 32174 38894 32226 38946
rect 32398 38894 32450 38946
rect 33294 38894 33346 38946
rect 35870 38894 35922 38946
rect 38446 38894 38498 38946
rect 45054 38894 45106 38946
rect 45390 38894 45442 38946
rect 46398 38894 46450 38946
rect 46622 38894 46674 38946
rect 47854 38894 47906 38946
rect 4622 38782 4674 38834
rect 5294 38782 5346 38834
rect 8878 38782 8930 38834
rect 11006 38782 11058 38834
rect 12014 38782 12066 38834
rect 12462 38782 12514 38834
rect 13582 38782 13634 38834
rect 16942 38782 16994 38834
rect 18398 38782 18450 38834
rect 19854 38782 19906 38834
rect 20526 38782 20578 38834
rect 21310 38782 21362 38834
rect 22542 38782 22594 38834
rect 23214 38782 23266 38834
rect 24446 38782 24498 38834
rect 26014 38782 26066 38834
rect 26238 38782 26290 38834
rect 27134 38782 27186 38834
rect 29150 38782 29202 38834
rect 33182 38782 33234 38834
rect 33742 38782 33794 38834
rect 34078 38782 34130 38834
rect 35198 38782 35250 38834
rect 36094 38782 36146 38834
rect 36990 38782 37042 38834
rect 37214 38782 37266 38834
rect 37550 38782 37602 38834
rect 37774 38782 37826 38834
rect 37998 38782 38050 38834
rect 38110 38782 38162 38834
rect 39678 38782 39730 38834
rect 39902 38782 39954 38834
rect 41134 38782 41186 38834
rect 42142 38782 42194 38834
rect 43038 38782 43090 38834
rect 43374 38782 43426 38834
rect 43710 38782 43762 38834
rect 44158 38782 44210 38834
rect 44942 38782 44994 38834
rect 45614 38782 45666 38834
rect 45726 38782 45778 38834
rect 45950 38782 46002 38834
rect 46958 38782 47010 38834
rect 47406 38782 47458 38834
rect 48190 38782 48242 38834
rect 1710 38670 1762 38722
rect 3838 38670 3890 38722
rect 8206 38670 8258 38722
rect 9550 38670 9602 38722
rect 9886 38670 9938 38722
rect 10782 38670 10834 38722
rect 11342 38670 11394 38722
rect 12686 38670 12738 38722
rect 14254 38670 14306 38722
rect 16382 38670 16434 38722
rect 17838 38670 17890 38722
rect 19966 38670 20018 38722
rect 20862 38670 20914 38722
rect 25342 38670 25394 38722
rect 26798 38670 26850 38722
rect 31390 38670 31442 38722
rect 36430 38670 36482 38722
rect 40126 38670 40178 38722
rect 40350 38670 40402 38722
rect 41358 38670 41410 38722
rect 41918 38670 41970 38722
rect 47518 38670 47570 38722
rect 18846 38558 18898 38610
rect 21758 38558 21810 38610
rect 32286 38558 32338 38610
rect 35086 38558 35138 38610
rect 42030 38558 42082 38610
rect 44382 38558 44434 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 19406 38222 19458 38274
rect 19630 38222 19682 38274
rect 20190 38222 20242 38274
rect 21422 38222 21474 38274
rect 22206 38222 22258 38274
rect 29150 38222 29202 38274
rect 30382 38222 30434 38274
rect 30830 38222 30882 38274
rect 32510 38222 32562 38274
rect 32958 38222 33010 38274
rect 2718 38110 2770 38162
rect 6078 38110 6130 38162
rect 10446 38110 10498 38162
rect 10894 38110 10946 38162
rect 11566 38110 11618 38162
rect 12462 38110 12514 38162
rect 17278 38110 17330 38162
rect 20302 38110 20354 38162
rect 29374 38110 29426 38162
rect 29710 38110 29762 38162
rect 32734 38110 32786 38162
rect 33182 38110 33234 38162
rect 34302 38110 34354 38162
rect 36430 38110 36482 38162
rect 39678 38110 39730 38162
rect 43150 38110 43202 38162
rect 43598 38110 43650 38162
rect 47406 38110 47458 38162
rect 3278 37998 3330 38050
rect 3838 37998 3890 38050
rect 7310 37998 7362 38050
rect 8094 37998 8146 38050
rect 8430 37998 8482 38050
rect 8766 37998 8818 38050
rect 9662 37998 9714 38050
rect 12238 37998 12290 38050
rect 13694 37998 13746 38050
rect 14366 37998 14418 38050
rect 18622 37998 18674 38050
rect 18846 37998 18898 38050
rect 19070 37998 19122 38050
rect 19742 37998 19794 38050
rect 21534 37998 21586 38050
rect 26574 37998 26626 38050
rect 29598 37998 29650 38050
rect 32062 37998 32114 38050
rect 32398 37998 32450 38050
rect 33630 37998 33682 38050
rect 40126 37998 40178 38050
rect 41246 37998 41298 38050
rect 41918 37998 41970 38050
rect 43038 37998 43090 38050
rect 43486 37998 43538 38050
rect 44158 37998 44210 38050
rect 44830 37998 44882 38050
rect 45726 37998 45778 38050
rect 46734 37998 46786 38050
rect 47518 37998 47570 38050
rect 2830 37886 2882 37938
rect 3166 37886 3218 37938
rect 6190 37886 6242 37938
rect 6414 37886 6466 37938
rect 7870 37886 7922 37938
rect 9214 37886 9266 37938
rect 9886 37886 9938 37938
rect 10334 37886 10386 37938
rect 12574 37886 12626 37938
rect 15150 37886 15202 37938
rect 17726 37886 17778 37938
rect 18398 37886 18450 37938
rect 19294 37886 19346 37938
rect 20414 37886 20466 37938
rect 21422 37886 21474 37938
rect 22094 37886 22146 37938
rect 22206 37886 22258 37938
rect 22990 37886 23042 37938
rect 30270 37886 30322 37938
rect 30382 37886 30434 37938
rect 30942 37886 30994 37938
rect 32174 37886 32226 37938
rect 45838 37886 45890 37938
rect 47630 37886 47682 37938
rect 2606 37774 2658 37826
rect 6974 37774 7026 37826
rect 7982 37774 8034 37826
rect 18062 37774 18114 37826
rect 28590 37774 28642 37826
rect 29822 37774 29874 37826
rect 31502 37774 31554 37826
rect 43710 37774 43762 37826
rect 45054 37774 45106 37826
rect 45166 37774 45218 37826
rect 46846 37774 46898 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 17838 37438 17890 37490
rect 19406 37438 19458 37490
rect 19630 37438 19682 37490
rect 23662 37438 23714 37490
rect 25678 37438 25730 37490
rect 27582 37438 27634 37490
rect 33742 37438 33794 37490
rect 34750 37438 34802 37490
rect 34862 37438 34914 37490
rect 35646 37438 35698 37490
rect 36094 37438 36146 37490
rect 41022 37438 41074 37490
rect 42590 37438 42642 37490
rect 46286 37438 46338 37490
rect 47070 37438 47122 37490
rect 5742 37326 5794 37378
rect 8542 37326 8594 37378
rect 15150 37326 15202 37378
rect 23886 37326 23938 37378
rect 23998 37326 24050 37378
rect 26574 37326 26626 37378
rect 34190 37326 34242 37378
rect 35198 37326 35250 37378
rect 43038 37326 43090 37378
rect 44494 37326 44546 37378
rect 46174 37326 46226 37378
rect 46958 37326 47010 37378
rect 47742 37326 47794 37378
rect 3054 37214 3106 37266
rect 3502 37214 3554 37266
rect 5070 37214 5122 37266
rect 8094 37214 8146 37266
rect 8766 37214 8818 37266
rect 9774 37214 9826 37266
rect 14142 37214 14194 37266
rect 14814 37214 14866 37266
rect 16494 37214 16546 37266
rect 16830 37214 16882 37266
rect 17502 37214 17554 37266
rect 18622 37214 18674 37266
rect 19070 37214 19122 37266
rect 19742 37214 19794 37266
rect 22990 37214 23042 37266
rect 25566 37214 25618 37266
rect 27582 37214 27634 37266
rect 27806 37214 27858 37266
rect 28590 37214 28642 37266
rect 28926 37214 28978 37266
rect 29150 37214 29202 37266
rect 33630 37214 33682 37266
rect 33966 37214 34018 37266
rect 34638 37214 34690 37266
rect 34974 37214 35026 37266
rect 37102 37214 37154 37266
rect 41918 37214 41970 37266
rect 43934 37214 43986 37266
rect 47070 37214 47122 37266
rect 47854 37214 47906 37266
rect 7870 37102 7922 37154
rect 8654 37102 8706 37154
rect 10558 37102 10610 37154
rect 12686 37102 12738 37154
rect 13918 37102 13970 37154
rect 14478 37102 14530 37154
rect 18174 37102 18226 37154
rect 20078 37102 20130 37154
rect 22206 37102 22258 37154
rect 23550 37102 23602 37154
rect 24670 37102 24722 37154
rect 29934 37102 29986 37154
rect 32062 37102 32114 37154
rect 33182 37102 33234 37154
rect 33854 37102 33906 37154
rect 37886 37102 37938 37154
rect 40014 37102 40066 37154
rect 40910 37102 40962 37154
rect 2942 36990 2994 37042
rect 3278 36990 3330 37042
rect 33070 36990 33122 37042
rect 46286 36990 46338 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 18510 36654 18562 36706
rect 19854 36654 19906 36706
rect 38110 36654 38162 36706
rect 40350 36654 40402 36706
rect 43038 36654 43090 36706
rect 1710 36542 1762 36594
rect 3838 36542 3890 36594
rect 14926 36542 14978 36594
rect 17054 36542 17106 36594
rect 18174 36542 18226 36594
rect 25342 36542 25394 36594
rect 25678 36542 25730 36594
rect 30606 36542 30658 36594
rect 32622 36542 32674 36594
rect 34750 36542 34802 36594
rect 37886 36542 37938 36594
rect 41358 36542 41410 36594
rect 43822 36542 43874 36594
rect 44942 36542 44994 36594
rect 48190 36542 48242 36594
rect 4622 36430 4674 36482
rect 12014 36430 12066 36482
rect 14142 36430 14194 36482
rect 18062 36430 18114 36482
rect 18846 36430 18898 36482
rect 19294 36430 19346 36482
rect 20526 36430 20578 36482
rect 20862 36430 20914 36482
rect 21534 36430 21586 36482
rect 22542 36430 22594 36482
rect 28590 36430 28642 36482
rect 29262 36430 29314 36482
rect 31054 36430 31106 36482
rect 31950 36430 32002 36482
rect 37662 36430 37714 36482
rect 38334 36430 38386 36482
rect 40574 36430 40626 36482
rect 43262 36430 43314 36482
rect 43934 36430 43986 36482
rect 45390 36430 45442 36482
rect 5742 36318 5794 36370
rect 9774 36318 9826 36370
rect 19966 36318 20018 36370
rect 23214 36318 23266 36370
rect 27806 36318 27858 36370
rect 29710 36318 29762 36370
rect 36990 36318 37042 36370
rect 37326 36318 37378 36370
rect 37550 36318 37602 36370
rect 39790 36318 39842 36370
rect 40014 36318 40066 36370
rect 40126 36318 40178 36370
rect 41022 36318 41074 36370
rect 46062 36318 46114 36370
rect 5630 36206 5682 36258
rect 12574 36206 12626 36258
rect 20638 36206 20690 36258
rect 21646 36206 21698 36258
rect 21758 36206 21810 36258
rect 21982 36206 22034 36258
rect 29486 36206 29538 36258
rect 29598 36206 29650 36258
rect 29822 36206 29874 36258
rect 30606 36206 30658 36258
rect 30718 36206 30770 36258
rect 30942 36206 30994 36258
rect 36430 36206 36482 36258
rect 37102 36206 37154 36258
rect 42254 36206 42306 36258
rect 42702 36206 42754 36258
rect 44830 36206 44882 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 3278 35870 3330 35922
rect 7086 35870 7138 35922
rect 7198 35870 7250 35922
rect 7310 35870 7362 35922
rect 8206 35870 8258 35922
rect 8878 35870 8930 35922
rect 18174 35870 18226 35922
rect 22654 35870 22706 35922
rect 23998 35870 24050 35922
rect 24558 35870 24610 35922
rect 26910 35870 26962 35922
rect 28142 35870 28194 35922
rect 28814 35870 28866 35922
rect 29150 35870 29202 35922
rect 29598 35870 29650 35922
rect 29934 35870 29986 35922
rect 30830 35870 30882 35922
rect 32062 35870 32114 35922
rect 33406 35870 33458 35922
rect 36094 35870 36146 35922
rect 39902 35870 39954 35922
rect 41694 35870 41746 35922
rect 41918 35870 41970 35922
rect 47518 35870 47570 35922
rect 48190 35870 48242 35922
rect 3726 35758 3778 35810
rect 4174 35758 4226 35810
rect 4398 35758 4450 35810
rect 8654 35758 8706 35810
rect 8990 35758 9042 35810
rect 21310 35758 21362 35810
rect 25566 35758 25618 35810
rect 27358 35758 27410 35810
rect 28254 35758 28306 35810
rect 30046 35758 30098 35810
rect 31390 35758 31442 35810
rect 46286 35758 46338 35810
rect 47070 35758 47122 35810
rect 47406 35758 47458 35810
rect 47854 35758 47906 35810
rect 3166 35646 3218 35698
rect 3502 35646 3554 35698
rect 4062 35646 4114 35698
rect 4846 35646 4898 35698
rect 6862 35646 6914 35698
rect 7982 35646 8034 35698
rect 8094 35646 8146 35698
rect 8430 35646 8482 35698
rect 13806 35646 13858 35698
rect 22094 35646 22146 35698
rect 22542 35646 22594 35698
rect 22766 35646 22818 35698
rect 23214 35646 23266 35698
rect 23774 35646 23826 35698
rect 24110 35646 24162 35698
rect 24446 35646 24498 35698
rect 24782 35646 24834 35698
rect 25230 35646 25282 35698
rect 25342 35646 25394 35698
rect 25790 35646 25842 35698
rect 26686 35646 26738 35698
rect 27694 35646 27746 35698
rect 30382 35646 30434 35698
rect 30606 35646 30658 35698
rect 30718 35646 30770 35698
rect 31054 35646 31106 35698
rect 31726 35646 31778 35698
rect 32174 35646 32226 35698
rect 33070 35646 33122 35698
rect 35982 35646 36034 35698
rect 36318 35646 36370 35698
rect 36542 35646 36594 35698
rect 39790 35646 39842 35698
rect 42030 35646 42082 35698
rect 42478 35646 42530 35698
rect 46062 35646 46114 35698
rect 46398 35646 46450 35698
rect 10894 35534 10946 35586
rect 13022 35534 13074 35586
rect 17726 35534 17778 35586
rect 18062 35534 18114 35586
rect 18734 35534 18786 35586
rect 19182 35534 19234 35586
rect 23662 35534 23714 35586
rect 26014 35534 26066 35586
rect 34078 35534 34130 35586
rect 34526 35534 34578 35586
rect 37326 35534 37378 35586
rect 39454 35534 39506 35586
rect 43150 35534 43202 35586
rect 45278 35534 45330 35586
rect 46958 35534 47010 35586
rect 5070 35422 5122 35474
rect 6638 35422 6690 35474
rect 33966 35422 34018 35474
rect 45838 35422 45890 35474
rect 46622 35422 46674 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 3950 35086 4002 35138
rect 11902 35086 11954 35138
rect 12238 35086 12290 35138
rect 12910 35086 12962 35138
rect 23774 35086 23826 35138
rect 25006 35086 25058 35138
rect 36990 35086 37042 35138
rect 37550 35086 37602 35138
rect 37774 35086 37826 35138
rect 43262 35086 43314 35138
rect 3054 34974 3106 35026
rect 8094 34974 8146 35026
rect 8878 34974 8930 35026
rect 9550 34974 9602 35026
rect 17950 34974 18002 35026
rect 19966 34974 20018 35026
rect 20302 34974 20354 35026
rect 23550 34974 23602 35026
rect 26350 34974 26402 35026
rect 29262 34974 29314 35026
rect 35422 34974 35474 35026
rect 37326 34974 37378 35026
rect 40462 34974 40514 35026
rect 42590 34974 42642 35026
rect 43486 34974 43538 35026
rect 44942 34974 44994 35026
rect 48190 34974 48242 35026
rect 2158 34862 2210 34914
rect 3614 34862 3666 34914
rect 4398 34862 4450 34914
rect 4622 34862 4674 34914
rect 6750 34862 6802 34914
rect 7086 34862 7138 34914
rect 7310 34862 7362 34914
rect 8766 34862 8818 34914
rect 9214 34862 9266 34914
rect 9998 34862 10050 34914
rect 11454 34862 11506 34914
rect 13470 34862 13522 34914
rect 14030 34862 14082 34914
rect 15150 34862 15202 34914
rect 18286 34862 18338 34914
rect 22094 34862 22146 34914
rect 22430 34862 22482 34914
rect 23438 34862 23490 34914
rect 34190 34862 34242 34914
rect 37102 34862 37154 34914
rect 38558 34862 38610 34914
rect 39790 34862 39842 34914
rect 43038 34862 43090 34914
rect 45390 34862 45442 34914
rect 2270 34750 2322 34802
rect 2606 34750 2658 34802
rect 2942 34750 2994 34802
rect 3166 34750 3218 34802
rect 4510 34750 4562 34802
rect 5630 34750 5682 34802
rect 5966 34750 6018 34802
rect 7758 34750 7810 34802
rect 7982 34750 8034 34802
rect 8206 34750 8258 34802
rect 11230 34750 11282 34802
rect 11566 34750 11618 34802
rect 12462 34750 12514 34802
rect 12798 34750 12850 34802
rect 13806 34750 13858 34802
rect 15822 34750 15874 34802
rect 19406 34750 19458 34802
rect 22206 34750 22258 34802
rect 24222 34750 24274 34802
rect 24558 34750 24610 34802
rect 24894 34750 24946 34802
rect 25790 34750 25842 34802
rect 27022 34750 27074 34802
rect 29934 34750 29986 34802
rect 38222 34750 38274 34802
rect 38334 34750 38386 34802
rect 43598 34750 43650 34802
rect 43822 34750 43874 34802
rect 46062 34750 46114 34802
rect 2494 34638 2546 34690
rect 6862 34638 6914 34690
rect 13694 34638 13746 34690
rect 13918 34638 13970 34690
rect 14702 34638 14754 34690
rect 18510 34638 18562 34690
rect 18622 34638 18674 34690
rect 18734 34638 18786 34690
rect 18846 34638 18898 34690
rect 19294 34638 19346 34690
rect 20862 34638 20914 34690
rect 21870 34638 21922 34690
rect 23214 34638 23266 34690
rect 25006 34638 25058 34690
rect 25454 34638 25506 34690
rect 25678 34638 25730 34690
rect 26910 34638 26962 34690
rect 27470 34638 27522 34690
rect 27918 34638 27970 34690
rect 29374 34638 29426 34690
rect 36094 34638 36146 34690
rect 36430 34638 36482 34690
rect 38894 34638 38946 34690
rect 39342 34638 39394 34690
rect 44270 34638 44322 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 13246 34302 13298 34354
rect 13582 34302 13634 34354
rect 16382 34302 16434 34354
rect 18398 34302 18450 34354
rect 19294 34302 19346 34354
rect 23998 34302 24050 34354
rect 32174 34302 32226 34354
rect 36654 34302 36706 34354
rect 41246 34302 41298 34354
rect 2494 34190 2546 34242
rect 5966 34190 6018 34242
rect 13470 34190 13522 34242
rect 14142 34190 14194 34242
rect 16494 34190 16546 34242
rect 17950 34190 18002 34242
rect 18958 34190 19010 34242
rect 23774 34190 23826 34242
rect 24110 34190 24162 34242
rect 26462 34190 26514 34242
rect 29710 34190 29762 34242
rect 33854 34190 33906 34242
rect 39678 34190 39730 34242
rect 40014 34190 40066 34242
rect 40350 34190 40402 34242
rect 40910 34190 40962 34242
rect 1822 34078 1874 34130
rect 5182 34078 5234 34130
rect 9774 34078 9826 34130
rect 13022 34078 13074 34130
rect 18174 34078 18226 34130
rect 18622 34078 18674 34130
rect 19182 34078 19234 34130
rect 19406 34078 19458 34130
rect 19630 34078 19682 34130
rect 20526 34078 20578 34130
rect 24334 34078 24386 34130
rect 25790 34078 25842 34130
rect 29038 34078 29090 34130
rect 32398 34078 32450 34130
rect 33070 34078 33122 34130
rect 36318 34078 36370 34130
rect 36542 34078 36594 34130
rect 36766 34078 36818 34130
rect 36990 34078 37042 34130
rect 42142 34078 42194 34130
rect 43150 34078 43202 34130
rect 4622 33966 4674 34018
rect 8094 33966 8146 34018
rect 10558 33966 10610 34018
rect 12686 33966 12738 34018
rect 13358 33966 13410 34018
rect 14478 33966 14530 34018
rect 15038 33966 15090 34018
rect 15822 33966 15874 34018
rect 18286 33966 18338 34018
rect 20078 33966 20130 34018
rect 21310 33966 21362 34018
rect 23438 33966 23490 34018
rect 25454 33966 25506 34018
rect 28590 33966 28642 34018
rect 31838 33966 31890 34018
rect 35982 33966 36034 34018
rect 37438 33966 37490 34018
rect 38670 33966 38722 34018
rect 39342 33966 39394 34018
rect 41694 33966 41746 34018
rect 42478 33966 42530 34018
rect 46958 33966 47010 34018
rect 14590 33854 14642 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 11118 33518 11170 33570
rect 30270 33518 30322 33570
rect 30718 33518 30770 33570
rect 31614 33518 31666 33570
rect 44158 33518 44210 33570
rect 46398 33518 46450 33570
rect 46622 33518 46674 33570
rect 48078 33518 48130 33570
rect 7982 33406 8034 33458
rect 9438 33406 9490 33458
rect 10334 33406 10386 33458
rect 11230 33406 11282 33458
rect 13582 33406 13634 33458
rect 15710 33406 15762 33458
rect 20414 33406 20466 33458
rect 22430 33406 22482 33458
rect 26910 33406 26962 33458
rect 29486 33406 29538 33458
rect 30718 33406 30770 33458
rect 31166 33406 31218 33458
rect 32062 33406 32114 33458
rect 33070 33406 33122 33458
rect 43710 33406 43762 33458
rect 44942 33406 44994 33458
rect 46062 33406 46114 33458
rect 7758 33294 7810 33346
rect 9886 33294 9938 33346
rect 16382 33294 16434 33346
rect 17502 33294 17554 33346
rect 21534 33294 21586 33346
rect 22318 33294 22370 33346
rect 22542 33294 22594 33346
rect 22878 33294 22930 33346
rect 23550 33294 23602 33346
rect 23886 33294 23938 33346
rect 24334 33294 24386 33346
rect 26014 33294 26066 33346
rect 27582 33294 27634 33346
rect 28254 33294 28306 33346
rect 29262 33294 29314 33346
rect 29374 33294 29426 33346
rect 29822 33294 29874 33346
rect 35982 33294 36034 33346
rect 37326 33294 37378 33346
rect 37550 33294 37602 33346
rect 38222 33294 38274 33346
rect 38782 33294 38834 33346
rect 39790 33294 39842 33346
rect 40014 33294 40066 33346
rect 40910 33294 40962 33346
rect 41582 33294 41634 33346
rect 44046 33294 44098 33346
rect 45502 33294 45554 33346
rect 47070 33294 47122 33346
rect 47630 33294 47682 33346
rect 7086 33182 7138 33234
rect 18286 33182 18338 33234
rect 21310 33182 21362 33234
rect 23214 33182 23266 33234
rect 24558 33182 24610 33234
rect 25230 33182 25282 33234
rect 32286 33182 32338 33234
rect 35198 33182 35250 33234
rect 37886 33182 37938 33234
rect 38558 33182 38610 33234
rect 39230 33182 39282 33234
rect 39454 33182 39506 33234
rect 39902 33182 39954 33234
rect 40350 33182 40402 33234
rect 45838 33182 45890 33234
rect 46062 33182 46114 33234
rect 6750 33070 6802 33122
rect 6974 33070 7026 33122
rect 8990 33070 9042 33122
rect 23550 33070 23602 33122
rect 24894 33070 24946 33122
rect 26238 33070 26290 33122
rect 27358 33070 27410 33122
rect 27694 33070 27746 33122
rect 27918 33070 27970 33122
rect 28590 33070 28642 33122
rect 29598 33070 29650 33122
rect 30382 33070 30434 33122
rect 31614 33070 31666 33122
rect 32062 33070 32114 33122
rect 36430 33070 36482 33122
rect 37438 33070 37490 33122
rect 39118 33070 39170 33122
rect 44158 33070 44210 33122
rect 47966 33126 48018 33178
rect 48078 33182 48130 33234
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 14478 32734 14530 32786
rect 14590 32734 14642 32786
rect 15150 32734 15202 32786
rect 18174 32734 18226 32786
rect 30270 32734 30322 32786
rect 33966 32734 34018 32786
rect 34078 32734 34130 32786
rect 34862 32734 34914 32786
rect 39790 32734 39842 32786
rect 44494 32734 44546 32786
rect 4958 32622 5010 32674
rect 8766 32622 8818 32674
rect 14142 32622 14194 32674
rect 20190 32622 20242 32674
rect 24558 32622 24610 32674
rect 26686 32622 26738 32674
rect 27918 32622 27970 32674
rect 29822 32622 29874 32674
rect 33406 32622 33458 32674
rect 33742 32622 33794 32674
rect 34750 32622 34802 32674
rect 37214 32622 37266 32674
rect 40238 32622 40290 32674
rect 44942 32622 44994 32674
rect 48078 32622 48130 32674
rect 8318 32510 8370 32562
rect 8878 32510 8930 32562
rect 10446 32510 10498 32562
rect 13918 32510 13970 32562
rect 14366 32510 14418 32562
rect 14814 32510 14866 32562
rect 15374 32510 15426 32562
rect 16830 32510 16882 32562
rect 17950 32510 18002 32562
rect 18398 32510 18450 32562
rect 18622 32510 18674 32562
rect 23550 32510 23602 32562
rect 24670 32510 24722 32562
rect 25230 32510 25282 32562
rect 28478 32510 28530 32562
rect 28814 32510 28866 32562
rect 29038 32510 29090 32562
rect 29374 32510 29426 32562
rect 33070 32510 33122 32562
rect 34190 32510 34242 32562
rect 34302 32510 34354 32562
rect 35422 32510 35474 32562
rect 36542 32510 36594 32562
rect 39678 32510 39730 32562
rect 39902 32510 39954 32562
rect 41134 32510 41186 32562
rect 45950 32510 46002 32562
rect 48190 32510 48242 32562
rect 9662 32398 9714 32450
rect 11118 32398 11170 32450
rect 13246 32398 13298 32450
rect 16046 32398 16098 32450
rect 16382 32398 16434 32450
rect 17502 32398 17554 32450
rect 18286 32398 18338 32450
rect 28030 32398 28082 32450
rect 29262 32398 29314 32450
rect 35982 32398 36034 32450
rect 39342 32398 39394 32450
rect 41918 32398 41970 32450
rect 44046 32398 44098 32450
rect 8766 32286 8818 32338
rect 17390 32286 17442 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 43374 31950 43426 32002
rect 44046 31950 44098 32002
rect 4622 31838 4674 31890
rect 7758 31838 7810 31890
rect 15374 31838 15426 31890
rect 17502 31838 17554 31890
rect 17838 31838 17890 31890
rect 22878 31838 22930 31890
rect 25006 31838 25058 31890
rect 26014 31838 26066 31890
rect 29934 31838 29986 31890
rect 32062 31838 32114 31890
rect 33966 31838 34018 31890
rect 38334 31838 38386 31890
rect 42366 31838 42418 31890
rect 43038 31838 43090 31890
rect 44270 31838 44322 31890
rect 1822 31726 1874 31778
rect 5966 31726 6018 31778
rect 6414 31726 6466 31778
rect 10558 31726 10610 31778
rect 13470 31726 13522 31778
rect 13918 31726 13970 31778
rect 14142 31726 14194 31778
rect 14590 31726 14642 31778
rect 20638 31726 20690 31778
rect 22094 31726 22146 31778
rect 25902 31726 25954 31778
rect 26126 31726 26178 31778
rect 26798 31726 26850 31778
rect 26910 31726 26962 31778
rect 27358 31726 27410 31778
rect 27694 31726 27746 31778
rect 27918 31726 27970 31778
rect 29150 31726 29202 31778
rect 39566 31726 39618 31778
rect 44830 31726 44882 31778
rect 45054 31726 45106 31778
rect 45390 31726 45442 31778
rect 45726 31726 45778 31778
rect 46062 31726 46114 31778
rect 47406 31726 47458 31778
rect 2494 31614 2546 31666
rect 5630 31614 5682 31666
rect 5742 31614 5794 31666
rect 6190 31614 6242 31666
rect 6862 31614 6914 31666
rect 7086 31614 7138 31666
rect 9886 31614 9938 31666
rect 11790 31614 11842 31666
rect 11902 31614 11954 31666
rect 13806 31614 13858 31666
rect 19966 31614 20018 31666
rect 21310 31614 21362 31666
rect 21646 31614 21698 31666
rect 38670 31614 38722 31666
rect 40238 31614 40290 31666
rect 43150 31614 43202 31666
rect 43710 31614 43762 31666
rect 45166 31614 45218 31666
rect 45950 31614 46002 31666
rect 46398 31614 46450 31666
rect 46846 31614 46898 31666
rect 6638 31502 6690 31554
rect 13694 31502 13746 31554
rect 25678 31502 25730 31554
rect 26574 31502 26626 31554
rect 27022 31502 27074 31554
rect 27806 31502 27858 31554
rect 28366 31502 28418 31554
rect 33182 31502 33234 31554
rect 33518 31502 33570 31554
rect 34638 31502 34690 31554
rect 35198 31502 35250 31554
rect 35982 31502 36034 31554
rect 36542 31502 36594 31554
rect 37102 31502 37154 31554
rect 37438 31502 37490 31554
rect 37774 31502 37826 31554
rect 38782 31502 38834 31554
rect 45278 31502 45330 31554
rect 46510 31502 46562 31554
rect 46958 31502 47010 31554
rect 47966 31502 48018 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 6974 31166 7026 31218
rect 7198 31166 7250 31218
rect 8094 31166 8146 31218
rect 8654 31166 8706 31218
rect 16270 31166 16322 31218
rect 20638 31166 20690 31218
rect 21422 31166 21474 31218
rect 22654 31166 22706 31218
rect 25566 31166 25618 31218
rect 25902 31166 25954 31218
rect 26574 31166 26626 31218
rect 26798 31166 26850 31218
rect 27134 31166 27186 31218
rect 27358 31166 27410 31218
rect 32286 31166 32338 31218
rect 41358 31166 41410 31218
rect 41918 31166 41970 31218
rect 43038 31166 43090 31218
rect 43150 31166 43202 31218
rect 43262 31166 43314 31218
rect 44046 31166 44098 31218
rect 44158 31166 44210 31218
rect 4398 31054 4450 31106
rect 7310 31054 7362 31106
rect 7758 31054 7810 31106
rect 7870 31054 7922 31106
rect 8542 31054 8594 31106
rect 8878 31054 8930 31106
rect 10782 31054 10834 31106
rect 14926 31054 14978 31106
rect 20750 31054 20802 31106
rect 27582 31054 27634 31106
rect 29038 31054 29090 31106
rect 31614 31054 31666 31106
rect 44270 31054 44322 31106
rect 47182 31054 47234 31106
rect 3726 30942 3778 30994
rect 8318 30942 8370 30994
rect 11118 30942 11170 30994
rect 11566 30942 11618 30994
rect 12126 30942 12178 30994
rect 15486 30942 15538 30994
rect 17390 30942 17442 30994
rect 21870 30942 21922 30994
rect 23662 30942 23714 30994
rect 26126 30942 26178 30994
rect 6526 30830 6578 30882
rect 12574 30830 12626 30882
rect 14142 30830 14194 30882
rect 14590 30830 14642 30882
rect 15150 30830 15202 30882
rect 16718 30830 16770 30882
rect 18174 30830 18226 30882
rect 20302 30830 20354 30882
rect 22318 30830 22370 30882
rect 23102 30830 23154 30882
rect 24222 30830 24274 30882
rect 24670 30830 24722 30882
rect 26686 30830 26738 30882
rect 27246 30830 27298 30882
rect 27694 30830 27746 30882
rect 28030 30942 28082 30994
rect 28254 30942 28306 30994
rect 31726 30942 31778 30994
rect 31838 30942 31890 30994
rect 34862 30942 34914 30994
rect 35310 30942 35362 30994
rect 36542 30942 36594 30994
rect 37438 30942 37490 30994
rect 40910 30942 40962 30994
rect 41134 30942 41186 30994
rect 41582 30942 41634 30994
rect 42814 30942 42866 30994
rect 43374 30942 43426 30994
rect 43934 30942 43986 30994
rect 44494 30942 44546 30994
rect 47966 30942 48018 30994
rect 31166 30830 31218 30882
rect 33406 30830 33458 30882
rect 34302 30830 34354 30882
rect 35758 30830 35810 30882
rect 36206 30830 36258 30882
rect 38110 30830 38162 30882
rect 40238 30830 40290 30882
rect 41246 30830 41298 30882
rect 42030 30830 42082 30882
rect 42478 30830 42530 30882
rect 45054 30830 45106 30882
rect 23998 30718 24050 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 25454 30382 25506 30434
rect 27918 30382 27970 30434
rect 31390 30382 31442 30434
rect 34078 30382 34130 30434
rect 4622 30270 4674 30322
rect 13806 30270 13858 30322
rect 22542 30270 22594 30322
rect 30270 30270 30322 30322
rect 32062 30270 32114 30322
rect 45278 30270 45330 30322
rect 1822 30158 1874 30210
rect 5630 30158 5682 30210
rect 6190 30158 6242 30210
rect 6414 30158 6466 30210
rect 7310 30158 7362 30210
rect 8542 30158 8594 30210
rect 9214 30158 9266 30210
rect 20750 30158 20802 30210
rect 22990 30158 23042 30210
rect 25566 30158 25618 30210
rect 26462 30158 26514 30210
rect 26798 30158 26850 30210
rect 27134 30158 27186 30210
rect 27470 30158 27522 30210
rect 30718 30158 30770 30210
rect 31054 30158 31106 30210
rect 34078 30158 34130 30210
rect 34750 30158 34802 30210
rect 36430 30158 36482 30210
rect 36990 30158 37042 30210
rect 43486 30158 43538 30210
rect 47406 30158 47458 30210
rect 48078 30158 48130 30210
rect 2494 30046 2546 30098
rect 5742 30046 5794 30098
rect 5966 30046 6018 30098
rect 6638 30046 6690 30098
rect 6750 30046 6802 30098
rect 6974 30046 7026 30098
rect 7534 30046 7586 30098
rect 7870 30046 7922 30098
rect 8430 30046 8482 30098
rect 14926 30046 14978 30098
rect 18734 30046 18786 30098
rect 25902 30046 25954 30098
rect 26238 30046 26290 30098
rect 27694 30046 27746 30098
rect 30382 30046 30434 30098
rect 31502 30046 31554 30098
rect 31726 30046 31778 30098
rect 33406 30046 33458 30098
rect 33742 30046 33794 30098
rect 35086 30046 35138 30098
rect 35422 30046 35474 30098
rect 41806 30046 41858 30098
rect 7198 29934 7250 29986
rect 7758 29934 7810 29986
rect 8206 29934 8258 29986
rect 11342 29934 11394 29986
rect 12910 29934 12962 29986
rect 13694 29934 13746 29986
rect 13918 29934 13970 29986
rect 14142 29934 14194 29986
rect 14590 29934 14642 29986
rect 21422 29934 21474 29986
rect 24110 29934 24162 29986
rect 24558 29934 24610 29986
rect 25006 29934 25058 29986
rect 25454 29934 25506 29986
rect 26014 29934 26066 29986
rect 27246 29934 27298 29986
rect 28254 29934 28306 29986
rect 30830 29934 30882 29986
rect 32174 29934 32226 29986
rect 33070 29934 33122 29986
rect 34414 29934 34466 29986
rect 35870 29934 35922 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 5070 29598 5122 29650
rect 5966 29598 6018 29650
rect 6190 29598 6242 29650
rect 6974 29598 7026 29650
rect 16830 29598 16882 29650
rect 17726 29598 17778 29650
rect 18958 29598 19010 29650
rect 32286 29598 32338 29650
rect 33630 29598 33682 29650
rect 33854 29598 33906 29650
rect 5630 29486 5682 29538
rect 5742 29486 5794 29538
rect 6302 29486 6354 29538
rect 8990 29486 9042 29538
rect 12798 29486 12850 29538
rect 27358 29486 27410 29538
rect 33742 29486 33794 29538
rect 39790 29486 39842 29538
rect 40350 29486 40402 29538
rect 40910 29486 40962 29538
rect 41246 29486 41298 29538
rect 42702 29486 42754 29538
rect 1822 29374 1874 29426
rect 4846 29374 4898 29426
rect 5182 29374 5234 29426
rect 6750 29374 6802 29426
rect 7310 29374 7362 29426
rect 7534 29374 7586 29426
rect 7758 29374 7810 29426
rect 7982 29374 8034 29426
rect 8318 29374 8370 29426
rect 8654 29374 8706 29426
rect 12462 29374 12514 29426
rect 13134 29374 13186 29426
rect 13582 29374 13634 29426
rect 17726 29374 17778 29426
rect 17950 29374 18002 29426
rect 23214 29374 23266 29426
rect 24222 29374 24274 29426
rect 25342 29374 25394 29426
rect 33406 29374 33458 29426
rect 34078 29374 34130 29426
rect 34526 29374 34578 29426
rect 38782 29374 38834 29426
rect 42590 29374 42642 29426
rect 42926 29374 42978 29426
rect 43262 29374 43314 29426
rect 43710 29374 43762 29426
rect 45390 29374 45442 29426
rect 2494 29262 2546 29314
rect 4622 29262 4674 29314
rect 8542 29262 8594 29314
rect 9550 29262 9602 29314
rect 11678 29262 11730 29314
rect 14254 29262 14306 29314
rect 16382 29262 16434 29314
rect 17502 29262 17554 29314
rect 19070 29262 19122 29314
rect 20302 29262 20354 29314
rect 22430 29262 22482 29314
rect 24446 29262 24498 29314
rect 31726 29262 31778 29314
rect 35198 29262 35250 29314
rect 37326 29262 37378 29314
rect 37886 29262 37938 29314
rect 38334 29262 38386 29314
rect 39230 29262 39282 29314
rect 39566 29262 39618 29314
rect 39902 29262 39954 29314
rect 40238 29262 40290 29314
rect 41694 29262 41746 29314
rect 44158 29262 44210 29314
rect 46062 29262 46114 29314
rect 48190 29262 48242 29314
rect 5630 29150 5682 29202
rect 8094 29150 8146 29202
rect 23886 29150 23938 29202
rect 31950 29150 32002 29202
rect 41582 29150 41634 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 19070 28814 19122 28866
rect 19294 28814 19346 28866
rect 33518 28814 33570 28866
rect 33854 28814 33906 28866
rect 35198 28814 35250 28866
rect 43710 28814 43762 28866
rect 44046 28814 44098 28866
rect 45726 28814 45778 28866
rect 46062 28814 46114 28866
rect 3726 28702 3778 28754
rect 11678 28702 11730 28754
rect 12798 28702 12850 28754
rect 17390 28702 17442 28754
rect 19182 28702 19234 28754
rect 19630 28702 19682 28754
rect 20638 28702 20690 28754
rect 21534 28702 21586 28754
rect 22430 28702 22482 28754
rect 23998 28702 24050 28754
rect 26126 28702 26178 28754
rect 27470 28702 27522 28754
rect 35982 28702 36034 28754
rect 43710 28702 43762 28754
rect 44158 28702 44210 28754
rect 47630 28702 47682 28754
rect 3614 28590 3666 28642
rect 4062 28590 4114 28642
rect 4622 28590 4674 28642
rect 4734 28590 4786 28642
rect 5070 28590 5122 28642
rect 6190 28590 6242 28642
rect 7310 28590 7362 28642
rect 8654 28590 8706 28642
rect 11790 28590 11842 28642
rect 12014 28590 12066 28642
rect 12350 28590 12402 28642
rect 12686 28590 12738 28642
rect 13022 28590 13074 28642
rect 14926 28590 14978 28642
rect 19518 28590 19570 28642
rect 20190 28590 20242 28642
rect 22094 28590 22146 28642
rect 22542 28590 22594 28642
rect 23214 28602 23266 28654
rect 27134 28590 27186 28642
rect 27582 28590 27634 28642
rect 28478 28590 28530 28642
rect 29150 28590 29202 28642
rect 31166 28590 31218 28642
rect 33294 28590 33346 28642
rect 34190 28590 34242 28642
rect 34750 28590 34802 28642
rect 35086 28590 35138 28642
rect 36430 28590 36482 28642
rect 41806 28590 41858 28642
rect 43374 28590 43426 28642
rect 44830 28590 44882 28642
rect 45054 28590 45106 28642
rect 46062 28590 46114 28642
rect 47406 28590 47458 28642
rect 48190 28590 48242 28642
rect 3054 28478 3106 28530
rect 3166 28478 3218 28530
rect 3390 28478 3442 28530
rect 3950 28478 4002 28530
rect 4510 28478 4562 28530
rect 5630 28478 5682 28530
rect 7198 28478 7250 28530
rect 7982 28478 8034 28530
rect 8318 28478 8370 28530
rect 8430 28478 8482 28530
rect 9102 28478 9154 28530
rect 19742 28478 19794 28530
rect 19966 28478 20018 28530
rect 21422 28478 21474 28530
rect 21646 28478 21698 28530
rect 22318 28478 22370 28530
rect 22878 28478 22930 28530
rect 28590 28478 28642 28530
rect 29262 28478 29314 28530
rect 32286 28478 32338 28530
rect 38670 28478 38722 28530
rect 42814 28478 42866 28530
rect 6638 28366 6690 28418
rect 7646 28366 7698 28418
rect 8766 28366 8818 28418
rect 8990 28366 9042 28418
rect 10782 28366 10834 28418
rect 27918 28366 27970 28418
rect 30606 28366 30658 28418
rect 43038 28366 43090 28418
rect 43262 28366 43314 28418
rect 45390 28366 45442 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 9662 28030 9714 28082
rect 10558 28030 10610 28082
rect 15822 28030 15874 28082
rect 18846 28030 18898 28082
rect 22878 28030 22930 28082
rect 23438 28030 23490 28082
rect 26238 28030 26290 28082
rect 26574 28030 26626 28082
rect 28030 28030 28082 28082
rect 29374 28030 29426 28082
rect 30046 28030 30098 28082
rect 31278 28030 31330 28082
rect 40350 28030 40402 28082
rect 41246 28030 41298 28082
rect 41470 28030 41522 28082
rect 41582 28030 41634 28082
rect 42142 28030 42194 28082
rect 42478 28030 42530 28082
rect 11678 27918 11730 27970
rect 14814 27918 14866 27970
rect 14926 27918 14978 27970
rect 26686 27918 26738 27970
rect 29486 27918 29538 27970
rect 29822 27918 29874 27970
rect 40238 27918 40290 27970
rect 8654 27806 8706 27858
rect 10334 27806 10386 27858
rect 11006 27806 11058 27858
rect 14590 27806 14642 27858
rect 15710 27806 15762 27858
rect 18622 27806 18674 27858
rect 19070 27806 19122 27858
rect 19182 27806 19234 27858
rect 20078 27806 20130 27858
rect 20302 27806 20354 27858
rect 21086 27806 21138 27858
rect 21758 27806 21810 27858
rect 22654 27806 22706 27858
rect 22990 27806 23042 27858
rect 27582 27806 27634 27858
rect 27806 27806 27858 27858
rect 29150 27806 29202 27858
rect 30718 27806 30770 27858
rect 31166 27806 31218 27858
rect 31726 27806 31778 27858
rect 31950 27806 32002 27858
rect 33742 27806 33794 27858
rect 36990 27806 37042 27858
rect 41134 27806 41186 27858
rect 43598 27806 43650 27858
rect 6078 27694 6130 27746
rect 13806 27694 13858 27746
rect 16158 27694 16210 27746
rect 16830 27694 16882 27746
rect 17502 27694 17554 27746
rect 18958 27694 19010 27746
rect 20638 27694 20690 27746
rect 22430 27694 22482 27746
rect 24334 27694 24386 27746
rect 25342 27694 25394 27746
rect 27694 27694 27746 27746
rect 30158 27694 30210 27746
rect 33182 27694 33234 27746
rect 33294 27694 33346 27746
rect 34414 27694 34466 27746
rect 36542 27694 36594 27746
rect 37662 27694 37714 27746
rect 39790 27694 39842 27746
rect 41582 27694 41634 27746
rect 45390 27694 45442 27746
rect 15374 27582 15426 27634
rect 15934 27582 15986 27634
rect 17390 27582 17442 27634
rect 20750 27582 20802 27634
rect 21870 27582 21922 27634
rect 25230 27582 25282 27634
rect 32286 27582 32338 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 30158 27246 30210 27298
rect 37438 27246 37490 27298
rect 37774 27246 37826 27298
rect 2494 27134 2546 27186
rect 4622 27134 4674 27186
rect 8990 27134 9042 27186
rect 9326 27134 9378 27186
rect 14366 27134 14418 27186
rect 16718 27134 16770 27186
rect 18846 27134 18898 27186
rect 19630 27134 19682 27186
rect 20414 27134 20466 27186
rect 21310 27134 21362 27186
rect 25678 27134 25730 27186
rect 27358 27134 27410 27186
rect 30382 27134 30434 27186
rect 31502 27134 31554 27186
rect 32286 27134 32338 27186
rect 32734 27134 32786 27186
rect 33966 27134 34018 27186
rect 34974 27134 35026 27186
rect 35422 27134 35474 27186
rect 38446 27134 38498 27186
rect 40686 27134 40738 27186
rect 42478 27134 42530 27186
rect 48078 27134 48130 27186
rect 1822 27022 1874 27074
rect 6078 27022 6130 27074
rect 12238 27022 12290 27074
rect 14814 27022 14866 27074
rect 16046 27022 16098 27074
rect 24222 27022 24274 27074
rect 26014 27022 26066 27074
rect 32622 27022 32674 27074
rect 32846 27022 32898 27074
rect 33182 27022 33234 27074
rect 33854 27022 33906 27074
rect 34078 27022 34130 27074
rect 34302 27022 34354 27074
rect 34526 27022 34578 27074
rect 37550 27022 37602 27074
rect 37998 27022 38050 27074
rect 38670 27022 38722 27074
rect 39230 27022 39282 27074
rect 39342 27022 39394 27074
rect 39566 27022 39618 27074
rect 40350 27022 40402 27074
rect 41358 27022 41410 27074
rect 42254 27022 42306 27074
rect 42702 27022 42754 27074
rect 43150 27022 43202 27074
rect 43598 27022 43650 27074
rect 43934 27022 43986 27074
rect 45278 27022 45330 27074
rect 6862 26910 6914 26962
rect 11454 26910 11506 26962
rect 14254 26910 14306 26962
rect 14590 26910 14642 26962
rect 19854 26910 19906 26962
rect 23438 26910 23490 26962
rect 24558 26910 24610 26962
rect 24894 26910 24946 26962
rect 25678 26910 25730 26962
rect 26238 26910 26290 26962
rect 26574 26910 26626 26962
rect 29822 26910 29874 26962
rect 38334 26910 38386 26962
rect 40126 26910 40178 26962
rect 41022 26910 41074 26962
rect 42030 26910 42082 26962
rect 42926 26910 42978 26962
rect 43822 26910 43874 26962
rect 45950 26910 46002 26962
rect 19966 26798 20018 26850
rect 25790 26798 25842 26850
rect 26910 26798 26962 26850
rect 31390 26798 31442 26850
rect 33070 26798 33122 26850
rect 39454 26798 39506 26850
rect 39678 26798 39730 26850
rect 42478 26798 42530 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 5966 26462 6018 26514
rect 6302 26462 6354 26514
rect 7758 26462 7810 26514
rect 7870 26462 7922 26514
rect 8430 26462 8482 26514
rect 10558 26462 10610 26514
rect 16270 26462 16322 26514
rect 16606 26462 16658 26514
rect 18062 26462 18114 26514
rect 25790 26462 25842 26514
rect 29598 26462 29650 26514
rect 33854 26462 33906 26514
rect 34638 26462 34690 26514
rect 37550 26462 37602 26514
rect 38446 26462 38498 26514
rect 39790 26462 39842 26514
rect 43934 26462 43986 26514
rect 44382 26462 44434 26514
rect 44942 26462 44994 26514
rect 8318 26350 8370 26402
rect 8542 26350 8594 26402
rect 9886 26350 9938 26402
rect 10110 26350 10162 26402
rect 13694 26350 13746 26402
rect 16382 26350 16434 26402
rect 17614 26350 17666 26402
rect 21422 26350 21474 26402
rect 22318 26350 22370 26402
rect 24558 26350 24610 26402
rect 27358 26350 27410 26402
rect 39230 26350 39282 26402
rect 40910 26350 40962 26402
rect 41806 26350 41858 26402
rect 42030 26350 42082 26402
rect 42814 26350 42866 26402
rect 43038 26350 43090 26402
rect 43486 26350 43538 26402
rect 44046 26350 44098 26402
rect 44494 26350 44546 26402
rect 47630 26350 47682 26402
rect 48078 26350 48130 26402
rect 4622 26238 4674 26290
rect 4846 26238 4898 26290
rect 5182 26238 5234 26290
rect 5406 26238 5458 26290
rect 7086 26238 7138 26290
rect 7310 26238 7362 26290
rect 7982 26238 8034 26290
rect 9774 26238 9826 26290
rect 10222 26238 10274 26290
rect 10670 26238 10722 26290
rect 10782 26238 10834 26290
rect 12910 26238 12962 26290
rect 16830 26238 16882 26290
rect 18622 26238 18674 26290
rect 19070 26238 19122 26290
rect 19630 26238 19682 26290
rect 20638 26238 20690 26290
rect 22206 26238 22258 26290
rect 23998 26238 24050 26290
rect 25230 26238 25282 26290
rect 25678 26238 25730 26290
rect 25902 26238 25954 26290
rect 26686 26238 26738 26290
rect 33406 26238 33458 26290
rect 33630 26238 33682 26290
rect 34078 26238 34130 26290
rect 38334 26238 38386 26290
rect 38782 26238 38834 26290
rect 39006 26238 39058 26290
rect 39342 26238 39394 26290
rect 41022 26238 41074 26290
rect 41694 26238 41746 26290
rect 42142 26238 42194 26290
rect 42590 26238 42642 26290
rect 43598 26238 43650 26290
rect 44830 26238 44882 26290
rect 45054 26238 45106 26290
rect 46510 26238 46562 26290
rect 46622 26238 46674 26290
rect 46958 26238 47010 26290
rect 47182 26238 47234 26290
rect 47406 26238 47458 26290
rect 1710 26126 1762 26178
rect 3838 26126 3890 26178
rect 5070 26126 5122 26178
rect 15822 26126 15874 26178
rect 16494 26126 16546 26178
rect 19406 26126 19458 26178
rect 25454 26126 25506 26178
rect 33518 26126 33570 26178
rect 37886 26126 37938 26178
rect 42702 26126 42754 26178
rect 47070 26126 47122 26178
rect 47966 26126 48018 26178
rect 19518 26014 19570 26066
rect 37998 26014 38050 26066
rect 41246 26014 41298 26066
rect 45278 26014 45330 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 3502 25678 3554 25730
rect 28030 25678 28082 25730
rect 38782 25678 38834 25730
rect 7310 25566 7362 25618
rect 16382 25566 16434 25618
rect 20302 25566 20354 25618
rect 20638 25566 20690 25618
rect 30830 25566 30882 25618
rect 32958 25566 33010 25618
rect 33294 25566 33346 25618
rect 33742 25566 33794 25618
rect 39118 25566 39170 25618
rect 48190 25566 48242 25618
rect 3054 25454 3106 25506
rect 3950 25454 4002 25506
rect 4286 25454 4338 25506
rect 4398 25454 4450 25506
rect 4734 25454 4786 25506
rect 7086 25454 7138 25506
rect 10670 25454 10722 25506
rect 13470 25454 13522 25506
rect 17502 25454 17554 25506
rect 25118 25454 25170 25506
rect 27246 25454 27298 25506
rect 30158 25454 30210 25506
rect 36430 25454 36482 25506
rect 36990 25454 37042 25506
rect 37214 25454 37266 25506
rect 37326 25454 37378 25506
rect 39790 25454 39842 25506
rect 40238 25454 40290 25506
rect 40686 25454 40738 25506
rect 41022 25454 41074 25506
rect 41358 25454 41410 25506
rect 42030 25454 42082 25506
rect 43150 25454 43202 25506
rect 43598 25454 43650 25506
rect 44046 25454 44098 25506
rect 45390 25454 45442 25506
rect 3614 25342 3666 25394
rect 4622 25342 4674 25394
rect 5630 25342 5682 25394
rect 6750 25342 6802 25394
rect 7422 25342 7474 25394
rect 8430 25342 8482 25394
rect 8654 25342 8706 25394
rect 8878 25342 8930 25394
rect 8990 25342 9042 25394
rect 9774 25342 9826 25394
rect 10334 25342 10386 25394
rect 10446 25342 10498 25394
rect 11118 25342 11170 25394
rect 14254 25342 14306 25394
rect 18174 25342 18226 25394
rect 21982 25342 22034 25394
rect 27022 25342 27074 25394
rect 27806 25342 27858 25394
rect 28478 25342 28530 25394
rect 38110 25342 38162 25394
rect 38446 25342 38498 25394
rect 39006 25342 39058 25394
rect 39678 25342 39730 25394
rect 42366 25342 42418 25394
rect 42590 25342 42642 25394
rect 44270 25342 44322 25394
rect 44830 25342 44882 25394
rect 44942 25342 44994 25394
rect 46062 25342 46114 25394
rect 2718 25230 2770 25282
rect 2942 25230 2994 25282
rect 3502 25230 3554 25282
rect 4062 25230 4114 25282
rect 5966 25230 6018 25282
rect 6414 25230 6466 25282
rect 7758 25230 7810 25282
rect 8094 25230 8146 25282
rect 9886 25230 9938 25282
rect 10110 25230 10162 25282
rect 11230 25230 11282 25282
rect 11454 25230 11506 25282
rect 20750 25230 20802 25282
rect 27918 25230 27970 25282
rect 29710 25230 29762 25282
rect 33406 25230 33458 25282
rect 33854 25230 33906 25282
rect 37774 25230 37826 25282
rect 39566 25230 39618 25282
rect 41022 25230 41074 25282
rect 42254 25230 42306 25282
rect 42814 25230 42866 25282
rect 43038 25230 43090 25282
rect 43822 25230 43874 25282
rect 43934 25230 43986 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 5966 24894 6018 24946
rect 8206 24894 8258 24946
rect 10222 24894 10274 24946
rect 11790 24894 11842 24946
rect 16382 24894 16434 24946
rect 24446 24894 24498 24946
rect 32510 24894 32562 24946
rect 39790 24894 39842 24946
rect 42590 24894 42642 24946
rect 44046 24894 44098 24946
rect 45950 24894 46002 24946
rect 9886 24782 9938 24834
rect 9998 24782 10050 24834
rect 11342 24782 11394 24834
rect 11566 24782 11618 24834
rect 12238 24782 12290 24834
rect 12350 24782 12402 24834
rect 16718 24782 16770 24834
rect 24334 24782 24386 24834
rect 28590 24782 28642 24834
rect 33854 24782 33906 24834
rect 39902 24782 39954 24834
rect 42478 24782 42530 24834
rect 43150 24782 43202 24834
rect 46062 24782 46114 24834
rect 1822 24670 1874 24722
rect 4846 24670 4898 24722
rect 5182 24670 5234 24722
rect 5406 24670 5458 24722
rect 6302 24670 6354 24722
rect 8318 24670 8370 24722
rect 8542 24670 8594 24722
rect 8766 24670 8818 24722
rect 10334 24670 10386 24722
rect 10670 24670 10722 24722
rect 10894 24670 10946 24722
rect 12014 24670 12066 24722
rect 20190 24670 20242 24722
rect 23550 24670 23602 24722
rect 25342 24670 25394 24722
rect 25790 24670 25842 24722
rect 31278 24670 31330 24722
rect 31502 24670 31554 24722
rect 33070 24670 33122 24722
rect 36318 24670 36370 24722
rect 39454 24670 39506 24722
rect 40014 24670 40066 24722
rect 44830 24670 44882 24722
rect 2494 24558 2546 24610
rect 4622 24558 4674 24610
rect 5070 24558 5122 24610
rect 6750 24558 6802 24610
rect 10558 24558 10610 24610
rect 16830 24558 16882 24610
rect 17390 24558 17442 24610
rect 19518 24558 19570 24610
rect 20750 24558 20802 24610
rect 22878 24558 22930 24610
rect 35982 24558 36034 24610
rect 37102 24558 37154 24610
rect 39230 24558 39282 24610
rect 44158 24558 44210 24610
rect 45054 24558 45106 24610
rect 45502 24558 45554 24610
rect 45838 24558 45890 24610
rect 8094 24446 8146 24498
rect 12350 24446 12402 24498
rect 24446 24446 24498 24498
rect 31838 24446 31890 24498
rect 43038 24446 43090 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 21310 24110 21362 24162
rect 30494 24110 30546 24162
rect 9998 23998 10050 24050
rect 12126 23998 12178 24050
rect 16382 23998 16434 24050
rect 19742 23998 19794 24050
rect 21534 23998 21586 24050
rect 24558 23998 24610 24050
rect 26686 23998 26738 24050
rect 30270 23998 30322 24050
rect 37998 23998 38050 24050
rect 38334 23998 38386 24050
rect 42590 23998 42642 24050
rect 45278 23998 45330 24050
rect 4510 23886 4562 23938
rect 5966 23886 6018 23938
rect 8206 23886 8258 23938
rect 8654 23886 8706 23938
rect 8990 23886 9042 23938
rect 12798 23886 12850 23938
rect 13582 23886 13634 23938
rect 16830 23886 16882 23938
rect 20750 23886 20802 23938
rect 21870 23886 21922 23938
rect 21982 23886 22034 23938
rect 22542 23886 22594 23938
rect 22766 23886 22818 23938
rect 22990 23886 23042 23938
rect 23886 23886 23938 23938
rect 27246 23886 27298 23938
rect 27694 23886 27746 23938
rect 28142 23886 28194 23938
rect 29150 23886 29202 23938
rect 29374 23886 29426 23938
rect 29598 23886 29650 23938
rect 29822 23886 29874 23938
rect 36430 23886 36482 23938
rect 37886 23886 37938 23938
rect 39342 23886 39394 23938
rect 40014 23886 40066 23938
rect 41246 23886 41298 23938
rect 41806 23886 41858 23938
rect 42030 23886 42082 23938
rect 43150 23886 43202 23938
rect 43598 23886 43650 23938
rect 48078 23886 48130 23938
rect 4174 23774 4226 23826
rect 6750 23774 6802 23826
rect 7086 23774 7138 23826
rect 7758 23774 7810 23826
rect 8430 23774 8482 23826
rect 14254 23774 14306 23826
rect 17614 23774 17666 23826
rect 20414 23774 20466 23826
rect 23102 23774 23154 23826
rect 27022 23774 27074 23826
rect 28478 23774 28530 23826
rect 29486 23774 29538 23826
rect 31950 23774 32002 23826
rect 41694 23774 41746 23826
rect 42926 23774 42978 23826
rect 43710 23774 43762 23826
rect 43822 23774 43874 23826
rect 47406 23774 47458 23826
rect 4286 23662 4338 23714
rect 5630 23662 5682 23714
rect 7422 23662 7474 23714
rect 8542 23662 8594 23714
rect 20190 23662 20242 23714
rect 21758 23662 21810 23714
rect 23214 23662 23266 23714
rect 27358 23662 27410 23714
rect 27470 23662 27522 23714
rect 28030 23662 28082 23714
rect 28590 23662 28642 23714
rect 30830 23662 30882 23714
rect 38782 23662 38834 23714
rect 39454 23662 39506 23714
rect 39566 23662 39618 23714
rect 41022 23662 41074 23714
rect 42590 23662 42642 23714
rect 42702 23662 42754 23714
rect 44270 23662 44322 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 3950 23326 4002 23378
rect 5854 23326 5906 23378
rect 13582 23326 13634 23378
rect 14366 23326 14418 23378
rect 14590 23326 14642 23378
rect 17950 23326 18002 23378
rect 24558 23326 24610 23378
rect 36990 23326 37042 23378
rect 38446 23326 38498 23378
rect 41806 23326 41858 23378
rect 42254 23326 42306 23378
rect 42702 23326 42754 23378
rect 44494 23326 44546 23378
rect 47854 23326 47906 23378
rect 3278 23214 3330 23266
rect 3390 23214 3442 23266
rect 4510 23214 4562 23266
rect 5966 23214 6018 23266
rect 6526 23214 6578 23266
rect 6862 23214 6914 23266
rect 8654 23214 8706 23266
rect 8766 23214 8818 23266
rect 13470 23214 13522 23266
rect 14142 23214 14194 23266
rect 14926 23214 14978 23266
rect 16158 23214 16210 23266
rect 18622 23214 18674 23266
rect 20526 23214 20578 23266
rect 23102 23214 23154 23266
rect 23998 23214 24050 23266
rect 24110 23214 24162 23266
rect 24670 23214 24722 23266
rect 25230 23214 25282 23266
rect 25790 23214 25842 23266
rect 26238 23214 26290 23266
rect 26462 23214 26514 23266
rect 29598 23214 29650 23266
rect 36542 23214 36594 23266
rect 39454 23214 39506 23266
rect 44942 23214 44994 23266
rect 46398 23214 46450 23266
rect 3614 23102 3666 23154
rect 4062 23102 4114 23154
rect 4398 23102 4450 23154
rect 5406 23102 5458 23154
rect 15262 23102 15314 23154
rect 15934 23102 15986 23154
rect 18958 23102 19010 23154
rect 20302 23102 20354 23154
rect 21310 23102 21362 23154
rect 22766 23102 22818 23154
rect 27134 23102 27186 23154
rect 30270 23102 30322 23154
rect 30718 23102 30770 23154
rect 31278 23102 31330 23154
rect 31614 23102 31666 23154
rect 31838 23102 31890 23154
rect 33070 23102 33122 23154
rect 33294 23102 33346 23154
rect 34302 23102 34354 23154
rect 34974 23102 35026 23154
rect 35422 23102 35474 23154
rect 35534 23102 35586 23154
rect 35646 23102 35698 23154
rect 35982 23102 36034 23154
rect 36318 23102 36370 23154
rect 36878 23102 36930 23154
rect 37326 23102 37378 23154
rect 38782 23102 38834 23154
rect 39118 23102 39170 23154
rect 41470 23102 41522 23154
rect 41694 23102 41746 23154
rect 41918 23102 41970 23154
rect 42478 23102 42530 23154
rect 45166 23102 45218 23154
rect 45390 23102 45442 23154
rect 45838 23102 45890 23154
rect 48190 23102 48242 23154
rect 14478 22990 14530 23042
rect 15486 22990 15538 23042
rect 16830 22990 16882 23042
rect 17502 22990 17554 23042
rect 26350 22990 26402 23042
rect 27470 22990 27522 23042
rect 33854 22990 33906 23042
rect 34750 22990 34802 23042
rect 36094 22990 36146 23042
rect 37102 22990 37154 23042
rect 37886 22990 37938 23042
rect 42366 22990 42418 23042
rect 45054 22990 45106 23042
rect 47630 22990 47682 23042
rect 3950 22878 4002 22930
rect 8654 22878 8706 22930
rect 13694 22878 13746 22930
rect 23214 22878 23266 22930
rect 23998 22878 24050 22930
rect 24558 22878 24610 22930
rect 25342 22878 25394 22930
rect 25678 22878 25730 22930
rect 32174 22878 32226 22930
rect 44270 22878 44322 22930
rect 44606 22878 44658 22930
rect 46062 22878 46114 22930
rect 46286 22878 46338 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 17390 22542 17442 22594
rect 43934 22542 43986 22594
rect 4622 22430 4674 22482
rect 10894 22430 10946 22482
rect 15710 22430 15762 22482
rect 16270 22430 16322 22482
rect 17838 22430 17890 22482
rect 21646 22430 21698 22482
rect 21982 22430 22034 22482
rect 24558 22430 24610 22482
rect 26686 22430 26738 22482
rect 29150 22430 29202 22482
rect 36094 22430 36146 22482
rect 39902 22430 39954 22482
rect 43710 22430 43762 22482
rect 45278 22430 45330 22482
rect 1710 22318 1762 22370
rect 5630 22318 5682 22370
rect 6414 22318 6466 22370
rect 7422 22318 7474 22370
rect 8094 22318 8146 22370
rect 14478 22318 14530 22370
rect 16942 22318 16994 22370
rect 17166 22318 17218 22370
rect 20750 22318 20802 22370
rect 21422 22318 21474 22370
rect 22990 22318 23042 22370
rect 23102 22318 23154 22370
rect 23438 22318 23490 22370
rect 23774 22318 23826 22370
rect 31950 22318 32002 22370
rect 33182 22318 33234 22370
rect 36990 22318 37042 22370
rect 40462 22318 40514 22370
rect 41358 22318 41410 22370
rect 42030 22318 42082 22370
rect 42814 22318 42866 22370
rect 43262 22318 43314 22370
rect 48078 22318 48130 22370
rect 2494 22206 2546 22258
rect 6302 22206 6354 22258
rect 7534 22206 7586 22258
rect 8766 22206 8818 22258
rect 17502 22206 17554 22258
rect 19966 22206 20018 22258
rect 22878 22206 22930 22258
rect 31278 22206 31330 22258
rect 32286 22206 32338 22258
rect 32846 22206 32898 22258
rect 33966 22206 34018 22258
rect 37774 22206 37826 22258
rect 40238 22206 40290 22258
rect 42366 22206 42418 22258
rect 42926 22206 42978 22258
rect 43374 22206 43426 22258
rect 47406 22206 47458 22258
rect 5742 22094 5794 22146
rect 5966 22094 6018 22146
rect 6078 22094 6130 22146
rect 7758 22094 7810 22146
rect 14590 22094 14642 22146
rect 14702 22094 14754 22146
rect 14926 22094 14978 22146
rect 16718 22094 16770 22146
rect 21870 22094 21922 22146
rect 22094 22094 22146 22146
rect 22766 22094 22818 22146
rect 27358 22094 27410 22146
rect 27470 22094 27522 22146
rect 27582 22094 27634 22146
rect 27806 22094 27858 22146
rect 28478 22094 28530 22146
rect 32398 22094 32450 22146
rect 32622 22094 32674 22146
rect 41470 22094 41522 22146
rect 44270 22094 44322 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 3838 21758 3890 21810
rect 6862 21758 6914 21810
rect 8654 21758 8706 21810
rect 16718 21758 16770 21810
rect 23102 21758 23154 21810
rect 23326 21758 23378 21810
rect 24334 21758 24386 21810
rect 24446 21758 24498 21810
rect 28814 21758 28866 21810
rect 29486 21758 29538 21810
rect 30158 21758 30210 21810
rect 31726 21758 31778 21810
rect 32398 21758 32450 21810
rect 33070 21758 33122 21810
rect 35534 21758 35586 21810
rect 38110 21758 38162 21810
rect 38782 21758 38834 21810
rect 41806 21758 41858 21810
rect 41918 21758 41970 21810
rect 47966 21758 48018 21810
rect 3166 21646 3218 21698
rect 3278 21646 3330 21698
rect 3502 21646 3554 21698
rect 4958 21646 5010 21698
rect 6078 21646 6130 21698
rect 6750 21646 6802 21698
rect 7534 21646 7586 21698
rect 8430 21646 8482 21698
rect 14030 21646 14082 21698
rect 14254 21646 14306 21698
rect 18062 21646 18114 21698
rect 23438 21646 23490 21698
rect 27358 21646 27410 21698
rect 30494 21646 30546 21698
rect 33406 21646 33458 21698
rect 34190 21646 34242 21698
rect 34638 21646 34690 21698
rect 39118 21646 39170 21698
rect 44494 21646 44546 21698
rect 44606 21646 44658 21698
rect 45614 21646 45666 21698
rect 3614 21534 3666 21586
rect 3950 21534 4002 21586
rect 4286 21534 4338 21586
rect 4510 21534 4562 21586
rect 5182 21534 5234 21586
rect 5854 21534 5906 21586
rect 6526 21534 6578 21586
rect 7870 21534 7922 21586
rect 8206 21534 8258 21586
rect 8878 21534 8930 21586
rect 10782 21534 10834 21586
rect 14814 21534 14866 21586
rect 15822 21534 15874 21586
rect 16382 21534 16434 21586
rect 16606 21534 16658 21586
rect 16942 21534 16994 21586
rect 22430 21534 22482 21586
rect 23998 21534 24050 21586
rect 24222 21534 24274 21586
rect 28030 21534 28082 21586
rect 28478 21534 28530 21586
rect 28814 21534 28866 21586
rect 29038 21534 29090 21586
rect 30830 21534 30882 21586
rect 31278 21534 31330 21586
rect 31838 21534 31890 21586
rect 32286 21534 32338 21586
rect 32510 21534 32562 21586
rect 33966 21534 34018 21586
rect 34414 21534 34466 21586
rect 35086 21534 35138 21586
rect 36318 21534 36370 21586
rect 37438 21534 37490 21586
rect 38334 21534 38386 21586
rect 41470 21534 41522 21586
rect 41694 21534 41746 21586
rect 42142 21534 42194 21586
rect 43038 21534 43090 21586
rect 44830 21534 44882 21586
rect 45054 21534 45106 21586
rect 45502 21534 45554 21586
rect 46062 21534 46114 21586
rect 46398 21534 46450 21586
rect 46734 21534 46786 21586
rect 47182 21534 47234 21586
rect 47294 21534 47346 21586
rect 4734 21422 4786 21474
rect 6302 21422 6354 21474
rect 9662 21422 9714 21474
rect 11454 21422 11506 21474
rect 13582 21422 13634 21474
rect 13918 21422 13970 21474
rect 14590 21422 14642 21474
rect 15598 21422 15650 21474
rect 25230 21422 25282 21474
rect 31054 21422 31106 21474
rect 34302 21422 34354 21474
rect 35982 21422 36034 21474
rect 36878 21422 36930 21474
rect 37214 21422 37266 21474
rect 37774 21422 37826 21474
rect 42478 21422 42530 21474
rect 42590 21422 42642 21474
rect 45278 21422 45330 21474
rect 46958 21422 47010 21474
rect 47742 21422 47794 21474
rect 47854 21422 47906 21474
rect 6862 21310 6914 21362
rect 15150 21310 15202 21362
rect 15486 21310 15538 21362
rect 23774 21310 23826 21362
rect 34974 21310 35026 21362
rect 42926 21310 42978 21362
rect 45950 21310 46002 21362
rect 46286 21310 46338 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 10782 20974 10834 21026
rect 19294 20974 19346 21026
rect 27134 20974 27186 21026
rect 29486 20974 29538 21026
rect 43934 20974 43986 21026
rect 44270 20974 44322 21026
rect 2494 20862 2546 20914
rect 4622 20862 4674 20914
rect 6414 20862 6466 20914
rect 8542 20862 8594 20914
rect 9662 20862 9714 20914
rect 11454 20862 11506 20914
rect 14702 20862 14754 20914
rect 18398 20862 18450 20914
rect 20638 20862 20690 20914
rect 32062 20862 32114 20914
rect 41806 20862 41858 20914
rect 42926 20862 42978 20914
rect 43710 20862 43762 20914
rect 46062 20862 46114 20914
rect 48190 20862 48242 20914
rect 1710 20750 1762 20802
rect 5742 20750 5794 20802
rect 11006 20750 11058 20802
rect 14142 20750 14194 20802
rect 14814 20750 14866 20802
rect 15150 20750 15202 20802
rect 17166 20750 17218 20802
rect 19966 20750 20018 20802
rect 21646 20750 21698 20802
rect 21982 20750 22034 20802
rect 23214 20750 23266 20802
rect 25118 20750 25170 20802
rect 26462 20750 26514 20802
rect 27806 20750 27858 20802
rect 33966 20750 34018 20802
rect 41694 20750 41746 20802
rect 45390 20750 45442 20802
rect 9214 20638 9266 20690
rect 9550 20638 9602 20690
rect 9998 20638 10050 20690
rect 15262 20638 15314 20690
rect 18286 20638 18338 20690
rect 19742 20638 19794 20690
rect 19854 20638 19906 20690
rect 21310 20638 21362 20690
rect 21422 20638 21474 20690
rect 21870 20638 21922 20690
rect 23550 20638 23602 20690
rect 25902 20638 25954 20690
rect 27582 20638 27634 20690
rect 27694 20638 27746 20690
rect 29598 20638 29650 20690
rect 29934 20638 29986 20690
rect 41246 20638 41298 20690
rect 41358 20638 41410 20690
rect 42142 20638 42194 20690
rect 42814 20638 42866 20690
rect 8990 20526 9042 20578
rect 9774 20526 9826 20578
rect 10446 20526 10498 20578
rect 14590 20526 14642 20578
rect 20750 20526 20802 20578
rect 22878 20526 22930 20578
rect 28366 20526 28418 20578
rect 30270 20526 30322 20578
rect 30718 20526 30770 20578
rect 31166 20526 31218 20578
rect 35534 20526 35586 20578
rect 36094 20526 36146 20578
rect 37214 20526 37266 20578
rect 41022 20526 41074 20578
rect 42254 20526 42306 20578
rect 42366 20526 42418 20578
rect 43374 20526 43426 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 9886 20190 9938 20242
rect 16270 20190 16322 20242
rect 33294 20190 33346 20242
rect 33630 20190 33682 20242
rect 41246 20190 41298 20242
rect 9774 20078 9826 20130
rect 12798 20078 12850 20130
rect 23102 20078 23154 20130
rect 23886 20078 23938 20130
rect 25902 20078 25954 20130
rect 30382 20078 30434 20130
rect 31838 20078 31890 20130
rect 33854 20078 33906 20130
rect 35310 20078 35362 20130
rect 41918 20078 41970 20130
rect 8206 19966 8258 20018
rect 9998 19966 10050 20018
rect 10446 19966 10498 20018
rect 15934 19966 15986 20018
rect 16606 19966 16658 20018
rect 16830 19966 16882 20018
rect 18846 19966 18898 20018
rect 23550 19966 23602 20018
rect 25566 19966 25618 20018
rect 26798 19966 26850 20018
rect 28366 19966 28418 20018
rect 33406 19966 33458 20018
rect 34302 19966 34354 20018
rect 36542 19966 36594 20018
rect 40014 19966 40066 20018
rect 40350 19966 40402 20018
rect 40910 19966 40962 20018
rect 41134 19966 41186 20018
rect 41358 19966 41410 20018
rect 41582 19966 41634 20018
rect 42142 19966 42194 20018
rect 43374 19966 43426 20018
rect 3390 19854 3442 19906
rect 8878 19854 8930 19906
rect 22430 19854 22482 19906
rect 24334 19854 24386 19906
rect 26350 19854 26402 19906
rect 29486 19854 29538 19906
rect 31502 19854 31554 19906
rect 32398 19854 32450 19906
rect 33518 19854 33570 19906
rect 34974 19854 35026 19906
rect 35982 19854 36034 19906
rect 36094 19854 36146 19906
rect 37214 19854 37266 19906
rect 39342 19854 39394 19906
rect 40238 19854 40290 19906
rect 42478 19854 42530 19906
rect 46846 19854 46898 19906
rect 8766 19742 8818 19794
rect 31950 19742 32002 19794
rect 32510 19742 32562 19794
rect 34638 19742 34690 19794
rect 35310 19742 35362 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 7086 19406 7138 19458
rect 7422 19406 7474 19458
rect 20750 19406 20802 19458
rect 31054 19406 31106 19458
rect 42590 19406 42642 19458
rect 4622 19294 4674 19346
rect 8990 19294 9042 19346
rect 11118 19294 11170 19346
rect 13470 19294 13522 19346
rect 15710 19294 15762 19346
rect 16382 19294 16434 19346
rect 18174 19294 18226 19346
rect 20302 19294 20354 19346
rect 20638 19294 20690 19346
rect 21422 19294 21474 19346
rect 23550 19294 23602 19346
rect 25678 19294 25730 19346
rect 27806 19294 27858 19346
rect 32622 19294 32674 19346
rect 34750 19294 34802 19346
rect 42030 19294 42082 19346
rect 44158 19294 44210 19346
rect 44942 19294 44994 19346
rect 46062 19294 46114 19346
rect 48190 19294 48242 19346
rect 1822 19182 1874 19234
rect 6526 19182 6578 19234
rect 6862 19182 6914 19234
rect 7646 19182 7698 19234
rect 8318 19182 8370 19234
rect 15262 19182 15314 19234
rect 17502 19182 17554 19234
rect 24334 19170 24386 19222
rect 24894 19182 24946 19234
rect 30046 19182 30098 19234
rect 30382 19182 30434 19234
rect 30718 19182 30770 19234
rect 31950 19182 32002 19234
rect 35422 19182 35474 19234
rect 37326 19182 37378 19234
rect 43934 19182 43986 19234
rect 44830 19182 44882 19234
rect 45390 19182 45442 19234
rect 2494 19070 2546 19122
rect 5630 19070 5682 19122
rect 13806 19070 13858 19122
rect 14814 19070 14866 19122
rect 29150 19070 29202 19122
rect 29710 19070 29762 19122
rect 30158 19070 30210 19122
rect 35534 19070 35586 19122
rect 35758 19070 35810 19122
rect 36206 19070 36258 19122
rect 42814 19070 42866 19122
rect 43262 19070 43314 19122
rect 5742 18958 5794 19010
rect 5854 18958 5906 19010
rect 6638 18958 6690 19010
rect 13582 18958 13634 19010
rect 14366 18958 14418 19010
rect 29262 18958 29314 19010
rect 29934 18958 29986 19010
rect 30942 18958 30994 19010
rect 31502 18958 31554 19010
rect 35198 18958 35250 19010
rect 35310 18958 35362 19010
rect 36318 18958 36370 19010
rect 42702 18958 42754 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 4398 18622 4450 18674
rect 4622 18622 4674 18674
rect 21870 18622 21922 18674
rect 24670 18622 24722 18674
rect 35646 18622 35698 18674
rect 36542 18622 36594 18674
rect 47518 18622 47570 18674
rect 17502 18510 17554 18562
rect 20974 18510 21026 18562
rect 28030 18510 28082 18562
rect 31166 18510 31218 18562
rect 31502 18510 31554 18562
rect 33630 18510 33682 18562
rect 33854 18510 33906 18562
rect 35422 18510 35474 18562
rect 35870 18510 35922 18562
rect 36430 18510 36482 18562
rect 47630 18510 47682 18562
rect 3166 18398 3218 18450
rect 3502 18398 3554 18450
rect 3726 18398 3778 18450
rect 4062 18398 4114 18450
rect 4510 18398 4562 18450
rect 5294 18398 5346 18450
rect 10670 18398 10722 18450
rect 11454 18398 11506 18450
rect 12126 18398 12178 18450
rect 17838 18398 17890 18450
rect 18622 18398 18674 18450
rect 20078 18398 20130 18450
rect 21310 18398 21362 18450
rect 22206 18398 22258 18450
rect 22654 18398 22706 18450
rect 23214 18398 23266 18450
rect 23550 18398 23602 18450
rect 25230 18398 25282 18450
rect 30942 18398 30994 18450
rect 31726 18398 31778 18450
rect 32286 18398 32338 18450
rect 34862 18398 34914 18450
rect 35198 18398 35250 18450
rect 35534 18398 35586 18450
rect 36766 18398 36818 18450
rect 37102 18398 37154 18450
rect 40910 18398 40962 18450
rect 44270 18398 44322 18450
rect 6078 18286 6130 18338
rect 8206 18286 8258 18338
rect 8654 18286 8706 18338
rect 14254 18286 14306 18338
rect 15710 18286 15762 18338
rect 16942 18286 16994 18338
rect 19966 18286 20018 18338
rect 24110 18286 24162 18338
rect 33182 18286 33234 18338
rect 34302 18286 34354 18338
rect 37774 18286 37826 18338
rect 39902 18286 39954 18338
rect 40238 18286 40290 18338
rect 41694 18286 41746 18338
rect 43822 18286 43874 18338
rect 44942 18286 44994 18338
rect 47070 18286 47122 18338
rect 48190 18286 48242 18338
rect 10670 18174 10722 18226
rect 11006 18174 11058 18226
rect 15934 18174 15986 18226
rect 16270 18174 16322 18226
rect 18286 18174 18338 18226
rect 33966 18174 34018 18226
rect 40350 18174 40402 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 23326 17838 23378 17890
rect 23662 17838 23714 17890
rect 24222 17838 24274 17890
rect 25342 17838 25394 17890
rect 43710 17838 43762 17890
rect 4622 17726 4674 17778
rect 10558 17726 10610 17778
rect 12686 17726 12738 17778
rect 14142 17726 14194 17778
rect 20862 17726 20914 17778
rect 23438 17726 23490 17778
rect 23886 17726 23938 17778
rect 24334 17726 24386 17778
rect 25342 17726 25394 17778
rect 28030 17726 28082 17778
rect 29150 17726 29202 17778
rect 33518 17726 33570 17778
rect 34526 17726 34578 17778
rect 37214 17726 37266 17778
rect 40910 17726 40962 17778
rect 43598 17726 43650 17778
rect 45726 17726 45778 17778
rect 46174 17726 46226 17778
rect 47182 17726 47234 17778
rect 1822 17614 1874 17666
rect 8878 17614 8930 17666
rect 9886 17614 9938 17666
rect 17054 17614 17106 17666
rect 19070 17614 19122 17666
rect 19630 17614 19682 17666
rect 25790 17614 25842 17666
rect 26350 17614 26402 17666
rect 27134 17614 27186 17666
rect 27694 17614 27746 17666
rect 32062 17614 32114 17666
rect 32398 17614 32450 17666
rect 33182 17614 33234 17666
rect 34862 17614 34914 17666
rect 35422 17614 35474 17666
rect 37886 17614 37938 17666
rect 43374 17614 43426 17666
rect 45278 17614 45330 17666
rect 45614 17614 45666 17666
rect 2494 17502 2546 17554
rect 9214 17502 9266 17554
rect 16270 17502 16322 17554
rect 17390 17502 17442 17554
rect 17502 17502 17554 17554
rect 17614 17502 17666 17554
rect 19966 17502 20018 17554
rect 21870 17502 21922 17554
rect 22430 17502 22482 17554
rect 22766 17502 22818 17554
rect 22990 17502 23042 17554
rect 25678 17502 25730 17554
rect 27246 17502 27298 17554
rect 28590 17502 28642 17554
rect 31278 17502 31330 17554
rect 36430 17502 36482 17554
rect 44158 17502 44210 17554
rect 46622 17502 46674 17554
rect 47854 17502 47906 17554
rect 48190 17502 48242 17554
rect 5630 17390 5682 17442
rect 5966 17390 6018 17442
rect 6974 17390 7026 17442
rect 9102 17390 9154 17442
rect 18174 17390 18226 17442
rect 18622 17390 18674 17442
rect 19630 17390 19682 17442
rect 21310 17390 21362 17442
rect 22654 17390 22706 17442
rect 24894 17390 24946 17442
rect 27358 17390 27410 17442
rect 28254 17390 28306 17442
rect 28478 17390 28530 17442
rect 32734 17390 32786 17442
rect 33966 17390 34018 17442
rect 36094 17390 36146 17442
rect 44046 17390 44098 17442
rect 45390 17390 45442 17442
rect 45726 17390 45778 17442
rect 46286 17390 46338 17442
rect 46734 17390 46786 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 9662 17054 9714 17106
rect 12014 17054 12066 17106
rect 16046 17054 16098 17106
rect 16270 17054 16322 17106
rect 20638 17054 20690 17106
rect 26910 17054 26962 17106
rect 31054 17054 31106 17106
rect 31838 17054 31890 17106
rect 40350 17054 40402 17106
rect 41134 17054 41186 17106
rect 42142 17054 42194 17106
rect 42590 17054 42642 17106
rect 3390 16942 3442 16994
rect 4062 16942 4114 16994
rect 4846 16942 4898 16994
rect 6862 16942 6914 16994
rect 13134 16942 13186 16994
rect 23662 16942 23714 16994
rect 29486 16942 29538 16994
rect 30830 16942 30882 16994
rect 31166 16942 31218 16994
rect 31950 16942 32002 16994
rect 32286 16942 32338 16994
rect 38670 16942 38722 16994
rect 39902 16942 39954 16994
rect 41582 16942 41634 16994
rect 4286 16830 4338 16882
rect 4510 16830 4562 16882
rect 5406 16830 5458 16882
rect 6078 16830 6130 16882
rect 9550 16830 9602 16882
rect 9774 16830 9826 16882
rect 10222 16830 10274 16882
rect 11342 16830 11394 16882
rect 11790 16830 11842 16882
rect 12350 16830 12402 16882
rect 15598 16830 15650 16882
rect 18062 16830 18114 16882
rect 18398 16830 18450 16882
rect 18622 16830 18674 16882
rect 19966 16830 20018 16882
rect 24446 16830 24498 16882
rect 25342 16830 25394 16882
rect 26014 16830 26066 16882
rect 30270 16830 30322 16882
rect 31278 16830 31330 16882
rect 31502 16830 31554 16882
rect 37886 16830 37938 16882
rect 38894 16830 38946 16882
rect 39566 16830 39618 16882
rect 40910 16830 40962 16882
rect 41358 16830 41410 16882
rect 42926 16830 42978 16882
rect 3278 16718 3330 16770
rect 4398 16718 4450 16770
rect 8990 16718 9042 16770
rect 11902 16718 11954 16770
rect 15262 16718 15314 16770
rect 16158 16718 16210 16770
rect 19518 16718 19570 16770
rect 21086 16718 21138 16770
rect 21534 16718 21586 16770
rect 26238 16718 26290 16770
rect 27358 16718 27410 16770
rect 35086 16718 35138 16770
rect 41022 16718 41074 16770
rect 44942 16718 44994 16770
rect 3614 16606 3666 16658
rect 5182 16606 5234 16658
rect 19070 16606 19122 16658
rect 19742 16606 19794 16658
rect 20414 16606 20466 16658
rect 25678 16606 25730 16658
rect 32398 16606 32450 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 9550 16270 9602 16322
rect 10110 16270 10162 16322
rect 34974 16270 35026 16322
rect 35310 16270 35362 16322
rect 3054 16158 3106 16210
rect 4846 16158 4898 16210
rect 5854 16158 5906 16210
rect 8990 16158 9042 16210
rect 9214 16158 9266 16210
rect 11118 16158 11170 16210
rect 12350 16158 12402 16210
rect 12910 16158 12962 16210
rect 19630 16158 19682 16210
rect 21982 16158 22034 16210
rect 23214 16158 23266 16210
rect 28142 16158 28194 16210
rect 29150 16158 29202 16210
rect 29374 16158 29426 16210
rect 29710 16158 29762 16210
rect 30382 16158 30434 16210
rect 30718 16158 30770 16210
rect 32846 16158 32898 16210
rect 34974 16158 35026 16210
rect 35870 16158 35922 16210
rect 36430 16158 36482 16210
rect 37774 16158 37826 16210
rect 39902 16184 39954 16236
rect 41134 16158 41186 16210
rect 41358 16158 41410 16210
rect 43486 16158 43538 16210
rect 44942 16158 44994 16210
rect 45278 16158 45330 16210
rect 47406 16158 47458 16210
rect 3390 16046 3442 16098
rect 3838 16046 3890 16098
rect 4398 16046 4450 16098
rect 6414 16046 6466 16098
rect 9886 16046 9938 16098
rect 11790 16046 11842 16098
rect 12686 16046 12738 16098
rect 13582 16046 13634 16098
rect 14478 16046 14530 16098
rect 15150 16046 15202 16098
rect 18174 16046 18226 16098
rect 18398 16046 18450 16098
rect 19070 16046 19122 16098
rect 19406 16046 19458 16098
rect 21198 16046 21250 16098
rect 21534 16046 21586 16098
rect 22318 16046 22370 16098
rect 23102 16046 23154 16098
rect 23326 16046 23378 16098
rect 23774 16046 23826 16098
rect 24558 16046 24610 16098
rect 25230 16046 25282 16098
rect 28590 16046 28642 16098
rect 33630 16046 33682 16098
rect 35422 16046 35474 16098
rect 35646 16046 35698 16098
rect 37102 16046 37154 16098
rect 44270 16046 44322 16098
rect 48078 16046 48130 16098
rect 3726 15934 3778 15986
rect 6190 15934 6242 15986
rect 12014 15934 12066 15986
rect 13918 15934 13970 15986
rect 14254 15934 14306 15986
rect 14814 15934 14866 15986
rect 20302 15934 20354 15986
rect 20526 15934 20578 15986
rect 21422 15934 21474 15986
rect 26014 15934 26066 15986
rect 28478 15934 28530 15986
rect 34526 15934 34578 15986
rect 35982 15934 36034 15986
rect 40574 15934 40626 15986
rect 3166 15822 3218 15874
rect 3950 15822 4002 15874
rect 10446 15822 10498 15874
rect 14478 15822 14530 15874
rect 15486 15822 15538 15874
rect 17950 15822 18002 15874
rect 18286 15822 18338 15874
rect 19070 15822 19122 15874
rect 20414 15822 20466 15874
rect 23998 15822 24050 15874
rect 29598 15822 29650 15874
rect 29822 15822 29874 15874
rect 30270 15822 30322 15874
rect 33966 15822 34018 15874
rect 40238 15822 40290 15874
rect 44830 15822 44882 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 5742 15486 5794 15538
rect 9550 15486 9602 15538
rect 9774 15486 9826 15538
rect 10670 15486 10722 15538
rect 11342 15486 11394 15538
rect 11790 15486 11842 15538
rect 18398 15486 18450 15538
rect 18846 15486 18898 15538
rect 20974 15486 21026 15538
rect 21870 15486 21922 15538
rect 22878 15486 22930 15538
rect 23438 15486 23490 15538
rect 24110 15486 24162 15538
rect 24446 15486 24498 15538
rect 29038 15486 29090 15538
rect 29262 15486 29314 15538
rect 31614 15486 31666 15538
rect 31838 15486 31890 15538
rect 33854 15486 33906 15538
rect 35422 15486 35474 15538
rect 36542 15486 36594 15538
rect 39118 15486 39170 15538
rect 40014 15486 40066 15538
rect 2494 15374 2546 15426
rect 15710 15374 15762 15426
rect 19742 15374 19794 15426
rect 19966 15374 20018 15426
rect 20750 15374 20802 15426
rect 26126 15374 26178 15426
rect 26910 15374 26962 15426
rect 27022 15374 27074 15426
rect 27134 15374 27186 15426
rect 28702 15374 28754 15426
rect 29374 15374 29426 15426
rect 31278 15374 31330 15426
rect 31726 15374 31778 15426
rect 33518 15374 33570 15426
rect 35086 15374 35138 15426
rect 36094 15374 36146 15426
rect 36990 15374 37042 15426
rect 38334 15374 38386 15426
rect 47406 15374 47458 15426
rect 1822 15262 1874 15314
rect 5518 15262 5570 15314
rect 6078 15262 6130 15314
rect 6862 15262 6914 15314
rect 10222 15262 10274 15314
rect 10558 15262 10610 15314
rect 11566 15262 11618 15314
rect 16382 15262 16434 15314
rect 19518 15262 19570 15314
rect 20190 15262 20242 15314
rect 20638 15262 20690 15314
rect 21198 15262 21250 15314
rect 22430 15262 22482 15314
rect 23550 15262 23602 15314
rect 25566 15262 25618 15314
rect 26014 15262 26066 15314
rect 27694 15262 27746 15314
rect 27918 15262 27970 15314
rect 28142 15262 28194 15314
rect 28590 15262 28642 15314
rect 30046 15262 30098 15314
rect 30606 15262 30658 15314
rect 31502 15262 31554 15314
rect 34190 15262 34242 15314
rect 34750 15262 34802 15314
rect 35870 15262 35922 15314
rect 37438 15262 37490 15314
rect 38558 15262 38610 15314
rect 43822 15262 43874 15314
rect 48078 15262 48130 15314
rect 4622 15150 4674 15202
rect 8990 15150 9042 15202
rect 9662 15150 9714 15202
rect 10446 15150 10498 15202
rect 11678 15150 11730 15202
rect 13582 15150 13634 15202
rect 18734 15150 18786 15202
rect 20862 15150 20914 15202
rect 25790 15150 25842 15202
rect 26462 15150 26514 15202
rect 28478 15150 28530 15202
rect 37774 15150 37826 15202
rect 39566 15150 39618 15202
rect 40910 15150 40962 15202
rect 43038 15150 43090 15202
rect 44718 15150 44770 15202
rect 45278 15150 45330 15202
rect 19182 15038 19234 15090
rect 23438 15038 23490 15090
rect 27582 15038 27634 15090
rect 39454 15038 39506 15090
rect 44606 15038 44658 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 3502 14702 3554 14754
rect 3838 14702 3890 14754
rect 11790 14702 11842 14754
rect 19630 14702 19682 14754
rect 28254 14702 28306 14754
rect 4062 14590 4114 14642
rect 6078 14590 6130 14642
rect 14926 14590 14978 14642
rect 18734 14590 18786 14642
rect 21310 14590 21362 14642
rect 23438 14590 23490 14642
rect 24670 14590 24722 14642
rect 25006 14590 25058 14642
rect 27134 14590 27186 14642
rect 29710 14590 29762 14642
rect 34750 14590 34802 14642
rect 38222 14590 38274 14642
rect 42590 14590 42642 14642
rect 43374 14590 43426 14642
rect 45726 14590 45778 14642
rect 4398 14478 4450 14530
rect 10894 14478 10946 14530
rect 11566 14478 11618 14530
rect 15038 14478 15090 14530
rect 15486 14478 15538 14530
rect 15934 14478 15986 14530
rect 19406 14478 19458 14530
rect 19854 14478 19906 14530
rect 24110 14478 24162 14530
rect 27806 14478 27858 14530
rect 29374 14478 29426 14530
rect 30606 14478 30658 14530
rect 35310 14478 35362 14530
rect 35870 14478 35922 14530
rect 36542 14478 36594 14530
rect 37214 14478 37266 14530
rect 37998 14478 38050 14530
rect 38334 14478 38386 14530
rect 39006 14478 39058 14530
rect 39342 14478 39394 14530
rect 39902 14478 39954 14530
rect 40238 14478 40290 14530
rect 40462 14478 40514 14530
rect 42926 14478 42978 14530
rect 43150 14478 43202 14530
rect 43486 14478 43538 14530
rect 45278 14478 45330 14530
rect 45390 14478 45442 14530
rect 45614 14478 45666 14530
rect 46958 14478 47010 14530
rect 4846 14366 4898 14418
rect 12126 14366 12178 14418
rect 12574 14366 12626 14418
rect 13470 14366 13522 14418
rect 13582 14366 13634 14418
rect 14814 14366 14866 14418
rect 16606 14366 16658 14418
rect 4510 14254 4562 14306
rect 4622 14254 4674 14306
rect 10894 14254 10946 14306
rect 11342 14254 11394 14306
rect 12910 14254 12962 14306
rect 19182 14366 19234 14418
rect 19406 14366 19458 14418
rect 20302 14366 20354 14418
rect 29486 14366 29538 14418
rect 30158 14366 30210 14418
rect 35982 14366 36034 14418
rect 37102 14366 37154 14418
rect 37326 14366 37378 14418
rect 40798 14366 40850 14418
rect 41134 14366 41186 14418
rect 41470 14366 41522 14418
rect 43934 14366 43986 14418
rect 46174 14366 46226 14418
rect 13806 14254 13858 14306
rect 18958 14254 19010 14306
rect 19518 14254 19570 14306
rect 20414 14254 20466 14306
rect 20526 14254 20578 14306
rect 28366 14254 28418 14306
rect 28478 14254 28530 14306
rect 35086 14254 35138 14306
rect 36094 14254 36146 14306
rect 37774 14254 37826 14306
rect 38558 14254 38610 14306
rect 42030 14254 42082 14306
rect 43374 14254 43426 14306
rect 44046 14254 44098 14306
rect 44270 14254 44322 14306
rect 45726 14254 45778 14306
rect 46510 14254 46562 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 6526 13918 6578 13970
rect 10894 13918 10946 13970
rect 15710 13918 15762 13970
rect 18398 13918 18450 13970
rect 25902 13918 25954 13970
rect 27470 13918 27522 13970
rect 28030 13918 28082 13970
rect 28366 13918 28418 13970
rect 28702 13918 28754 13970
rect 31950 13918 32002 13970
rect 41022 13918 41074 13970
rect 42590 13918 42642 13970
rect 44494 13918 44546 13970
rect 11902 13806 11954 13858
rect 14030 13806 14082 13858
rect 17950 13806 18002 13858
rect 18958 13806 19010 13858
rect 21758 13806 21810 13858
rect 27806 13806 27858 13858
rect 28254 13806 28306 13858
rect 29934 13806 29986 13858
rect 30606 13806 30658 13858
rect 36318 13806 36370 13858
rect 39230 13806 39282 13858
rect 39454 13806 39506 13858
rect 47406 13806 47458 13858
rect 1822 13694 1874 13746
rect 4958 13694 5010 13746
rect 5182 13694 5234 13746
rect 7086 13694 7138 13746
rect 7534 13694 7586 13746
rect 10222 13694 10274 13746
rect 11230 13694 11282 13746
rect 12238 13694 12290 13746
rect 14142 13694 14194 13746
rect 14590 13694 14642 13746
rect 17838 13694 17890 13746
rect 23886 13694 23938 13746
rect 26238 13694 26290 13746
rect 26462 13694 26514 13746
rect 27694 13694 27746 13746
rect 28590 13694 28642 13746
rect 28814 13694 28866 13746
rect 30158 13694 30210 13746
rect 30718 13694 30770 13746
rect 31390 13694 31442 13746
rect 31614 13694 31666 13746
rect 31838 13694 31890 13746
rect 33182 13694 33234 13746
rect 35534 13694 35586 13746
rect 39118 13694 39170 13746
rect 39678 13694 39730 13746
rect 42814 13694 42866 13746
rect 43822 13694 43874 13746
rect 43934 13694 43986 13746
rect 44046 13694 44098 13746
rect 48078 13694 48130 13746
rect 2494 13582 2546 13634
rect 4622 13582 4674 13634
rect 12014 13582 12066 13634
rect 13806 13582 13858 13634
rect 25342 13582 25394 13634
rect 31726 13582 31778 13634
rect 32398 13582 32450 13634
rect 34302 13582 34354 13634
rect 38446 13582 38498 13634
rect 40126 13582 40178 13634
rect 41694 13582 41746 13634
rect 43038 13582 43090 13634
rect 43374 13582 43426 13634
rect 45278 13582 45330 13634
rect 5518 13470 5570 13522
rect 6862 13470 6914 13522
rect 10334 13470 10386 13522
rect 14814 13470 14866 13522
rect 17950 13470 18002 13522
rect 18734 13470 18786 13522
rect 32510 13470 32562 13522
rect 34190 13470 34242 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 3726 13134 3778 13186
rect 4062 13134 4114 13186
rect 38110 13134 38162 13186
rect 7086 13022 7138 13074
rect 7758 13022 7810 13074
rect 9102 13022 9154 13074
rect 11230 13022 11282 13074
rect 12126 13022 12178 13074
rect 13694 13022 13746 13074
rect 15150 13022 15202 13074
rect 16270 13022 16322 13074
rect 18734 13022 18786 13074
rect 21310 13022 21362 13074
rect 22430 13022 22482 13074
rect 23326 13022 23378 13074
rect 23774 13022 23826 13074
rect 29374 13022 29426 13074
rect 29710 13022 29762 13074
rect 31054 13022 31106 13074
rect 33182 13022 33234 13074
rect 34414 13022 34466 13074
rect 38894 13022 38946 13074
rect 40462 13022 40514 13074
rect 6302 12910 6354 12962
rect 6750 12910 6802 12962
rect 6862 12910 6914 12962
rect 8318 12910 8370 12962
rect 11678 12910 11730 12962
rect 12686 12910 12738 12962
rect 14030 12910 14082 12962
rect 17726 12910 17778 12962
rect 17950 12910 18002 12962
rect 18286 12910 18338 12962
rect 18958 12910 19010 12962
rect 19854 12910 19906 12962
rect 20302 12910 20354 12962
rect 23102 12910 23154 12962
rect 24334 12910 24386 12962
rect 26014 12910 26066 12962
rect 26238 12910 26290 12962
rect 26574 12910 26626 12962
rect 29150 12910 29202 12962
rect 33854 12910 33906 12962
rect 34750 12910 34802 12962
rect 38222 12910 38274 12962
rect 40574 12910 40626 12962
rect 41918 12910 41970 12962
rect 42478 12910 42530 12962
rect 42702 12910 42754 12962
rect 43598 12910 43650 12962
rect 44046 12910 44098 12962
rect 44270 12910 44322 12962
rect 45166 12910 45218 12962
rect 45390 12910 45442 12962
rect 3838 12798 3890 12850
rect 4734 12798 4786 12850
rect 5070 12798 5122 12850
rect 5630 12798 5682 12850
rect 7198 12798 7250 12850
rect 14478 12798 14530 12850
rect 14814 12798 14866 12850
rect 15038 12798 15090 12850
rect 18174 12798 18226 12850
rect 19070 12798 19122 12850
rect 26910 12798 26962 12850
rect 27022 12798 27074 12850
rect 34974 12798 35026 12850
rect 40014 12798 40066 12850
rect 45726 12798 45778 12850
rect 46062 12798 46114 12850
rect 47854 12798 47906 12850
rect 5742 12686 5794 12738
rect 5854 12686 5906 12738
rect 12462 12686 12514 12738
rect 15598 12686 15650 12738
rect 17614 12686 17666 12738
rect 20862 12686 20914 12738
rect 21870 12686 21922 12738
rect 24110 12686 24162 12738
rect 25454 12686 25506 12738
rect 25678 12686 25730 12738
rect 25902 12686 25954 12738
rect 26462 12686 26514 12738
rect 29598 12686 29650 12738
rect 29822 12686 29874 12738
rect 34414 12686 34466 12738
rect 34526 12686 34578 12738
rect 40126 12686 40178 12738
rect 42142 12686 42194 12738
rect 42926 12686 42978 12738
rect 43038 12686 43090 12738
rect 46398 12686 46450 12738
rect 47630 12686 47682 12738
rect 48190 12686 48242 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 5294 12350 5346 12402
rect 9886 12350 9938 12402
rect 11342 12350 11394 12402
rect 16718 12350 16770 12402
rect 31166 12350 31218 12402
rect 31390 12350 31442 12402
rect 32062 12350 32114 12402
rect 41134 12350 41186 12402
rect 41358 12350 41410 12402
rect 42254 12350 42306 12402
rect 42478 12350 42530 12402
rect 5406 12238 5458 12290
rect 8094 12238 8146 12290
rect 9550 12238 9602 12290
rect 11678 12238 11730 12290
rect 12014 12238 12066 12290
rect 15486 12238 15538 12290
rect 17614 12238 17666 12290
rect 17950 12238 18002 12290
rect 22542 12238 22594 12290
rect 25790 12238 25842 12290
rect 26686 12238 26738 12290
rect 29038 12238 29090 12290
rect 31278 12238 31330 12290
rect 40126 12238 40178 12290
rect 43598 12238 43650 12290
rect 47406 12238 47458 12290
rect 1822 12126 1874 12178
rect 4958 12126 5010 12178
rect 5630 12126 5682 12178
rect 8766 12126 8818 12178
rect 10334 12126 10386 12178
rect 10782 12126 10834 12178
rect 12350 12126 12402 12178
rect 16270 12126 16322 12178
rect 16606 12126 16658 12178
rect 16942 12126 16994 12178
rect 17390 12126 17442 12178
rect 21422 12126 21474 12178
rect 21758 12126 21810 12178
rect 25566 12126 25618 12178
rect 26238 12126 26290 12178
rect 26798 12126 26850 12178
rect 30382 12126 30434 12178
rect 30942 12126 30994 12178
rect 31614 12126 31666 12178
rect 33294 12126 33346 12178
rect 34078 12126 34130 12178
rect 37326 12126 37378 12178
rect 37774 12126 37826 12178
rect 37998 12126 38050 12178
rect 39006 12126 39058 12178
rect 39230 12126 39282 12178
rect 39454 12126 39506 12178
rect 39678 12126 39730 12178
rect 40014 12126 40066 12178
rect 40910 12126 40962 12178
rect 41582 12126 41634 12178
rect 42702 12126 42754 12178
rect 43486 12126 43538 12178
rect 43934 12126 43986 12178
rect 44158 12126 44210 12178
rect 48078 12126 48130 12178
rect 2494 12014 2546 12066
rect 4622 12014 4674 12066
rect 5966 12014 6018 12066
rect 12798 12014 12850 12066
rect 13358 12014 13410 12066
rect 17838 12014 17890 12066
rect 18510 12014 18562 12066
rect 20638 12014 20690 12066
rect 24670 12014 24722 12066
rect 26462 12014 26514 12066
rect 28926 12014 28978 12066
rect 36206 12014 36258 12066
rect 36654 12014 36706 12066
rect 37550 12014 37602 12066
rect 37886 12014 37938 12066
rect 39342 12014 39394 12066
rect 41022 12014 41074 12066
rect 44942 12014 44994 12066
rect 45278 12014 45330 12066
rect 25230 11902 25282 11954
rect 30494 11902 30546 11954
rect 36542 11902 36594 11954
rect 44494 11902 44546 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 3614 11566 3666 11618
rect 6414 11566 6466 11618
rect 24110 11566 24162 11618
rect 42254 11566 42306 11618
rect 43822 11566 43874 11618
rect 45054 11566 45106 11618
rect 4398 11454 4450 11506
rect 10222 11454 10274 11506
rect 16718 11454 16770 11506
rect 18846 11454 18898 11506
rect 22206 11454 22258 11506
rect 26462 11454 26514 11506
rect 28590 11454 28642 11506
rect 29598 11454 29650 11506
rect 30270 11454 30322 11506
rect 42142 11454 42194 11506
rect 3390 11342 3442 11394
rect 4286 11342 4338 11394
rect 4622 11342 4674 11394
rect 4846 11342 4898 11394
rect 5630 11342 5682 11394
rect 5854 11342 5906 11394
rect 5966 11342 6018 11394
rect 7310 11342 7362 11394
rect 10894 11342 10946 11394
rect 11118 11342 11170 11394
rect 12126 11342 12178 11394
rect 15374 11342 15426 11394
rect 16046 11342 16098 11394
rect 21870 11342 21922 11394
rect 23214 11342 23266 11394
rect 23326 11342 23378 11394
rect 23438 11342 23490 11394
rect 23774 11342 23826 11394
rect 25790 11342 25842 11394
rect 30494 11342 30546 11394
rect 36430 11342 36482 11394
rect 36990 11342 37042 11394
rect 37774 11342 37826 11394
rect 38446 11342 38498 11394
rect 39342 11342 39394 11394
rect 40798 11342 40850 11394
rect 42702 11342 42754 11394
rect 42814 11342 42866 11394
rect 43150 11342 43202 11394
rect 44830 11342 44882 11394
rect 45278 11342 45330 11394
rect 45502 11342 45554 11394
rect 46734 11342 46786 11394
rect 8094 11230 8146 11282
rect 11566 11230 11618 11282
rect 11678 11230 11730 11282
rect 12238 11230 12290 11282
rect 15598 11230 15650 11282
rect 29934 11230 29986 11282
rect 31950 11230 32002 11282
rect 37102 11230 37154 11282
rect 37662 11230 37714 11282
rect 38670 11230 38722 11282
rect 40238 11230 40290 11282
rect 43038 11230 43090 11282
rect 43934 11230 43986 11282
rect 45614 11230 45666 11282
rect 45950 11230 46002 11282
rect 3950 11118 4002 11170
rect 10670 11118 10722 11170
rect 11006 11118 11058 11170
rect 11902 11118 11954 11170
rect 12350 11118 12402 11170
rect 12574 11118 12626 11170
rect 22766 11118 22818 11170
rect 30830 11118 30882 11170
rect 37326 11118 37378 11170
rect 38222 11118 38274 11170
rect 40126 11118 40178 11170
rect 40350 11118 40402 11170
rect 41806 11118 41858 11170
rect 43598 11118 43650 11170
rect 46286 11118 46338 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 6526 10782 6578 10834
rect 9662 10782 9714 10834
rect 12574 10782 12626 10834
rect 21534 10782 21586 10834
rect 33406 10782 33458 10834
rect 33630 10782 33682 10834
rect 33742 10782 33794 10834
rect 37662 10782 37714 10834
rect 38334 10782 38386 10834
rect 39230 10782 39282 10834
rect 39790 10782 39842 10834
rect 42030 10782 42082 10834
rect 5182 10670 5234 10722
rect 9550 10670 9602 10722
rect 9886 10670 9938 10722
rect 10110 10670 10162 10722
rect 15038 10670 15090 10722
rect 31278 10670 31330 10722
rect 32510 10670 32562 10722
rect 33966 10670 34018 10722
rect 39902 10670 39954 10722
rect 40238 10670 40290 10722
rect 40910 10670 40962 10722
rect 41470 10670 41522 10722
rect 42478 10670 42530 10722
rect 47966 10670 48018 10722
rect 4622 10558 4674 10610
rect 6750 10558 6802 10610
rect 7198 10558 7250 10610
rect 12238 10558 12290 10610
rect 12686 10558 12738 10610
rect 15262 10558 15314 10610
rect 18174 10558 18226 10610
rect 21310 10558 21362 10610
rect 25342 10558 25394 10610
rect 25566 10558 25618 10610
rect 25790 10558 25842 10610
rect 31950 10558 32002 10610
rect 33518 10558 33570 10610
rect 36430 10558 36482 10610
rect 37102 10558 37154 10610
rect 37998 10558 38050 10610
rect 38334 10558 38386 10610
rect 38670 10558 38722 10610
rect 39566 10558 39618 10610
rect 41246 10558 41298 10610
rect 43486 10558 43538 10610
rect 1710 10446 1762 10498
rect 3838 10446 3890 10498
rect 5070 10446 5122 10498
rect 6638 10446 6690 10498
rect 18846 10446 18898 10498
rect 20974 10446 21026 10498
rect 21422 10446 21474 10498
rect 25678 10446 25730 10498
rect 29150 10446 29202 10498
rect 34302 10446 34354 10498
rect 37438 10446 37490 10498
rect 39006 10446 39058 10498
rect 4958 10334 5010 10386
rect 12462 10334 12514 10386
rect 32398 10334 32450 10386
rect 39118 10446 39170 10498
rect 40350 10446 40402 10498
rect 41022 10446 41074 10498
rect 42142 10446 42194 10498
rect 37886 10334 37938 10386
rect 41582 10334 41634 10386
rect 41806 10334 41858 10386
rect 42590 10334 42642 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 12238 9998 12290 10050
rect 13582 9998 13634 10050
rect 18846 9998 18898 10050
rect 27918 9998 27970 10050
rect 37214 9998 37266 10050
rect 37550 9998 37602 10050
rect 39342 9998 39394 10050
rect 41582 9998 41634 10050
rect 3502 9886 3554 9938
rect 4398 9886 4450 9938
rect 8542 9886 8594 9938
rect 11342 9886 11394 9938
rect 13694 9886 13746 9938
rect 14814 9886 14866 9938
rect 16942 9886 16994 9938
rect 23438 9886 23490 9938
rect 23886 9886 23938 9938
rect 25006 9886 25058 9938
rect 27134 9886 27186 9938
rect 31502 9886 31554 9938
rect 33630 9886 33682 9938
rect 35086 9886 35138 9938
rect 37550 9886 37602 9938
rect 38894 9886 38946 9938
rect 45054 9886 45106 9938
rect 45278 9886 45330 9938
rect 47406 9886 47458 9938
rect 3390 9774 3442 9826
rect 3614 9774 3666 9826
rect 4062 9774 4114 9826
rect 5630 9774 5682 9826
rect 10446 9774 10498 9826
rect 10670 9774 10722 9826
rect 11006 9774 11058 9826
rect 12574 9774 12626 9826
rect 14142 9774 14194 9826
rect 17502 9774 17554 9826
rect 18062 9774 18114 9826
rect 18846 9774 18898 9826
rect 21310 9774 21362 9826
rect 21870 9774 21922 9826
rect 24222 9774 24274 9826
rect 27582 9774 27634 9826
rect 27806 9774 27858 9826
rect 30718 9774 30770 9826
rect 34862 9774 34914 9826
rect 34974 9774 35026 9826
rect 35422 9774 35474 9826
rect 35758 9774 35810 9826
rect 35982 9774 36034 9826
rect 36206 9774 36258 9826
rect 36430 9774 36482 9826
rect 39118 9774 39170 9826
rect 40798 9774 40850 9826
rect 41470 9774 41522 9826
rect 42030 9774 42082 9826
rect 43374 9774 43426 9826
rect 44270 9774 44322 9826
rect 48078 9774 48130 9826
rect 6414 9662 6466 9714
rect 19182 9662 19234 9714
rect 22654 9662 22706 9714
rect 27470 9662 27522 9714
rect 41022 9662 41074 9714
rect 43822 9662 43874 9714
rect 10782 9550 10834 9602
rect 12350 9550 12402 9602
rect 17278 9550 17330 9602
rect 21534 9550 21586 9602
rect 21646 9550 21698 9602
rect 21758 9550 21810 9602
rect 22766 9550 22818 9602
rect 34414 9550 34466 9602
rect 35198 9550 35250 9602
rect 36094 9550 36146 9602
rect 37102 9550 37154 9602
rect 39790 9550 39842 9602
rect 42926 9550 42978 9602
rect 43150 9550 43202 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 6302 9214 6354 9266
rect 9662 9214 9714 9266
rect 10782 9214 10834 9266
rect 10894 9214 10946 9266
rect 16270 9214 16322 9266
rect 16830 9214 16882 9266
rect 24782 9214 24834 9266
rect 25790 9214 25842 9266
rect 26014 9214 26066 9266
rect 32510 9214 32562 9266
rect 39566 9214 39618 9266
rect 40238 9214 40290 9266
rect 40910 9214 40962 9266
rect 42926 9214 42978 9266
rect 6078 9102 6130 9154
rect 6414 9102 6466 9154
rect 6638 9102 6690 9154
rect 7198 9102 7250 9154
rect 7310 9102 7362 9154
rect 12350 9102 12402 9154
rect 15934 9102 15986 9154
rect 25678 9046 25730 9098
rect 25902 9102 25954 9154
rect 28702 9102 28754 9154
rect 35198 9102 35250 9154
rect 35310 9102 35362 9154
rect 36430 9102 36482 9154
rect 40350 9102 40402 9154
rect 41134 9102 41186 9154
rect 41358 9102 41410 9154
rect 43038 9102 43090 9154
rect 6974 8990 7026 9042
rect 10334 8990 10386 9042
rect 10670 8990 10722 9042
rect 11566 8990 11618 9042
rect 17390 8990 17442 9042
rect 24110 8990 24162 9042
rect 25230 8990 25282 9042
rect 26798 8990 26850 9042
rect 27022 8990 27074 9042
rect 27134 8990 27186 9042
rect 27918 8990 27970 9042
rect 33294 8990 33346 9042
rect 33518 8990 33570 9042
rect 35646 8990 35698 9042
rect 39678 8990 39730 9042
rect 40014 8990 40066 9042
rect 41918 8990 41970 9042
rect 42030 8990 42082 9042
rect 42142 8990 42194 9042
rect 42254 8990 42306 9042
rect 42478 8990 42530 9042
rect 43150 8990 43202 9042
rect 43374 8990 43426 9042
rect 44270 8990 44322 9042
rect 48078 8990 48130 9042
rect 4062 8878 4114 8930
rect 14478 8878 14530 8930
rect 18174 8878 18226 8930
rect 20302 8878 20354 8930
rect 20862 8878 20914 8930
rect 21198 8878 21250 8930
rect 23326 8878 23378 8930
rect 30830 8878 30882 8930
rect 34078 8878 34130 8930
rect 34750 8878 34802 8930
rect 38558 8878 38610 8930
rect 41022 8878 41074 8930
rect 44158 8878 44210 8930
rect 44942 8878 44994 8930
rect 45278 8878 45330 8930
rect 47406 8878 47458 8930
rect 3502 8766 3554 8818
rect 3838 8766 3890 8818
rect 7758 8766 7810 8818
rect 27582 8766 27634 8818
rect 34862 8766 34914 8818
rect 43598 8766 43650 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 13582 8430 13634 8482
rect 18398 8430 18450 8482
rect 40350 8430 40402 8482
rect 44158 8430 44210 8482
rect 47182 8430 47234 8482
rect 4622 8318 4674 8370
rect 5854 8318 5906 8370
rect 12126 8318 12178 8370
rect 16718 8318 16770 8370
rect 18734 8318 18786 8370
rect 20190 8318 20242 8370
rect 21422 8318 21474 8370
rect 23774 8318 23826 8370
rect 24110 8318 24162 8370
rect 24558 8318 24610 8370
rect 27470 8318 27522 8370
rect 29262 8318 29314 8370
rect 30382 8318 30434 8370
rect 34302 8318 34354 8370
rect 35646 8318 35698 8370
rect 37214 8318 37266 8370
rect 37438 8318 37490 8370
rect 38334 8318 38386 8370
rect 40238 8318 40290 8370
rect 41582 8318 41634 8370
rect 43822 8318 43874 8370
rect 1822 8206 1874 8258
rect 10894 8206 10946 8258
rect 11902 8206 11954 8258
rect 12910 8206 12962 8258
rect 13694 8206 13746 8258
rect 16270 8206 16322 8258
rect 18062 8206 18114 8258
rect 18398 8206 18450 8258
rect 19630 8206 19682 8258
rect 20638 8206 20690 8258
rect 21534 8206 21586 8258
rect 21982 8206 22034 8258
rect 22766 8206 22818 8258
rect 22990 8206 23042 8258
rect 23214 8206 23266 8258
rect 25902 8206 25954 8258
rect 26238 8206 26290 8258
rect 27694 8206 27746 8258
rect 29150 8206 29202 8258
rect 29598 8206 29650 8258
rect 31502 8206 31554 8258
rect 35086 8206 35138 8258
rect 35198 8206 35250 8258
rect 36430 8206 36482 8258
rect 36990 8206 37042 8258
rect 38782 8206 38834 8258
rect 40126 8206 40178 8258
rect 40910 8206 40962 8258
rect 41246 8206 41298 8258
rect 42142 8206 42194 8258
rect 43598 8206 43650 8258
rect 45278 8262 45330 8314
rect 45502 8318 45554 8370
rect 46846 8318 46898 8370
rect 2494 8094 2546 8146
rect 11230 8094 11282 8146
rect 17278 8094 17330 8146
rect 20302 8094 20354 8146
rect 21422 8094 21474 8146
rect 22542 8094 22594 8146
rect 23886 8094 23938 8146
rect 25230 8094 25282 8146
rect 25566 8094 25618 8146
rect 25678 8094 25730 8146
rect 26798 8094 26850 8146
rect 28478 8094 28530 8146
rect 28590 8094 28642 8146
rect 29486 8094 29538 8146
rect 30046 8094 30098 8146
rect 32174 8094 32226 8146
rect 37662 8094 37714 8146
rect 37886 8094 37938 8146
rect 42366 8094 42418 8146
rect 42590 8094 42642 8146
rect 42814 8094 42866 8146
rect 43150 8094 43202 8146
rect 43262 8094 43314 8146
rect 45838 8094 45890 8146
rect 46174 8094 46226 8146
rect 46510 8094 46562 8146
rect 47854 8094 47906 8146
rect 5070 7982 5122 8034
rect 12574 7982 12626 8034
rect 13582 7982 13634 8034
rect 16046 7982 16098 8034
rect 16158 7982 16210 8034
rect 16718 7982 16770 8034
rect 16830 7982 16882 8034
rect 17054 7982 17106 8034
rect 17838 7982 17890 8034
rect 17950 7982 18002 8034
rect 19406 7982 19458 8034
rect 20190 7982 20242 8034
rect 20526 7982 20578 8034
rect 21758 7982 21810 8034
rect 23326 7982 23378 8034
rect 26462 7982 26514 8034
rect 28254 7982 28306 8034
rect 30270 7982 30322 8034
rect 34750 7982 34802 8034
rect 34862 7982 34914 8034
rect 34974 7982 35026 8034
rect 35758 7982 35810 8034
rect 36094 7982 36146 8034
rect 37550 7982 37602 8034
rect 44942 7982 44994 8034
rect 47070 7982 47122 8034
rect 47518 7982 47570 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 3502 7646 3554 7698
rect 3726 7646 3778 7698
rect 4622 7646 4674 7698
rect 22990 7646 23042 7698
rect 32398 7646 32450 7698
rect 39454 7646 39506 7698
rect 41470 7646 41522 7698
rect 42478 7646 42530 7698
rect 42814 7646 42866 7698
rect 44718 7646 44770 7698
rect 2942 7534 2994 7586
rect 8990 7534 9042 7586
rect 12798 7534 12850 7586
rect 14590 7534 14642 7586
rect 17614 7534 17666 7586
rect 23774 7534 23826 7586
rect 24110 7534 24162 7586
rect 31166 7534 31218 7586
rect 32510 7534 32562 7586
rect 33518 7534 33570 7586
rect 35534 7534 35586 7586
rect 43374 7534 43426 7586
rect 47406 7534 47458 7586
rect 4174 7422 4226 7474
rect 4398 7422 4450 7474
rect 5070 7422 5122 7474
rect 5518 7422 5570 7474
rect 8654 7422 8706 7474
rect 9662 7422 9714 7474
rect 13022 7422 13074 7474
rect 13806 7422 13858 7474
rect 22654 7422 22706 7474
rect 23326 7422 23378 7474
rect 23998 7422 24050 7474
rect 25566 7422 25618 7474
rect 31950 7422 32002 7474
rect 33294 7422 33346 7474
rect 37662 7422 37714 7474
rect 41358 7422 41410 7474
rect 41582 7422 41634 7474
rect 41694 7422 41746 7474
rect 43262 7422 43314 7474
rect 43598 7422 43650 7474
rect 43822 7422 43874 7474
rect 44382 7422 44434 7474
rect 44830 7422 44882 7474
rect 48078 7422 48130 7474
rect 2830 7310 2882 7362
rect 3614 7310 3666 7362
rect 4510 7310 4562 7362
rect 6190 7310 6242 7362
rect 8318 7310 8370 7362
rect 8878 7310 8930 7362
rect 10334 7310 10386 7362
rect 12462 7310 12514 7362
rect 16718 7310 16770 7362
rect 26238 7310 26290 7362
rect 28366 7310 28418 7362
rect 29038 7310 29090 7362
rect 39566 7310 39618 7362
rect 40014 7310 40066 7362
rect 44606 7310 44658 7362
rect 45278 7310 45330 7362
rect 3166 7198 3218 7250
rect 24334 7198 24386 7250
rect 24558 7198 24610 7250
rect 42030 7198 42082 7250
rect 44158 7198 44210 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 13022 6862 13074 6914
rect 30270 6862 30322 6914
rect 40238 6862 40290 6914
rect 41022 6862 41074 6914
rect 42254 6862 42306 6914
rect 45054 6862 45106 6914
rect 45278 6862 45330 6914
rect 45502 6862 45554 6914
rect 4622 6750 4674 6802
rect 5182 6750 5234 6802
rect 6414 6750 6466 6802
rect 11118 6750 11170 6802
rect 12014 6750 12066 6802
rect 16382 6750 16434 6802
rect 17054 6750 17106 6802
rect 17838 6750 17890 6802
rect 29262 6750 29314 6802
rect 33854 6750 33906 6802
rect 37774 6750 37826 6802
rect 39902 6750 39954 6802
rect 46734 6750 46786 6802
rect 1822 6638 1874 6690
rect 6862 6638 6914 6690
rect 7310 6638 7362 6690
rect 7870 6638 7922 6690
rect 8206 6638 8258 6690
rect 8990 6638 9042 6690
rect 12574 6638 12626 6690
rect 13582 6638 13634 6690
rect 16718 6638 16770 6690
rect 17390 6638 17442 6690
rect 20750 6638 20802 6690
rect 26014 6638 26066 6690
rect 29374 6638 29426 6690
rect 29598 6638 29650 6690
rect 30046 6638 30098 6690
rect 30942 6638 30994 6690
rect 32174 6638 32226 6690
rect 33294 6638 33346 6690
rect 35758 6638 35810 6690
rect 36990 6638 37042 6690
rect 40238 6638 40290 6690
rect 43710 6638 43762 6690
rect 43822 6638 43874 6690
rect 44046 6638 44098 6690
rect 44830 6638 44882 6690
rect 47630 6638 47682 6690
rect 48190 6638 48242 6690
rect 2494 6526 2546 6578
rect 5630 6526 5682 6578
rect 6302 6526 6354 6578
rect 6638 6526 6690 6578
rect 12126 6526 12178 6578
rect 12462 6526 12514 6578
rect 14254 6526 14306 6578
rect 19966 6526 20018 6578
rect 21310 6526 21362 6578
rect 24222 6526 24274 6578
rect 28254 6526 28306 6578
rect 29150 6526 29202 6578
rect 32958 6526 33010 6578
rect 40574 6526 40626 6578
rect 41134 6526 41186 6578
rect 42366 6526 42418 6578
rect 42926 6526 42978 6578
rect 43262 6526 43314 6578
rect 44158 6526 44210 6578
rect 44382 6526 44434 6578
rect 45614 6526 45666 6578
rect 45950 6526 46002 6578
rect 47854 6526 47906 6578
rect 5966 6414 6018 6466
rect 7198 6414 7250 6466
rect 7422 6414 7474 6466
rect 16942 6414 16994 6466
rect 17166 6414 17218 6466
rect 21422 6414 21474 6466
rect 21534 6414 21586 6466
rect 28590 6414 28642 6466
rect 30606 6414 30658 6466
rect 31054 6414 31106 6466
rect 31278 6414 31330 6466
rect 31614 6414 31666 6466
rect 32510 6414 32562 6466
rect 41022 6414 41074 6466
rect 41582 6414 41634 6466
rect 41918 6414 41970 6466
rect 42142 6414 42194 6466
rect 42590 6414 42642 6466
rect 42814 6414 42866 6466
rect 46286 6414 46338 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4734 6078 4786 6130
rect 5182 6078 5234 6130
rect 8766 6078 8818 6130
rect 15598 6078 15650 6130
rect 16270 6078 16322 6130
rect 20862 6078 20914 6130
rect 26574 6078 26626 6130
rect 33742 6078 33794 6130
rect 33966 6078 34018 6130
rect 38670 6078 38722 6130
rect 39342 6078 39394 6130
rect 39454 6078 39506 6130
rect 41246 6078 41298 6130
rect 44606 6078 44658 6130
rect 45054 6078 45106 6130
rect 5070 5966 5122 6018
rect 7982 5966 8034 6018
rect 16158 5966 16210 6018
rect 16382 5966 16434 6018
rect 25230 5966 25282 6018
rect 26462 5966 26514 6018
rect 26686 5966 26738 6018
rect 34974 5966 35026 6018
rect 36094 5966 36146 6018
rect 41134 5966 41186 6018
rect 47406 5966 47458 6018
rect 4174 5854 4226 5906
rect 5406 5854 5458 5906
rect 6526 5854 6578 5906
rect 7422 5854 7474 5906
rect 7870 5854 7922 5906
rect 8094 5854 8146 5906
rect 15150 5854 15202 5906
rect 17950 5854 18002 5906
rect 21198 5854 21250 5906
rect 21758 5854 21810 5906
rect 25454 5854 25506 5906
rect 32286 5854 32338 5906
rect 33630 5854 33682 5906
rect 34190 5854 34242 5906
rect 34862 5854 34914 5906
rect 35422 5854 35474 5906
rect 39230 5854 39282 5906
rect 39566 5854 39618 5906
rect 39790 5854 39842 5906
rect 40798 5854 40850 5906
rect 41806 5854 41858 5906
rect 42702 5854 42754 5906
rect 42814 5854 42866 5906
rect 43038 5854 43090 5906
rect 43486 5854 43538 5906
rect 48078 5854 48130 5906
rect 6190 5742 6242 5794
rect 6974 5742 7026 5794
rect 10110 5742 10162 5794
rect 17614 5742 17666 5794
rect 22430 5742 22482 5794
rect 24558 5742 24610 5794
rect 26014 5742 26066 5794
rect 29262 5742 29314 5794
rect 33182 5742 33234 5794
rect 33854 5742 33906 5794
rect 38222 5742 38274 5794
rect 40126 5742 40178 5794
rect 40238 5742 40290 5794
rect 41582 5742 41634 5794
rect 45278 5742 45330 5794
rect 4398 5630 4450 5682
rect 7198 5630 7250 5682
rect 18958 5630 19010 5682
rect 25902 5630 25954 5682
rect 33070 5630 33122 5682
rect 41358 5630 41410 5682
rect 42254 5630 42306 5682
rect 43710 5630 43762 5682
rect 44046 5630 44098 5682
rect 44382 5630 44434 5682
rect 45054 5630 45106 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 22542 5294 22594 5346
rect 30270 5294 30322 5346
rect 39902 5294 39954 5346
rect 40238 5294 40290 5346
rect 41582 5294 41634 5346
rect 41918 5294 41970 5346
rect 9662 5182 9714 5234
rect 10782 5182 10834 5234
rect 12910 5182 12962 5234
rect 14926 5182 14978 5234
rect 15262 5182 15314 5234
rect 15710 5182 15762 5234
rect 19518 5182 19570 5234
rect 20414 5182 20466 5234
rect 21534 5182 21586 5234
rect 23550 5182 23602 5234
rect 24670 5182 24722 5234
rect 25118 5182 25170 5234
rect 26462 5182 26514 5234
rect 26910 5182 26962 5234
rect 29150 5182 29202 5234
rect 29598 5182 29650 5234
rect 31054 5182 31106 5234
rect 32174 5182 32226 5234
rect 34302 5182 34354 5234
rect 34750 5182 34802 5234
rect 35870 5182 35922 5234
rect 42702 5182 42754 5234
rect 43486 5182 43538 5234
rect 44382 5182 44434 5234
rect 44830 5182 44882 5234
rect 5854 5070 5906 5122
rect 6190 5070 6242 5122
rect 6750 5070 6802 5122
rect 10110 5070 10162 5122
rect 16158 5070 16210 5122
rect 16606 5070 16658 5122
rect 19854 5070 19906 5122
rect 20526 5070 20578 5122
rect 21310 5070 21362 5122
rect 21646 5070 21698 5122
rect 22318 5070 22370 5122
rect 22766 5070 22818 5122
rect 23438 5070 23490 5122
rect 23998 5070 24050 5122
rect 24782 5070 24834 5122
rect 29486 5070 29538 5122
rect 31502 5070 31554 5122
rect 34638 5070 34690 5122
rect 35086 5070 35138 5122
rect 35646 5070 35698 5122
rect 36318 5070 36370 5122
rect 36990 5070 37042 5122
rect 40238 5070 40290 5122
rect 40686 5070 40738 5122
rect 41358 5070 41410 5122
rect 42814 5070 42866 5122
rect 46958 5070 47010 5122
rect 47630 5070 47682 5122
rect 5966 4958 6018 5010
rect 7534 4958 7586 5010
rect 15038 4958 15090 5010
rect 15710 4958 15762 5010
rect 15822 4958 15874 5010
rect 17390 4958 17442 5010
rect 20078 4958 20130 5010
rect 21982 4958 22034 5010
rect 23774 4958 23826 5010
rect 27806 4958 27858 5010
rect 30494 4958 30546 5010
rect 35310 4958 35362 5010
rect 35870 4958 35922 5010
rect 41022 4958 41074 5010
rect 16046 4846 16098 4898
rect 20302 4846 20354 4898
rect 22430 4846 22482 4898
rect 23550 4846 23602 4898
rect 25678 4846 25730 4898
rect 26014 4846 26066 4898
rect 28142 4846 28194 4898
rect 28590 4846 28642 4898
rect 30382 4846 30434 4898
rect 34862 4846 34914 4898
rect 36094 4846 36146 4898
rect 37998 4846 38050 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 7758 4510 7810 4562
rect 17614 4510 17666 4562
rect 17838 4510 17890 4562
rect 17950 4510 18002 4562
rect 33294 4510 33346 4562
rect 7422 4398 7474 4450
rect 8654 4398 8706 4450
rect 8990 4398 9042 4450
rect 11006 4398 11058 4450
rect 14254 4398 14306 4450
rect 17390 4398 17442 4450
rect 19294 4398 19346 4450
rect 22542 4398 22594 4450
rect 25230 4398 25282 4450
rect 30046 4398 30098 4450
rect 33518 4398 33570 4450
rect 39566 4398 39618 4450
rect 40910 4398 40962 4450
rect 41246 4398 41298 4450
rect 41582 4398 41634 4450
rect 42142 4398 42194 4450
rect 45390 4398 45442 4450
rect 4174 4286 4226 4338
rect 10222 4286 10274 4338
rect 13582 4286 13634 4338
rect 18510 4286 18562 4338
rect 21870 4286 21922 4338
rect 25790 4286 25842 4338
rect 29262 4286 29314 4338
rect 34078 4286 34130 4338
rect 40350 4286 40402 4338
rect 43598 4286 43650 4338
rect 4958 4174 5010 4226
rect 7086 4174 7138 4226
rect 13134 4174 13186 4226
rect 16382 4174 16434 4226
rect 17726 4174 17778 4226
rect 21422 4174 21474 4226
rect 24670 4174 24722 4226
rect 26574 4174 26626 4226
rect 28702 4174 28754 4226
rect 32174 4174 32226 4226
rect 34750 4174 34802 4226
rect 36878 4174 36930 4226
rect 37438 4174 37490 4226
rect 42030 4174 42082 4226
rect 33630 4062 33682 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 7422 3726 7474 3778
rect 17278 3726 17330 3778
rect 24558 3726 24610 3778
rect 24894 3726 24946 3778
rect 26574 3726 26626 3778
rect 26910 3726 26962 3778
rect 28702 3726 28754 3778
rect 40014 3726 40066 3778
rect 7534 3614 7586 3666
rect 17166 3614 17218 3666
rect 22094 3614 22146 3666
rect 28590 3614 28642 3666
rect 30270 3614 30322 3666
rect 32958 3614 33010 3666
rect 35086 3614 35138 3666
rect 36990 3614 37042 3666
rect 45502 3614 45554 3666
rect 7758 3502 7810 3554
rect 16382 3502 16434 3554
rect 17614 3502 17666 3554
rect 21086 3502 21138 3554
rect 26574 3502 26626 3554
rect 29038 3502 29090 3554
rect 32286 3502 32338 3554
rect 35982 3502 36034 3554
rect 42366 3502 42418 3554
rect 43934 3502 43986 3554
rect 47630 3502 47682 3554
rect 8206 3390 8258 3442
rect 17054 3390 17106 3442
rect 19294 3390 19346 3442
rect 24670 3390 24722 3442
rect 44158 3390 44210 3442
rect 47854 3390 47906 3442
rect 48190 3390 48242 3442
rect 3838 3278 3890 3330
rect 5518 3278 5570 3330
rect 6974 3278 7026 3330
rect 8542 3278 8594 3330
rect 10110 3278 10162 3330
rect 11678 3278 11730 3330
rect 12574 3278 12626 3330
rect 13470 3278 13522 3330
rect 15374 3278 15426 3330
rect 25230 3278 25282 3330
rect 25790 3278 25842 3330
rect 27358 3278 27410 3330
rect 38894 3278 38946 3330
rect 42702 3278 42754 3330
rect 44494 3278 44546 3330
rect 44942 3278 44994 3330
rect 46174 3278 46226 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 13470 1710 13522 1762
rect 14590 1710 14642 1762
<< metal2 >>
rect 6272 49200 6384 50000
rect 18592 49200 18704 50000
rect 30912 49200 31024 50000
rect 43232 49200 43344 50000
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 5964 43538 6020 43550
rect 5964 43486 5966 43538
rect 6018 43486 6020 43538
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 5964 41972 6020 43486
rect 6076 41972 6132 41982
rect 5964 41970 6132 41972
rect 5964 41918 6078 41970
rect 6130 41918 6132 41970
rect 5964 41916 6132 41918
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 4620 41300 4676 41310
rect 4620 40404 4676 41244
rect 6076 41300 6132 41916
rect 6076 41206 6132 41244
rect 4620 40402 4900 40404
rect 4620 40350 4622 40402
rect 4674 40350 4900 40402
rect 4620 40348 4900 40350
rect 4620 40338 4676 40348
rect 1708 40290 1764 40302
rect 1708 40238 1710 40290
rect 1762 40238 1764 40290
rect 1708 39508 1764 40238
rect 3836 40292 3892 40302
rect 3836 40290 4004 40292
rect 3836 40238 3838 40290
rect 3890 40238 4004 40290
rect 3836 40236 4004 40238
rect 3836 40226 3892 40236
rect 2716 39620 2772 39630
rect 2716 39618 3220 39620
rect 2716 39566 2718 39618
rect 2770 39566 3220 39618
rect 2716 39564 3220 39566
rect 2716 39554 2772 39564
rect 1708 39442 1764 39452
rect 2828 39394 2884 39406
rect 2828 39342 2830 39394
rect 2882 39342 2884 39394
rect 2828 38836 2884 39342
rect 3052 39396 3108 39406
rect 3052 39302 3108 39340
rect 3164 39396 3220 39564
rect 3388 39508 3444 39518
rect 3388 39414 3444 39452
rect 3500 39508 3556 39518
rect 3836 39508 3892 39518
rect 3500 39506 3892 39508
rect 3500 39454 3502 39506
rect 3554 39454 3838 39506
rect 3890 39454 3892 39506
rect 3500 39452 3892 39454
rect 3164 39394 3332 39396
rect 3164 39342 3166 39394
rect 3218 39342 3332 39394
rect 3164 39340 3332 39342
rect 3164 39330 3220 39340
rect 2828 38770 2884 38780
rect 1708 38722 1764 38734
rect 1708 38670 1710 38722
rect 1762 38670 1764 38722
rect 1708 38052 1764 38670
rect 2716 38724 2772 38734
rect 2716 38162 2772 38668
rect 2716 38110 2718 38162
rect 2770 38110 2772 38162
rect 2716 38098 2772 38110
rect 1708 37986 1764 37996
rect 3276 38050 3332 39340
rect 3276 37998 3278 38050
rect 3330 37998 3332 38050
rect 3276 37986 3332 37998
rect 3388 38836 3444 38846
rect 2828 37940 2884 37950
rect 3164 37940 3220 37950
rect 2828 37938 3220 37940
rect 2828 37886 2830 37938
rect 2882 37886 3166 37938
rect 3218 37886 3220 37938
rect 2828 37884 3220 37886
rect 2828 37874 2884 37884
rect 3164 37874 3220 37884
rect 2604 37828 2660 37838
rect 2604 37734 2660 37772
rect 3276 37828 3332 37838
rect 3052 37268 3108 37278
rect 3276 37268 3332 37772
rect 3052 37266 3332 37268
rect 3052 37214 3054 37266
rect 3106 37214 3332 37266
rect 3052 37212 3332 37214
rect 3052 37202 3108 37212
rect 2940 37042 2996 37054
rect 2940 36990 2942 37042
rect 2994 36990 2996 37042
rect 1708 36594 1764 36606
rect 1708 36542 1710 36594
rect 1762 36542 1764 36594
rect 1708 35812 1764 36542
rect 2940 36596 2996 36990
rect 2940 36530 2996 36540
rect 3276 37042 3332 37054
rect 3276 36990 3278 37042
rect 3330 36990 3332 37042
rect 3276 35922 3332 36990
rect 3276 35870 3278 35922
rect 3330 35870 3332 35922
rect 3276 35858 3332 35870
rect 1708 35746 1764 35756
rect 3164 35700 3220 35710
rect 3164 35698 3332 35700
rect 3164 35646 3166 35698
rect 3218 35646 3332 35698
rect 3164 35644 3332 35646
rect 3164 35634 3220 35644
rect 3052 35028 3108 35038
rect 2156 35026 3108 35028
rect 2156 34974 3054 35026
rect 3106 34974 3108 35026
rect 2156 34972 3108 34974
rect 2156 34914 2212 34972
rect 3052 34962 3108 34972
rect 2156 34862 2158 34914
rect 2210 34862 2212 34914
rect 2156 34850 2212 34862
rect 3276 34916 3332 35644
rect 3276 34850 3332 34860
rect 2268 34804 2324 34814
rect 2604 34804 2660 34814
rect 2940 34804 2996 34814
rect 2268 34802 2436 34804
rect 2268 34750 2270 34802
rect 2322 34750 2436 34802
rect 2268 34748 2436 34750
rect 2268 34738 2324 34748
rect 2380 34692 2436 34748
rect 2604 34802 2940 34804
rect 2604 34750 2606 34802
rect 2658 34750 2940 34802
rect 2604 34748 2940 34750
rect 2604 34738 2660 34748
rect 2940 34710 2996 34748
rect 3164 34802 3220 34814
rect 3164 34750 3166 34802
rect 3218 34750 3220 34802
rect 2380 34626 2436 34636
rect 2492 34690 2548 34702
rect 2492 34638 2494 34690
rect 2546 34638 2548 34690
rect 2492 34242 2548 34638
rect 3164 34692 3220 34750
rect 3276 34692 3332 34702
rect 3164 34636 3276 34692
rect 3276 34626 3332 34636
rect 3388 34468 3444 38780
rect 3500 37268 3556 39452
rect 3836 39442 3892 39452
rect 3948 39284 4004 40236
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4172 39732 4228 39742
rect 4172 39730 4788 39732
rect 4172 39678 4174 39730
rect 4226 39678 4788 39730
rect 4172 39676 4788 39678
rect 4172 39666 4228 39676
rect 4060 39508 4116 39518
rect 4060 39396 4116 39452
rect 4508 39506 4564 39518
rect 4508 39454 4510 39506
rect 4562 39454 4564 39506
rect 4508 39396 4564 39454
rect 4732 39506 4788 39676
rect 4732 39454 4734 39506
rect 4786 39454 4788 39506
rect 4732 39442 4788 39454
rect 4060 39394 4228 39396
rect 4060 39342 4062 39394
rect 4114 39342 4228 39394
rect 4060 39340 4228 39342
rect 4060 39330 4116 39340
rect 3948 39218 4004 39228
rect 3836 38724 3892 38734
rect 3836 38630 3892 38668
rect 3836 38052 3892 38062
rect 3892 37996 4004 38052
rect 3836 37958 3892 37996
rect 3500 37266 3668 37268
rect 3500 37214 3502 37266
rect 3554 37214 3668 37266
rect 3500 37212 3668 37214
rect 3500 37202 3556 37212
rect 3500 35698 3556 35710
rect 3500 35646 3502 35698
rect 3554 35646 3556 35698
rect 3500 35140 3556 35646
rect 3612 35140 3668 37212
rect 3836 36596 3892 36606
rect 3836 36502 3892 36540
rect 3724 35812 3780 35822
rect 3724 35718 3780 35756
rect 3948 35700 4004 37996
rect 4172 35810 4228 39340
rect 4508 39330 4564 39340
rect 4620 39394 4676 39406
rect 4620 39342 4622 39394
rect 4674 39342 4676 39394
rect 4620 39284 4676 39342
rect 4620 39218 4676 39228
rect 4620 38836 4676 38846
rect 4844 38836 4900 40348
rect 6076 38948 6132 38958
rect 6076 38854 6132 38892
rect 5292 38836 5348 38846
rect 4620 38834 5348 38836
rect 4620 38782 4622 38834
rect 4674 38782 5294 38834
rect 5346 38782 5348 38834
rect 4620 38780 5348 38782
rect 4620 38770 4676 38780
rect 5292 38770 5348 38780
rect 6300 38668 6356 49200
rect 18620 46116 18676 49200
rect 30940 46450 30996 49200
rect 30940 46398 30942 46450
rect 30994 46398 30996 46450
rect 30940 46386 30996 46398
rect 32620 46450 32676 46462
rect 32620 46398 32622 46450
rect 32674 46398 32676 46450
rect 18620 46060 18900 46116
rect 18508 46004 18564 46014
rect 18620 46004 18676 46060
rect 18508 46002 18676 46004
rect 18508 45950 18510 46002
rect 18562 45950 18676 46002
rect 18508 45948 18676 45950
rect 18508 45938 18564 45948
rect 11340 45890 11396 45902
rect 11340 45838 11342 45890
rect 11394 45838 11396 45890
rect 10668 45778 10724 45790
rect 10668 45726 10670 45778
rect 10722 45726 10724 45778
rect 10668 45220 10724 45726
rect 10444 45164 10724 45220
rect 10892 45778 10948 45790
rect 10892 45726 10894 45778
rect 10946 45726 10948 45778
rect 10444 44548 10500 45164
rect 10444 44482 10500 44492
rect 10556 44996 10612 45006
rect 10892 44996 10948 45726
rect 10556 44994 10948 44996
rect 10556 44942 10558 44994
rect 10610 44942 10948 44994
rect 10556 44940 10948 44942
rect 11116 45666 11172 45678
rect 11116 45614 11118 45666
rect 11170 45614 11172 45666
rect 7644 44436 7700 44446
rect 7644 44342 7700 44380
rect 10444 44324 10500 44334
rect 9996 44322 10500 44324
rect 9996 44270 10446 44322
rect 10498 44270 10500 44322
rect 9996 44268 10500 44270
rect 9772 44210 9828 44222
rect 9772 44158 9774 44210
rect 9826 44158 9828 44210
rect 9772 43540 9828 44158
rect 9772 43474 9828 43484
rect 9884 43652 9940 43662
rect 6636 43428 6692 43438
rect 6636 43334 6692 43372
rect 8876 43426 8932 43438
rect 8876 43374 8878 43426
rect 8930 43374 8932 43426
rect 8876 43204 8932 43374
rect 8876 43138 8932 43148
rect 9548 43426 9604 43438
rect 9548 43374 9550 43426
rect 9602 43374 9604 43426
rect 9548 43204 9604 43374
rect 9772 43316 9828 43326
rect 9884 43316 9940 43596
rect 9772 43314 9940 43316
rect 9772 43262 9774 43314
rect 9826 43262 9940 43314
rect 9772 43260 9940 43262
rect 9772 43250 9828 43260
rect 9548 43138 9604 43148
rect 9996 42868 10052 44268
rect 10444 44258 10500 44268
rect 10556 44212 10612 44940
rect 10780 44212 10836 44222
rect 10556 44156 10780 44212
rect 10780 44146 10836 44156
rect 10892 44098 10948 44110
rect 10892 44046 10894 44098
rect 10946 44046 10948 44098
rect 10892 43652 10948 44046
rect 11116 43708 11172 45614
rect 11340 44210 11396 45838
rect 17500 45892 17556 45902
rect 17500 45330 17556 45836
rect 17500 45278 17502 45330
rect 17554 45278 17556 45330
rect 13468 45108 13524 45118
rect 13804 45108 13860 45118
rect 13468 45106 13860 45108
rect 13468 45054 13470 45106
rect 13522 45054 13806 45106
rect 13858 45054 13860 45106
rect 13468 45052 13860 45054
rect 13468 45042 13524 45052
rect 12684 44994 12740 45006
rect 12684 44942 12686 44994
rect 12738 44942 12740 44994
rect 11564 44436 11620 44446
rect 11564 44322 11620 44380
rect 12012 44436 12068 44446
rect 12012 44342 12068 44380
rect 12684 44434 12740 44942
rect 12684 44382 12686 44434
rect 12738 44382 12740 44434
rect 12684 44370 12740 44382
rect 11564 44270 11566 44322
rect 11618 44270 11620 44322
rect 11564 44258 11620 44270
rect 11340 44158 11342 44210
rect 11394 44158 11396 44210
rect 11340 44100 11396 44158
rect 11340 44034 11396 44044
rect 11452 44212 11508 44222
rect 11452 43764 11508 44156
rect 12908 44212 12964 44222
rect 13468 44212 13524 44222
rect 12908 44210 13524 44212
rect 12908 44158 12910 44210
rect 12962 44158 13470 44210
rect 13522 44158 13524 44210
rect 12908 44156 13524 44158
rect 12908 44146 12964 44156
rect 13468 44146 13524 44156
rect 12124 44098 12180 44110
rect 12124 44046 12126 44098
rect 12178 44046 12180 44098
rect 11676 43764 11732 43774
rect 11452 43708 11676 43764
rect 11116 43652 11396 43708
rect 11676 43698 11732 43708
rect 10948 43596 11060 43652
rect 10892 43586 10948 43596
rect 10444 43428 10500 43438
rect 10444 43334 10500 43372
rect 11004 43428 11060 43596
rect 11340 43538 11396 43652
rect 11340 43486 11342 43538
rect 11394 43486 11396 43538
rect 11340 43474 11396 43486
rect 11900 43540 11956 43550
rect 11900 43446 11956 43484
rect 11004 43362 11060 43372
rect 11564 43428 11620 43438
rect 11564 43334 11620 43372
rect 9660 42866 10052 42868
rect 9660 42814 9998 42866
rect 10050 42814 10052 42866
rect 9660 42812 10052 42814
rect 6860 42084 6916 42094
rect 6860 41970 6916 42028
rect 6860 41918 6862 41970
rect 6914 41918 6916 41970
rect 6860 41906 6916 41918
rect 8988 41858 9044 41870
rect 8988 41806 8990 41858
rect 9042 41806 9044 41858
rect 8988 41636 9044 41806
rect 8988 41570 9044 41580
rect 9660 40402 9716 42812
rect 9996 42802 10052 42812
rect 10108 43314 10164 43326
rect 10108 43262 10110 43314
rect 10162 43262 10164 43314
rect 10108 41972 10164 43262
rect 10556 43314 10612 43326
rect 10556 43262 10558 43314
rect 10610 43262 10612 43314
rect 10556 43092 10612 43262
rect 10780 43316 10836 43326
rect 10780 43222 10836 43260
rect 10892 43314 10948 43326
rect 10892 43262 10894 43314
rect 10946 43262 10948 43314
rect 10332 41972 10388 41982
rect 10108 41970 10332 41972
rect 10108 41918 10110 41970
rect 10162 41918 10332 41970
rect 10108 41916 10332 41918
rect 10108 41906 10164 41916
rect 10332 41906 10388 41916
rect 9884 41858 9940 41870
rect 9884 41806 9886 41858
rect 9938 41806 9940 41858
rect 9884 41636 9940 41806
rect 10444 41860 10500 41870
rect 10444 41766 10500 41804
rect 10556 41748 10612 43036
rect 10780 42084 10836 42094
rect 10780 41990 10836 42028
rect 10892 41972 10948 43262
rect 11788 43314 11844 43326
rect 11788 43262 11790 43314
rect 11842 43262 11844 43314
rect 11788 43092 11844 43262
rect 11788 43026 11844 43036
rect 12124 43092 12180 44046
rect 12684 44098 12740 44110
rect 12684 44046 12686 44098
rect 12738 44046 12740 44098
rect 12572 43538 12628 43550
rect 12572 43486 12574 43538
rect 12626 43486 12628 43538
rect 12236 43428 12292 43438
rect 12236 43334 12292 43372
rect 12348 43426 12404 43438
rect 12348 43374 12350 43426
rect 12402 43374 12404 43426
rect 12348 43316 12404 43374
rect 12572 43428 12628 43486
rect 12572 43362 12628 43372
rect 12348 43250 12404 43260
rect 12124 43026 12180 43036
rect 12684 42308 12740 44046
rect 13804 43708 13860 45052
rect 14588 44994 14644 45006
rect 16716 44996 16772 45006
rect 14588 44942 14590 44994
rect 14642 44942 14644 44994
rect 14588 44548 14644 44942
rect 16604 44940 16716 44996
rect 14588 44482 14644 44492
rect 16156 44548 16212 44558
rect 16156 44454 16212 44492
rect 15148 44436 15204 44446
rect 15148 44434 15428 44436
rect 15148 44382 15150 44434
rect 15202 44382 15428 44434
rect 15148 44380 15428 44382
rect 15148 44370 15204 44380
rect 13580 43652 13636 43662
rect 13580 43558 13636 43596
rect 13692 43652 13860 43708
rect 14140 44322 14196 44334
rect 14140 44270 14142 44322
rect 14194 44270 14196 44322
rect 12684 42242 12740 42252
rect 12908 42754 12964 42766
rect 12908 42702 12910 42754
rect 12962 42702 12964 42754
rect 11900 42082 11956 42094
rect 11900 42030 11902 42082
rect 11954 42030 11956 42082
rect 10892 41906 10948 41916
rect 11676 41972 11732 41982
rect 11676 41878 11732 41916
rect 11228 41860 11284 41870
rect 11228 41766 11284 41804
rect 11788 41858 11844 41870
rect 11788 41806 11790 41858
rect 11842 41806 11844 41858
rect 10892 41748 10948 41758
rect 10556 41746 10948 41748
rect 10556 41694 10894 41746
rect 10946 41694 10948 41746
rect 10556 41692 10948 41694
rect 9884 41570 9940 41580
rect 10332 41188 10388 41198
rect 10332 40514 10388 41132
rect 10332 40462 10334 40514
rect 10386 40462 10388 40514
rect 10332 40450 10388 40462
rect 9660 40350 9662 40402
rect 9714 40350 9716 40402
rect 9660 40338 9716 40350
rect 10780 40292 10836 41692
rect 10892 41682 10948 41692
rect 11116 41748 11172 41758
rect 11116 41654 11172 41692
rect 11788 41748 11844 41806
rect 11788 41682 11844 41692
rect 11900 41636 11956 42030
rect 12572 42084 12628 42094
rect 12572 42082 12852 42084
rect 12572 42030 12574 42082
rect 12626 42030 12852 42082
rect 12572 42028 12852 42030
rect 12572 42018 12628 42028
rect 12460 41970 12516 41982
rect 12460 41918 12462 41970
rect 12514 41918 12516 41970
rect 11900 41570 11956 41580
rect 12012 41860 12068 41870
rect 12012 41298 12068 41804
rect 12460 41860 12516 41918
rect 12460 41794 12516 41804
rect 12012 41246 12014 41298
rect 12066 41246 12068 41298
rect 12012 41234 12068 41246
rect 12572 41746 12628 41758
rect 12572 41694 12574 41746
rect 12626 41694 12628 41746
rect 10892 41186 10948 41198
rect 10892 41134 10894 41186
rect 10946 41134 10948 41186
rect 10892 40964 10948 41134
rect 12348 41186 12404 41198
rect 12348 41134 12350 41186
rect 12402 41134 12404 41186
rect 11340 40964 11396 40974
rect 10892 40908 11340 40964
rect 11340 40404 11396 40908
rect 12348 40628 12404 41134
rect 12572 40628 12628 41694
rect 12348 40562 12404 40572
rect 12460 40572 12628 40628
rect 12460 40404 12516 40572
rect 12796 40516 12852 42028
rect 12908 41860 12964 42702
rect 13580 42756 13636 42766
rect 13692 42756 13748 43652
rect 13916 43428 13972 43438
rect 14140 43428 14196 44270
rect 14364 44322 14420 44334
rect 14364 44270 14366 44322
rect 14418 44270 14420 44322
rect 14364 44100 14420 44270
rect 15372 44324 15428 44380
rect 15596 44324 15652 44334
rect 15372 44322 15652 44324
rect 15372 44270 15598 44322
rect 15650 44270 15652 44322
rect 15372 44268 15652 44270
rect 15596 44258 15652 44268
rect 15820 44324 15876 44334
rect 15036 44212 15092 44222
rect 15036 44118 15092 44156
rect 15260 44210 15316 44222
rect 15260 44158 15262 44210
rect 15314 44158 15316 44210
rect 14364 44034 14420 44044
rect 15260 43764 15316 44158
rect 15820 44100 15876 44268
rect 15820 44034 15876 44044
rect 16044 44322 16100 44334
rect 16044 44270 16046 44322
rect 16098 44270 16100 44322
rect 16044 44100 16100 44270
rect 16044 44034 16100 44044
rect 16492 44322 16548 44334
rect 16492 44270 16494 44322
rect 16546 44270 16548 44322
rect 15260 43698 15316 43708
rect 16044 43764 16100 43774
rect 16492 43764 16548 44270
rect 16604 44212 16660 44940
rect 16716 44902 16772 44940
rect 17388 44436 17444 44446
rect 17388 44342 17444 44380
rect 16604 44146 16660 44156
rect 16716 44322 16772 44334
rect 16716 44270 16718 44322
rect 16770 44270 16772 44322
rect 16100 43708 16548 43764
rect 16716 43764 16772 44270
rect 16940 44322 16996 44334
rect 16940 44270 16942 44322
rect 16994 44270 16996 44322
rect 16940 44100 16996 44270
rect 17276 44324 17332 44334
rect 17052 44212 17108 44222
rect 17052 44118 17108 44156
rect 16940 44034 16996 44044
rect 16716 43708 16884 43764
rect 16044 43670 16100 43708
rect 16604 43652 16660 43662
rect 13916 43426 14196 43428
rect 13916 43374 13918 43426
rect 13970 43374 14196 43426
rect 13916 43372 14196 43374
rect 13916 43362 13972 43372
rect 14140 43316 14196 43372
rect 14140 43250 14196 43260
rect 16492 43538 16548 43550
rect 16492 43486 16494 43538
rect 16546 43486 16548 43538
rect 16492 43092 16548 43486
rect 13580 42754 13748 42756
rect 13580 42702 13582 42754
rect 13634 42702 13748 42754
rect 13580 42700 13748 42702
rect 13580 42690 13636 42700
rect 13132 41860 13188 41870
rect 12908 41804 13132 41860
rect 12908 41076 12964 41086
rect 12908 40982 12964 41020
rect 13132 40964 13188 41804
rect 13692 41300 13748 42700
rect 16268 43036 16548 43092
rect 14252 42644 14308 42654
rect 14028 42642 14308 42644
rect 14028 42590 14254 42642
rect 14306 42590 14308 42642
rect 14028 42588 14308 42590
rect 13804 42308 13860 42318
rect 13804 41972 13860 42252
rect 14028 42194 14084 42588
rect 14252 42578 14308 42588
rect 14028 42142 14030 42194
rect 14082 42142 14084 42194
rect 14028 42130 14084 42142
rect 16044 42084 16100 42094
rect 14140 41972 14196 41982
rect 13804 41970 13972 41972
rect 13804 41918 13806 41970
rect 13858 41918 13972 41970
rect 13804 41916 13972 41918
rect 13804 41906 13860 41916
rect 13692 41234 13748 41244
rect 13580 41188 13636 41198
rect 13580 41094 13636 41132
rect 13468 41076 13524 41086
rect 13468 40982 13524 41020
rect 13692 41076 13748 41086
rect 13916 41076 13972 41916
rect 14140 41878 14196 41916
rect 15372 41972 15428 41982
rect 15372 41878 15428 41916
rect 16044 41970 16100 42028
rect 16044 41918 16046 41970
rect 16098 41918 16100 41970
rect 16044 41906 16100 41918
rect 16268 41860 16324 43036
rect 16380 42868 16436 42878
rect 16604 42868 16660 43596
rect 16716 43540 16772 43550
rect 16716 43446 16772 43484
rect 16380 42866 16660 42868
rect 16380 42814 16382 42866
rect 16434 42814 16660 42866
rect 16380 42812 16660 42814
rect 16828 42866 16884 43708
rect 17276 43762 17332 44268
rect 17276 43710 17278 43762
rect 17330 43710 17332 43762
rect 17276 43698 17332 43710
rect 16828 42814 16830 42866
rect 16882 42814 16884 42866
rect 16380 42802 16436 42812
rect 16828 42802 16884 42814
rect 16940 43652 16996 43662
rect 16940 42754 16996 43596
rect 17500 43540 17556 45278
rect 18060 45892 18116 45902
rect 17836 45106 17892 45118
rect 17836 45054 17838 45106
rect 17890 45054 17892 45106
rect 17836 44436 17892 45054
rect 17836 44370 17892 44380
rect 17836 43652 17892 43662
rect 17836 43558 17892 43596
rect 18060 43650 18116 45836
rect 18732 45890 18788 45902
rect 18732 45838 18734 45890
rect 18786 45838 18788 45890
rect 18060 43598 18062 43650
rect 18114 43598 18116 43650
rect 18060 43586 18116 43598
rect 18172 45106 18228 45118
rect 18172 45054 18174 45106
rect 18226 45054 18228 45106
rect 18172 44996 18228 45054
rect 18396 45108 18452 45118
rect 18396 45014 18452 45052
rect 16940 42702 16942 42754
rect 16994 42702 16996 42754
rect 16716 42644 16772 42654
rect 16604 42588 16716 42644
rect 16604 41860 16660 42588
rect 16716 42550 16772 42588
rect 16716 42084 16772 42094
rect 16716 41970 16772 42028
rect 16828 42084 16884 42094
rect 16940 42084 16996 42702
rect 17276 42756 17332 42766
rect 17500 42756 17556 43484
rect 17276 42754 17556 42756
rect 17276 42702 17278 42754
rect 17330 42702 17556 42754
rect 17276 42700 17556 42702
rect 17724 43538 17780 43550
rect 17724 43486 17726 43538
rect 17778 43486 17780 43538
rect 17276 42690 17332 42700
rect 17612 42644 17668 42654
rect 17612 42550 17668 42588
rect 17724 42532 17780 43486
rect 18172 43538 18228 44940
rect 18172 43486 18174 43538
rect 18226 43486 18228 43538
rect 18172 43474 18228 43486
rect 18508 44884 18564 44894
rect 18732 44884 18788 45838
rect 18844 45330 18900 46060
rect 20748 46060 21028 46116
rect 19628 45892 19684 45902
rect 19628 45798 19684 45836
rect 18844 45278 18846 45330
rect 18898 45278 18900 45330
rect 18844 45266 18900 45278
rect 19068 45778 19124 45790
rect 19068 45726 19070 45778
rect 19122 45726 19124 45778
rect 19068 44996 19124 45726
rect 19852 45668 19908 45678
rect 19628 45666 19908 45668
rect 19628 45614 19854 45666
rect 19906 45614 19908 45666
rect 19628 45612 19908 45614
rect 19628 45108 19684 45612
rect 19852 45602 19908 45612
rect 20076 45668 20132 45678
rect 20076 45666 20244 45668
rect 20076 45614 20078 45666
rect 20130 45614 20244 45666
rect 20076 45612 20244 45614
rect 20076 45602 20132 45612
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 20188 45332 20244 45612
rect 20076 45276 20244 45332
rect 19740 45108 19796 45118
rect 19628 45106 19796 45108
rect 19628 45054 19742 45106
rect 19794 45054 19796 45106
rect 19628 45052 19796 45054
rect 19740 45042 19796 45052
rect 19068 44930 19124 44940
rect 19404 44994 19460 45006
rect 19404 44942 19406 44994
rect 19458 44942 19460 44994
rect 18508 44882 18788 44884
rect 18508 44830 18510 44882
rect 18562 44830 18788 44882
rect 18508 44828 18788 44830
rect 18172 42756 18228 42766
rect 17948 42532 18004 42542
rect 17724 42530 18004 42532
rect 17724 42478 17950 42530
rect 18002 42478 18004 42530
rect 17724 42476 18004 42478
rect 16828 42082 16996 42084
rect 16828 42030 16830 42082
rect 16882 42030 16996 42082
rect 16828 42028 16996 42030
rect 17164 42196 17220 42206
rect 16828 42018 16884 42028
rect 16716 41918 16718 41970
rect 16770 41918 16772 41970
rect 16716 41906 16772 41918
rect 16268 41858 16660 41860
rect 16268 41806 16270 41858
rect 16322 41806 16660 41858
rect 16268 41804 16660 41806
rect 14476 41300 14532 41310
rect 14476 41206 14532 41244
rect 13692 41074 13972 41076
rect 13692 41022 13694 41074
rect 13746 41022 13972 41074
rect 13692 41020 13972 41022
rect 13692 41010 13748 41020
rect 13132 40898 13188 40908
rect 13580 40964 13636 40974
rect 11340 40348 11844 40404
rect 10892 40292 10948 40302
rect 10780 40236 10892 40292
rect 10892 40226 10948 40236
rect 9660 39732 9716 39742
rect 9660 39730 9828 39732
rect 9660 39678 9662 39730
rect 9714 39678 9828 39730
rect 9660 39676 9828 39678
rect 9660 39666 9716 39676
rect 6748 39618 6804 39630
rect 6748 39566 6750 39618
rect 6802 39566 6804 39618
rect 6300 38612 6580 38668
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 6076 38164 6132 38174
rect 5740 38162 6132 38164
rect 5740 38110 6078 38162
rect 6130 38110 6132 38162
rect 5740 38108 6132 38110
rect 5740 37378 5796 38108
rect 6076 38098 6132 38108
rect 6188 37940 6244 37950
rect 6076 37938 6244 37940
rect 6076 37886 6190 37938
rect 6242 37886 6244 37938
rect 6076 37884 6244 37886
rect 6076 37828 6132 37884
rect 6188 37874 6244 37884
rect 6412 37938 6468 37950
rect 6412 37886 6414 37938
rect 6466 37886 6468 37938
rect 6076 37762 6132 37772
rect 5740 37326 5742 37378
rect 5794 37326 5796 37378
rect 5740 37314 5796 37326
rect 5068 37268 5124 37278
rect 4844 37212 5068 37268
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4620 36484 4676 36494
rect 4844 36484 4900 37212
rect 5068 37174 5124 37212
rect 4620 36482 4900 36484
rect 4620 36430 4622 36482
rect 4674 36430 4900 36482
rect 4620 36428 4900 36430
rect 4620 36418 4676 36428
rect 5740 36372 5796 36382
rect 5740 36278 5796 36316
rect 5628 36258 5684 36270
rect 5628 36206 5630 36258
rect 5682 36206 5684 36258
rect 4396 35812 4452 35822
rect 4172 35758 4174 35810
rect 4226 35758 4228 35810
rect 4172 35746 4228 35758
rect 4284 35756 4396 35812
rect 4060 35700 4116 35710
rect 3948 35698 4116 35700
rect 3948 35646 4062 35698
rect 4114 35646 4116 35698
rect 3948 35644 4116 35646
rect 4060 35634 4116 35644
rect 3948 35140 4004 35150
rect 3612 35138 4004 35140
rect 3612 35086 3950 35138
rect 4002 35086 4004 35138
rect 3612 35084 4004 35086
rect 4284 35140 4340 35756
rect 4396 35718 4452 35756
rect 4844 35698 4900 35710
rect 4844 35646 4846 35698
rect 4898 35646 4900 35698
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4732 35140 4788 35150
rect 4844 35140 4900 35646
rect 4284 35084 4676 35140
rect 3500 34692 3556 35084
rect 3948 35074 4004 35084
rect 3500 34626 3556 34636
rect 3612 34914 3668 34926
rect 3612 34862 3614 34914
rect 3666 34862 3668 34914
rect 3612 34804 3668 34862
rect 4396 34916 4452 34926
rect 4396 34822 4452 34860
rect 4620 34914 4676 35084
rect 4788 35084 4900 35140
rect 5068 35474 5124 35486
rect 5068 35422 5070 35474
rect 5122 35422 5124 35474
rect 4732 35074 4788 35084
rect 4620 34862 4622 34914
rect 4674 34862 4676 34914
rect 4620 34850 4676 34862
rect 5068 34916 5124 35422
rect 5404 35140 5460 35150
rect 5460 35084 5572 35140
rect 5404 35074 5460 35084
rect 5068 34850 5124 34860
rect 3612 34468 3668 34748
rect 3388 34412 3668 34468
rect 4508 34802 4564 34814
rect 4508 34750 4510 34802
rect 4562 34750 4564 34802
rect 4508 34468 4564 34750
rect 5516 34804 5572 35084
rect 5628 35028 5684 36206
rect 6412 35924 6468 37886
rect 6412 35858 6468 35868
rect 5628 34962 5684 34972
rect 5628 34804 5684 34814
rect 5516 34802 5684 34804
rect 5516 34750 5630 34802
rect 5682 34750 5684 34802
rect 5516 34748 5684 34750
rect 5628 34738 5684 34748
rect 5964 34802 6020 34814
rect 5964 34750 5966 34802
rect 6018 34750 6020 34802
rect 4620 34468 4676 34478
rect 4508 34412 4620 34468
rect 2492 34190 2494 34242
rect 2546 34190 2548 34242
rect 2492 34178 2548 34190
rect 1820 34130 1876 34142
rect 1820 34078 1822 34130
rect 1874 34078 1876 34130
rect 1820 31778 1876 34078
rect 4620 34018 4676 34412
rect 5964 34468 6020 34750
rect 5964 34402 6020 34412
rect 5964 34244 6020 34254
rect 5964 34150 6020 34188
rect 5180 34132 5236 34142
rect 4620 33966 4622 34018
rect 4674 33966 4676 34018
rect 4620 33954 4676 33966
rect 4956 34130 5236 34132
rect 4956 34078 5182 34130
rect 5234 34078 5236 34130
rect 4956 34076 5236 34078
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4956 32674 5012 34076
rect 5180 34066 5236 34076
rect 4956 32622 4958 32674
rect 5010 32622 5012 32674
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 1820 31726 1822 31778
rect 1874 31726 1876 31778
rect 1820 31332 1876 31726
rect 3724 31892 3780 31902
rect 2492 31668 2548 31678
rect 2492 31574 2548 31612
rect 1820 30210 1876 31276
rect 3724 31332 3780 31836
rect 4620 31892 4676 31902
rect 4956 31892 5012 32622
rect 4620 31890 4900 31892
rect 4620 31838 4622 31890
rect 4674 31838 4900 31890
rect 4620 31836 4900 31838
rect 4620 31826 4676 31836
rect 3724 30994 3780 31276
rect 4396 31556 4452 31566
rect 4396 31106 4452 31500
rect 4396 31054 4398 31106
rect 4450 31054 4452 31106
rect 4396 31042 4452 31054
rect 3724 30942 3726 30994
rect 3778 30942 3780 30994
rect 3724 30930 3780 30942
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 1820 30158 1822 30210
rect 1874 30158 1876 30210
rect 1820 30146 1876 30158
rect 4620 30322 4676 30334
rect 4620 30270 4622 30322
rect 4674 30270 4676 30322
rect 2492 30100 2548 30110
rect 2492 30006 2548 30044
rect 4620 29652 4676 30270
rect 4844 29988 4900 31836
rect 4956 31826 5012 31836
rect 5964 33124 6020 33134
rect 5964 31778 6020 33068
rect 6524 31892 6580 38612
rect 6748 37268 6804 39566
rect 7532 39508 7588 39518
rect 7532 39414 7588 39452
rect 8540 39396 8596 39406
rect 8540 39060 8596 39340
rect 8540 38966 8596 39004
rect 9660 38946 9716 38958
rect 9660 38894 9662 38946
rect 9714 38894 9716 38946
rect 8876 38834 8932 38846
rect 8876 38782 8878 38834
rect 8930 38782 8932 38834
rect 8204 38724 8260 38734
rect 8092 38722 8260 38724
rect 8092 38670 8206 38722
rect 8258 38670 8260 38722
rect 8092 38668 8260 38670
rect 8876 38724 8932 38782
rect 9548 38724 9604 38734
rect 8876 38722 9604 38724
rect 8876 38670 9550 38722
rect 9602 38670 9604 38722
rect 8876 38668 9604 38670
rect 7308 38164 7364 38174
rect 7308 38050 7364 38108
rect 7308 37998 7310 38050
rect 7362 37998 7364 38050
rect 7308 37986 7364 37998
rect 8092 38052 8148 38668
rect 8204 38658 8260 38668
rect 9548 38658 9604 38668
rect 9660 38668 9716 38894
rect 9772 38948 9828 39676
rect 10220 39620 10276 39630
rect 10220 39618 10612 39620
rect 10220 39566 10222 39618
rect 10274 39566 10612 39618
rect 10220 39564 10612 39566
rect 10220 39554 10276 39564
rect 10108 39508 10164 39518
rect 10108 39414 10164 39452
rect 9996 39396 10052 39406
rect 10444 39396 10500 39406
rect 9996 39302 10052 39340
rect 10220 39394 10500 39396
rect 10220 39342 10446 39394
rect 10498 39342 10500 39394
rect 10220 39340 10500 39342
rect 10220 39284 10276 39340
rect 10444 39330 10500 39340
rect 10108 39228 10276 39284
rect 10108 39058 10164 39228
rect 10108 39006 10110 39058
rect 10162 39006 10164 39058
rect 10108 38994 10164 39006
rect 10444 39060 10500 39070
rect 9772 38882 9828 38892
rect 10332 38948 10388 38958
rect 9884 38722 9940 38734
rect 9884 38670 9886 38722
rect 9938 38670 9940 38722
rect 9660 38612 9828 38668
rect 8092 37958 8148 37996
rect 8428 38050 8484 38062
rect 8428 37998 8430 38050
rect 8482 37998 8484 38050
rect 7868 37940 7924 37950
rect 7868 37846 7924 37884
rect 8428 37940 8484 37998
rect 8764 38052 8820 38062
rect 8764 37958 8820 37996
rect 9660 38050 9716 38062
rect 9660 37998 9662 38050
rect 9714 37998 9716 38050
rect 8428 37874 8484 37884
rect 9212 37938 9268 37950
rect 9212 37886 9214 37938
rect 9266 37886 9268 37938
rect 6748 37202 6804 37212
rect 6972 37828 7028 37838
rect 6860 36372 6916 36382
rect 6860 35812 6916 36316
rect 6860 35698 6916 35756
rect 6860 35646 6862 35698
rect 6914 35646 6916 35698
rect 6860 35634 6916 35646
rect 6636 35474 6692 35486
rect 6636 35422 6638 35474
rect 6690 35422 6692 35474
rect 6636 34916 6692 35422
rect 6636 34850 6692 34860
rect 6748 34916 6804 34926
rect 6972 34916 7028 37772
rect 7980 37828 8036 37838
rect 7980 37826 8260 37828
rect 7980 37774 7982 37826
rect 8034 37774 8260 37826
rect 7980 37772 8260 37774
rect 7980 37762 8036 37772
rect 8092 37266 8148 37278
rect 8092 37214 8094 37266
rect 8146 37214 8148 37266
rect 7868 37156 7924 37166
rect 8092 37156 8148 37214
rect 7868 37154 8148 37156
rect 7868 37102 7870 37154
rect 7922 37102 8148 37154
rect 7868 37100 8148 37102
rect 7868 36708 7924 37100
rect 7084 36652 7924 36708
rect 7084 35922 7140 36652
rect 7308 36484 7364 36494
rect 7084 35870 7086 35922
rect 7138 35870 7140 35922
rect 7084 35858 7140 35870
rect 7196 35924 7252 35934
rect 7196 35830 7252 35868
rect 7308 35922 7364 36428
rect 8204 36484 8260 37772
rect 8540 37380 8596 37390
rect 8540 37286 8596 37324
rect 8764 37268 8820 37278
rect 8764 37266 9156 37268
rect 8764 37214 8766 37266
rect 8818 37214 9156 37266
rect 8764 37212 9156 37214
rect 8764 37202 8820 37212
rect 8652 37154 8708 37166
rect 8652 37102 8654 37154
rect 8706 37102 8708 37154
rect 8652 36484 8708 37102
rect 8652 36428 9044 36484
rect 8204 36418 8260 36428
rect 8876 36260 8932 36270
rect 7308 35870 7310 35922
rect 7362 35870 7364 35922
rect 7308 35858 7364 35870
rect 7420 35980 8148 36036
rect 6748 34914 7028 34916
rect 6748 34862 6750 34914
rect 6802 34862 7028 34914
rect 6748 34860 7028 34862
rect 7084 35252 7140 35262
rect 7084 34914 7140 35196
rect 7084 34862 7086 34914
rect 7138 34862 7140 34914
rect 6748 34850 6804 34860
rect 7084 34850 7140 34862
rect 7308 34916 7364 34926
rect 7420 34916 7476 35980
rect 8092 35924 8148 35980
rect 8204 35924 8260 35934
rect 8092 35922 8260 35924
rect 8092 35870 8206 35922
rect 8258 35870 8260 35922
rect 8092 35868 8260 35870
rect 8204 35858 8260 35868
rect 8876 35922 8932 36204
rect 8876 35870 8878 35922
rect 8930 35870 8932 35922
rect 8876 35858 8932 35870
rect 8652 35812 8708 35822
rect 8652 35718 8708 35756
rect 8988 35810 9044 36428
rect 8988 35758 8990 35810
rect 9042 35758 9044 35810
rect 8988 35746 9044 35758
rect 7980 35698 8036 35710
rect 7980 35646 7982 35698
rect 8034 35646 8036 35698
rect 7980 35476 8036 35646
rect 8092 35700 8148 35710
rect 8092 35698 8260 35700
rect 8092 35646 8094 35698
rect 8146 35646 8260 35698
rect 8092 35644 8260 35646
rect 8092 35634 8148 35644
rect 7980 35420 8148 35476
rect 7868 35364 7924 35374
rect 7308 34914 7476 34916
rect 7308 34862 7310 34914
rect 7362 34862 7476 34914
rect 7308 34860 7476 34862
rect 7756 35140 7812 35150
rect 7308 34850 7364 34860
rect 7756 34804 7812 35084
rect 7868 34804 7924 35308
rect 8092 35026 8148 35420
rect 8204 35364 8260 35644
rect 8204 35298 8260 35308
rect 8428 35698 8484 35710
rect 8428 35646 8430 35698
rect 8482 35646 8484 35698
rect 8092 34974 8094 35026
rect 8146 34974 8148 35026
rect 8092 34962 8148 34974
rect 7980 34804 8036 34814
rect 7868 34802 8036 34804
rect 7868 34750 7982 34802
rect 8034 34750 8036 34802
rect 7868 34748 8036 34750
rect 7756 34710 7812 34748
rect 6860 34690 6916 34702
rect 6860 34638 6862 34690
rect 6914 34638 6916 34690
rect 6860 34244 6916 34638
rect 6860 34178 6916 34188
rect 7756 34468 7812 34478
rect 7756 33346 7812 34412
rect 7980 34020 8036 34748
rect 8204 34804 8260 34814
rect 8428 34804 8484 35646
rect 8876 35026 8932 35038
rect 8876 34974 8878 35026
rect 8930 34974 8932 35026
rect 8764 34916 8820 34926
rect 8764 34822 8820 34860
rect 8260 34748 8484 34804
rect 8876 34804 8932 34974
rect 8204 34710 8260 34748
rect 8876 34738 8932 34748
rect 9100 34692 9156 37212
rect 9212 34914 9268 37886
rect 9660 35588 9716 37998
rect 9772 37940 9828 38612
rect 9884 38164 9940 38670
rect 10332 38164 10388 38892
rect 10444 38946 10500 39004
rect 10444 38894 10446 38946
rect 10498 38894 10500 38946
rect 10444 38882 10500 38894
rect 10556 38612 10612 39564
rect 11004 39060 11060 39070
rect 11004 38836 11060 39004
rect 10892 38834 11060 38836
rect 10892 38782 11006 38834
rect 11058 38782 11060 38834
rect 10892 38780 11060 38782
rect 10556 38546 10612 38556
rect 10780 38724 10836 38734
rect 10444 38164 10500 38174
rect 10332 38162 10500 38164
rect 10332 38110 10446 38162
rect 10498 38110 10500 38162
rect 10332 38108 10500 38110
rect 9884 38098 9940 38108
rect 10444 38098 10500 38108
rect 9772 37874 9828 37884
rect 9884 37938 9940 37950
rect 9884 37886 9886 37938
rect 9938 37886 9940 37938
rect 9884 37380 9940 37886
rect 10332 37940 10388 37950
rect 10332 37846 10388 37884
rect 9660 35252 9716 35532
rect 9660 35186 9716 35196
rect 9772 37268 9828 37278
rect 9772 36370 9828 37212
rect 9772 36318 9774 36370
rect 9826 36318 9828 36370
rect 9548 35028 9604 35038
rect 9212 34862 9214 34914
rect 9266 34862 9268 34914
rect 9212 34850 9268 34862
rect 9436 35026 9604 35028
rect 9436 34974 9550 35026
rect 9602 34974 9604 35026
rect 9436 34972 9604 34974
rect 9100 34626 9156 34636
rect 8092 34020 8148 34030
rect 7980 34018 8148 34020
rect 7980 33966 8094 34018
rect 8146 33966 8148 34018
rect 7980 33964 8148 33966
rect 7980 33458 8036 33964
rect 8092 33954 8148 33964
rect 7980 33406 7982 33458
rect 8034 33406 8036 33458
rect 7980 33394 8036 33406
rect 9436 33458 9492 34972
rect 9548 34962 9604 34972
rect 9772 34130 9828 36318
rect 9884 34916 9940 37324
rect 10556 37154 10612 37166
rect 10556 37102 10558 37154
rect 10610 37102 10612 37154
rect 10556 35364 10612 37102
rect 10556 35298 10612 35308
rect 10780 35140 10836 38668
rect 10892 38162 10948 38780
rect 11004 38770 11060 38780
rect 11564 39060 11620 39070
rect 10892 38110 10894 38162
rect 10946 38110 10948 38162
rect 10892 38098 10948 38110
rect 11340 38722 11396 38734
rect 11340 38670 11342 38722
rect 11394 38670 11396 38722
rect 11340 38612 11396 38670
rect 11340 37380 11396 38556
rect 11564 38162 11620 39004
rect 11676 38946 11732 38958
rect 11676 38894 11678 38946
rect 11730 38894 11732 38946
rect 11676 38724 11732 38894
rect 11676 38658 11732 38668
rect 11788 38388 11844 40348
rect 12348 40348 12516 40404
rect 12684 40514 12852 40516
rect 12684 40462 12798 40514
rect 12850 40462 12852 40514
rect 12684 40460 12852 40462
rect 12348 40068 12404 40348
rect 12460 40234 12516 40246
rect 12460 40182 12462 40234
rect 12514 40182 12516 40234
rect 12460 40180 12516 40182
rect 12684 40180 12740 40460
rect 12796 40450 12852 40460
rect 13132 40628 13188 40638
rect 13132 40514 13188 40572
rect 13132 40462 13134 40514
rect 13186 40462 13188 40514
rect 13132 40450 13188 40462
rect 12460 40124 12740 40180
rect 12348 40012 12516 40068
rect 12348 39394 12404 39406
rect 12348 39342 12350 39394
rect 12402 39342 12404 39394
rect 12012 38836 12068 38846
rect 12348 38836 12404 39342
rect 12012 38834 12404 38836
rect 12012 38782 12014 38834
rect 12066 38782 12404 38834
rect 12012 38780 12404 38782
rect 12460 38834 12516 40012
rect 12908 39396 12964 39406
rect 12908 38946 12964 39340
rect 12908 38894 12910 38946
rect 12962 38894 12964 38946
rect 12908 38882 12964 38894
rect 13132 38948 13188 38958
rect 13132 38854 13188 38892
rect 12460 38782 12462 38834
rect 12514 38782 12516 38834
rect 12012 38668 12068 38780
rect 12460 38770 12516 38782
rect 13580 38836 13636 40908
rect 13804 40516 13860 40526
rect 13916 40516 13972 41020
rect 13804 40514 13972 40516
rect 13804 40462 13806 40514
rect 13858 40462 13972 40514
rect 13804 40460 13972 40462
rect 14140 40516 14196 40526
rect 13804 38948 13860 40460
rect 14140 40422 14196 40460
rect 14476 40516 14532 40526
rect 13804 38882 13860 38892
rect 14140 40292 14196 40302
rect 14140 39394 14196 40236
rect 14476 39618 14532 40460
rect 15932 40516 15988 40526
rect 15932 40422 15988 40460
rect 15708 40404 15764 40414
rect 15708 40310 15764 40348
rect 16268 40402 16324 41804
rect 16268 40350 16270 40402
rect 16322 40350 16324 40402
rect 16268 40338 16324 40350
rect 16604 40516 16660 40526
rect 16492 40178 16548 40190
rect 16492 40126 16494 40178
rect 16546 40126 16548 40178
rect 14476 39566 14478 39618
rect 14530 39566 14532 39618
rect 14476 39554 14532 39566
rect 15932 39618 15988 39630
rect 15932 39566 15934 39618
rect 15986 39566 15988 39618
rect 15484 39508 15540 39518
rect 15484 39506 15876 39508
rect 15484 39454 15486 39506
rect 15538 39454 15876 39506
rect 15484 39452 15876 39454
rect 15484 39442 15540 39452
rect 14140 39342 14142 39394
rect 14194 39342 14196 39394
rect 13580 38742 13636 38780
rect 12684 38724 12740 38734
rect 12012 38612 12516 38668
rect 12684 38630 12740 38668
rect 11788 38332 12068 38388
rect 11564 38110 11566 38162
rect 11618 38110 11620 38162
rect 11564 38098 11620 38110
rect 11900 38164 11956 38174
rect 11340 37314 11396 37324
rect 10892 35588 10948 35598
rect 10892 35252 10948 35532
rect 10892 35186 10948 35196
rect 10780 35074 10836 35084
rect 11676 35140 11732 35150
rect 9996 34916 10052 34926
rect 9884 34860 9996 34916
rect 9996 34822 10052 34860
rect 11452 34916 11508 34926
rect 11452 34822 11508 34860
rect 11228 34804 11284 34814
rect 11228 34710 11284 34748
rect 11564 34802 11620 34814
rect 11564 34750 11566 34802
rect 11618 34750 11620 34802
rect 9772 34078 9774 34130
rect 9826 34078 9828 34130
rect 9772 34066 9828 34078
rect 9884 34692 9940 34702
rect 9436 33406 9438 33458
rect 9490 33406 9492 33458
rect 9436 33394 9492 33406
rect 9884 33908 9940 34636
rect 10556 34020 10612 34030
rect 11228 34020 11284 34030
rect 10556 34018 11172 34020
rect 10556 33966 10558 34018
rect 10610 33966 11172 34018
rect 10556 33964 11172 33966
rect 10556 33954 10612 33964
rect 7756 33294 7758 33346
rect 7810 33294 7812 33346
rect 7756 33282 7812 33294
rect 9884 33346 9940 33852
rect 11116 33570 11172 33964
rect 11116 33518 11118 33570
rect 11170 33518 11172 33570
rect 11116 33506 11172 33518
rect 10332 33460 10388 33470
rect 10332 33366 10388 33404
rect 11228 33458 11284 33964
rect 11228 33406 11230 33458
rect 11282 33406 11284 33458
rect 11228 33394 11284 33406
rect 9884 33294 9886 33346
rect 9938 33294 9940 33346
rect 9884 33282 9940 33294
rect 7084 33236 7140 33246
rect 7084 33234 7364 33236
rect 7084 33182 7086 33234
rect 7138 33182 7364 33234
rect 7084 33180 7364 33182
rect 7084 33170 7140 33180
rect 6748 33124 6804 33134
rect 6972 33124 7028 33134
rect 6748 33030 6804 33068
rect 6860 33122 7028 33124
rect 6860 33070 6974 33122
rect 7026 33070 7028 33122
rect 6860 33068 7028 33070
rect 6860 32004 6916 33068
rect 6972 33058 7028 33068
rect 6748 31948 6916 32004
rect 6636 31892 6692 31902
rect 6524 31836 6636 31892
rect 6636 31826 6692 31836
rect 5964 31726 5966 31778
rect 6018 31726 6020 31778
rect 5964 31714 6020 31726
rect 6412 31778 6468 31790
rect 6412 31726 6414 31778
rect 6466 31726 6468 31778
rect 5628 31666 5684 31678
rect 5628 31614 5630 31666
rect 5682 31614 5684 31666
rect 5628 30436 5684 31614
rect 5740 31668 5796 31678
rect 5740 31574 5796 31612
rect 6188 31668 6244 31678
rect 5628 30380 5908 30436
rect 5628 30212 5684 30222
rect 5628 30118 5684 30156
rect 5740 30100 5796 30110
rect 5740 30006 5796 30044
rect 4844 29922 4900 29932
rect 5740 29876 5796 29886
rect 4620 29586 4676 29596
rect 5068 29652 5124 29662
rect 5068 29558 5124 29596
rect 5628 29538 5684 29550
rect 5628 29486 5630 29538
rect 5682 29486 5684 29538
rect 1820 29426 1876 29438
rect 1820 29374 1822 29426
rect 1874 29374 1876 29426
rect 1820 27748 1876 29374
rect 3164 29428 3220 29438
rect 2492 29316 2548 29326
rect 2492 29222 2548 29260
rect 3052 28868 3108 28878
rect 1820 27074 1876 27692
rect 2492 28644 2548 28654
rect 2492 27186 2548 28588
rect 2492 27134 2494 27186
rect 2546 27134 2548 27186
rect 2492 27122 2548 27134
rect 3052 28530 3108 28812
rect 3052 28478 3054 28530
rect 3106 28478 3108 28530
rect 1820 27022 1822 27074
rect 1874 27022 1876 27074
rect 1708 26178 1764 26190
rect 1708 26126 1710 26178
rect 1762 26126 1764 26178
rect 1708 25284 1764 26126
rect 1708 25218 1764 25228
rect 1820 24722 1876 27022
rect 3052 25508 3108 28478
rect 3164 28530 3220 29372
rect 4620 29428 4676 29438
rect 3724 29316 3780 29326
rect 3612 29204 3668 29214
rect 3500 28644 3556 28654
rect 3164 28478 3166 28530
rect 3218 28478 3220 28530
rect 3164 28466 3220 28478
rect 3388 28588 3500 28644
rect 3388 28530 3444 28588
rect 3500 28578 3556 28588
rect 3612 28642 3668 29148
rect 3724 28754 3780 29260
rect 4620 29314 4676 29372
rect 4620 29262 4622 29314
rect 4674 29262 4676 29314
rect 4620 29250 4676 29262
rect 4844 29426 4900 29438
rect 4844 29374 4846 29426
rect 4898 29374 4900 29426
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4844 28868 4900 29374
rect 4172 28812 4900 28868
rect 5180 29426 5236 29438
rect 5180 29374 5182 29426
rect 5234 29374 5236 29426
rect 5180 28868 5236 29374
rect 5628 29428 5684 29486
rect 5740 29540 5796 29820
rect 5852 29652 5908 30380
rect 6188 30210 6244 31612
rect 6188 30158 6190 30210
rect 6242 30158 6244 30210
rect 6188 30146 6244 30158
rect 6412 30210 6468 31726
rect 6636 31556 6692 31566
rect 6636 31462 6692 31500
rect 6748 31332 6804 31948
rect 6524 31276 6804 31332
rect 6860 31666 6916 31678
rect 6860 31614 6862 31666
rect 6914 31614 6916 31666
rect 6524 30884 6580 31276
rect 6860 31220 6916 31614
rect 7084 31668 7140 31678
rect 6972 31220 7028 31230
rect 6860 31218 7028 31220
rect 6860 31166 6974 31218
rect 7026 31166 7028 31218
rect 6860 31164 7028 31166
rect 6972 31154 7028 31164
rect 7084 30996 7140 31612
rect 7084 30930 7140 30940
rect 7196 31332 7252 31342
rect 7196 31218 7252 31276
rect 7196 31166 7198 31218
rect 7250 31166 7252 31218
rect 6524 30882 6692 30884
rect 6524 30830 6526 30882
rect 6578 30830 6692 30882
rect 6524 30828 6692 30830
rect 6524 30818 6580 30828
rect 6412 30158 6414 30210
rect 6466 30158 6468 30210
rect 6412 30146 6468 30158
rect 5964 30100 6020 30110
rect 5964 30006 6020 30044
rect 6636 30098 6692 30828
rect 7196 30772 7252 31166
rect 7196 30706 7252 30716
rect 7308 31108 7364 33180
rect 8988 33124 9044 33134
rect 8988 33122 9380 33124
rect 8988 33070 8990 33122
rect 9042 33070 9380 33122
rect 8988 33068 9380 33070
rect 8988 33058 9044 33068
rect 7756 32676 7812 32686
rect 7756 31890 7812 32620
rect 8764 32676 8820 32686
rect 8764 32582 8820 32620
rect 8316 32562 8372 32574
rect 8316 32510 8318 32562
rect 8370 32510 8372 32562
rect 8316 32452 8372 32510
rect 8876 32564 8932 32574
rect 8876 32562 9044 32564
rect 8876 32510 8878 32562
rect 8930 32510 9044 32562
rect 8876 32508 9044 32510
rect 8876 32498 8932 32508
rect 8316 32386 8372 32396
rect 7756 31838 7758 31890
rect 7810 31838 7812 31890
rect 7756 31332 7812 31838
rect 8764 32338 8820 32350
rect 8764 32286 8766 32338
rect 8818 32286 8820 32338
rect 7756 31266 7812 31276
rect 8652 31668 8708 31678
rect 8092 31220 8148 31230
rect 8092 31218 8484 31220
rect 8092 31166 8094 31218
rect 8146 31166 8484 31218
rect 8092 31164 8484 31166
rect 8092 31154 8148 31164
rect 7756 31108 7812 31118
rect 7308 31106 7812 31108
rect 7308 31054 7310 31106
rect 7362 31054 7758 31106
rect 7810 31054 7812 31106
rect 7308 31052 7812 31054
rect 7308 30212 7364 31052
rect 7756 31042 7812 31052
rect 7868 31108 7924 31118
rect 8428 31108 8484 31164
rect 8652 31218 8708 31612
rect 8652 31166 8654 31218
rect 8706 31166 8708 31218
rect 8652 31154 8708 31166
rect 8540 31108 8596 31118
rect 7868 31106 8036 31108
rect 7868 31054 7870 31106
rect 7922 31054 8036 31106
rect 7868 31052 8036 31054
rect 8428 31106 8596 31108
rect 8428 31054 8542 31106
rect 8594 31054 8596 31106
rect 8428 31052 8596 31054
rect 8764 31108 8820 32286
rect 8876 31108 8932 31118
rect 8764 31106 8932 31108
rect 8764 31054 8878 31106
rect 8930 31054 8932 31106
rect 8764 31052 8932 31054
rect 7868 31042 7924 31052
rect 7084 30210 7364 30212
rect 7084 30158 7310 30210
rect 7362 30158 7364 30210
rect 7084 30156 7364 30158
rect 6636 30046 6638 30098
rect 6690 30046 6692 30098
rect 6188 29988 6244 29998
rect 6188 29764 6244 29932
rect 6636 29988 6692 30046
rect 6748 30100 6804 30110
rect 6972 30100 7028 30110
rect 6748 30098 6916 30100
rect 6748 30046 6750 30098
rect 6802 30046 6916 30098
rect 6748 30044 6916 30046
rect 6748 30034 6804 30044
rect 6636 29922 6692 29932
rect 5964 29652 6020 29662
rect 5852 29650 6020 29652
rect 5852 29598 5966 29650
rect 6018 29598 6020 29650
rect 5852 29596 6020 29598
rect 5964 29586 6020 29596
rect 6188 29650 6244 29708
rect 6188 29598 6190 29650
rect 6242 29598 6244 29650
rect 6188 29586 6244 29598
rect 6300 29540 6356 29550
rect 5740 29538 5908 29540
rect 5740 29486 5742 29538
rect 5794 29486 5908 29538
rect 5740 29484 5908 29486
rect 5740 29474 5796 29484
rect 5628 29362 5684 29372
rect 5628 29204 5684 29214
rect 5628 29110 5684 29148
rect 3724 28702 3726 28754
rect 3778 28702 3780 28754
rect 3724 28690 3780 28702
rect 3836 28756 3892 28766
rect 3892 28700 4116 28756
rect 3836 28690 3892 28700
rect 3612 28590 3614 28642
rect 3666 28590 3668 28642
rect 3612 28578 3668 28590
rect 4060 28642 4116 28700
rect 4060 28590 4062 28642
rect 4114 28590 4116 28642
rect 4060 28578 4116 28590
rect 3388 28478 3390 28530
rect 3442 28478 3444 28530
rect 3388 28466 3444 28478
rect 3948 28530 4004 28542
rect 3948 28478 3950 28530
rect 4002 28478 4004 28530
rect 3948 28420 4004 28478
rect 4172 28420 4228 28812
rect 5068 28756 5124 28766
rect 4620 28642 4676 28654
rect 4620 28590 4622 28642
rect 4674 28590 4676 28642
rect 4508 28532 4564 28542
rect 3948 28364 4228 28420
rect 4284 28530 4564 28532
rect 4284 28478 4510 28530
rect 4562 28478 4564 28530
rect 4284 28476 4564 28478
rect 4172 27748 4228 27758
rect 4172 26964 4228 27692
rect 4172 26898 4228 26908
rect 3724 26292 3780 26302
rect 3500 26236 3724 26292
rect 3500 25730 3556 26236
rect 3724 26226 3780 26236
rect 3836 26180 3892 26190
rect 3836 26086 3892 26124
rect 3500 25678 3502 25730
rect 3554 25678 3556 25730
rect 3500 25666 3556 25678
rect 4172 25732 4228 25742
rect 4284 25732 4340 28476
rect 4508 28466 4564 28476
rect 4620 28532 4676 28590
rect 4732 28644 4788 28654
rect 4732 28550 4788 28588
rect 5068 28642 5124 28700
rect 5068 28590 5070 28642
rect 5122 28590 5124 28642
rect 4620 28466 4676 28476
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4620 27300 4676 27310
rect 4620 27188 4676 27244
rect 4620 27186 4788 27188
rect 4620 27134 4622 27186
rect 4674 27134 4788 27186
rect 4620 27132 4788 27134
rect 4620 27122 4676 27132
rect 4620 26964 4676 26974
rect 4620 26290 4676 26908
rect 4620 26238 4622 26290
rect 4674 26238 4676 26290
rect 4620 26226 4676 26238
rect 4732 26068 4788 27132
rect 5068 26908 5124 28590
rect 5180 28420 5236 28812
rect 5628 28530 5684 28542
rect 5628 28478 5630 28530
rect 5682 28478 5684 28530
rect 5404 28420 5460 28430
rect 5180 28364 5404 28420
rect 5404 28354 5460 28364
rect 5628 27300 5684 28478
rect 5628 27234 5684 27244
rect 5852 26908 5908 29484
rect 6300 29446 6356 29484
rect 6860 29540 6916 30044
rect 6972 30006 7028 30044
rect 6972 29652 7028 29662
rect 7084 29652 7140 30156
rect 7308 30146 7364 30156
rect 7420 30772 7476 30782
rect 6972 29650 7140 29652
rect 6972 29598 6974 29650
rect 7026 29598 7140 29650
rect 6972 29596 7140 29598
rect 7196 29986 7252 29998
rect 7196 29934 7198 29986
rect 7250 29934 7252 29986
rect 7196 29764 7252 29934
rect 6972 29586 7028 29596
rect 6860 29474 6916 29484
rect 6076 29428 6132 29438
rect 6076 28644 6132 29372
rect 6748 29426 6804 29438
rect 6748 29374 6750 29426
rect 6802 29374 6804 29426
rect 6188 28644 6244 28654
rect 6076 28642 6244 28644
rect 6076 28590 6190 28642
rect 6242 28590 6244 28642
rect 6076 28588 6244 28590
rect 6188 28578 6244 28588
rect 5068 26852 5460 26908
rect 4844 26292 4900 26302
rect 4844 26198 4900 26236
rect 5180 26290 5236 26302
rect 5180 26238 5182 26290
rect 5234 26238 5236 26290
rect 5068 26180 5124 26190
rect 5068 26086 5124 26124
rect 4732 26012 4900 26068
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4844 25732 4900 26012
rect 4284 25676 4452 25732
rect 4172 25620 4228 25676
rect 4172 25564 4340 25620
rect 3052 25414 3108 25452
rect 3948 25508 4004 25518
rect 3948 25414 4004 25452
rect 4284 25506 4340 25564
rect 4284 25454 4286 25506
rect 4338 25454 4340 25506
rect 4284 25442 4340 25454
rect 4396 25506 4452 25676
rect 4396 25454 4398 25506
rect 4450 25454 4452 25506
rect 4396 25442 4452 25454
rect 4620 25676 4900 25732
rect 5180 25732 5236 26238
rect 3612 25396 3668 25406
rect 3612 25302 3668 25340
rect 4620 25394 4676 25676
rect 5180 25666 5236 25676
rect 5404 26290 5460 26852
rect 5404 26238 5406 26290
rect 5458 26238 5460 26290
rect 4732 25508 4788 25518
rect 4732 25414 4788 25452
rect 4620 25342 4622 25394
rect 4674 25342 4676 25394
rect 2716 25282 2772 25294
rect 2716 25230 2718 25282
rect 2770 25230 2772 25282
rect 2716 24836 2772 25230
rect 2940 25284 2996 25294
rect 2940 25190 2996 25228
rect 3500 25284 3556 25294
rect 2716 24770 2772 24780
rect 1820 24670 1822 24722
rect 1874 24670 1876 24722
rect 1820 24658 1876 24670
rect 2492 24612 2548 24622
rect 2492 24518 2548 24556
rect 3276 23716 3332 23726
rect 3276 23268 3332 23660
rect 3500 23604 3556 25228
rect 4060 25284 4116 25294
rect 4620 25284 4676 25342
rect 4060 25282 4228 25284
rect 4060 25230 4062 25282
rect 4114 25230 4228 25282
rect 4060 25228 4228 25230
rect 4060 25218 4116 25228
rect 4172 25172 4228 25228
rect 4396 25228 4676 25284
rect 4396 25172 4452 25228
rect 4172 25116 4452 25172
rect 5404 24948 5460 26238
rect 5628 26852 5908 26908
rect 5964 28420 6020 28430
rect 5628 25508 5684 26852
rect 5964 26514 6020 28364
rect 6636 28420 6692 28430
rect 6636 28326 6692 28364
rect 6748 28308 6804 29374
rect 7196 28530 7252 29708
rect 7308 29988 7364 29998
rect 7308 29426 7364 29932
rect 7308 29374 7310 29426
rect 7362 29374 7364 29426
rect 7308 29362 7364 29374
rect 7420 29428 7476 30716
rect 7980 30212 8036 31052
rect 8540 31042 8596 31052
rect 8876 31042 8932 31052
rect 8316 30996 8372 31006
rect 8316 30902 8372 30940
rect 8988 30324 9044 32508
rect 8540 30268 9044 30324
rect 7980 30156 8484 30212
rect 7532 30100 7588 30110
rect 7532 30006 7588 30044
rect 7868 30098 7924 30110
rect 7868 30046 7870 30098
rect 7922 30046 7924 30098
rect 7756 29988 7812 29998
rect 7644 29986 7812 29988
rect 7644 29934 7758 29986
rect 7810 29934 7812 29986
rect 7644 29932 7812 29934
rect 7644 29652 7700 29932
rect 7756 29922 7812 29932
rect 7868 29988 7924 30046
rect 7868 29922 7924 29932
rect 7980 29764 8036 30156
rect 8428 30100 8484 30156
rect 8428 30006 8484 30044
rect 8540 30210 8596 30268
rect 9212 30212 9268 30222
rect 8540 30158 8542 30210
rect 8594 30158 8596 30210
rect 8204 29988 8260 29998
rect 8204 29986 8372 29988
rect 8204 29934 8206 29986
rect 8258 29934 8372 29986
rect 8204 29932 8372 29934
rect 8204 29922 8260 29932
rect 7532 29428 7588 29438
rect 7420 29426 7588 29428
rect 7420 29374 7534 29426
rect 7586 29374 7588 29426
rect 7420 29372 7588 29374
rect 7532 29362 7588 29372
rect 7308 28644 7364 28654
rect 7644 28644 7700 29596
rect 7756 29708 8036 29764
rect 7756 29426 7812 29708
rect 7756 29374 7758 29426
rect 7810 29374 7812 29426
rect 7756 29362 7812 29374
rect 7868 29540 7924 29550
rect 7868 29204 7924 29484
rect 7980 29428 8036 29438
rect 7980 29426 8260 29428
rect 7980 29374 7982 29426
rect 8034 29374 8260 29426
rect 7980 29372 8260 29374
rect 7980 29362 8036 29372
rect 7868 29148 8036 29204
rect 7308 28642 7700 28644
rect 7308 28590 7310 28642
rect 7362 28590 7700 28642
rect 7308 28588 7700 28590
rect 7308 28578 7364 28588
rect 7196 28478 7198 28530
rect 7250 28478 7252 28530
rect 7196 28466 7252 28478
rect 7980 28530 8036 29148
rect 7980 28478 7982 28530
rect 8034 28478 8036 28530
rect 7980 28466 8036 28478
rect 8092 29202 8148 29214
rect 8092 29150 8094 29202
rect 8146 29150 8148 29202
rect 8092 28532 8148 29150
rect 8092 28466 8148 28476
rect 8204 28756 8260 29372
rect 8316 29426 8372 29932
rect 8540 29540 8596 30158
rect 8540 29474 8596 29484
rect 8988 30156 9212 30212
rect 8988 29538 9044 30156
rect 8988 29486 8990 29538
rect 9042 29486 9044 29538
rect 8988 29474 9044 29486
rect 8316 29374 8318 29426
rect 8370 29374 8372 29426
rect 8316 29362 8372 29374
rect 8652 29426 8708 29438
rect 8652 29374 8654 29426
rect 8706 29374 8708 29426
rect 8540 29316 8596 29326
rect 8540 29222 8596 29260
rect 8204 28700 8484 28756
rect 7644 28418 7700 28430
rect 7644 28366 7646 28418
rect 7698 28366 7700 28418
rect 7084 28308 7140 28318
rect 6748 28252 7084 28308
rect 6076 27746 6132 27758
rect 6076 27694 6078 27746
rect 6130 27694 6132 27746
rect 6076 27074 6132 27694
rect 6076 27022 6078 27074
rect 6130 27022 6132 27074
rect 6076 26964 6132 27022
rect 6748 26908 6804 28252
rect 7084 28242 7140 28252
rect 6076 26898 6132 26908
rect 5964 26462 5966 26514
rect 6018 26462 6020 26514
rect 5964 26450 6020 26462
rect 6300 26852 6804 26908
rect 6300 26514 6356 26852
rect 6300 26462 6302 26514
rect 6354 26462 6356 26514
rect 6300 26450 6356 26462
rect 6748 25620 6804 26852
rect 6860 26962 6916 26974
rect 6860 26910 6862 26962
rect 6914 26910 6916 26962
rect 6860 26516 6916 26910
rect 6860 26450 6916 26460
rect 7084 26292 7140 26302
rect 7308 26292 7364 26302
rect 7084 26290 7364 26292
rect 7084 26238 7086 26290
rect 7138 26238 7310 26290
rect 7362 26238 7364 26290
rect 7084 26236 7364 26238
rect 7084 26226 7140 26236
rect 6748 25564 6916 25620
rect 5628 25394 5684 25452
rect 5628 25342 5630 25394
rect 5682 25342 5684 25394
rect 5628 25330 5684 25342
rect 6748 25396 6804 25406
rect 6748 25302 6804 25340
rect 5964 25284 6020 25294
rect 6412 25284 6468 25294
rect 5964 25282 6412 25284
rect 5964 25230 5966 25282
rect 6018 25230 6412 25282
rect 5964 25228 6412 25230
rect 5964 25218 6020 25228
rect 5964 24948 6020 24958
rect 5404 24946 6020 24948
rect 5404 24894 5966 24946
rect 6018 24894 6020 24946
rect 5404 24892 6020 24894
rect 5180 24836 5236 24846
rect 4844 24722 4900 24734
rect 4844 24670 4846 24722
rect 4898 24670 4900 24722
rect 4620 24612 4676 24622
rect 4284 24610 4676 24612
rect 4284 24558 4622 24610
rect 4674 24558 4676 24610
rect 4284 24556 4676 24558
rect 4172 23826 4228 23838
rect 4172 23774 4174 23826
rect 4226 23774 4228 23826
rect 4172 23716 4228 23774
rect 4172 23650 4228 23660
rect 4284 23714 4340 24556
rect 4620 24546 4676 24556
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4844 24164 4900 24670
rect 5180 24722 5236 24780
rect 5180 24670 5182 24722
rect 5234 24670 5236 24722
rect 5180 24658 5236 24670
rect 5404 24722 5460 24892
rect 5964 24882 6020 24892
rect 5404 24670 5406 24722
rect 5458 24670 5460 24722
rect 5404 24658 5460 24670
rect 5068 24612 5124 24622
rect 5068 24518 5124 24556
rect 4508 24108 4900 24164
rect 4508 23938 4564 24108
rect 4508 23886 4510 23938
rect 4562 23886 4564 23938
rect 4508 23874 4564 23886
rect 5964 23940 6020 23950
rect 6076 23940 6132 25228
rect 6412 25190 6468 25228
rect 6300 24722 6356 24734
rect 6300 24670 6302 24722
rect 6354 24670 6356 24722
rect 6300 24612 6356 24670
rect 6748 24612 6804 24622
rect 6300 24610 6804 24612
rect 6300 24558 6750 24610
rect 6802 24558 6804 24610
rect 6300 24556 6804 24558
rect 6748 24052 6804 24556
rect 6748 23986 6804 23996
rect 5964 23938 6132 23940
rect 5964 23886 5966 23938
rect 6018 23886 6132 23938
rect 5964 23884 6132 23886
rect 6188 23940 6244 23950
rect 5964 23874 6020 23884
rect 5852 23828 5908 23838
rect 4284 23662 4286 23714
rect 4338 23662 4340 23714
rect 3612 23604 3668 23614
rect 3500 23548 3612 23604
rect 3612 23538 3668 23548
rect 3948 23380 4004 23390
rect 4284 23380 4340 23662
rect 5628 23714 5684 23726
rect 5628 23662 5630 23714
rect 5682 23662 5684 23714
rect 4508 23604 4564 23614
rect 3948 23378 4452 23380
rect 3948 23326 3950 23378
rect 4002 23326 4452 23378
rect 3948 23324 4452 23326
rect 3948 23314 4004 23324
rect 3164 23266 3332 23268
rect 3164 23214 3278 23266
rect 3330 23214 3332 23266
rect 3164 23212 3332 23214
rect 1708 22370 1764 22382
rect 1708 22318 1710 22370
rect 1762 22318 1764 22370
rect 1708 20802 1764 22318
rect 2492 22258 2548 22270
rect 2492 22206 2494 22258
rect 2546 22206 2548 22258
rect 2492 21812 2548 22206
rect 2492 21746 2548 21756
rect 3164 21698 3220 23212
rect 3276 23202 3332 23212
rect 3388 23266 3444 23278
rect 3388 23214 3390 23266
rect 3442 23214 3444 23266
rect 3388 22596 3444 23214
rect 3388 22530 3444 22540
rect 3612 23154 3668 23166
rect 3612 23102 3614 23154
rect 3666 23102 3668 23154
rect 3164 21646 3166 21698
rect 3218 21646 3220 21698
rect 3164 21634 3220 21646
rect 3276 21698 3332 21710
rect 3276 21646 3278 21698
rect 3330 21646 3332 21698
rect 2492 21476 2548 21486
rect 2492 20914 2548 21420
rect 3276 21028 3332 21646
rect 3500 21700 3556 21710
rect 3500 21606 3556 21644
rect 3612 21586 3668 23102
rect 4060 23156 4116 23166
rect 4060 23062 4116 23100
rect 4396 23154 4452 23324
rect 4508 23266 4564 23548
rect 5628 23604 5684 23662
rect 5628 23538 5684 23548
rect 5852 23378 5908 23772
rect 5852 23326 5854 23378
rect 5906 23326 5908 23378
rect 5852 23314 5908 23326
rect 4508 23214 4510 23266
rect 4562 23214 4564 23266
rect 4508 23202 4564 23214
rect 5964 23266 6020 23278
rect 5964 23214 5966 23266
rect 6018 23214 6020 23266
rect 4396 23102 4398 23154
rect 4450 23102 4452 23154
rect 4396 23090 4452 23102
rect 5404 23154 5460 23166
rect 5404 23102 5406 23154
rect 5458 23102 5460 23154
rect 3948 22930 4004 22942
rect 3948 22878 3950 22930
rect 4002 22878 4004 22930
rect 3836 21812 3892 21822
rect 3836 21718 3892 21756
rect 3612 21534 3614 21586
rect 3666 21534 3668 21586
rect 3612 21522 3668 21534
rect 3948 21586 4004 22878
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4620 22596 4676 22606
rect 4620 22482 4676 22540
rect 5404 22596 5460 23102
rect 5404 22530 5460 22540
rect 5628 23156 5684 23166
rect 4620 22430 4622 22482
rect 4674 22430 4676 22482
rect 4620 22418 4676 22430
rect 5628 22372 5684 23100
rect 5964 22372 6020 23214
rect 5628 22278 5684 22316
rect 5852 22316 6020 22372
rect 4956 22148 5012 22158
rect 4396 21700 4452 21710
rect 4452 21644 4564 21700
rect 4396 21634 4452 21644
rect 3948 21534 3950 21586
rect 4002 21534 4004 21586
rect 3948 21522 4004 21534
rect 4284 21588 4340 21598
rect 4284 21494 4340 21532
rect 4508 21586 4564 21644
rect 4956 21698 5012 22092
rect 4956 21646 4958 21698
rect 5010 21646 5012 21698
rect 4956 21634 5012 21646
rect 5740 22148 5796 22158
rect 5852 22148 5908 22316
rect 5740 22146 5908 22148
rect 5740 22094 5742 22146
rect 5794 22094 5908 22146
rect 5740 22092 5908 22094
rect 5964 22146 6020 22158
rect 5964 22094 5966 22146
rect 6018 22094 6020 22146
rect 4508 21534 4510 21586
rect 4562 21534 4564 21586
rect 4508 21522 4564 21534
rect 5180 21588 5236 21598
rect 5180 21494 5236 21532
rect 4732 21476 4788 21486
rect 4732 21382 4788 21420
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 3276 20962 3332 20972
rect 4620 21028 4676 21038
rect 2492 20862 2494 20914
rect 2546 20862 2548 20914
rect 2492 20850 2548 20862
rect 4620 20914 4676 20972
rect 5740 21028 5796 22092
rect 5964 21700 6020 22094
rect 6076 22148 6132 22158
rect 6076 22054 6132 22092
rect 6076 21700 6132 21710
rect 5964 21698 6132 21700
rect 5964 21646 6078 21698
rect 6130 21646 6132 21698
rect 5964 21644 6132 21646
rect 6076 21634 6132 21644
rect 5852 21588 5908 21598
rect 5852 21494 5908 21532
rect 5740 20962 5796 20972
rect 4620 20862 4622 20914
rect 4674 20862 4676 20914
rect 4620 20850 4676 20862
rect 1708 20750 1710 20802
rect 1762 20750 1764 20802
rect 1708 20188 1764 20750
rect 5740 20802 5796 20814
rect 5740 20750 5742 20802
rect 5794 20750 5796 20802
rect 4956 20580 5012 20590
rect 4844 20524 4956 20580
rect 1708 20132 1876 20188
rect 1820 19236 1876 20132
rect 1820 17666 1876 19180
rect 3388 19906 3444 19918
rect 3388 19854 3390 19906
rect 3442 19854 3444 19906
rect 3388 19236 3444 19854
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4620 19348 4676 19358
rect 3388 19170 3444 19180
rect 4396 19346 4676 19348
rect 4396 19294 4622 19346
rect 4674 19294 4676 19346
rect 4396 19292 4676 19294
rect 2492 19124 2548 19134
rect 2492 19030 2548 19068
rect 3612 18676 3668 18686
rect 4396 18676 4452 19292
rect 4620 19282 4676 19292
rect 3164 18452 3220 18462
rect 3164 18358 3220 18396
rect 3500 18452 3556 18462
rect 3612 18452 3668 18620
rect 3500 18450 3668 18452
rect 3500 18398 3502 18450
rect 3554 18398 3668 18450
rect 3500 18396 3668 18398
rect 3724 18674 4452 18676
rect 3724 18622 4398 18674
rect 4450 18622 4452 18674
rect 3724 18620 4452 18622
rect 3724 18450 3780 18620
rect 4396 18610 4452 18620
rect 4508 19124 4564 19134
rect 3724 18398 3726 18450
rect 3778 18398 3780 18450
rect 3500 18386 3556 18396
rect 3724 18386 3780 18398
rect 4060 18450 4116 18462
rect 4060 18398 4062 18450
rect 4114 18398 4116 18450
rect 1820 17614 1822 17666
rect 1874 17614 1876 17666
rect 1820 17602 1876 17614
rect 2492 17556 2548 17566
rect 2492 17554 3332 17556
rect 2492 17502 2494 17554
rect 2546 17502 3332 17554
rect 2492 17500 3332 17502
rect 2492 17490 2548 17500
rect 3276 16770 3332 17500
rect 4060 17444 4116 18398
rect 4508 18450 4564 19068
rect 4620 18676 4676 18686
rect 4844 18676 4900 20524
rect 4956 20514 5012 20524
rect 4676 18620 4900 18676
rect 5292 19236 5348 19246
rect 4620 18582 4676 18620
rect 4508 18398 4510 18450
rect 4562 18398 4564 18450
rect 4508 18386 4564 18398
rect 4956 18452 5012 18462
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 3388 16996 3444 17006
rect 3444 16940 3556 16996
rect 3388 16902 3444 16940
rect 3276 16718 3278 16770
rect 3330 16718 3332 16770
rect 3276 16706 3332 16718
rect 3052 16212 3108 16222
rect 2492 16210 3108 16212
rect 2492 16158 3054 16210
rect 3106 16158 3108 16210
rect 2492 16156 3108 16158
rect 3500 16212 3556 16940
rect 4060 16994 4116 17388
rect 4060 16942 4062 16994
rect 4114 16942 4116 16994
rect 3724 16772 3780 16782
rect 3612 16716 3724 16772
rect 3612 16658 3668 16716
rect 3724 16706 3780 16716
rect 3612 16606 3614 16658
rect 3666 16606 3668 16658
rect 3612 16594 3668 16606
rect 4060 16548 4116 16942
rect 4620 17778 4676 17790
rect 4620 17726 4622 17778
rect 4674 17726 4676 17778
rect 4284 16884 4340 16894
rect 4284 16790 4340 16828
rect 4508 16882 4564 16894
rect 4508 16830 4510 16882
rect 4562 16830 4564 16882
rect 4396 16772 4452 16782
rect 4396 16678 4452 16716
rect 4508 16660 4564 16830
rect 4620 16884 4676 17726
rect 4844 16996 4900 17006
rect 4844 16902 4900 16940
rect 4620 16818 4676 16828
rect 4508 16604 4900 16660
rect 4060 16492 4340 16548
rect 3500 16156 3668 16212
rect 2492 15426 2548 16156
rect 3052 16146 3108 16156
rect 3388 16100 3444 16110
rect 3388 16006 3444 16044
rect 3612 15988 3668 16156
rect 3836 16100 3892 16110
rect 4284 16100 4340 16492
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4844 16436 4900 16604
rect 4844 16210 4900 16380
rect 4844 16158 4846 16210
rect 4898 16158 4900 16210
rect 4844 16146 4900 16158
rect 4396 16100 4452 16110
rect 4284 16098 4452 16100
rect 4284 16046 4398 16098
rect 4450 16046 4452 16098
rect 4284 16044 4452 16046
rect 3836 16006 3892 16044
rect 3724 15988 3780 15998
rect 3612 15986 3780 15988
rect 3612 15934 3726 15986
rect 3778 15934 3780 15986
rect 3612 15932 3780 15934
rect 3164 15876 3220 15886
rect 3164 15874 3332 15876
rect 3164 15822 3166 15874
rect 3218 15822 3332 15874
rect 3164 15820 3332 15822
rect 3164 15810 3220 15820
rect 2492 15374 2494 15426
rect 2546 15374 2548 15426
rect 2492 15362 2548 15374
rect 1820 15314 1876 15326
rect 1820 15262 1822 15314
rect 1874 15262 1876 15314
rect 1820 15204 1876 15262
rect 1820 13746 1876 15148
rect 3276 14756 3332 15820
rect 3724 15148 3780 15932
rect 3948 15874 4004 15886
rect 3948 15822 3950 15874
rect 4002 15822 4004 15874
rect 3948 15148 4004 15822
rect 4396 15764 4452 16044
rect 4396 15708 4788 15764
rect 4620 15202 4676 15214
rect 4620 15150 4622 15202
rect 4674 15150 4676 15202
rect 4620 15148 4676 15150
rect 3724 15092 3892 15148
rect 3948 15092 4676 15148
rect 4732 15148 4788 15708
rect 4732 15092 4900 15148
rect 3500 14756 3556 14766
rect 3276 14754 3668 14756
rect 3276 14702 3502 14754
rect 3554 14702 3668 14754
rect 3276 14700 3668 14702
rect 3500 14690 3556 14700
rect 1820 13694 1822 13746
rect 1874 13694 1876 13746
rect 1820 12178 1876 13694
rect 2492 13634 2548 13646
rect 2492 13582 2494 13634
rect 2546 13582 2548 13634
rect 2492 13188 2548 13582
rect 2492 13122 2548 13132
rect 1820 12126 1822 12178
rect 1874 12126 1876 12178
rect 1820 12114 1876 12126
rect 2492 12066 2548 12078
rect 2492 12014 2494 12066
rect 2546 12014 2548 12066
rect 2492 11508 2548 12014
rect 3612 11620 3668 14700
rect 3836 14754 3892 15092
rect 3836 14702 3838 14754
rect 3890 14702 3892 14754
rect 3836 14690 3892 14702
rect 4060 14642 4116 15092
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4060 14590 4062 14642
rect 4114 14590 4116 14642
rect 4060 14578 4116 14590
rect 4396 14532 4452 14542
rect 4396 14438 4452 14476
rect 4844 14418 4900 15092
rect 4956 14532 5012 18396
rect 5292 18450 5348 19180
rect 5740 19236 5796 20750
rect 5740 19170 5796 19180
rect 5628 19124 5684 19134
rect 5628 19030 5684 19068
rect 5740 19012 5796 19022
rect 5740 18918 5796 18956
rect 5852 19010 5908 19022
rect 5852 18958 5854 19010
rect 5906 18958 5908 19010
rect 5292 18398 5294 18450
rect 5346 18398 5348 18450
rect 5292 18386 5348 18398
rect 5628 18452 5684 18462
rect 5852 18452 5908 18958
rect 5684 18396 5908 18452
rect 5628 18386 5684 18396
rect 6076 18340 6132 18350
rect 5740 18338 6132 18340
rect 5740 18286 6078 18338
rect 6130 18286 6132 18338
rect 5740 18284 6132 18286
rect 5628 17444 5684 17454
rect 5628 17350 5684 17388
rect 5404 16884 5460 16894
rect 5404 16790 5460 16828
rect 5180 16658 5236 16670
rect 5180 16606 5182 16658
rect 5234 16606 5236 16658
rect 5180 16436 5236 16606
rect 5180 16370 5236 16380
rect 5740 15538 5796 18284
rect 6076 18274 6132 18284
rect 5964 17442 6020 17454
rect 5964 17390 5966 17442
rect 6018 17390 6020 17442
rect 5852 16436 5908 16446
rect 5852 16210 5908 16380
rect 5852 16158 5854 16210
rect 5906 16158 5908 16210
rect 5852 16146 5908 16158
rect 5964 16100 6020 17390
rect 5964 16034 6020 16044
rect 6076 16882 6132 16894
rect 6076 16830 6078 16882
rect 6130 16830 6132 16882
rect 5740 15486 5742 15538
rect 5794 15486 5796 15538
rect 5740 15474 5796 15486
rect 5516 15316 5572 15326
rect 5516 15222 5572 15260
rect 6076 15314 6132 16830
rect 6188 15988 6244 23884
rect 6748 23828 6804 23838
rect 6860 23828 6916 25564
rect 7084 25506 7140 25518
rect 7084 25454 7086 25506
rect 7138 25454 7140 25506
rect 6748 23826 6916 23828
rect 6748 23774 6750 23826
rect 6802 23774 6916 23826
rect 6748 23772 6916 23774
rect 6748 23762 6804 23772
rect 6748 23604 6804 23614
rect 6524 23266 6580 23278
rect 6524 23214 6526 23266
rect 6578 23214 6580 23266
rect 6300 22596 6356 22606
rect 6300 22258 6356 22540
rect 6412 22372 6468 22382
rect 6524 22372 6580 23214
rect 6468 22316 6580 22372
rect 6412 22278 6468 22316
rect 6300 22206 6302 22258
rect 6354 22206 6356 22258
rect 6300 22194 6356 22206
rect 6748 21698 6804 23548
rect 6860 23266 6916 23772
rect 6860 23214 6862 23266
rect 6914 23214 6916 23266
rect 6860 23202 6916 23214
rect 6972 25396 7028 25406
rect 6860 21812 6916 21822
rect 6860 21718 6916 21756
rect 6748 21646 6750 21698
rect 6802 21646 6804 21698
rect 6748 21634 6804 21646
rect 6524 21586 6580 21598
rect 6524 21534 6526 21586
rect 6578 21534 6580 21586
rect 6300 21474 6356 21486
rect 6300 21422 6302 21474
rect 6354 21422 6356 21474
rect 6300 20916 6356 21422
rect 6524 21364 6580 21534
rect 6860 21364 6916 21374
rect 6524 21362 6916 21364
rect 6524 21310 6862 21362
rect 6914 21310 6916 21362
rect 6524 21308 6916 21310
rect 6860 21298 6916 21308
rect 6412 20916 6468 20926
rect 6300 20914 6468 20916
rect 6300 20862 6414 20914
rect 6466 20862 6468 20914
rect 6300 20860 6468 20862
rect 6412 20850 6468 20860
rect 6524 19796 6580 19806
rect 6524 19234 6580 19740
rect 6524 19182 6526 19234
rect 6578 19182 6580 19234
rect 6524 19170 6580 19182
rect 6860 19236 6916 19246
rect 6972 19236 7028 25340
rect 7084 25284 7140 25454
rect 7084 25218 7140 25228
rect 7196 23940 7252 26236
rect 7308 26226 7364 26236
rect 7308 25732 7364 25742
rect 7308 25618 7364 25676
rect 7308 25566 7310 25618
rect 7362 25566 7364 25618
rect 7308 25554 7364 25566
rect 7644 25508 7700 28366
rect 8204 27188 8260 28700
rect 8316 28530 8372 28542
rect 8316 28478 8318 28530
rect 8370 28478 8372 28530
rect 8316 28308 8372 28478
rect 8428 28530 8484 28700
rect 8652 28642 8708 29374
rect 8652 28590 8654 28642
rect 8706 28590 8708 28642
rect 8652 28578 8708 28590
rect 8428 28478 8430 28530
rect 8482 28478 8484 28530
rect 8428 28466 8484 28478
rect 9100 28532 9156 28542
rect 9100 28438 9156 28476
rect 8316 28242 8372 28252
rect 8764 28418 8820 28430
rect 8764 28366 8766 28418
rect 8818 28366 8820 28418
rect 8652 28084 8708 28094
rect 8652 27858 8708 28028
rect 8652 27806 8654 27858
rect 8706 27806 8708 27858
rect 8652 27794 8708 27806
rect 8204 26908 8260 27132
rect 7756 26852 8260 26908
rect 7756 26514 7812 26852
rect 7756 26462 7758 26514
rect 7810 26462 7812 26514
rect 7756 26450 7812 26462
rect 7868 26516 7924 26526
rect 8428 26516 8484 26526
rect 7868 26514 8372 26516
rect 7868 26462 7870 26514
rect 7922 26462 8372 26514
rect 7868 26460 8372 26462
rect 7868 26450 7924 26460
rect 8316 26402 8372 26460
rect 8428 26422 8484 26460
rect 8316 26350 8318 26402
rect 8370 26350 8372 26402
rect 8316 26338 8372 26350
rect 8540 26402 8596 26414
rect 8540 26350 8542 26402
rect 8594 26350 8596 26402
rect 7980 26292 8036 26302
rect 7644 25442 7700 25452
rect 7868 26290 8036 26292
rect 7868 26238 7982 26290
rect 8034 26238 8036 26290
rect 7868 26236 8036 26238
rect 7420 25396 7476 25406
rect 7420 25302 7476 25340
rect 7756 25284 7812 25294
rect 7756 25190 7812 25228
rect 7196 23874 7252 23884
rect 7868 24836 7924 26236
rect 7980 26226 8036 26236
rect 8540 25732 8596 26350
rect 8540 25666 8596 25676
rect 8652 25508 8708 25518
rect 8428 25394 8484 25406
rect 8428 25342 8430 25394
rect 8482 25342 8484 25394
rect 8092 25284 8148 25294
rect 8092 25190 8148 25228
rect 7084 23826 7140 23838
rect 7084 23774 7086 23826
rect 7138 23774 7140 23826
rect 7084 23716 7140 23774
rect 7756 23828 7812 23838
rect 7868 23828 7924 24780
rect 8204 24946 8260 24958
rect 8204 24894 8206 24946
rect 8258 24894 8260 24946
rect 7756 23826 7924 23828
rect 7756 23774 7758 23826
rect 7810 23774 7924 23826
rect 7756 23772 7924 23774
rect 8092 24498 8148 24510
rect 8092 24446 8094 24498
rect 8146 24446 8148 24498
rect 7756 23762 7812 23772
rect 7420 23716 7476 23726
rect 7084 23714 7476 23716
rect 7084 23662 7422 23714
rect 7474 23662 7476 23714
rect 7084 23660 7476 23662
rect 7084 19458 7140 23660
rect 7420 23650 7476 23660
rect 8092 22596 8148 24446
rect 8204 23938 8260 24894
rect 8316 24724 8372 24734
rect 8316 24630 8372 24668
rect 8428 24276 8484 25342
rect 8652 25394 8708 25452
rect 8652 25342 8654 25394
rect 8706 25342 8708 25394
rect 8540 25284 8596 25294
rect 8540 24722 8596 25228
rect 8540 24670 8542 24722
rect 8594 24670 8596 24722
rect 8540 24658 8596 24670
rect 8428 24220 8596 24276
rect 8204 23886 8206 23938
rect 8258 23886 8260 23938
rect 8204 23874 8260 23886
rect 8316 24052 8372 24062
rect 7532 22540 8148 22596
rect 7420 22372 7476 22382
rect 7420 22278 7476 22316
rect 7532 22258 7588 22540
rect 7532 22206 7534 22258
rect 7586 22206 7588 22258
rect 7532 22036 7588 22206
rect 8092 22370 8148 22382
rect 8092 22318 8094 22370
rect 8146 22318 8148 22370
rect 7420 21980 7588 22036
rect 7756 22146 7812 22158
rect 7756 22094 7758 22146
rect 7810 22094 7812 22146
rect 7420 21812 7476 21980
rect 7420 21746 7476 21756
rect 7532 21698 7588 21710
rect 7532 21646 7534 21698
rect 7586 21646 7588 21698
rect 7532 21588 7588 21646
rect 7756 21700 7812 22094
rect 7756 21634 7812 21644
rect 7532 21522 7588 21532
rect 7868 21586 7924 21598
rect 7868 21534 7870 21586
rect 7922 21534 7924 21586
rect 7868 21364 7924 21534
rect 7868 21298 7924 21308
rect 7084 19406 7086 19458
rect 7138 19406 7140 19458
rect 7084 19394 7140 19406
rect 7420 19796 7476 19806
rect 7420 19458 7476 19740
rect 7420 19406 7422 19458
rect 7474 19406 7476 19458
rect 7420 19394 7476 19406
rect 6860 19234 7028 19236
rect 6860 19182 6862 19234
rect 6914 19182 7028 19234
rect 6860 19180 7028 19182
rect 7644 19234 7700 19246
rect 7644 19182 7646 19234
rect 7698 19182 7700 19234
rect 6860 19170 6916 19180
rect 6636 19012 6692 19022
rect 6636 18564 6692 18956
rect 7644 19012 7700 19182
rect 8092 19236 8148 22318
rect 8204 21588 8260 21598
rect 8204 21494 8260 21532
rect 8204 21364 8260 21374
rect 8316 21364 8372 23996
rect 8428 23828 8484 23838
rect 8428 23734 8484 23772
rect 8540 23714 8596 24220
rect 8540 23662 8542 23714
rect 8594 23662 8596 23714
rect 8540 23650 8596 23662
rect 8652 23938 8708 25342
rect 8764 24722 8820 28366
rect 8988 28420 9044 28430
rect 8988 28326 9044 28364
rect 8988 27188 9044 27198
rect 8988 27094 9044 27132
rect 8876 25396 8932 25406
rect 8876 25302 8932 25340
rect 8988 25394 9044 25406
rect 8988 25342 8990 25394
rect 9042 25342 9044 25394
rect 8764 24670 8766 24722
rect 8818 24670 8820 24722
rect 8764 24658 8820 24670
rect 8876 25172 8932 25182
rect 8652 23886 8654 23938
rect 8706 23886 8708 23938
rect 8652 23268 8708 23886
rect 8652 23174 8708 23212
rect 8764 23268 8820 23278
rect 8876 23268 8932 25116
rect 8988 23940 9044 25342
rect 8988 23846 9044 23884
rect 8764 23266 8932 23268
rect 8764 23214 8766 23266
rect 8818 23214 8932 23266
rect 8764 23212 8932 23214
rect 8764 23202 8820 23212
rect 8652 22932 8708 22942
rect 8652 22930 8932 22932
rect 8652 22878 8654 22930
rect 8706 22878 8932 22930
rect 8652 22876 8932 22878
rect 8652 22866 8708 22876
rect 8764 22258 8820 22270
rect 8764 22206 8766 22258
rect 8818 22206 8820 22258
rect 8540 21812 8596 21822
rect 8428 21700 8484 21710
rect 8428 21606 8484 21644
rect 8260 21308 8372 21364
rect 8204 21298 8260 21308
rect 8540 20914 8596 21756
rect 8652 21812 8708 21822
rect 8764 21812 8820 22206
rect 8652 21810 8820 21812
rect 8652 21758 8654 21810
rect 8706 21758 8820 21810
rect 8652 21756 8820 21758
rect 8652 21746 8708 21756
rect 8876 21586 8932 22876
rect 8876 21534 8878 21586
rect 8930 21534 8932 21586
rect 8876 21522 8932 21534
rect 9212 21028 9268 30156
rect 9324 27860 9380 33068
rect 10444 32564 10500 32574
rect 10444 32562 10612 32564
rect 10444 32510 10446 32562
rect 10498 32510 10612 32562
rect 10444 32508 10612 32510
rect 10444 32498 10500 32508
rect 9660 32452 9716 32462
rect 9548 30100 9604 30110
rect 9548 29314 9604 30044
rect 9548 29262 9550 29314
rect 9602 29262 9604 29314
rect 9548 29250 9604 29262
rect 9660 28644 9716 32396
rect 10556 31780 10612 32508
rect 10556 31686 10612 31724
rect 11116 32450 11172 32462
rect 11116 32398 11118 32450
rect 11170 32398 11172 32450
rect 9884 31668 9940 31678
rect 9884 31574 9940 31612
rect 11116 31668 11172 32398
rect 11564 32452 11620 34750
rect 11564 32386 11620 32396
rect 11116 31602 11172 31612
rect 10780 31106 10836 31118
rect 10780 31054 10782 31106
rect 10834 31054 10836 31106
rect 10780 30996 10836 31054
rect 10780 30930 10836 30940
rect 11116 30996 11172 31006
rect 11564 30996 11620 31006
rect 11116 30994 11620 30996
rect 11116 30942 11118 30994
rect 11170 30942 11566 30994
rect 11618 30942 11620 30994
rect 11116 30940 11620 30942
rect 11116 30930 11172 30940
rect 11564 30884 11620 30940
rect 11340 29988 11396 29998
rect 11564 29988 11620 30828
rect 11340 29986 11620 29988
rect 11340 29934 11342 29986
rect 11394 29934 11620 29986
rect 11340 29932 11620 29934
rect 10780 28756 10836 28766
rect 9660 28084 9716 28588
rect 10556 28700 10780 28756
rect 9660 27990 9716 28028
rect 10332 28196 10388 28206
rect 9324 27794 9380 27804
rect 10332 27858 10388 28140
rect 10332 27806 10334 27858
rect 10386 27806 10388 27858
rect 10332 27794 10388 27806
rect 10556 28082 10612 28700
rect 10780 28690 10836 28700
rect 11004 28532 11060 28542
rect 10780 28418 10836 28430
rect 10780 28366 10782 28418
rect 10834 28366 10836 28418
rect 10780 28196 10836 28366
rect 10780 28130 10836 28140
rect 10556 28030 10558 28082
rect 10610 28030 10612 28082
rect 9324 27186 9380 27198
rect 9324 27134 9326 27186
rect 9378 27134 9380 27186
rect 9324 26908 9380 27134
rect 10556 26908 10612 28030
rect 11004 27858 11060 28476
rect 11340 28196 11396 29932
rect 11676 29540 11732 35084
rect 11900 35138 11956 38108
rect 12012 36482 12068 38332
rect 12460 38164 12516 38612
rect 12460 38070 12516 38108
rect 12236 38052 12292 38062
rect 12012 36430 12014 36482
rect 12066 36430 12068 36482
rect 12012 36260 12068 36430
rect 12012 36194 12068 36204
rect 12124 37996 12236 38052
rect 11900 35086 11902 35138
rect 11954 35086 11956 35138
rect 11900 35074 11956 35086
rect 12124 34804 12180 37996
rect 12236 37958 12292 37996
rect 13692 38052 13748 38062
rect 13692 37958 13748 37996
rect 12572 37938 12628 37950
rect 12572 37886 12574 37938
rect 12626 37886 12628 37938
rect 12572 37156 12628 37886
rect 14140 37266 14196 39342
rect 15372 39396 15428 39406
rect 15372 39060 15428 39340
rect 15372 38994 15428 39004
rect 14364 38836 14420 38846
rect 14252 38724 14308 38734
rect 14252 38630 14308 38668
rect 14140 37214 14142 37266
rect 14194 37214 14196 37266
rect 14140 37202 14196 37214
rect 14364 38050 14420 38780
rect 15820 38668 15876 39452
rect 15932 38836 15988 39566
rect 15932 38770 15988 38780
rect 16380 38722 16436 38734
rect 16380 38670 16382 38722
rect 16434 38670 16436 38722
rect 16380 38668 16436 38670
rect 15820 38612 16436 38668
rect 16492 38388 16548 40126
rect 16492 38322 16548 38332
rect 16604 40180 16660 40460
rect 16716 40180 16772 40190
rect 16604 40178 16772 40180
rect 16604 40126 16718 40178
rect 16770 40126 16772 40178
rect 16604 40124 16772 40126
rect 16604 38276 16660 40124
rect 16716 40114 16772 40124
rect 16828 40178 16884 40190
rect 16828 40126 16830 40178
rect 16882 40126 16884 40178
rect 16828 39956 16884 40126
rect 16716 39900 16884 39956
rect 16716 39730 16772 39900
rect 16716 39678 16718 39730
rect 16770 39678 16772 39730
rect 16716 39666 16772 39678
rect 16940 38836 16996 38846
rect 16828 38834 16996 38836
rect 16828 38782 16942 38834
rect 16994 38782 16996 38834
rect 16828 38780 16996 38782
rect 16828 38500 16884 38780
rect 16940 38770 16996 38780
rect 17164 38668 17220 42140
rect 17836 41860 17892 41870
rect 17836 41188 17892 41804
rect 17836 41122 17892 41132
rect 17948 40964 18004 42476
rect 17948 40898 18004 40908
rect 18060 41412 18116 41422
rect 18060 40514 18116 41356
rect 18060 40462 18062 40514
rect 18114 40462 18116 40514
rect 18060 40450 18116 40462
rect 18172 40404 18228 42700
rect 18508 42532 18564 44828
rect 19404 43764 19460 44942
rect 19516 44212 19572 44222
rect 19516 44118 19572 44156
rect 20076 44100 20132 45276
rect 20524 45218 20580 45230
rect 20524 45166 20526 45218
rect 20578 45166 20580 45218
rect 20300 44322 20356 44334
rect 20300 44270 20302 44322
rect 20354 44270 20356 44322
rect 20300 44212 20356 44270
rect 20300 44146 20356 44156
rect 20076 44044 20244 44100
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 20188 43764 20244 44044
rect 20188 43708 20356 43764
rect 19404 43698 19460 43708
rect 18732 43426 18788 43438
rect 18732 43374 18734 43426
rect 18786 43374 18788 43426
rect 18732 42980 18788 43374
rect 20076 43428 20132 43438
rect 18732 42924 19348 42980
rect 19180 42756 19236 42766
rect 18508 42466 18564 42476
rect 18844 42754 19236 42756
rect 18844 42702 19182 42754
rect 19234 42702 19236 42754
rect 18844 42700 19236 42702
rect 18396 42196 18452 42206
rect 18452 42140 18676 42196
rect 18396 42130 18452 42140
rect 18620 42082 18676 42140
rect 18620 42030 18622 42082
rect 18674 42030 18676 42082
rect 18620 42018 18676 42030
rect 18732 42084 18788 42094
rect 18844 42084 18900 42700
rect 19180 42690 19236 42700
rect 18788 42028 18900 42084
rect 18732 41990 18788 42028
rect 18956 41972 19012 41982
rect 19180 41972 19236 41982
rect 18956 41878 19012 41916
rect 19068 41970 19236 41972
rect 19068 41918 19182 41970
rect 19234 41918 19236 41970
rect 19068 41916 19236 41918
rect 18396 41858 18452 41870
rect 18396 41806 18398 41858
rect 18450 41806 18452 41858
rect 18396 40628 18452 41806
rect 19068 41188 19124 41916
rect 19180 41906 19236 41916
rect 18732 41132 19124 41188
rect 19292 41188 19348 42924
rect 19404 42866 19460 42878
rect 19404 42814 19406 42866
rect 19458 42814 19460 42866
rect 19404 42196 19460 42814
rect 19404 42130 19460 42140
rect 19628 42642 19684 42654
rect 19628 42590 19630 42642
rect 19682 42590 19684 42642
rect 19628 41970 19684 42590
rect 20076 42644 20132 43372
rect 20300 42868 20356 43708
rect 20412 43538 20468 43550
rect 20412 43486 20414 43538
rect 20466 43486 20468 43538
rect 20412 43092 20468 43486
rect 20524 43204 20580 45166
rect 20748 44546 20804 46060
rect 20972 46004 21028 46060
rect 21532 46004 21588 46014
rect 20972 46002 21588 46004
rect 20972 45950 21534 46002
rect 21586 45950 21588 46002
rect 20972 45948 21588 45950
rect 21532 45938 21588 45948
rect 23660 46004 23716 46014
rect 24556 46004 24612 46014
rect 23660 46002 23940 46004
rect 23660 45950 23662 46002
rect 23714 45950 23940 46002
rect 23660 45948 23940 45950
rect 23660 45938 23716 45948
rect 20748 44494 20750 44546
rect 20802 44494 20804 44546
rect 20748 44482 20804 44494
rect 20860 45890 20916 45902
rect 20860 45838 20862 45890
rect 20914 45838 20916 45890
rect 20636 44210 20692 44222
rect 20636 44158 20638 44210
rect 20690 44158 20692 44210
rect 20636 43428 20692 44158
rect 20860 44212 20916 45838
rect 21980 45218 22036 45230
rect 21980 45166 21982 45218
rect 22034 45166 22036 45218
rect 21420 45108 21476 45118
rect 21420 45014 21476 45052
rect 20860 44146 20916 44156
rect 21420 43764 21476 43774
rect 21476 43708 21588 43764
rect 21420 43698 21476 43708
rect 20636 43362 20692 43372
rect 20524 43148 20804 43204
rect 20412 43036 20692 43092
rect 20300 42802 20356 42812
rect 20412 42866 20468 42878
rect 20412 42814 20414 42866
rect 20466 42814 20468 42866
rect 20188 42756 20244 42766
rect 20188 42662 20244 42700
rect 20076 42578 20132 42588
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19628 41918 19630 41970
rect 19682 41918 19684 41970
rect 19628 41906 19684 41918
rect 20412 41524 20468 42814
rect 19852 41468 20468 41524
rect 20524 41636 20580 41646
rect 19852 41412 19908 41468
rect 19852 41318 19908 41356
rect 19516 41188 19572 41198
rect 19292 41132 19516 41188
rect 18396 40572 18676 40628
rect 18172 40402 18452 40404
rect 18172 40350 18174 40402
rect 18226 40350 18452 40402
rect 18172 40348 18452 40350
rect 18172 40338 18228 40348
rect 18284 39508 18340 39518
rect 18172 39396 18228 39406
rect 18172 38946 18228 39340
rect 18172 38894 18174 38946
rect 18226 38894 18228 38946
rect 16828 38434 16884 38444
rect 16940 38612 17220 38668
rect 17836 38724 17892 38762
rect 18172 38668 18228 38894
rect 18284 38946 18340 39452
rect 18396 39284 18452 40348
rect 18396 39218 18452 39228
rect 18508 40402 18564 40414
rect 18508 40350 18510 40402
rect 18562 40350 18564 40402
rect 18284 38894 18286 38946
rect 18338 38894 18340 38946
rect 18284 38882 18340 38894
rect 18396 38834 18452 38846
rect 18396 38782 18398 38834
rect 18450 38782 18452 38834
rect 18396 38668 18452 38782
rect 17836 38658 17892 38668
rect 18060 38612 18228 38668
rect 18284 38612 18452 38668
rect 16716 38276 16772 38286
rect 16604 38220 16716 38276
rect 16716 38210 16772 38220
rect 14364 37998 14366 38050
rect 14418 37998 14420 38050
rect 12684 37156 12740 37166
rect 12572 37154 12740 37156
rect 12572 37102 12686 37154
rect 12738 37102 12740 37154
rect 12572 37100 12740 37102
rect 12572 36260 12628 36270
rect 12572 36166 12628 36204
rect 12236 35140 12292 35150
rect 12684 35140 12740 37100
rect 13916 37156 13972 37166
rect 13916 37062 13972 37100
rect 14140 36484 14196 36494
rect 14364 36484 14420 37998
rect 15148 37940 15204 37950
rect 15148 37846 15204 37884
rect 15148 37380 15204 37390
rect 14924 37378 15204 37380
rect 14924 37326 15150 37378
rect 15202 37326 15204 37378
rect 14924 37324 15204 37326
rect 14812 37266 14868 37278
rect 14812 37214 14814 37266
rect 14866 37214 14868 37266
rect 14476 37156 14532 37166
rect 14812 37156 14868 37214
rect 14476 37154 14868 37156
rect 14476 37102 14478 37154
rect 14530 37102 14868 37154
rect 14476 37100 14868 37102
rect 14476 37090 14532 37100
rect 14924 36594 14980 37324
rect 15148 37314 15204 37324
rect 16492 37268 16548 37278
rect 16828 37268 16884 37278
rect 16492 37266 16828 37268
rect 16492 37214 16494 37266
rect 16546 37214 16828 37266
rect 16492 37212 16828 37214
rect 16492 37202 16548 37212
rect 16828 37174 16884 37212
rect 14924 36542 14926 36594
rect 14978 36542 14980 36594
rect 14924 36530 14980 36542
rect 14140 36482 14420 36484
rect 14140 36430 14142 36482
rect 14194 36430 14420 36482
rect 14140 36428 14420 36430
rect 13804 35700 13860 35710
rect 14140 35700 14196 36428
rect 13804 35698 14196 35700
rect 13804 35646 13806 35698
rect 13858 35646 14196 35698
rect 13804 35644 14196 35646
rect 16604 36260 16660 36270
rect 13804 35634 13860 35644
rect 13020 35586 13076 35598
rect 13020 35534 13022 35586
rect 13074 35534 13076 35586
rect 12236 35138 12740 35140
rect 12236 35086 12238 35138
rect 12290 35086 12740 35138
rect 12236 35084 12740 35086
rect 12908 35140 12964 35150
rect 13020 35140 13076 35534
rect 13580 35364 13636 35374
rect 12908 35138 13076 35140
rect 12908 35086 12910 35138
rect 12962 35086 13076 35138
rect 12908 35084 13076 35086
rect 13468 35252 13524 35262
rect 12236 35074 12292 35084
rect 12908 35074 12964 35084
rect 13468 34914 13524 35196
rect 13468 34862 13470 34914
rect 13522 34862 13524 34914
rect 13468 34850 13524 34862
rect 12124 34738 12180 34748
rect 12460 34804 12516 34814
rect 12460 33796 12516 34748
rect 12796 34804 12852 34814
rect 12796 34710 12852 34748
rect 13244 34356 13300 34366
rect 13244 34262 13300 34300
rect 13580 34354 13636 35308
rect 14028 35364 14084 35374
rect 14028 34914 14084 35308
rect 14028 34862 14030 34914
rect 14082 34862 14084 34914
rect 13804 34804 13860 34814
rect 13804 34710 13860 34748
rect 13580 34302 13582 34354
rect 13634 34302 13636 34354
rect 13580 34290 13636 34302
rect 13692 34690 13748 34702
rect 13692 34638 13694 34690
rect 13746 34638 13748 34690
rect 13692 34356 13748 34638
rect 13916 34692 13972 34702
rect 13916 34598 13972 34636
rect 13692 34290 13748 34300
rect 13468 34244 13524 34254
rect 13468 34150 13524 34188
rect 13020 34130 13076 34142
rect 13020 34078 13022 34130
rect 13074 34078 13076 34130
rect 12684 34020 12740 34030
rect 13020 34020 13076 34078
rect 12684 34018 13076 34020
rect 12684 33966 12686 34018
rect 12738 33966 13076 34018
rect 12684 33964 13076 33966
rect 13356 34020 13412 34030
rect 12684 33908 12740 33964
rect 13356 33926 13412 33964
rect 12684 33842 12740 33852
rect 12460 33730 12516 33740
rect 13580 33460 13636 33470
rect 13580 33366 13636 33404
rect 14028 32788 14084 34862
rect 15148 34914 15204 34926
rect 15148 34862 15150 34914
rect 15202 34862 15204 34914
rect 14700 34692 14756 34702
rect 14756 34636 14868 34692
rect 14700 34598 14756 34636
rect 14364 34356 14420 34366
rect 14140 34244 14196 34254
rect 14140 34150 14196 34188
rect 14028 32722 14084 32732
rect 14140 33460 14196 33470
rect 14140 32674 14196 33404
rect 14140 32622 14142 32674
rect 14194 32622 14196 32674
rect 14140 32610 14196 32622
rect 13916 32564 13972 32574
rect 13244 32452 13300 32462
rect 13300 32396 13524 32452
rect 13244 32358 13300 32396
rect 13356 31892 13412 31902
rect 11788 31668 11844 31678
rect 11788 31574 11844 31612
rect 11900 31668 11956 31678
rect 12124 31668 12180 31678
rect 11900 31666 12124 31668
rect 11900 31614 11902 31666
rect 11954 31614 12124 31666
rect 11900 31612 12124 31614
rect 11900 31602 11956 31612
rect 12124 31602 12180 31612
rect 12124 30996 12180 31006
rect 12124 30212 12180 30940
rect 12572 30884 12628 30894
rect 12572 30790 12628 30828
rect 12460 30324 12516 30334
rect 12124 30146 12180 30156
rect 12348 30268 12460 30324
rect 11340 28130 11396 28140
rect 11564 29484 11732 29540
rect 11004 27806 11006 27858
rect 11058 27806 11060 27858
rect 11004 27794 11060 27806
rect 11452 26962 11508 26974
rect 11452 26910 11454 26962
rect 11506 26910 11508 26962
rect 9324 26852 9940 26908
rect 10556 26852 10836 26908
rect 9884 26404 9940 26852
rect 10556 26516 10612 26526
rect 10556 26422 10612 26460
rect 10108 26404 10164 26414
rect 9884 26402 10052 26404
rect 9884 26350 9886 26402
rect 9938 26350 10052 26402
rect 9884 26348 10052 26350
rect 9884 26338 9940 26348
rect 9772 26290 9828 26302
rect 9772 26238 9774 26290
rect 9826 26238 9828 26290
rect 9772 25396 9828 26238
rect 9548 25394 9828 25396
rect 9548 25342 9774 25394
rect 9826 25342 9828 25394
rect 9548 25340 9828 25342
rect 9324 25284 9380 25294
rect 9324 24500 9380 25228
rect 9436 25172 9492 25182
rect 9548 25172 9604 25340
rect 9772 25330 9828 25340
rect 9884 25284 9940 25294
rect 9884 25190 9940 25228
rect 9492 25116 9604 25172
rect 9772 25172 9828 25182
rect 9436 25106 9492 25116
rect 9772 25060 9828 25116
rect 9772 25004 9940 25060
rect 9884 24836 9940 25004
rect 9884 24770 9940 24780
rect 9996 24834 10052 26348
rect 10108 26402 10276 26404
rect 10108 26350 10110 26402
rect 10162 26350 10276 26402
rect 10108 26348 10276 26350
rect 10108 26338 10164 26348
rect 10220 26290 10276 26348
rect 10220 26238 10222 26290
rect 10274 26238 10276 26290
rect 10220 26226 10276 26238
rect 10668 26290 10724 26302
rect 10668 26238 10670 26290
rect 10722 26238 10724 26290
rect 10444 25508 10500 25518
rect 10332 25394 10388 25406
rect 10332 25342 10334 25394
rect 10386 25342 10388 25394
rect 9996 24782 9998 24834
rect 10050 24782 10052 24834
rect 9996 24724 10052 24782
rect 10108 25282 10164 25294
rect 10108 25230 10110 25282
rect 10162 25230 10164 25282
rect 10108 24724 10164 25230
rect 10332 25172 10388 25342
rect 10444 25394 10500 25452
rect 10668 25506 10724 26238
rect 10780 26292 10836 26852
rect 11452 26516 11508 26910
rect 11564 26908 11620 29484
rect 11676 29316 11732 29326
rect 11676 29222 11732 29260
rect 12012 28868 12068 28878
rect 11676 28756 11732 28766
rect 11676 28662 11732 28700
rect 11788 28642 11844 28654
rect 11788 28590 11790 28642
rect 11842 28590 11844 28642
rect 11788 28308 11844 28590
rect 12012 28642 12068 28812
rect 12012 28590 12014 28642
rect 12066 28590 12068 28642
rect 12012 28578 12068 28590
rect 12348 28642 12404 30268
rect 12460 30258 12516 30268
rect 12908 29986 12964 29998
rect 12908 29934 12910 29986
rect 12962 29934 12964 29986
rect 12908 29876 12964 29934
rect 12796 29540 12852 29550
rect 12684 29538 12852 29540
rect 12684 29486 12798 29538
rect 12850 29486 12852 29538
rect 12684 29484 12852 29486
rect 12348 28590 12350 28642
rect 12402 28590 12404 28642
rect 12348 28578 12404 28590
rect 12460 29428 12516 29438
rect 11676 28252 11844 28308
rect 12460 28532 12516 29372
rect 12684 28868 12740 29484
rect 12796 29474 12852 29484
rect 12684 28642 12740 28812
rect 12796 29316 12852 29326
rect 12796 28754 12852 29260
rect 12796 28702 12798 28754
rect 12850 28702 12852 28754
rect 12796 28690 12852 28702
rect 12684 28590 12686 28642
rect 12738 28590 12740 28642
rect 12684 28578 12740 28590
rect 11676 27970 11732 28252
rect 11676 27918 11678 27970
rect 11730 27918 11732 27970
rect 11676 27906 11732 27918
rect 12236 27074 12292 27086
rect 12236 27022 12238 27074
rect 12290 27022 12292 27074
rect 12236 26964 12292 27022
rect 12460 26964 12516 28476
rect 12236 26908 12516 26964
rect 12908 26908 12964 29820
rect 13020 29988 13076 29998
rect 13020 28642 13076 29932
rect 13132 29426 13188 29438
rect 13132 29374 13134 29426
rect 13186 29374 13188 29426
rect 13132 28756 13188 29374
rect 13132 28690 13188 28700
rect 13020 28590 13022 28642
rect 13074 28590 13076 28642
rect 13020 28578 13076 28590
rect 11564 26852 11732 26908
rect 11452 26450 11508 26460
rect 10780 26290 10948 26292
rect 10780 26238 10782 26290
rect 10834 26238 10948 26290
rect 10780 26236 10948 26238
rect 10780 26226 10836 26236
rect 10668 25454 10670 25506
rect 10722 25454 10724 25506
rect 10668 25442 10724 25454
rect 10444 25342 10446 25394
rect 10498 25342 10500 25394
rect 10444 25330 10500 25342
rect 10332 25106 10388 25116
rect 10220 24948 10276 24958
rect 10220 24946 10724 24948
rect 10220 24894 10222 24946
rect 10274 24894 10724 24946
rect 10220 24892 10724 24894
rect 10220 24882 10276 24892
rect 10332 24724 10388 24734
rect 10108 24722 10388 24724
rect 10108 24670 10334 24722
rect 10386 24670 10388 24722
rect 10108 24668 10388 24670
rect 9996 24658 10052 24668
rect 10332 24658 10388 24668
rect 10668 24722 10724 24892
rect 10668 24670 10670 24722
rect 10722 24670 10724 24722
rect 10668 24658 10724 24670
rect 10892 24836 10948 26236
rect 11116 25394 11172 25406
rect 11116 25342 11118 25394
rect 11170 25342 11172 25394
rect 11116 25172 11172 25342
rect 11228 25284 11284 25294
rect 11228 25190 11284 25228
rect 11452 25284 11508 25294
rect 11452 25282 11620 25284
rect 11452 25230 11454 25282
rect 11506 25230 11620 25282
rect 11452 25228 11620 25230
rect 11452 25218 11508 25228
rect 11116 25106 11172 25116
rect 11340 24836 11396 24846
rect 10892 24834 11396 24836
rect 10892 24782 11342 24834
rect 11394 24782 11396 24834
rect 10892 24780 11396 24782
rect 10892 24722 10948 24780
rect 11340 24770 11396 24780
rect 11564 24834 11620 25228
rect 11564 24782 11566 24834
rect 11618 24782 11620 24834
rect 11564 24770 11620 24782
rect 10892 24670 10894 24722
rect 10946 24670 10948 24722
rect 10892 24658 10948 24670
rect 10556 24610 10612 24622
rect 10556 24558 10558 24610
rect 10610 24558 10612 24610
rect 9324 24444 10052 24500
rect 9996 24050 10052 24444
rect 9996 23998 9998 24050
rect 10050 23998 10052 24050
rect 9996 23986 10052 23998
rect 10556 24052 10612 24558
rect 10556 23986 10612 23996
rect 10892 23268 10948 23278
rect 10892 22482 10948 23212
rect 10892 22430 10894 22482
rect 10946 22430 10948 22482
rect 10892 22418 10948 22430
rect 10780 21588 10836 21598
rect 10780 21494 10836 21532
rect 9660 21474 9716 21486
rect 9660 21422 9662 21474
rect 9714 21422 9716 21474
rect 9660 21364 9716 21422
rect 11452 21476 11508 21486
rect 11452 21382 11508 21420
rect 9660 21298 9716 21308
rect 10780 21028 10836 21038
rect 9212 20972 9380 21028
rect 8540 20862 8542 20914
rect 8594 20862 8596 20914
rect 8540 20850 8596 20862
rect 9212 20692 9268 20702
rect 9100 20690 9268 20692
rect 9100 20638 9214 20690
rect 9266 20638 9268 20690
rect 9100 20636 9268 20638
rect 8988 20578 9044 20590
rect 8988 20526 8990 20578
rect 9042 20526 9044 20578
rect 8204 20018 8260 20030
rect 8204 19966 8206 20018
rect 8258 19966 8260 20018
rect 8204 19908 8260 19966
rect 8204 19842 8260 19852
rect 8876 19906 8932 19918
rect 8876 19854 8878 19906
rect 8930 19854 8932 19906
rect 8764 19796 8820 19806
rect 8764 19702 8820 19740
rect 8316 19236 8372 19246
rect 8092 19234 8372 19236
rect 8092 19182 8318 19234
rect 8370 19182 8372 19234
rect 8092 19180 8372 19182
rect 7644 18946 7700 18956
rect 8204 19012 8260 19022
rect 6636 18508 7028 18564
rect 6972 18340 7028 18508
rect 6860 17444 6916 17454
rect 6860 16994 6916 17388
rect 6860 16942 6862 16994
rect 6914 16942 6916 16994
rect 6860 16930 6916 16942
rect 6972 17442 7028 18284
rect 8204 18338 8260 18956
rect 8316 18452 8372 19180
rect 8876 19012 8932 19854
rect 8988 19908 9044 20526
rect 8988 19842 9044 19852
rect 8988 19348 9044 19358
rect 9100 19348 9156 20636
rect 9212 20626 9268 20636
rect 8988 19346 9156 19348
rect 8988 19294 8990 19346
rect 9042 19294 9156 19346
rect 8988 19292 9156 19294
rect 8988 19282 9044 19292
rect 9324 19124 9380 20972
rect 9660 20916 9716 20926
rect 9548 20914 9716 20916
rect 9548 20862 9662 20914
rect 9714 20862 9716 20914
rect 9548 20860 9716 20862
rect 9548 20690 9604 20860
rect 9660 20850 9716 20860
rect 9548 20638 9550 20690
rect 9602 20638 9604 20690
rect 9548 20626 9604 20638
rect 9996 20690 10052 20702
rect 9996 20638 9998 20690
rect 10050 20638 10052 20690
rect 9772 20580 9828 20590
rect 9772 20486 9828 20524
rect 9884 20244 9940 20254
rect 9996 20244 10052 20638
rect 10444 20580 10500 20590
rect 10444 20486 10500 20524
rect 9884 20242 10052 20244
rect 9884 20190 9886 20242
rect 9938 20190 10052 20242
rect 9884 20188 10052 20190
rect 9884 20178 9940 20188
rect 9772 20132 9828 20142
rect 9772 20038 9828 20076
rect 10780 20132 10836 20972
rect 11452 20916 11508 20926
rect 11676 20916 11732 26852
rect 12236 26292 12292 26908
rect 12908 26852 13076 26908
rect 12236 26226 12292 26236
rect 12908 26292 12964 26302
rect 12908 26198 12964 26236
rect 11788 25396 11844 25406
rect 11788 24946 11844 25340
rect 11788 24894 11790 24946
rect 11842 24894 11844 24946
rect 11788 24882 11844 24894
rect 12236 25060 12292 25070
rect 12236 24834 12292 25004
rect 12236 24782 12238 24834
rect 12290 24782 12292 24834
rect 12236 24770 12292 24782
rect 12348 24836 12404 24846
rect 12348 24834 12516 24836
rect 12348 24782 12350 24834
rect 12402 24782 12516 24834
rect 12348 24780 12516 24782
rect 12348 24770 12404 24780
rect 12012 24722 12068 24734
rect 12012 24670 12014 24722
rect 12066 24670 12068 24722
rect 12012 24500 12068 24670
rect 12348 24500 12404 24510
rect 12012 24498 12404 24500
rect 12012 24446 12350 24498
rect 12402 24446 12404 24498
rect 12012 24444 12404 24446
rect 12348 24434 12404 24444
rect 12124 24052 12180 24062
rect 12124 23958 12180 23996
rect 12460 23940 12516 24780
rect 12460 23156 12516 23884
rect 12460 23090 12516 23100
rect 12796 23938 12852 23950
rect 12796 23886 12798 23938
rect 12850 23886 12852 23938
rect 11452 20914 11732 20916
rect 11452 20862 11454 20914
rect 11506 20862 11732 20914
rect 11452 20860 11732 20862
rect 12796 21588 12852 23886
rect 10780 20066 10836 20076
rect 11004 20802 11060 20814
rect 11004 20750 11006 20802
rect 11058 20750 11060 20802
rect 9996 20020 10052 20030
rect 9996 19926 10052 19964
rect 10444 20018 10500 20030
rect 10444 19966 10446 20018
rect 10498 19966 10500 20018
rect 10444 19796 10500 19966
rect 11004 20020 11060 20750
rect 10444 19730 10500 19740
rect 10892 19908 10948 19918
rect 8876 18946 8932 18956
rect 8988 19068 9380 19124
rect 10556 19684 10612 19694
rect 8316 18386 8372 18396
rect 8204 18286 8206 18338
rect 8258 18286 8260 18338
rect 8204 18274 8260 18286
rect 8652 18340 8708 18350
rect 8652 18246 8708 18284
rect 6972 17390 6974 17442
rect 7026 17390 7028 17442
rect 6412 16100 6468 16110
rect 6412 16006 6468 16044
rect 6188 15986 6356 15988
rect 6188 15934 6190 15986
rect 6242 15934 6356 15986
rect 6188 15932 6356 15934
rect 6188 15922 6244 15932
rect 6076 15262 6078 15314
rect 6130 15262 6132 15314
rect 6076 15204 6132 15262
rect 6300 15148 6356 15932
rect 6076 14642 6132 15148
rect 6076 14590 6078 14642
rect 6130 14590 6132 14642
rect 6076 14578 6132 14590
rect 6188 15092 6356 15148
rect 6412 15316 6468 15326
rect 6412 15148 6468 15260
rect 6860 15316 6916 15326
rect 6860 15222 6916 15260
rect 6412 15092 6580 15148
rect 5012 14476 5236 14532
rect 4956 14466 5012 14476
rect 4844 14366 4846 14418
rect 4898 14366 4900 14418
rect 4844 14354 4900 14366
rect 4508 14306 4564 14318
rect 4508 14254 4510 14306
rect 4562 14254 4564 14306
rect 4508 13524 4564 14254
rect 4620 14306 4676 14318
rect 4620 14254 4622 14306
rect 4674 14254 4676 14306
rect 4620 13748 4676 14254
rect 4956 13748 5012 13758
rect 4620 13746 5012 13748
rect 4620 13694 4958 13746
rect 5010 13694 5012 13746
rect 4620 13692 5012 13694
rect 4620 13634 4676 13692
rect 4956 13682 5012 13692
rect 5180 13746 5236 14476
rect 5180 13694 5182 13746
rect 5234 13694 5236 13746
rect 5180 13682 5236 13694
rect 4620 13582 4622 13634
rect 4674 13582 4676 13634
rect 4620 13570 4676 13582
rect 4060 13468 4564 13524
rect 5516 13522 5572 13534
rect 5516 13470 5518 13522
rect 5570 13470 5572 13522
rect 3724 13188 3780 13198
rect 3724 13094 3780 13132
rect 4060 13186 4116 13468
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 5516 13300 5572 13470
rect 4476 13290 4740 13300
rect 4060 13134 4062 13186
rect 4114 13134 4116 13186
rect 4060 13122 4116 13134
rect 5068 13244 5572 13300
rect 4732 12908 5012 12964
rect 3836 12852 3892 12862
rect 3836 12758 3892 12796
rect 4284 12852 4340 12862
rect 3612 11618 3780 11620
rect 3612 11566 3614 11618
rect 3666 11566 3780 11618
rect 3612 11564 3780 11566
rect 3612 11554 3668 11564
rect 2492 11442 2548 11452
rect 3388 11396 3444 11406
rect 3388 11394 3668 11396
rect 3388 11342 3390 11394
rect 3442 11342 3668 11394
rect 3388 11340 3668 11342
rect 3388 11330 3444 11340
rect 1708 10500 1764 10510
rect 1708 10406 1764 10444
rect 3612 10500 3668 11340
rect 3500 10388 3556 10398
rect 3500 9938 3556 10332
rect 3500 9886 3502 9938
rect 3554 9886 3556 9938
rect 3500 9874 3556 9886
rect 3388 9828 3444 9866
rect 3388 9762 3444 9772
rect 3612 9826 3668 10444
rect 3612 9774 3614 9826
rect 3666 9774 3668 9826
rect 3612 9762 3668 9774
rect 3724 9828 3780 11564
rect 4284 11394 4340 12796
rect 4732 12852 4788 12908
rect 4732 12758 4788 12796
rect 4844 12740 4900 12750
rect 4620 12068 4676 12078
rect 4620 11974 4676 12012
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4396 11508 4452 11518
rect 4396 11414 4452 11452
rect 4284 11342 4286 11394
rect 4338 11342 4340 11394
rect 4284 11330 4340 11342
rect 4620 11396 4676 11406
rect 4620 11302 4676 11340
rect 4844 11394 4900 12684
rect 4956 12178 5012 12908
rect 4956 12126 4958 12178
rect 5010 12126 5012 12178
rect 4956 12114 5012 12126
rect 5068 12850 5124 13244
rect 5068 12798 5070 12850
rect 5122 12798 5124 12850
rect 5068 11844 5124 12798
rect 5292 12964 5348 12974
rect 5292 12402 5348 12908
rect 5628 12852 5684 12862
rect 5628 12758 5684 12796
rect 5740 12740 5796 12750
rect 5740 12646 5796 12684
rect 5852 12738 5908 12750
rect 5852 12686 5854 12738
rect 5906 12686 5908 12738
rect 5852 12404 5908 12686
rect 5292 12350 5294 12402
rect 5346 12350 5348 12402
rect 5292 12338 5348 12350
rect 5404 12348 5908 12404
rect 5404 12290 5460 12348
rect 5404 12238 5406 12290
rect 5458 12238 5460 12290
rect 5404 12226 5460 12238
rect 5068 11778 5124 11788
rect 5516 12068 5572 12348
rect 5628 12180 5684 12190
rect 5628 12178 6020 12180
rect 5628 12126 5630 12178
rect 5682 12126 6020 12178
rect 5628 12124 6020 12126
rect 5628 12114 5684 12124
rect 4844 11342 4846 11394
rect 4898 11342 4900 11394
rect 4844 11330 4900 11342
rect 5516 11396 5572 12012
rect 5628 11396 5684 11406
rect 5572 11394 5684 11396
rect 5572 11342 5630 11394
rect 5682 11342 5684 11394
rect 5572 11340 5684 11342
rect 5516 11302 5572 11340
rect 5628 11330 5684 11340
rect 5852 11394 5908 12124
rect 5964 12066 6020 12124
rect 5964 12014 5966 12066
rect 6018 12014 6020 12066
rect 5964 12002 6020 12014
rect 5852 11342 5854 11394
rect 5906 11342 5908 11394
rect 5852 11330 5908 11342
rect 5964 11844 6020 11854
rect 5964 11394 6020 11788
rect 5964 11342 5966 11394
rect 6018 11342 6020 11394
rect 5964 11330 6020 11342
rect 3948 11170 4004 11182
rect 6188 11172 6244 15092
rect 6524 13970 6580 15092
rect 6524 13918 6526 13970
rect 6578 13918 6580 13970
rect 6524 13906 6580 13918
rect 6972 13748 7028 17390
rect 8876 17666 8932 17678
rect 8876 17614 8878 17666
rect 8930 17614 8932 17666
rect 8876 16324 8932 17614
rect 8988 17220 9044 19068
rect 9884 18452 9940 18462
rect 9884 17666 9940 18396
rect 10556 18340 10612 19628
rect 10668 18452 10724 18462
rect 10668 18450 10836 18452
rect 10668 18398 10670 18450
rect 10722 18398 10836 18450
rect 10668 18396 10836 18398
rect 10668 18386 10724 18396
rect 9884 17614 9886 17666
rect 9938 17614 9940 17666
rect 9884 17602 9940 17614
rect 10444 18284 10612 18340
rect 9212 17554 9268 17566
rect 9212 17502 9214 17554
rect 9266 17502 9268 17554
rect 9100 17444 9156 17454
rect 9100 17350 9156 17388
rect 9212 17332 9268 17502
rect 9212 17276 9716 17332
rect 8988 17164 9380 17220
rect 9212 16884 9268 16894
rect 8876 16258 8932 16268
rect 8988 16828 9212 16884
rect 8988 16770 9044 16828
rect 9212 16818 9268 16828
rect 8988 16718 8990 16770
rect 9042 16718 9044 16770
rect 8988 16210 9044 16718
rect 8988 16158 8990 16210
rect 9042 16158 9044 16210
rect 8988 16146 9044 16158
rect 9212 16212 9268 16222
rect 9212 16118 9268 16156
rect 9212 15540 9268 15550
rect 8988 15484 9212 15540
rect 7308 15204 7364 15214
rect 7084 13748 7140 13758
rect 6972 13692 7084 13748
rect 7084 13654 7140 13692
rect 6860 13524 6916 13534
rect 6860 13522 7028 13524
rect 6860 13470 6862 13522
rect 6914 13470 7028 13522
rect 6860 13468 7028 13470
rect 6860 13458 6916 13468
rect 6300 12962 6356 12974
rect 6300 12910 6302 12962
rect 6354 12910 6356 12962
rect 6300 12404 6356 12910
rect 6300 12338 6356 12348
rect 6748 12962 6804 12974
rect 6748 12910 6750 12962
rect 6802 12910 6804 12962
rect 6748 11732 6804 12910
rect 6860 12964 6916 12974
rect 6860 12870 6916 12908
rect 6412 11676 6804 11732
rect 6972 12292 7028 13468
rect 7084 13076 7140 13086
rect 7084 12982 7140 13020
rect 7308 12964 7364 15148
rect 8988 15202 9044 15484
rect 9212 15474 9268 15484
rect 8988 15150 8990 15202
rect 9042 15150 9044 15202
rect 8988 15138 9044 15150
rect 9324 15148 9380 17164
rect 9660 17106 9716 17276
rect 9660 17054 9662 17106
rect 9714 17054 9716 17106
rect 9660 17042 9716 17054
rect 9548 16884 9604 16894
rect 9772 16884 9828 16894
rect 9548 16882 9716 16884
rect 9548 16830 9550 16882
rect 9602 16830 9716 16882
rect 9548 16828 9716 16830
rect 9548 16818 9604 16828
rect 9548 16324 9604 16334
rect 9548 15538 9604 16268
rect 9660 16212 9716 16828
rect 9772 16790 9828 16828
rect 10220 16884 10276 16894
rect 10108 16324 10164 16334
rect 10108 16230 10164 16268
rect 9660 16146 9716 16156
rect 9884 16098 9940 16110
rect 9884 16046 9886 16098
rect 9938 16046 9940 16098
rect 9548 15486 9550 15538
rect 9602 15486 9604 15538
rect 9548 15474 9604 15486
rect 9772 15540 9828 15550
rect 9884 15540 9940 16046
rect 9828 15484 9940 15540
rect 9772 15446 9828 15484
rect 10220 15314 10276 16828
rect 10444 16100 10500 18284
rect 10668 18228 10724 18238
rect 10556 18226 10724 18228
rect 10556 18174 10670 18226
rect 10722 18174 10724 18226
rect 10556 18172 10724 18174
rect 10556 17778 10612 18172
rect 10668 18162 10724 18172
rect 10556 17726 10558 17778
rect 10610 17726 10612 17778
rect 10556 17714 10612 17726
rect 10780 16212 10836 18396
rect 10892 18004 10948 19852
rect 11004 19348 11060 19964
rect 11452 19796 11508 20860
rect 12124 20132 12180 20142
rect 11452 19730 11508 19740
rect 12012 19796 12068 19806
rect 11116 19348 11172 19358
rect 11004 19346 11172 19348
rect 11004 19294 11118 19346
rect 11170 19294 11172 19346
rect 11004 19292 11172 19294
rect 11116 19282 11172 19292
rect 11452 18452 11508 18462
rect 11452 18358 11508 18396
rect 11004 18228 11060 18238
rect 11004 18226 11284 18228
rect 11004 18174 11006 18226
rect 11058 18174 11284 18226
rect 11004 18172 11284 18174
rect 11004 18162 11060 18172
rect 10892 17948 11172 18004
rect 11116 16212 11172 17948
rect 11228 16772 11284 18172
rect 12012 17892 12068 19740
rect 12124 18450 12180 20076
rect 12796 20130 12852 21532
rect 12796 20078 12798 20130
rect 12850 20078 12852 20130
rect 12124 18398 12126 18450
rect 12178 18398 12180 18450
rect 12124 18386 12180 18398
rect 12348 18452 12404 18462
rect 12012 17836 12180 17892
rect 12012 17668 12068 17678
rect 12012 17106 12068 17612
rect 12012 17054 12014 17106
rect 12066 17054 12068 17106
rect 12012 17042 12068 17054
rect 11900 16996 11956 17006
rect 11788 16940 11900 16996
rect 11228 16706 11284 16716
rect 11340 16884 11396 16894
rect 10780 16146 10836 16156
rect 10892 16210 11172 16212
rect 10892 16158 11118 16210
rect 11170 16158 11172 16210
rect 10892 16156 11172 16158
rect 10444 16044 10724 16100
rect 10668 15988 10724 16044
rect 10668 15932 10836 15988
rect 10444 15876 10500 15886
rect 10444 15874 10724 15876
rect 10444 15822 10446 15874
rect 10498 15822 10724 15874
rect 10444 15820 10724 15822
rect 10444 15810 10500 15820
rect 10668 15540 10724 15820
rect 10668 15446 10724 15484
rect 10220 15262 10222 15314
rect 10274 15262 10276 15314
rect 10220 15250 10276 15262
rect 10556 15316 10612 15326
rect 9660 15204 9716 15242
rect 9324 15092 9492 15148
rect 9660 15138 9716 15148
rect 10444 15204 10500 15242
rect 10556 15222 10612 15260
rect 10444 15138 10500 15148
rect 7532 13748 7588 13758
rect 7532 13654 7588 13692
rect 9100 13636 9156 13646
rect 7756 13076 7812 13086
rect 7756 12982 7812 13020
rect 9100 13074 9156 13580
rect 9100 13022 9102 13074
rect 9154 13022 9156 13074
rect 9100 13010 9156 13022
rect 7196 12850 7252 12862
rect 7196 12798 7198 12850
rect 7250 12798 7252 12850
rect 7196 12740 7252 12798
rect 7196 12674 7252 12684
rect 6412 11618 6468 11676
rect 6412 11566 6414 11618
rect 6466 11566 6468 11618
rect 6412 11554 6468 11566
rect 3948 11118 3950 11170
rect 4002 11118 4004 11170
rect 3948 10612 4004 11118
rect 5964 11116 6244 11172
rect 5180 10722 5236 10734
rect 5180 10670 5182 10722
rect 5234 10670 5236 10722
rect 3836 10500 3892 10510
rect 3836 10406 3892 10444
rect 3724 9762 3780 9772
rect 3500 8818 3556 8830
rect 3500 8766 3502 8818
rect 3554 8766 3556 8818
rect 3500 8428 3556 8766
rect 3836 8820 3892 8830
rect 3948 8820 4004 10556
rect 4620 10612 4676 10622
rect 5180 10612 5236 10670
rect 4620 10610 4900 10612
rect 4620 10558 4622 10610
rect 4674 10558 4900 10610
rect 4620 10556 4900 10558
rect 4620 10546 4676 10556
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4396 10052 4452 10062
rect 4396 9940 4452 9996
rect 4060 9938 4452 9940
rect 4060 9886 4398 9938
rect 4450 9886 4452 9938
rect 4060 9884 4452 9886
rect 4060 9826 4116 9884
rect 4396 9874 4452 9884
rect 4844 9940 4900 10556
rect 5180 10546 5236 10556
rect 5068 10500 5124 10510
rect 5068 10406 5124 10444
rect 4956 10388 5012 10398
rect 4956 10294 5012 10332
rect 4844 9874 4900 9884
rect 5068 10052 5124 10062
rect 4060 9774 4062 9826
rect 4114 9774 4116 9826
rect 4060 9762 4116 9774
rect 3836 8818 4004 8820
rect 3836 8766 3838 8818
rect 3890 8766 4004 8818
rect 3836 8764 4004 8766
rect 4060 8930 4116 8942
rect 4060 8878 4062 8930
rect 4114 8878 4116 8930
rect 3836 8708 3892 8764
rect 3388 8372 3556 8428
rect 3612 8652 3892 8708
rect 1820 8260 1876 8270
rect 1820 6690 1876 8204
rect 2492 8148 2548 8158
rect 2492 8146 2884 8148
rect 2492 8094 2494 8146
rect 2546 8094 2884 8146
rect 2492 8092 2884 8094
rect 2492 8082 2548 8092
rect 2828 7362 2884 8092
rect 2940 7586 2996 7598
rect 2940 7534 2942 7586
rect 2994 7534 2996 7586
rect 2940 7476 2996 7534
rect 2940 7410 2996 7420
rect 3388 7476 3444 8372
rect 3500 7700 3556 7710
rect 3612 7700 3668 8652
rect 4060 8428 4116 8878
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 3500 7698 3668 7700
rect 3500 7646 3502 7698
rect 3554 7646 3668 7698
rect 3500 7644 3668 7646
rect 3724 8372 4676 8428
rect 3724 7698 3780 8372
rect 4620 8370 4676 8372
rect 4620 8318 4622 8370
rect 4674 8318 4676 8370
rect 4620 8306 4676 8318
rect 5068 8034 5124 9996
rect 5964 10052 6020 11116
rect 6524 10836 6580 11676
rect 5964 9986 6020 9996
rect 6076 10834 6580 10836
rect 6076 10782 6526 10834
rect 6578 10782 6580 10834
rect 6076 10780 6580 10782
rect 5628 9940 5684 9950
rect 5628 9826 5684 9884
rect 5628 9774 5630 9826
rect 5682 9774 5684 9826
rect 5628 8428 5684 9774
rect 6076 9268 6132 10780
rect 6524 10770 6580 10780
rect 6748 10610 6804 10622
rect 6748 10558 6750 10610
rect 6802 10558 6804 10610
rect 6636 10498 6692 10510
rect 6636 10446 6638 10498
rect 6690 10446 6692 10498
rect 6412 9716 6468 9726
rect 6076 9154 6132 9212
rect 6300 9714 6468 9716
rect 6300 9662 6414 9714
rect 6466 9662 6468 9714
rect 6300 9660 6468 9662
rect 6300 9266 6356 9660
rect 6412 9650 6468 9660
rect 6300 9214 6302 9266
rect 6354 9214 6356 9266
rect 6300 9202 6356 9214
rect 6076 9102 6078 9154
rect 6130 9102 6132 9154
rect 6076 9090 6132 9102
rect 6412 9156 6468 9166
rect 6412 9062 6468 9100
rect 6636 9154 6692 10446
rect 6748 9940 6804 10558
rect 6748 9874 6804 9884
rect 6636 9102 6638 9154
rect 6690 9102 6692 9154
rect 6636 9090 6692 9102
rect 6972 9042 7028 12236
rect 7308 11394 7364 12908
rect 8316 12964 8372 12974
rect 8316 12870 8372 12908
rect 8764 12964 8820 12974
rect 8092 12740 8148 12750
rect 8092 12290 8148 12684
rect 8092 12238 8094 12290
rect 8146 12238 8148 12290
rect 8092 12226 8148 12238
rect 8764 12178 8820 12908
rect 8764 12126 8766 12178
rect 8818 12126 8820 12178
rect 8764 12114 8820 12126
rect 7308 11342 7310 11394
rect 7362 11342 7364 11394
rect 7308 11330 7364 11342
rect 8092 11284 8148 11294
rect 8092 11190 8148 11228
rect 7196 10612 7252 10622
rect 7196 10518 7252 10556
rect 9436 10500 9492 15092
rect 10220 13748 10276 13758
rect 10108 13746 10276 13748
rect 10108 13694 10222 13746
rect 10274 13694 10276 13746
rect 10108 13692 10276 13694
rect 9884 12404 9940 12414
rect 9884 12310 9940 12348
rect 9548 12292 9604 12302
rect 9548 11172 9604 12236
rect 9884 11620 9940 11630
rect 9548 11106 9604 11116
rect 9660 11284 9716 11294
rect 9660 10834 9716 11228
rect 9660 10782 9662 10834
rect 9714 10782 9716 10834
rect 9660 10770 9716 10782
rect 9548 10724 9604 10734
rect 9548 10630 9604 10668
rect 9884 10722 9940 11564
rect 10108 11508 10164 13692
rect 10220 13682 10276 13692
rect 10332 13524 10388 13534
rect 10332 13522 10500 13524
rect 10332 13470 10334 13522
rect 10386 13470 10500 13522
rect 10332 13468 10500 13470
rect 10332 13458 10388 13468
rect 10332 12404 10388 12414
rect 10332 12178 10388 12348
rect 10332 12126 10334 12178
rect 10386 12126 10388 12178
rect 10332 12114 10388 12126
rect 10444 11620 10500 13468
rect 10444 11554 10500 11564
rect 10780 12178 10836 15932
rect 10892 14532 10948 16156
rect 11116 16146 11172 16156
rect 11340 15538 11396 16828
rect 11788 16882 11844 16940
rect 11900 16930 11956 16940
rect 11788 16830 11790 16882
rect 11842 16830 11844 16882
rect 11788 16818 11844 16830
rect 11900 16772 11956 16782
rect 11900 16678 11956 16716
rect 11788 16324 11844 16334
rect 11788 16098 11844 16268
rect 11788 16046 11790 16098
rect 11842 16046 11844 16098
rect 11788 16034 11844 16046
rect 12012 16100 12068 16110
rect 12012 15986 12068 16044
rect 12012 15934 12014 15986
rect 12066 15934 12068 15986
rect 12012 15922 12068 15934
rect 11340 15486 11342 15538
rect 11394 15486 11396 15538
rect 10892 14530 11172 14532
rect 10892 14478 10894 14530
rect 10946 14478 11172 14530
rect 10892 14476 11172 14478
rect 10892 14466 10948 14476
rect 10892 14306 10948 14318
rect 10892 14254 10894 14306
rect 10946 14254 10948 14306
rect 10892 13970 10948 14254
rect 10892 13918 10894 13970
rect 10946 13918 10948 13970
rect 10892 13906 10948 13918
rect 11116 12852 11172 14476
rect 11340 14306 11396 15486
rect 11788 15540 11844 15550
rect 11340 14254 11342 14306
rect 11394 14254 11396 14306
rect 11340 14242 11396 14254
rect 11564 15314 11620 15326
rect 11564 15262 11566 15314
rect 11618 15262 11620 15314
rect 11564 14530 11620 15262
rect 11564 14478 11566 14530
rect 11618 14478 11620 14530
rect 11228 13746 11284 13758
rect 11228 13694 11230 13746
rect 11282 13694 11284 13746
rect 11228 13300 11284 13694
rect 11228 13234 11284 13244
rect 11228 13076 11284 13086
rect 11564 13076 11620 14478
rect 11676 15202 11732 15214
rect 11676 15150 11678 15202
rect 11730 15150 11732 15202
rect 11676 13860 11732 15150
rect 11788 14754 11844 15484
rect 12124 15148 12180 17836
rect 12348 16882 12404 18396
rect 12796 18452 12852 20078
rect 13020 19684 13076 26852
rect 13356 24724 13412 31836
rect 13468 31778 13524 32396
rect 13468 31726 13470 31778
rect 13522 31726 13524 31778
rect 13468 31714 13524 31726
rect 13580 31780 13636 31790
rect 13580 29428 13636 31724
rect 13916 31778 13972 32508
rect 14364 32562 14420 34300
rect 14476 34018 14532 34030
rect 14476 33966 14478 34018
rect 14530 33966 14532 34018
rect 14476 32786 14532 33966
rect 14700 34020 14756 34030
rect 14588 33906 14644 33918
rect 14588 33854 14590 33906
rect 14642 33854 14644 33906
rect 14588 33572 14644 33854
rect 14588 33506 14644 33516
rect 14476 32734 14478 32786
rect 14530 32734 14532 32786
rect 14476 32722 14532 32734
rect 14588 32788 14644 32798
rect 14700 32788 14756 33964
rect 14812 33908 14868 34636
rect 15036 34020 15092 34030
rect 15036 33926 15092 33964
rect 14812 33842 14868 33852
rect 15148 33460 15204 34862
rect 15820 34804 15876 34814
rect 15820 34802 16436 34804
rect 15820 34750 15822 34802
rect 15874 34750 16436 34802
rect 15820 34748 16436 34750
rect 15820 34738 15876 34748
rect 16380 34354 16436 34748
rect 16380 34302 16382 34354
rect 16434 34302 16436 34354
rect 16380 34290 16436 34302
rect 16492 34692 16548 34702
rect 16492 34242 16548 34636
rect 16492 34190 16494 34242
rect 16546 34190 16548 34242
rect 16492 34178 16548 34190
rect 15820 34018 15876 34030
rect 15820 33966 15822 34018
rect 15874 33966 15876 34018
rect 15148 33394 15204 33404
rect 15708 33572 15764 33582
rect 15708 33458 15764 33516
rect 15708 33406 15710 33458
rect 15762 33406 15764 33458
rect 15708 33394 15764 33406
rect 14588 32786 14756 32788
rect 14588 32734 14590 32786
rect 14642 32734 14756 32786
rect 14588 32732 14756 32734
rect 14812 32788 14868 32798
rect 14588 32722 14644 32732
rect 14364 32510 14366 32562
rect 14418 32510 14420 32562
rect 13916 31726 13918 31778
rect 13970 31726 13972 31778
rect 13916 31714 13972 31726
rect 14140 31778 14196 31790
rect 14140 31726 14142 31778
rect 14194 31726 14196 31778
rect 13804 31668 13860 31678
rect 13804 31574 13860 31612
rect 13692 31554 13748 31566
rect 13692 31502 13694 31554
rect 13746 31502 13748 31554
rect 13692 31108 13748 31502
rect 13692 31042 13748 31052
rect 14140 30884 14196 31726
rect 14364 31108 14420 32510
rect 14812 32562 14868 32732
rect 15148 32788 15204 32798
rect 15148 32694 15204 32732
rect 15372 32564 15428 32574
rect 15820 32564 15876 33966
rect 14812 32510 14814 32562
rect 14866 32510 14868 32562
rect 14812 32498 14868 32510
rect 15260 32562 15876 32564
rect 15260 32510 15374 32562
rect 15426 32510 15876 32562
rect 15260 32508 15876 32510
rect 16156 33796 16212 33806
rect 14588 31780 14644 31790
rect 14588 31686 14644 31724
rect 14364 31042 14420 31052
rect 14924 31108 14980 31118
rect 14924 31014 14980 31052
rect 14140 30790 14196 30828
rect 14588 30884 14644 30894
rect 14588 30790 14644 30828
rect 15148 30884 15204 30894
rect 15260 30884 15316 32508
rect 15372 32498 15428 32508
rect 16044 32450 16100 32462
rect 16044 32398 16046 32450
rect 16098 32398 16100 32450
rect 15372 32340 15428 32350
rect 15372 31890 15428 32284
rect 15372 31838 15374 31890
rect 15426 31838 15428 31890
rect 15372 31826 15428 31838
rect 15204 30828 15316 30884
rect 15484 30994 15540 31006
rect 15484 30942 15486 30994
rect 15538 30942 15540 30994
rect 15484 30884 15540 30942
rect 15596 30884 15652 30894
rect 15484 30828 15596 30884
rect 13804 30324 13860 30334
rect 13804 30230 13860 30268
rect 14924 30098 14980 30110
rect 14924 30046 14926 30098
rect 14978 30046 14980 30098
rect 13692 29988 13748 29998
rect 13692 29894 13748 29932
rect 13916 29986 13972 29998
rect 13916 29934 13918 29986
rect 13970 29934 13972 29986
rect 13580 29334 13636 29372
rect 13916 28980 13972 29934
rect 14140 29986 14196 29998
rect 14140 29934 14142 29986
rect 14194 29934 14196 29986
rect 14140 29876 14196 29934
rect 14588 29988 14644 29998
rect 14644 29932 14868 29988
rect 14588 29894 14644 29932
rect 14140 29810 14196 29820
rect 14252 29316 14308 29326
rect 14252 29222 14308 29260
rect 13692 28924 13972 28980
rect 13580 28868 13636 28878
rect 13692 28868 13748 28924
rect 13636 28812 13748 28868
rect 13580 26964 13636 28812
rect 13804 28756 13860 28766
rect 13580 26898 13636 26908
rect 13692 28084 13748 28094
rect 13692 26402 13748 28028
rect 13804 27860 13860 28700
rect 14812 27972 14868 29932
rect 14924 29316 14980 30046
rect 14924 29250 14980 29260
rect 14924 28644 14980 28654
rect 14924 28550 14980 28588
rect 14700 27970 14868 27972
rect 14700 27918 14814 27970
rect 14866 27918 14868 27970
rect 14700 27916 14868 27918
rect 14588 27860 14644 27870
rect 13804 27858 14644 27860
rect 13804 27806 14590 27858
rect 14642 27806 14644 27858
rect 13804 27804 14644 27806
rect 13804 27746 13860 27804
rect 14588 27794 14644 27804
rect 13804 27694 13806 27746
rect 13858 27694 13860 27746
rect 13804 27682 13860 27694
rect 14364 27636 14420 27646
rect 14364 27186 14420 27580
rect 14700 27188 14756 27916
rect 14812 27906 14868 27916
rect 14924 27972 14980 27982
rect 14924 27878 14980 27916
rect 15148 27412 15204 30828
rect 15596 30818 15652 30828
rect 16044 30884 16100 32398
rect 16156 31220 16212 33740
rect 16380 33460 16436 33470
rect 16380 33346 16436 33404
rect 16380 33294 16382 33346
rect 16434 33294 16436 33346
rect 16380 33282 16436 33294
rect 16380 32452 16436 32462
rect 16604 32452 16660 36204
rect 16940 32676 16996 38612
rect 17276 38162 17332 38174
rect 17276 38110 17278 38162
rect 17330 38110 17332 38162
rect 17276 37940 17332 38110
rect 17724 37940 17780 37950
rect 17276 37938 17780 37940
rect 17276 37886 17726 37938
rect 17778 37886 17780 37938
rect 17276 37884 17780 37886
rect 17500 37266 17556 37278
rect 17500 37214 17502 37266
rect 17554 37214 17556 37266
rect 17052 36594 17108 36606
rect 17052 36542 17054 36594
rect 17106 36542 17108 36594
rect 17052 36484 17108 36542
rect 17500 36484 17556 37214
rect 17724 36932 17780 37884
rect 18060 37828 18116 38612
rect 18060 37734 18116 37772
rect 17836 37492 17892 37502
rect 17836 37398 17892 37436
rect 18284 37268 18340 38612
rect 18396 37938 18452 37950
rect 18396 37886 18398 37938
rect 18450 37886 18452 37938
rect 18396 37828 18452 37886
rect 18396 37762 18452 37772
rect 18396 37268 18452 37278
rect 18284 37212 18396 37268
rect 18396 37202 18452 37212
rect 18172 37156 18228 37166
rect 18172 37062 18228 37100
rect 17836 36932 17892 36942
rect 17724 36876 17836 36932
rect 17836 36866 17892 36876
rect 18508 36706 18564 40350
rect 18620 39844 18676 40572
rect 18732 40626 18788 41132
rect 19516 41094 19572 41132
rect 19964 41076 20020 41086
rect 19628 41074 20020 41076
rect 19628 41022 19966 41074
rect 20018 41022 20020 41074
rect 19628 41020 20020 41022
rect 19068 40964 19124 40974
rect 18732 40574 18734 40626
rect 18786 40574 18788 40626
rect 18732 40562 18788 40574
rect 18956 40626 19012 40638
rect 18956 40574 18958 40626
rect 19010 40574 19012 40626
rect 18732 39844 18788 39854
rect 18620 39788 18732 39844
rect 18732 39778 18788 39788
rect 18844 39730 18900 39742
rect 18844 39678 18846 39730
rect 18898 39678 18900 39730
rect 18844 39620 18900 39678
rect 18844 39554 18900 39564
rect 18620 39508 18676 39518
rect 18620 38050 18676 39452
rect 18844 39284 18900 39294
rect 18844 38948 18900 39228
rect 18956 39172 19012 40574
rect 19068 39842 19124 40908
rect 19628 40628 19684 41020
rect 19964 41010 20020 41020
rect 20524 41074 20580 41580
rect 20636 41300 20692 43036
rect 20748 41858 20804 43148
rect 21308 42868 21364 42878
rect 21308 42774 21364 42812
rect 21084 41972 21140 41982
rect 21084 41878 21140 41916
rect 20748 41806 20750 41858
rect 20802 41806 20804 41858
rect 20748 41794 20804 41806
rect 20636 41234 20692 41244
rect 21420 41188 21476 41198
rect 21420 41094 21476 41132
rect 20524 41022 20526 41074
rect 20578 41022 20580 41074
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 20524 40740 20580 41022
rect 20748 41076 20804 41086
rect 20748 41074 21364 41076
rect 20748 41022 20750 41074
rect 20802 41022 21364 41074
rect 20748 41020 21364 41022
rect 20748 41010 20804 41020
rect 20524 40674 20580 40684
rect 20636 40962 20692 40974
rect 20636 40910 20638 40962
rect 20690 40910 20692 40962
rect 20188 40628 20244 40638
rect 19628 40572 19796 40628
rect 19068 39790 19070 39842
rect 19122 39790 19124 39842
rect 19068 39778 19124 39790
rect 19516 39844 19572 39854
rect 19516 39618 19572 39788
rect 19516 39566 19518 39618
rect 19570 39566 19572 39618
rect 19516 39554 19572 39566
rect 19740 39620 19796 40572
rect 20636 40628 20692 40910
rect 20636 40572 21252 40628
rect 20188 40516 20244 40572
rect 20188 40514 20916 40516
rect 20188 40462 20190 40514
rect 20242 40462 20916 40514
rect 20188 40460 20916 40462
rect 20188 40450 20244 40460
rect 20076 40402 20132 40414
rect 20076 40350 20078 40402
rect 20130 40350 20132 40402
rect 20076 39844 20132 40350
rect 20748 40292 20804 40302
rect 20076 39788 20356 39844
rect 19740 39554 19796 39564
rect 20076 39620 20132 39630
rect 19628 39508 19684 39518
rect 19628 39414 19684 39452
rect 19852 39506 19908 39518
rect 19852 39454 19854 39506
rect 19906 39454 19908 39506
rect 19852 39396 19908 39454
rect 20076 39396 20132 39564
rect 20076 39340 20244 39396
rect 19852 39330 19908 39340
rect 19836 39228 20100 39238
rect 18956 39106 19012 39116
rect 19516 39172 19572 39182
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 18844 38892 19012 38948
rect 18844 38612 18900 38622
rect 18844 38518 18900 38556
rect 18620 37998 18622 38050
rect 18674 37998 18676 38050
rect 18620 37492 18676 37998
rect 18844 38052 18900 38062
rect 18844 37958 18900 37996
rect 18620 37266 18676 37436
rect 18620 37214 18622 37266
rect 18674 37214 18676 37266
rect 18620 37202 18676 37214
rect 18508 36654 18510 36706
rect 18562 36654 18564 36706
rect 18508 36642 18564 36654
rect 18844 36932 18900 36942
rect 18172 36594 18228 36606
rect 18172 36542 18174 36594
rect 18226 36542 18228 36594
rect 18060 36484 18116 36494
rect 17052 36482 18116 36484
rect 17052 36430 18062 36482
rect 18114 36430 18116 36482
rect 17052 36428 18116 36430
rect 18060 36418 18116 36428
rect 17836 36260 17892 36270
rect 17724 35588 17780 35598
rect 17724 35494 17780 35532
rect 16940 32610 16996 32620
rect 17276 35364 17332 35374
rect 16828 32564 16884 32574
rect 16828 32470 16884 32508
rect 16380 32450 16660 32452
rect 16380 32398 16382 32450
rect 16434 32398 16660 32450
rect 16380 32396 16660 32398
rect 16268 31220 16324 31230
rect 16156 31164 16268 31220
rect 16268 31126 16324 31164
rect 16044 30818 16100 30828
rect 16380 30100 16436 32396
rect 17276 31668 17332 35308
rect 17836 34244 17892 36204
rect 18172 35922 18228 36542
rect 18844 36482 18900 36876
rect 18844 36430 18846 36482
rect 18898 36430 18900 36482
rect 18844 36418 18900 36430
rect 18172 35870 18174 35922
rect 18226 35870 18228 35922
rect 18172 35858 18228 35870
rect 18060 35586 18116 35598
rect 18060 35534 18062 35586
rect 18114 35534 18116 35586
rect 17948 35028 18004 35038
rect 18060 35028 18116 35534
rect 18732 35586 18788 35598
rect 18732 35534 18734 35586
rect 18786 35534 18788 35586
rect 18396 35028 18452 35038
rect 17948 35026 18340 35028
rect 17948 34974 17950 35026
rect 18002 34974 18340 35026
rect 17948 34972 18340 34974
rect 17948 34962 18004 34972
rect 18284 34914 18340 34972
rect 18284 34862 18286 34914
rect 18338 34862 18340 34914
rect 18284 34850 18340 34862
rect 18396 34356 18452 34972
rect 18060 34354 18452 34356
rect 18060 34302 18398 34354
rect 18450 34302 18452 34354
rect 18060 34300 18452 34302
rect 17948 34244 18004 34254
rect 17836 34242 18004 34244
rect 17836 34190 17950 34242
rect 18002 34190 18004 34242
rect 17836 34188 18004 34190
rect 17724 33908 17780 33918
rect 17612 33852 17724 33908
rect 17500 33460 17556 33470
rect 17500 33346 17556 33404
rect 17500 33294 17502 33346
rect 17554 33294 17556 33346
rect 17500 33282 17556 33294
rect 17500 32452 17556 32462
rect 17612 32452 17668 33852
rect 17724 33842 17780 33852
rect 17836 32900 17892 34188
rect 17948 34178 18004 34188
rect 17500 32450 17668 32452
rect 17500 32398 17502 32450
rect 17554 32398 17668 32450
rect 17500 32396 17668 32398
rect 17724 32844 17892 32900
rect 18060 34020 18116 34300
rect 18396 34290 18452 34300
rect 18508 34690 18564 34702
rect 18508 34638 18510 34690
rect 18562 34638 18564 34690
rect 17500 32386 17556 32396
rect 17388 32340 17444 32350
rect 17388 32246 17444 32284
rect 17724 32228 17780 32844
rect 17500 32172 17780 32228
rect 17836 32676 17892 32686
rect 17892 32620 18004 32676
rect 17500 31890 17556 32172
rect 17500 31838 17502 31890
rect 17554 31838 17556 31890
rect 17500 31826 17556 31838
rect 17836 31890 17892 32620
rect 17948 32562 18004 32620
rect 17948 32510 17950 32562
rect 18002 32510 18004 32562
rect 17948 32498 18004 32510
rect 17836 31838 17838 31890
rect 17890 31838 17892 31890
rect 17836 31826 17892 31838
rect 18060 31668 18116 33964
rect 18172 34132 18228 34142
rect 18172 32786 18228 34076
rect 18508 34132 18564 34638
rect 18620 34692 18676 34702
rect 18620 34598 18676 34636
rect 18732 34690 18788 35534
rect 18732 34638 18734 34690
rect 18786 34638 18788 34690
rect 18508 34066 18564 34076
rect 18620 34130 18676 34142
rect 18620 34078 18622 34130
rect 18674 34078 18676 34130
rect 18284 34018 18340 34030
rect 18284 33966 18286 34018
rect 18338 33966 18340 34018
rect 18284 33908 18340 33966
rect 18284 33842 18340 33852
rect 18508 33796 18564 33806
rect 18396 33740 18508 33796
rect 18284 33236 18340 33246
rect 18396 33236 18452 33740
rect 18508 33730 18564 33740
rect 18620 33796 18676 34078
rect 18732 34132 18788 34638
rect 18732 34066 18788 34076
rect 18844 34690 18900 34702
rect 18844 34638 18846 34690
rect 18898 34638 18900 34690
rect 18844 33796 18900 34638
rect 18956 34242 19012 38892
rect 19404 38500 19460 38510
rect 19292 38444 19404 38500
rect 19292 38276 19348 38444
rect 19404 38434 19460 38444
rect 19068 38220 19348 38276
rect 19404 38276 19460 38286
rect 19068 38050 19124 38220
rect 19404 38182 19460 38220
rect 19068 37998 19070 38050
rect 19122 37998 19124 38050
rect 19068 37986 19124 37998
rect 19292 37940 19348 37950
rect 19292 37846 19348 37884
rect 19404 37492 19460 37502
rect 19516 37492 19572 39116
rect 19852 39060 19908 39070
rect 19852 38834 19908 39004
rect 19852 38782 19854 38834
rect 19906 38782 19908 38834
rect 19852 38770 19908 38782
rect 20076 38946 20132 38958
rect 20076 38894 20078 38946
rect 20130 38894 20132 38946
rect 20076 38836 20132 38894
rect 20076 38770 20132 38780
rect 19964 38722 20020 38734
rect 19964 38670 19966 38722
rect 20018 38670 20020 38722
rect 19628 38612 19684 38622
rect 19628 38274 19684 38556
rect 19628 38222 19630 38274
rect 19682 38222 19684 38274
rect 19628 38210 19684 38222
rect 19740 38052 19796 38062
rect 19740 37958 19796 37996
rect 19404 37490 19572 37492
rect 19404 37438 19406 37490
rect 19458 37438 19572 37490
rect 19404 37436 19572 37438
rect 19628 37828 19684 37838
rect 19964 37828 20020 38670
rect 20188 38668 20244 39340
rect 20300 39172 20356 39788
rect 20748 39506 20804 40236
rect 20748 39454 20750 39506
rect 20802 39454 20804 39506
rect 20748 39442 20804 39454
rect 20412 39396 20468 39406
rect 20412 39394 20692 39396
rect 20412 39342 20414 39394
rect 20466 39342 20692 39394
rect 20412 39340 20692 39342
rect 20412 39330 20468 39340
rect 20300 39116 20580 39172
rect 20524 38834 20580 39116
rect 20524 38782 20526 38834
rect 20578 38782 20580 38834
rect 20076 38612 20132 38622
rect 20188 38612 20468 38668
rect 20076 38276 20132 38556
rect 20300 38388 20356 38398
rect 20188 38276 20244 38286
rect 20076 38274 20244 38276
rect 20076 38222 20190 38274
rect 20242 38222 20244 38274
rect 20076 38220 20244 38222
rect 20188 38210 20244 38220
rect 20300 38162 20356 38332
rect 20300 38110 20302 38162
rect 20354 38110 20356 38162
rect 20300 38098 20356 38110
rect 20412 37938 20468 38612
rect 20412 37886 20414 37938
rect 20466 37886 20468 37938
rect 20412 37874 20468 37886
rect 19964 37772 20244 37828
rect 19628 37490 19684 37772
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20188 37492 20244 37772
rect 19628 37438 19630 37490
rect 19682 37438 19684 37490
rect 19404 37426 19460 37436
rect 19628 37426 19684 37438
rect 20076 37436 20244 37492
rect 19068 37268 19124 37278
rect 19068 37174 19124 37212
rect 19740 37266 19796 37278
rect 19740 37214 19742 37266
rect 19794 37214 19796 37266
rect 19740 36708 19796 37214
rect 20076 37156 20132 37436
rect 20076 37062 20132 37100
rect 19852 36708 19908 36718
rect 19292 36706 19908 36708
rect 19292 36654 19854 36706
rect 19906 36654 19908 36706
rect 19292 36652 19908 36654
rect 19180 36484 19236 36494
rect 19180 35586 19236 36428
rect 19292 36482 19348 36652
rect 19852 36642 19908 36652
rect 19292 36430 19294 36482
rect 19346 36430 19348 36482
rect 19292 36418 19348 36430
rect 20524 36484 20580 38782
rect 20636 38668 20692 39340
rect 20860 38722 20916 40460
rect 21196 40402 21252 40572
rect 21196 40350 21198 40402
rect 21250 40350 21252 40402
rect 21196 40338 21252 40350
rect 21196 40180 21252 40190
rect 20860 38670 20862 38722
rect 20914 38670 20916 38722
rect 20636 38612 20804 38668
rect 20860 38658 20916 38670
rect 20972 40124 21196 40180
rect 20524 36390 20580 36428
rect 19964 36370 20020 36382
rect 19964 36318 19966 36370
rect 20018 36318 20020 36370
rect 19964 36260 20020 36318
rect 19964 36194 20020 36204
rect 20636 36258 20692 36270
rect 20636 36206 20638 36258
rect 20690 36206 20692 36258
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19180 35534 19182 35586
rect 19234 35534 19236 35586
rect 19180 35522 19236 35534
rect 20300 35588 20356 35598
rect 20636 35588 20692 36206
rect 20356 35532 20692 35588
rect 19964 35028 20020 35038
rect 19964 34934 20020 34972
rect 20300 35028 20356 35532
rect 20748 35252 20804 38612
rect 20860 36484 20916 36494
rect 20860 36390 20916 36428
rect 20748 35186 20804 35196
rect 20300 34934 20356 34972
rect 19404 34802 19460 34814
rect 19404 34750 19406 34802
rect 19458 34750 19460 34802
rect 19292 34692 19348 34702
rect 18956 34190 18958 34242
rect 19010 34190 19012 34242
rect 18956 33908 19012 34190
rect 18956 33842 19012 33852
rect 19068 34690 19348 34692
rect 19068 34638 19294 34690
rect 19346 34638 19348 34690
rect 19068 34636 19348 34638
rect 18620 33740 18900 33796
rect 19068 33796 19124 34636
rect 19292 34626 19348 34636
rect 19292 34356 19348 34366
rect 19404 34356 19460 34750
rect 20860 34692 20916 34702
rect 20860 34598 20916 34636
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19292 34354 19460 34356
rect 19292 34302 19294 34354
rect 19346 34302 19460 34354
rect 19292 34300 19460 34302
rect 19292 34290 19348 34300
rect 18284 33234 18452 33236
rect 18284 33182 18286 33234
rect 18338 33182 18452 33234
rect 18284 33180 18452 33182
rect 18284 33170 18340 33180
rect 18172 32734 18174 32786
rect 18226 32734 18228 32786
rect 18172 32722 18228 32734
rect 18396 32564 18452 32574
rect 18452 32508 18564 32564
rect 18396 32470 18452 32508
rect 17276 31612 17556 31668
rect 16828 31220 16884 31230
rect 16380 30034 16436 30044
rect 16604 30884 16660 30894
rect 16716 30884 16772 30894
rect 16660 30882 16772 30884
rect 16660 30830 16718 30882
rect 16770 30830 16772 30882
rect 16660 30828 16772 30830
rect 16044 29428 16100 29438
rect 15820 28084 15876 28094
rect 15820 27990 15876 28028
rect 15932 27972 15988 27982
rect 15708 27858 15764 27870
rect 15932 27860 15988 27916
rect 15708 27806 15710 27858
rect 15762 27806 15764 27858
rect 15372 27636 15428 27646
rect 15708 27636 15764 27806
rect 15148 27346 15204 27356
rect 15260 27634 15764 27636
rect 15260 27582 15374 27634
rect 15426 27582 15764 27634
rect 15260 27580 15764 27582
rect 15820 27804 15988 27860
rect 14364 27134 14366 27186
rect 14418 27134 14420 27186
rect 14364 27122 14420 27134
rect 14476 27132 14756 27188
rect 14252 26964 14308 26974
rect 14476 26964 14532 27132
rect 14812 27076 14868 27086
rect 15148 27076 15204 27086
rect 14812 27074 15148 27076
rect 14812 27022 14814 27074
rect 14866 27022 15148 27074
rect 14812 27020 15148 27022
rect 14812 27010 14868 27020
rect 15148 27010 15204 27020
rect 14252 26962 14532 26964
rect 14252 26910 14254 26962
rect 14306 26910 14532 26962
rect 14252 26908 14532 26910
rect 14588 26964 14644 27002
rect 14252 26898 14308 26908
rect 14588 26898 14644 26908
rect 13692 26350 13694 26402
rect 13746 26350 13748 26402
rect 13692 26338 13748 26350
rect 13468 26292 13524 26302
rect 13468 25506 13524 26236
rect 13468 25454 13470 25506
rect 13522 25454 13524 25506
rect 13468 25442 13524 25454
rect 14252 25396 14308 25406
rect 14252 25302 14308 25340
rect 13356 24658 13412 24668
rect 13580 23940 13636 23950
rect 13580 23846 13636 23884
rect 14252 23828 14308 23838
rect 13692 23826 14308 23828
rect 13692 23774 14254 23826
rect 14306 23774 14308 23826
rect 13692 23772 14308 23774
rect 13580 23380 13636 23390
rect 13692 23380 13748 23772
rect 14252 23762 14308 23772
rect 13580 23378 13748 23380
rect 13580 23326 13582 23378
rect 13634 23326 13748 23378
rect 13580 23324 13748 23326
rect 14364 23492 14420 23502
rect 14364 23378 14420 23436
rect 14364 23326 14366 23378
rect 14418 23326 14420 23378
rect 13580 23314 13636 23324
rect 14364 23314 14420 23326
rect 14588 23380 14644 23390
rect 14588 23286 14644 23324
rect 15260 23380 15316 27580
rect 15372 27570 15428 27580
rect 15820 27076 15876 27804
rect 15932 27636 15988 27646
rect 15932 27542 15988 27580
rect 15820 26178 15876 27020
rect 16044 27074 16100 29372
rect 16380 29316 16436 29326
rect 16380 29222 16436 29260
rect 16156 27748 16212 27758
rect 16156 27654 16212 27692
rect 16044 27022 16046 27074
rect 16098 27022 16100 27074
rect 16044 27010 16100 27022
rect 16604 26908 16660 30828
rect 16716 30818 16772 30828
rect 16828 29650 16884 31164
rect 16828 29598 16830 29650
rect 16882 29598 16884 29650
rect 16828 29540 16884 29598
rect 16828 29474 16884 29484
rect 17388 30994 17444 31006
rect 17388 30942 17390 30994
rect 17442 30942 17444 30994
rect 17388 29428 17444 30942
rect 17500 29652 17556 31612
rect 17836 31612 18116 31668
rect 18284 32450 18340 32462
rect 18284 32398 18286 32450
rect 18338 32398 18340 32450
rect 17724 29652 17780 29662
rect 17500 29650 17780 29652
rect 17500 29598 17726 29650
rect 17778 29598 17780 29650
rect 17500 29596 17780 29598
rect 17724 29586 17780 29596
rect 17388 28754 17444 29372
rect 17724 29426 17780 29438
rect 17724 29374 17726 29426
rect 17778 29374 17780 29426
rect 17388 28702 17390 28754
rect 17442 28702 17444 28754
rect 17388 28690 17444 28702
rect 17500 29314 17556 29326
rect 17500 29262 17502 29314
rect 17554 29262 17556 29314
rect 17500 27972 17556 29262
rect 17724 29316 17780 29374
rect 17724 29250 17780 29260
rect 17500 27906 17556 27916
rect 16828 27748 16884 27758
rect 16716 27636 16772 27646
rect 16716 27186 16772 27580
rect 16716 27134 16718 27186
rect 16770 27134 16772 27186
rect 16716 27122 16772 27134
rect 15820 26126 15822 26178
rect 15874 26126 15876 26178
rect 15820 26114 15876 26126
rect 16156 26852 16660 26908
rect 16828 26908 16884 27692
rect 17500 27748 17556 27758
rect 17500 27654 17556 27692
rect 17388 27636 17444 27646
rect 17388 27542 17444 27580
rect 16828 26852 17332 26908
rect 16156 24948 16212 26852
rect 16268 26628 16324 26638
rect 16268 26514 16324 26572
rect 16268 26462 16270 26514
rect 16322 26462 16324 26514
rect 16268 26450 16324 26462
rect 16604 26516 16660 26526
rect 16604 26422 16660 26460
rect 16380 26404 16436 26414
rect 16380 26310 16436 26348
rect 16828 26292 16884 26302
rect 16828 26198 16884 26236
rect 16492 26178 16548 26190
rect 16492 26126 16494 26178
rect 16546 26126 16548 26178
rect 16380 25844 16436 25854
rect 16380 25618 16436 25788
rect 16380 25566 16382 25618
rect 16434 25566 16436 25618
rect 16380 25554 16436 25566
rect 16492 25508 16548 26126
rect 16492 25452 16772 25508
rect 16380 24948 16436 24958
rect 15932 24892 16380 24948
rect 13468 23268 13524 23278
rect 13468 23174 13524 23212
rect 14140 23266 14196 23278
rect 14924 23268 14980 23278
rect 14140 23214 14142 23266
rect 14194 23214 14196 23266
rect 13692 22932 13748 22942
rect 13692 22838 13748 22876
rect 14028 21698 14084 21710
rect 14028 21646 14030 21698
rect 14082 21646 14084 21698
rect 13580 21474 13636 21486
rect 13580 21422 13582 21474
rect 13634 21422 13636 21474
rect 13580 20916 13636 21422
rect 13916 21476 13972 21486
rect 13916 21382 13972 21420
rect 13580 20850 13636 20860
rect 14028 20804 14084 21646
rect 14028 20738 14084 20748
rect 14140 21140 14196 23214
rect 14700 23212 14924 23268
rect 14476 23042 14532 23054
rect 14476 22990 14478 23042
rect 14530 22990 14532 23042
rect 14476 22932 14532 22990
rect 14476 22866 14532 22876
rect 14476 22372 14532 22382
rect 14700 22372 14756 23212
rect 14924 23174 14980 23212
rect 15260 23154 15316 23324
rect 15260 23102 15262 23154
rect 15314 23102 15316 23154
rect 15260 23090 15316 23102
rect 15484 23492 15540 23502
rect 15484 23042 15540 23436
rect 15932 23154 15988 24892
rect 16380 24854 16436 24892
rect 16716 24834 16772 25452
rect 16716 24782 16718 24834
rect 16770 24782 16772 24834
rect 16716 24770 16772 24782
rect 16828 24612 16884 24622
rect 16828 24518 16884 24556
rect 16380 24050 16436 24062
rect 16380 23998 16382 24050
rect 16434 23998 16436 24050
rect 15932 23102 15934 23154
rect 15986 23102 15988 23154
rect 15932 23090 15988 23102
rect 16156 23266 16212 23278
rect 16156 23214 16158 23266
rect 16210 23214 16212 23266
rect 15484 22990 15486 23042
rect 15538 22990 15540 23042
rect 15484 22820 15540 22990
rect 15484 22754 15540 22764
rect 15708 22484 15764 22494
rect 15708 22390 15764 22428
rect 14476 22370 14868 22372
rect 14476 22318 14478 22370
rect 14530 22318 14868 22370
rect 14476 22316 14868 22318
rect 14476 22306 14532 22316
rect 14588 22146 14644 22158
rect 14588 22094 14590 22146
rect 14642 22094 14644 22146
rect 14588 21812 14644 22094
rect 14252 21756 14644 21812
rect 14700 22146 14756 22158
rect 14700 22094 14702 22146
rect 14754 22094 14756 22146
rect 14252 21698 14308 21756
rect 14252 21646 14254 21698
rect 14306 21646 14308 21698
rect 14252 21634 14308 21646
rect 14700 21588 14756 22094
rect 14140 20802 14196 21084
rect 14588 21532 14756 21588
rect 14812 21586 14868 22316
rect 14812 21534 14814 21586
rect 14866 21534 14868 21586
rect 14588 21474 14644 21532
rect 14812 21522 14868 21534
rect 14924 22146 14980 22158
rect 14924 22094 14926 22146
rect 14978 22094 14980 22146
rect 14588 21422 14590 21474
rect 14642 21422 14644 21474
rect 14588 20916 14644 21422
rect 14588 20850 14644 20860
rect 14700 21364 14756 21374
rect 14700 20914 14756 21308
rect 14812 21140 14868 21150
rect 14924 21140 14980 22094
rect 15820 21588 15876 21598
rect 15820 21586 16100 21588
rect 15820 21534 15822 21586
rect 15874 21534 16100 21586
rect 15820 21532 16100 21534
rect 15820 21522 15876 21532
rect 15596 21474 15652 21486
rect 15596 21422 15598 21474
rect 15650 21422 15652 21474
rect 15148 21364 15204 21374
rect 14868 21084 14980 21140
rect 15036 21362 15204 21364
rect 15036 21310 15150 21362
rect 15202 21310 15204 21362
rect 15036 21308 15204 21310
rect 14812 21074 14868 21084
rect 14700 20862 14702 20914
rect 14754 20862 14756 20914
rect 14700 20850 14756 20862
rect 14140 20750 14142 20802
rect 14194 20750 14196 20802
rect 14140 19684 14196 20750
rect 14812 20804 14868 20814
rect 15036 20804 15092 21308
rect 15148 21298 15204 21308
rect 15484 21364 15540 21374
rect 15484 21270 15540 21308
rect 14868 20748 15092 20804
rect 15148 20804 15204 20814
rect 14812 20710 14868 20748
rect 15148 20710 15204 20748
rect 15260 20690 15316 20702
rect 15260 20638 15262 20690
rect 15314 20638 15316 20690
rect 13020 19618 13076 19628
rect 13916 19628 14196 19684
rect 14588 20578 14644 20590
rect 14588 20526 14590 20578
rect 14642 20526 14644 20578
rect 14588 20244 14644 20526
rect 13468 19348 13524 19358
rect 12796 18386 12852 18396
rect 13132 19346 13524 19348
rect 13132 19294 13470 19346
rect 13522 19294 13524 19346
rect 13132 19292 13524 19294
rect 12684 17778 12740 17790
rect 12684 17726 12686 17778
rect 12738 17726 12740 17778
rect 12684 17668 12740 17726
rect 13020 17668 13076 17678
rect 12684 17612 12964 17668
rect 12348 16830 12350 16882
rect 12402 16830 12404 16882
rect 12348 16818 12404 16830
rect 12908 16996 12964 17612
rect 12572 16324 12628 16334
rect 12348 16212 12404 16222
rect 12348 16118 12404 16156
rect 11788 14702 11790 14754
rect 11842 14702 11844 14754
rect 11788 14690 11844 14702
rect 12012 15092 12180 15148
rect 12012 14196 12068 15092
rect 12572 14644 12628 16268
rect 12908 16210 12964 16940
rect 12908 16158 12910 16210
rect 12962 16158 12964 16210
rect 12908 16146 12964 16158
rect 12684 16098 12740 16110
rect 12684 16046 12686 16098
rect 12738 16046 12740 16098
rect 12684 15988 12740 16046
rect 13020 15988 13076 17612
rect 13132 16994 13188 19292
rect 13468 19282 13524 19292
rect 13804 19124 13860 19134
rect 13804 19030 13860 19068
rect 13580 19012 13636 19022
rect 13580 18918 13636 18956
rect 13132 16942 13134 16994
rect 13186 16942 13188 16994
rect 13132 16930 13188 16942
rect 13916 16884 13972 19628
rect 14364 19012 14420 19022
rect 14364 18918 14420 18956
rect 14252 18340 14308 18350
rect 14588 18340 14644 20188
rect 15260 19234 15316 20638
rect 15596 20132 15652 21422
rect 16044 20356 16100 21532
rect 16156 21476 16212 23214
rect 16380 22820 16436 23998
rect 16828 23940 16884 23950
rect 16828 23846 16884 23884
rect 16380 22754 16436 22764
rect 16828 23268 16884 23278
rect 16828 23042 16884 23212
rect 16828 22990 16830 23042
rect 16882 22990 16884 23042
rect 16268 22484 16324 22494
rect 16828 22484 16884 22990
rect 16268 22482 16884 22484
rect 16268 22430 16270 22482
rect 16322 22430 16884 22482
rect 16268 22428 16884 22430
rect 17276 22596 17332 26852
rect 17612 26404 17668 26414
rect 17836 26404 17892 31612
rect 18284 31108 18340 32398
rect 18508 31444 18564 32508
rect 18620 32562 18676 33740
rect 19068 33730 19124 33740
rect 19180 34130 19236 34142
rect 19180 34078 19182 34130
rect 19234 34078 19236 34130
rect 19180 34020 19236 34078
rect 19180 33236 19236 33964
rect 19404 34130 19460 34142
rect 19404 34078 19406 34130
rect 19458 34078 19460 34130
rect 19404 33684 19460 34078
rect 19404 33618 19460 33628
rect 19516 34132 19572 34142
rect 19180 33170 19236 33180
rect 18620 32510 18622 32562
rect 18674 32510 18676 32562
rect 18620 31668 18676 32510
rect 18620 31602 18676 31612
rect 18508 31388 18900 31444
rect 18284 31042 18340 31052
rect 18172 30882 18228 30894
rect 18172 30830 18174 30882
rect 18226 30830 18228 30882
rect 18172 29652 18228 30830
rect 18732 30100 18788 30110
rect 18732 30006 18788 30044
rect 18172 29586 18228 29596
rect 18508 29540 18564 29550
rect 17948 29426 18004 29438
rect 17948 29374 17950 29426
rect 18002 29374 18004 29426
rect 17948 28868 18004 29374
rect 17948 28802 18004 28812
rect 18060 28756 18116 28766
rect 18060 26514 18116 28700
rect 18060 26462 18062 26514
rect 18114 26462 18116 26514
rect 18060 26450 18116 26462
rect 17612 26402 17836 26404
rect 17612 26350 17614 26402
rect 17666 26350 17836 26402
rect 17612 26348 17836 26350
rect 17612 26338 17668 26348
rect 17836 26338 17892 26348
rect 17388 26292 17444 26302
rect 17388 24610 17444 26236
rect 17948 25844 18004 25854
rect 17500 25508 17556 25518
rect 17500 25414 17556 25452
rect 17388 24558 17390 24610
rect 17442 24558 17444 24610
rect 17388 24546 17444 24558
rect 17612 23828 17668 23838
rect 17612 23734 17668 23772
rect 17948 23378 18004 25788
rect 18172 25394 18228 25406
rect 18172 25342 18174 25394
rect 18226 25342 18228 25394
rect 18172 24052 18228 25342
rect 18172 23986 18228 23996
rect 17948 23326 17950 23378
rect 18002 23326 18004 23378
rect 17948 23314 18004 23326
rect 18060 23940 18116 23950
rect 17500 23156 17556 23166
rect 17500 23042 17556 23100
rect 17500 22990 17502 23042
rect 17554 22990 17556 23042
rect 17500 22978 17556 22990
rect 17388 22596 17444 22606
rect 17276 22594 17444 22596
rect 17276 22542 17390 22594
rect 17442 22542 17444 22594
rect 17276 22540 17444 22542
rect 17276 22484 17332 22540
rect 16268 22418 16324 22428
rect 17276 22418 17332 22428
rect 16940 22372 16996 22382
rect 16828 22370 16996 22372
rect 16828 22318 16942 22370
rect 16994 22318 16996 22370
rect 16828 22316 16996 22318
rect 16716 22148 16772 22158
rect 16716 22054 16772 22092
rect 16828 21924 16884 22316
rect 16940 22306 16996 22316
rect 17164 22370 17220 22382
rect 17164 22318 17166 22370
rect 17218 22318 17220 22370
rect 16716 21868 16884 21924
rect 16716 21810 16772 21868
rect 16716 21758 16718 21810
rect 16770 21758 16772 21810
rect 16716 21746 16772 21758
rect 16604 21700 16660 21710
rect 16380 21588 16436 21598
rect 16380 21494 16436 21532
rect 16604 21586 16660 21644
rect 16604 21534 16606 21586
rect 16658 21534 16660 21586
rect 16604 21522 16660 21534
rect 16940 21586 16996 21598
rect 16940 21534 16942 21586
rect 16994 21534 16996 21586
rect 16156 21410 16212 21420
rect 16492 21364 16548 21374
rect 15596 20066 15652 20076
rect 15708 20300 16324 20356
rect 15708 19346 15764 20300
rect 16268 20242 16324 20300
rect 16268 20190 16270 20242
rect 16322 20190 16324 20242
rect 16268 20178 16324 20190
rect 15932 20018 15988 20030
rect 15932 19966 15934 20018
rect 15986 19966 15988 20018
rect 15932 19908 15988 19966
rect 15932 19842 15988 19852
rect 16380 19908 16436 19918
rect 15708 19294 15710 19346
rect 15762 19294 15764 19346
rect 15708 19282 15764 19294
rect 16380 19346 16436 19852
rect 16380 19294 16382 19346
rect 16434 19294 16436 19346
rect 16380 19282 16436 19294
rect 15260 19182 15262 19234
rect 15314 19182 15316 19234
rect 14812 19124 14868 19134
rect 14812 19030 14868 19068
rect 14252 18338 14644 18340
rect 14252 18286 14254 18338
rect 14306 18286 14644 18338
rect 14252 18284 14644 18286
rect 14252 18274 14308 18284
rect 14140 17780 14196 17790
rect 14140 17686 14196 17724
rect 13580 16100 13636 16110
rect 13580 16006 13636 16044
rect 12684 15932 13076 15988
rect 13916 15986 13972 16828
rect 15260 16770 15316 19182
rect 15260 16718 15262 16770
rect 15314 16718 15316 16770
rect 15260 16706 15316 16718
rect 15484 19012 15540 19022
rect 15484 16660 15540 18956
rect 15708 18338 15764 18350
rect 15708 18286 15710 18338
rect 15762 18286 15764 18338
rect 15708 17780 15764 18286
rect 15708 17108 15764 17724
rect 15932 18228 15988 18238
rect 16268 18228 16324 18238
rect 15932 17332 15988 18172
rect 16156 18226 16324 18228
rect 16156 18174 16270 18226
rect 16322 18174 16324 18226
rect 16156 18172 16324 18174
rect 16156 17668 16212 18172
rect 16268 18162 16324 18172
rect 16156 17602 16212 17612
rect 16268 17556 16324 17566
rect 16268 17462 16324 17500
rect 15932 17276 16324 17332
rect 16044 17108 16100 17118
rect 15708 17106 16100 17108
rect 15708 17054 16046 17106
rect 16098 17054 16100 17106
rect 15708 17052 16100 17054
rect 16044 17042 16100 17052
rect 16156 17108 16212 17118
rect 15596 16884 15652 16894
rect 15596 16790 15652 16828
rect 16156 16770 16212 17052
rect 16268 17106 16324 17276
rect 16268 17054 16270 17106
rect 16322 17054 16324 17106
rect 16268 17042 16324 17054
rect 16156 16718 16158 16770
rect 16210 16718 16212 16770
rect 16156 16706 16212 16718
rect 15484 16604 15652 16660
rect 13916 15934 13918 15986
rect 13970 15934 13972 15986
rect 13916 15922 13972 15934
rect 14140 16156 14420 16212
rect 13580 15202 13636 15214
rect 13580 15150 13582 15202
rect 13634 15150 13636 15202
rect 13580 15148 13636 15150
rect 14140 15148 14196 16156
rect 14364 16100 14420 16156
rect 14476 16100 14532 16110
rect 14364 16098 14532 16100
rect 14364 16046 14478 16098
rect 14530 16046 14532 16098
rect 14364 16044 14532 16046
rect 14476 16034 14532 16044
rect 15148 16100 15204 16110
rect 15148 16006 15204 16044
rect 13580 15092 14196 15148
rect 14252 15986 14308 15998
rect 14252 15934 14254 15986
rect 14306 15934 14308 15986
rect 14252 15148 14308 15934
rect 14812 15986 14868 15998
rect 14812 15934 14814 15986
rect 14866 15934 14868 15986
rect 14476 15876 14532 15886
rect 14476 15782 14532 15820
rect 14252 15092 14756 15148
rect 12572 14588 12740 14644
rect 12124 14420 12180 14430
rect 12572 14420 12628 14430
rect 12124 14418 12572 14420
rect 12124 14366 12126 14418
rect 12178 14366 12572 14418
rect 12124 14364 12572 14366
rect 12124 14354 12180 14364
rect 12572 14326 12628 14364
rect 12236 14196 12292 14206
rect 12012 14140 12180 14196
rect 11900 13860 11956 13870
rect 11676 13858 11956 13860
rect 11676 13806 11902 13858
rect 11954 13806 11956 13858
rect 11676 13804 11956 13806
rect 11900 13794 11956 13804
rect 12012 13636 12068 13646
rect 12012 13542 12068 13580
rect 11228 13074 11620 13076
rect 11228 13022 11230 13074
rect 11282 13022 11620 13074
rect 11228 13020 11620 13022
rect 11676 13300 11732 13310
rect 11228 13010 11284 13020
rect 11676 12964 11732 13244
rect 12124 13076 12180 14140
rect 12236 13746 12292 14140
rect 12236 13694 12238 13746
rect 12290 13694 12292 13746
rect 12236 13682 12292 13694
rect 12124 12982 12180 13020
rect 11340 12962 11732 12964
rect 11340 12910 11678 12962
rect 11730 12910 11732 12962
rect 11340 12908 11732 12910
rect 11116 12796 11284 12852
rect 10780 12126 10782 12178
rect 10834 12126 10836 12178
rect 10220 11508 10276 11518
rect 10108 11506 10276 11508
rect 10108 11454 10222 11506
rect 10274 11454 10276 11506
rect 10108 11452 10276 11454
rect 10220 11442 10276 11452
rect 9884 10670 9886 10722
rect 9938 10670 9940 10722
rect 9884 10658 9940 10670
rect 9996 11172 10052 11182
rect 9996 10612 10052 11116
rect 10668 11172 10724 11182
rect 10668 11078 10724 11116
rect 10780 10948 10836 12126
rect 10220 10892 10836 10948
rect 10892 11620 10948 11630
rect 10892 11394 10948 11564
rect 10892 11342 10894 11394
rect 10946 11342 10948 11394
rect 10108 10836 10164 10846
rect 10108 10722 10164 10780
rect 10108 10670 10110 10722
rect 10162 10670 10164 10722
rect 10108 10658 10164 10670
rect 9996 10546 10052 10556
rect 9436 10444 9716 10500
rect 7196 9940 7252 9950
rect 7196 9156 7252 9884
rect 8540 9940 8596 9950
rect 8540 9846 8596 9884
rect 7196 9062 7252 9100
rect 7308 9268 7364 9278
rect 7308 9154 7364 9212
rect 7308 9102 7310 9154
rect 7362 9102 7364 9154
rect 7308 9090 7364 9102
rect 9660 9266 9716 10444
rect 9660 9214 9662 9266
rect 9714 9214 9716 9266
rect 6972 8990 6974 9042
rect 7026 8990 7028 9042
rect 6972 8428 7028 8990
rect 7756 8820 7812 8830
rect 7756 8726 7812 8764
rect 8540 8820 8596 8830
rect 5068 7982 5070 8034
rect 5122 7982 5124 8034
rect 4620 7700 4676 7710
rect 3724 7646 3726 7698
rect 3778 7646 3780 7698
rect 3500 7634 3556 7644
rect 3724 7634 3780 7646
rect 4284 7698 4676 7700
rect 4284 7646 4622 7698
rect 4674 7646 4676 7698
rect 4284 7644 4676 7646
rect 4172 7588 4228 7598
rect 3388 7410 3444 7420
rect 4060 7476 4116 7486
rect 2828 7310 2830 7362
rect 2882 7310 2884 7362
rect 2828 7298 2884 7310
rect 3612 7362 3668 7374
rect 3612 7310 3614 7362
rect 3666 7310 3668 7362
rect 3164 7252 3220 7262
rect 3612 7252 3668 7310
rect 3164 7250 3668 7252
rect 3164 7198 3166 7250
rect 3218 7198 3668 7250
rect 3164 7196 3668 7198
rect 3164 7186 3220 7196
rect 1820 6638 1822 6690
rect 1874 6638 1876 6690
rect 1820 5012 1876 6638
rect 2492 6578 2548 6590
rect 2492 6526 2494 6578
rect 2546 6526 2548 6578
rect 2492 6132 2548 6526
rect 2492 6066 2548 6076
rect 4060 5684 4116 7420
rect 4172 7474 4228 7532
rect 4172 7422 4174 7474
rect 4226 7422 4228 7474
rect 4172 7410 4228 7422
rect 4172 5908 4228 5918
rect 4284 5908 4340 7644
rect 4620 7634 4676 7644
rect 5068 7588 5124 7982
rect 4396 7476 4452 7486
rect 4396 7382 4452 7420
rect 5068 7474 5124 7532
rect 5068 7422 5070 7474
rect 5122 7422 5124 7474
rect 4508 7362 4564 7374
rect 4508 7310 4510 7362
rect 4562 7310 4564 7362
rect 4508 7252 4564 7310
rect 4508 7196 5012 7252
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4620 6802 4676 6814
rect 4620 6750 4622 6802
rect 4674 6750 4676 6802
rect 4620 5908 4676 6750
rect 4732 6580 4788 6590
rect 4732 6130 4788 6524
rect 4732 6078 4734 6130
rect 4786 6078 4788 6130
rect 4732 6066 4788 6078
rect 4956 6020 5012 7196
rect 5068 6804 5124 7422
rect 5516 8372 5908 8428
rect 6972 8372 8148 8428
rect 5516 8260 5572 8372
rect 5852 8370 5908 8372
rect 5852 8318 5854 8370
rect 5906 8318 5908 8370
rect 5852 8306 5908 8318
rect 5516 7474 5572 8204
rect 5516 7422 5518 7474
rect 5570 7422 5572 7474
rect 5516 7410 5572 7422
rect 6188 7364 6244 7374
rect 6188 7362 6468 7364
rect 6188 7310 6190 7362
rect 6242 7310 6468 7362
rect 6188 7308 6468 7310
rect 6188 7298 6244 7308
rect 5180 6804 5236 6814
rect 5068 6802 5236 6804
rect 5068 6750 5182 6802
rect 5234 6750 5236 6802
rect 5068 6748 5236 6750
rect 5180 6738 5236 6748
rect 6412 6802 6468 7308
rect 6412 6750 6414 6802
rect 6466 6750 6468 6802
rect 6412 6738 6468 6750
rect 6748 6804 6804 6814
rect 5628 6580 5684 6590
rect 5684 6524 5908 6580
rect 5628 6486 5684 6524
rect 5404 6468 5460 6478
rect 5180 6132 5236 6142
rect 5180 6038 5236 6076
rect 5068 6020 5124 6030
rect 4956 6018 5124 6020
rect 4956 5966 5070 6018
rect 5122 5966 5124 6018
rect 4956 5964 5124 5966
rect 5068 5954 5124 5964
rect 4172 5906 4676 5908
rect 4172 5854 4174 5906
rect 4226 5854 4676 5906
rect 4172 5852 4676 5854
rect 5404 5906 5460 6412
rect 5404 5854 5406 5906
rect 5458 5854 5460 5906
rect 4172 5842 4228 5852
rect 5404 5842 5460 5854
rect 4396 5684 4452 5694
rect 4060 5682 4452 5684
rect 4060 5630 4398 5682
rect 4450 5630 4452 5682
rect 4060 5628 4452 5630
rect 4396 5618 4452 5628
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 5852 5122 5908 6524
rect 6300 6578 6356 6590
rect 6300 6526 6302 6578
rect 6354 6526 6356 6578
rect 5964 6468 6020 6478
rect 6300 6468 6356 6526
rect 5964 6466 6300 6468
rect 5964 6414 5966 6466
rect 6018 6414 6300 6466
rect 5964 6412 6300 6414
rect 5964 6402 6020 6412
rect 6300 6402 6356 6412
rect 6636 6578 6692 6590
rect 6636 6526 6638 6578
rect 6690 6526 6692 6578
rect 5852 5070 5854 5122
rect 5906 5070 5908 5122
rect 5852 5058 5908 5070
rect 5964 6244 6020 6254
rect 1820 4946 1876 4956
rect 4172 5012 4228 5022
rect 4172 4338 4228 4956
rect 5964 5010 6020 6188
rect 6636 6244 6692 6526
rect 6636 6178 6692 6188
rect 6524 5908 6580 5918
rect 6524 5814 6580 5852
rect 6188 5794 6244 5806
rect 6188 5742 6190 5794
rect 6242 5742 6244 5794
rect 6188 5122 6244 5742
rect 6188 5070 6190 5122
rect 6242 5070 6244 5122
rect 6188 5058 6244 5070
rect 6748 5122 6804 6748
rect 6860 6692 6916 6702
rect 7308 6692 7364 6702
rect 6860 6690 7364 6692
rect 6860 6638 6862 6690
rect 6914 6638 7310 6690
rect 7362 6638 7364 6690
rect 6860 6636 7364 6638
rect 6860 6626 6916 6636
rect 7308 6626 7364 6636
rect 7868 6690 7924 6702
rect 7868 6638 7870 6690
rect 7922 6638 7924 6690
rect 7196 6468 7252 6478
rect 7084 5908 7140 5918
rect 7196 5908 7252 6412
rect 7420 6466 7476 6478
rect 7420 6414 7422 6466
rect 7474 6414 7476 6466
rect 7420 6244 7476 6414
rect 7420 6178 7476 6188
rect 7868 6132 7924 6638
rect 7868 6066 7924 6076
rect 7980 6244 8036 6254
rect 7980 6018 8036 6188
rect 7980 5966 7982 6018
rect 8034 5966 8036 6018
rect 7980 5954 8036 5966
rect 7420 5908 7476 5918
rect 7196 5906 7476 5908
rect 7196 5854 7422 5906
rect 7474 5854 7476 5906
rect 7196 5852 7476 5854
rect 6748 5070 6750 5122
rect 6802 5070 6804 5122
rect 6748 5058 6804 5070
rect 6972 5794 7028 5806
rect 6972 5742 6974 5794
rect 7026 5742 7028 5794
rect 5964 4958 5966 5010
rect 6018 4958 6020 5010
rect 5964 4946 6020 4958
rect 4172 4286 4174 4338
rect 4226 4286 4228 4338
rect 4172 4274 4228 4286
rect 4956 4228 5012 4238
rect 4956 4134 5012 4172
rect 6972 4004 7028 5742
rect 7084 4226 7140 5852
rect 7420 5842 7476 5852
rect 7868 5908 7924 5918
rect 7868 5814 7924 5852
rect 8092 5906 8148 8372
rect 8204 7476 8260 7486
rect 8204 6804 8260 7420
rect 8204 6690 8260 6748
rect 8204 6638 8206 6690
rect 8258 6638 8260 6690
rect 8204 6626 8260 6638
rect 8316 7362 8372 7374
rect 8316 7310 8318 7362
rect 8370 7310 8372 7362
rect 8316 6244 8372 7310
rect 8316 6178 8372 6188
rect 8092 5854 8094 5906
rect 8146 5854 8148 5906
rect 8092 5842 8148 5854
rect 7196 5684 7252 5694
rect 7196 5682 7476 5684
rect 7196 5630 7198 5682
rect 7250 5630 7476 5682
rect 7196 5628 7476 5630
rect 7196 5618 7252 5628
rect 7420 4450 7476 5628
rect 7532 5012 7588 5022
rect 7532 5010 7812 5012
rect 7532 4958 7534 5010
rect 7586 4958 7812 5010
rect 7532 4956 7812 4958
rect 7532 4946 7588 4956
rect 7756 4562 7812 4956
rect 7756 4510 7758 4562
rect 7810 4510 7812 4562
rect 7756 4498 7812 4510
rect 7420 4398 7422 4450
rect 7474 4398 7476 4450
rect 7420 4386 7476 4398
rect 8540 4452 8596 8764
rect 9660 8428 9716 9214
rect 8764 8372 9716 8428
rect 8652 7476 8708 7486
rect 8764 7476 8820 8372
rect 8988 8148 9044 8158
rect 8988 7586 9044 8092
rect 8988 7534 8990 7586
rect 9042 7534 9044 7586
rect 8988 7522 9044 7534
rect 8652 7474 8820 7476
rect 8652 7422 8654 7474
rect 8706 7422 8820 7474
rect 8652 7420 8820 7422
rect 9660 7476 9716 7486
rect 8652 5796 8708 7420
rect 8876 7364 8932 7374
rect 8876 7270 8932 7308
rect 8988 6804 9044 6814
rect 9660 6804 9716 7420
rect 9660 6748 10164 6804
rect 8988 6690 9044 6748
rect 8988 6638 8990 6690
rect 9042 6638 9044 6690
rect 8988 6626 9044 6638
rect 8764 6132 8820 6142
rect 8764 6038 8820 6076
rect 9660 5908 9716 5918
rect 8764 5796 8820 5806
rect 8652 5740 8764 5796
rect 8764 5730 8820 5740
rect 9660 5234 9716 5852
rect 9660 5182 9662 5234
rect 9714 5182 9716 5234
rect 9660 5170 9716 5182
rect 10108 5794 10164 6748
rect 10220 6132 10276 10892
rect 10332 10612 10388 10622
rect 10332 9042 10388 10556
rect 10892 10612 10948 11342
rect 11116 11396 11172 11406
rect 11004 11170 11060 11182
rect 11004 11118 11006 11170
rect 11058 11118 11060 11170
rect 11004 10836 11060 11118
rect 11004 10770 11060 10780
rect 11116 10724 11172 11340
rect 11116 10658 11172 10668
rect 10892 10546 10948 10556
rect 10892 9996 11172 10052
rect 10444 9828 10500 9838
rect 10668 9828 10724 9838
rect 10892 9828 10948 9996
rect 10444 9826 10612 9828
rect 10444 9774 10446 9826
rect 10498 9774 10612 9826
rect 10444 9772 10612 9774
rect 10444 9762 10500 9772
rect 10332 8990 10334 9042
rect 10386 8990 10388 9042
rect 10332 8978 10388 8990
rect 10444 9604 10500 9614
rect 10332 7364 10388 7374
rect 10332 7270 10388 7308
rect 10444 6804 10500 9548
rect 10556 9492 10612 9772
rect 10668 9826 10948 9828
rect 10668 9774 10670 9826
rect 10722 9774 10948 9826
rect 10668 9772 10948 9774
rect 11004 9826 11060 9838
rect 11004 9774 11006 9826
rect 11058 9774 11060 9826
rect 10668 9762 10724 9772
rect 11004 9716 11060 9774
rect 10892 9660 11004 9716
rect 10780 9604 10836 9614
rect 10780 9510 10836 9548
rect 10556 9436 10724 9492
rect 10668 9268 10724 9436
rect 10780 9268 10836 9278
rect 10668 9266 10836 9268
rect 10668 9214 10782 9266
rect 10834 9214 10836 9266
rect 10668 9212 10836 9214
rect 10780 9202 10836 9212
rect 10892 9266 10948 9660
rect 11004 9650 11060 9660
rect 10892 9214 10894 9266
rect 10946 9214 10948 9266
rect 10892 9202 10948 9214
rect 10668 9044 10724 9054
rect 11116 9044 11172 9996
rect 10668 9042 11172 9044
rect 10668 8990 10670 9042
rect 10722 8990 11172 9042
rect 10668 8988 11172 8990
rect 11228 9940 11284 12796
rect 11340 12404 11396 12908
rect 11676 12898 11732 12908
rect 12684 12962 12740 14588
rect 13468 14420 13524 14430
rect 13468 14326 13524 14364
rect 13580 14418 13636 15092
rect 13580 14366 13582 14418
rect 13634 14366 13636 14418
rect 13580 14354 13636 14366
rect 14028 14420 14084 15092
rect 12908 14308 12964 14318
rect 13804 14308 13860 14318
rect 12908 14214 12964 14252
rect 13692 14306 13860 14308
rect 13692 14254 13806 14306
rect 13858 14254 13860 14306
rect 13692 14252 13860 14254
rect 13692 13074 13748 14252
rect 13804 14242 13860 14252
rect 14028 13858 14084 14364
rect 14028 13806 14030 13858
rect 14082 13806 14084 13858
rect 14028 13794 14084 13806
rect 14700 14420 14756 15092
rect 14812 14644 14868 15934
rect 15484 15874 15540 15886
rect 15484 15822 15486 15874
rect 15538 15822 15540 15874
rect 15484 15148 15540 15822
rect 15260 15092 15540 15148
rect 14924 14644 14980 14654
rect 14812 14642 14980 14644
rect 14812 14590 14926 14642
rect 14978 14590 14980 14642
rect 14812 14588 14980 14590
rect 14924 14578 14980 14588
rect 15036 14530 15092 14542
rect 15036 14478 15038 14530
rect 15090 14478 15092 14530
rect 14812 14420 14868 14430
rect 14700 14418 14868 14420
rect 14700 14366 14814 14418
rect 14866 14366 14868 14418
rect 14700 14364 14868 14366
rect 14700 14308 14756 14364
rect 14812 14354 14868 14364
rect 14924 14420 14980 14430
rect 15036 14420 15092 14478
rect 14980 14364 15092 14420
rect 14924 14354 14980 14364
rect 14140 13746 14196 13758
rect 14140 13694 14142 13746
rect 14194 13694 14196 13746
rect 13692 13022 13694 13074
rect 13746 13022 13748 13074
rect 13692 13010 13748 13022
rect 13804 13636 13860 13646
rect 12684 12910 12686 12962
rect 12738 12910 12740 12962
rect 11340 12310 11396 12348
rect 12460 12738 12516 12750
rect 12460 12686 12462 12738
rect 12514 12686 12516 12738
rect 11676 12292 11732 12302
rect 11676 12198 11732 12236
rect 12012 12290 12068 12302
rect 12012 12238 12014 12290
rect 12066 12238 12068 12290
rect 12012 12180 12068 12238
rect 11788 12124 12012 12180
rect 11676 11732 11732 11742
rect 11564 11284 11620 11294
rect 11564 11190 11620 11228
rect 11676 11282 11732 11676
rect 11676 11230 11678 11282
rect 11730 11230 11732 11282
rect 11676 11218 11732 11230
rect 11340 9940 11396 9950
rect 11228 9938 11396 9940
rect 11228 9886 11342 9938
rect 11394 9886 11396 9938
rect 11228 9884 11396 9886
rect 10668 7812 10724 8988
rect 11228 8428 11284 9884
rect 11340 9874 11396 9884
rect 11116 8372 11284 8428
rect 11564 9042 11620 9054
rect 11564 8990 11566 9042
rect 11618 8990 11620 9042
rect 10892 8260 10948 8270
rect 11116 8260 11172 8372
rect 10892 8258 11172 8260
rect 10892 8206 10894 8258
rect 10946 8206 11172 8258
rect 10892 8204 11172 8206
rect 10892 8194 10948 8204
rect 10668 7756 11060 7812
rect 10444 6738 10500 6748
rect 10780 7588 10836 7598
rect 10220 6066 10276 6076
rect 10108 5742 10110 5794
rect 10162 5742 10164 5794
rect 10108 5122 10164 5742
rect 10780 5234 10836 7532
rect 11004 6804 11060 7756
rect 11116 7028 11172 8204
rect 11228 8148 11284 8158
rect 11228 8054 11284 8092
rect 11564 7476 11620 8990
rect 11788 8428 11844 12124
rect 12012 12114 12068 12124
rect 12348 12178 12404 12190
rect 12348 12126 12350 12178
rect 12402 12126 12404 12178
rect 12348 12068 12404 12126
rect 12460 12068 12516 12686
rect 12684 12292 12740 12910
rect 12684 12226 12740 12236
rect 12796 12068 12852 12078
rect 12348 12066 12852 12068
rect 12348 12014 12798 12066
rect 12850 12014 12852 12066
rect 12348 12012 12852 12014
rect 12796 11732 12852 12012
rect 13356 12068 13412 12078
rect 13356 11974 13412 12012
rect 13804 11732 13860 13580
rect 14028 12964 14084 12974
rect 14140 12964 14196 13694
rect 14588 13748 14644 13758
rect 14700 13748 14756 14252
rect 14588 13746 14756 13748
rect 14588 13694 14590 13746
rect 14642 13694 14756 13746
rect 14588 13692 14756 13694
rect 15260 13748 15316 15092
rect 15484 14644 15540 14654
rect 15484 14530 15540 14588
rect 15484 14478 15486 14530
rect 15538 14478 15540 14530
rect 15484 14466 15540 14478
rect 14588 13682 14644 13692
rect 15260 13682 15316 13692
rect 14812 13524 14868 13534
rect 14812 13522 14980 13524
rect 14812 13470 14814 13522
rect 14866 13470 14980 13522
rect 14812 13468 14980 13470
rect 14812 13458 14868 13468
rect 14028 12962 14196 12964
rect 14028 12910 14030 12962
rect 14082 12910 14196 12962
rect 14028 12908 14196 12910
rect 14028 12068 14084 12908
rect 14476 12852 14532 12862
rect 14812 12852 14868 12862
rect 14476 12850 14868 12852
rect 14476 12798 14478 12850
rect 14530 12798 14814 12850
rect 14866 12798 14868 12850
rect 14476 12796 14868 12798
rect 14476 12786 14532 12796
rect 14812 12786 14868 12796
rect 14924 12068 14980 13468
rect 15148 13076 15204 13086
rect 15148 13074 15540 13076
rect 15148 13022 15150 13074
rect 15202 13022 15540 13074
rect 15148 13020 15540 13022
rect 15148 13010 15204 13020
rect 15036 12852 15092 12862
rect 15260 12852 15316 12862
rect 15036 12850 15260 12852
rect 15036 12798 15038 12850
rect 15090 12798 15260 12850
rect 15036 12796 15260 12798
rect 15036 12786 15092 12796
rect 15260 12786 15316 12796
rect 15484 12290 15540 13020
rect 15484 12238 15486 12290
rect 15538 12238 15540 12290
rect 15484 12226 15540 12238
rect 15596 12852 15652 16604
rect 15708 15876 15764 15886
rect 15708 15426 15764 15820
rect 15708 15374 15710 15426
rect 15762 15374 15764 15426
rect 15708 15362 15764 15374
rect 16380 15314 16436 15326
rect 16380 15262 16382 15314
rect 16434 15262 16436 15314
rect 16380 15148 16436 15262
rect 15932 15092 16436 15148
rect 15708 14644 15764 14654
rect 15708 13970 15764 14588
rect 15708 13918 15710 13970
rect 15762 13918 15764 13970
rect 15708 13906 15764 13918
rect 15932 14530 15988 15092
rect 15932 14478 15934 14530
rect 15986 14478 15988 14530
rect 15596 12738 15652 12796
rect 15596 12686 15598 12738
rect 15650 12686 15652 12738
rect 14924 12012 15204 12068
rect 14028 12002 14084 12012
rect 12796 11676 13076 11732
rect 12124 11396 12180 11406
rect 12124 11302 12180 11340
rect 12236 11284 12292 11294
rect 12236 11190 12292 11228
rect 11900 11172 11956 11182
rect 11900 11170 12068 11172
rect 11900 11118 11902 11170
rect 11954 11118 12068 11170
rect 11900 11116 12068 11118
rect 11900 11106 11956 11116
rect 12012 10052 12068 11116
rect 12348 11170 12404 11182
rect 12572 11172 12628 11182
rect 12348 11118 12350 11170
rect 12402 11118 12404 11170
rect 12236 10612 12292 10622
rect 12348 10612 12404 11118
rect 12292 10556 12404 10612
rect 12460 11170 12628 11172
rect 12460 11118 12574 11170
rect 12626 11118 12628 11170
rect 12460 11116 12628 11118
rect 12236 10518 12292 10556
rect 12460 10386 12516 11116
rect 12572 11106 12628 11116
rect 12572 10836 12628 10846
rect 12572 10834 12964 10836
rect 12572 10782 12574 10834
rect 12626 10782 12964 10834
rect 12572 10780 12964 10782
rect 12572 10770 12628 10780
rect 12684 10612 12740 10622
rect 12684 10518 12740 10556
rect 12460 10334 12462 10386
rect 12514 10334 12516 10386
rect 12236 10052 12292 10062
rect 12012 10050 12292 10052
rect 12012 9998 12238 10050
rect 12290 9998 12292 10050
rect 12012 9996 12292 9998
rect 12236 9986 12292 9996
rect 12460 10052 12516 10334
rect 12460 9986 12516 9996
rect 12572 9826 12628 9838
rect 12572 9774 12574 9826
rect 12626 9774 12628 9826
rect 12572 9716 12628 9774
rect 12348 9602 12404 9614
rect 12348 9550 12350 9602
rect 12402 9550 12404 9602
rect 12348 9154 12404 9550
rect 12348 9102 12350 9154
rect 12402 9102 12404 9154
rect 12348 9090 12404 9102
rect 12124 8484 12180 8494
rect 11788 8372 12068 8428
rect 11900 8260 11956 8270
rect 11900 8166 11956 8204
rect 11564 7410 11620 7420
rect 11116 6972 11284 7028
rect 11116 6804 11172 6814
rect 11004 6748 11116 6804
rect 11116 6710 11172 6748
rect 11228 6692 11284 6972
rect 12012 6802 12068 8372
rect 12124 8370 12180 8428
rect 12124 8318 12126 8370
rect 12178 8318 12180 8370
rect 12124 8306 12180 8318
rect 12460 8260 12516 8270
rect 12460 7362 12516 8204
rect 12460 7310 12462 7362
rect 12514 7310 12516 7362
rect 12012 6750 12014 6802
rect 12066 6750 12068 6802
rect 12012 6738 12068 6750
rect 12124 6804 12180 6814
rect 11228 6626 11284 6636
rect 12124 6578 12180 6748
rect 12124 6526 12126 6578
rect 12178 6526 12180 6578
rect 12124 6514 12180 6526
rect 12460 6578 12516 7310
rect 12572 8034 12628 9660
rect 12908 8260 12964 10780
rect 13020 10164 13076 11676
rect 13804 11666 13860 11676
rect 15036 10724 15092 10734
rect 14812 10722 15092 10724
rect 14812 10670 15038 10722
rect 15090 10670 15092 10722
rect 14812 10668 15092 10670
rect 13132 10164 13188 10174
rect 13020 10108 13132 10164
rect 13132 10098 13188 10108
rect 13580 10052 13636 10062
rect 13580 9958 13636 9996
rect 13692 9996 14532 10052
rect 13692 9938 13748 9996
rect 13692 9886 13694 9938
rect 13746 9886 13748 9938
rect 13692 9874 13748 9886
rect 14140 9826 14196 9838
rect 14140 9774 14142 9826
rect 14194 9774 14196 9826
rect 13580 8484 13636 8522
rect 13580 8418 13636 8428
rect 13804 8484 13860 8494
rect 12908 8166 12964 8204
rect 13692 8260 13748 8270
rect 13692 8166 13748 8204
rect 13580 8036 13636 8046
rect 12572 7982 12574 8034
rect 12626 7982 12628 8034
rect 12572 6690 12628 7982
rect 13468 8034 13636 8036
rect 13468 7982 13582 8034
rect 13634 7982 13636 8034
rect 13468 7980 13636 7982
rect 12796 7588 12852 7598
rect 12796 7494 12852 7532
rect 13020 7474 13076 7486
rect 13020 7422 13022 7474
rect 13074 7422 13076 7474
rect 13020 6914 13076 7422
rect 13020 6862 13022 6914
rect 13074 6862 13076 6914
rect 13020 6850 13076 6862
rect 13356 6804 13412 6814
rect 13468 6804 13524 7980
rect 13580 7970 13636 7980
rect 13412 6748 13524 6804
rect 13804 7474 13860 8428
rect 14140 8484 14196 9774
rect 14476 8930 14532 9996
rect 14812 9938 14868 10668
rect 15036 10658 15092 10668
rect 15148 10612 15204 12012
rect 15596 11956 15652 12686
rect 15932 12180 15988 14478
rect 16268 13076 16324 13086
rect 16268 12982 16324 13020
rect 16268 12180 16324 12190
rect 15932 12178 16324 12180
rect 15932 12126 16270 12178
rect 16322 12126 16324 12178
rect 15932 12124 16324 12126
rect 15596 11890 15652 11900
rect 16268 11732 16324 12124
rect 16268 11666 16324 11676
rect 15372 11396 15428 11406
rect 15260 10612 15316 10622
rect 15148 10610 15316 10612
rect 15148 10558 15262 10610
rect 15314 10558 15316 10610
rect 15148 10556 15316 10558
rect 15260 10546 15316 10556
rect 15372 10612 15428 11340
rect 16044 11394 16100 11406
rect 16044 11342 16046 11394
rect 16098 11342 16100 11394
rect 15596 11284 15652 11294
rect 15596 11190 15652 11228
rect 15372 10546 15428 10556
rect 14812 9886 14814 9938
rect 14866 9886 14868 9938
rect 14812 9874 14868 9886
rect 14476 8878 14478 8930
rect 14530 8878 14532 8930
rect 14476 8866 14532 8878
rect 15932 9154 15988 9166
rect 15932 9102 15934 9154
rect 15986 9102 15988 9154
rect 14140 8418 14196 8428
rect 14588 8036 14644 8046
rect 14588 7586 14644 7980
rect 14588 7534 14590 7586
rect 14642 7534 14644 7586
rect 14588 7522 14644 7534
rect 13804 7422 13806 7474
rect 13858 7422 13860 7474
rect 13356 6738 13412 6748
rect 12572 6638 12574 6690
rect 12626 6638 12628 6690
rect 12572 6626 12628 6638
rect 13580 6692 13636 6702
rect 13804 6692 13860 7422
rect 13580 6690 13860 6692
rect 13580 6638 13582 6690
rect 13634 6638 13860 6690
rect 13580 6636 13860 6638
rect 15596 6692 15652 6702
rect 12460 6526 12462 6578
rect 12514 6526 12516 6578
rect 12460 6514 12516 6526
rect 10780 5182 10782 5234
rect 10834 5182 10836 5234
rect 10780 5170 10836 5182
rect 12908 5234 12964 5246
rect 12908 5182 12910 5234
rect 12962 5182 12964 5234
rect 10108 5070 10110 5122
rect 10162 5070 10164 5122
rect 8652 4452 8708 4462
rect 8540 4450 8708 4452
rect 8540 4398 8654 4450
rect 8706 4398 8708 4450
rect 8540 4396 8708 4398
rect 8652 4386 8708 4396
rect 8988 4452 9044 4462
rect 8988 4358 9044 4396
rect 10108 4340 10164 5070
rect 11004 4452 11060 4462
rect 11004 4358 11060 4396
rect 10220 4340 10276 4350
rect 10108 4338 10276 4340
rect 10108 4286 10222 4338
rect 10274 4286 10276 4338
rect 10108 4284 10276 4286
rect 10220 4274 10276 4284
rect 12908 4340 12964 5182
rect 12908 4274 12964 4284
rect 13580 4338 13636 6636
rect 14252 6580 14308 6590
rect 14252 6486 14308 6524
rect 15596 6132 15652 6636
rect 15148 6130 15652 6132
rect 15148 6078 15598 6130
rect 15650 6078 15652 6130
rect 15148 6076 15652 6078
rect 15036 6020 15092 6030
rect 14924 5236 14980 5246
rect 14252 5234 14980 5236
rect 14252 5182 14926 5234
rect 14978 5182 14980 5234
rect 14252 5180 14980 5182
rect 14252 4450 14308 5180
rect 14924 5170 14980 5180
rect 15036 5010 15092 5964
rect 15148 5906 15204 6076
rect 15596 6066 15652 6076
rect 15932 6020 15988 9102
rect 16044 9156 16100 11342
rect 16492 10500 16548 21308
rect 16940 21140 16996 21534
rect 16940 21074 16996 21084
rect 17164 21028 17220 22318
rect 17388 21476 17444 22540
rect 17836 22484 17892 22494
rect 17836 22390 17892 22428
rect 17500 22260 17556 22270
rect 17500 22258 17892 22260
rect 17500 22206 17502 22258
rect 17554 22206 17892 22258
rect 17500 22204 17892 22206
rect 17500 22194 17556 22204
rect 17388 21420 17780 21476
rect 17164 20962 17220 20972
rect 17500 21252 17556 21262
rect 17164 20804 17220 20814
rect 16828 20802 17220 20804
rect 16828 20750 17166 20802
rect 17218 20750 17220 20802
rect 16828 20748 17220 20750
rect 16604 20580 16660 20590
rect 16604 20018 16660 20524
rect 16604 19966 16606 20018
rect 16658 19966 16660 20018
rect 16604 19954 16660 19966
rect 16828 20244 16884 20748
rect 17164 20738 17220 20748
rect 16828 20018 16884 20188
rect 16828 19966 16830 20018
rect 16882 19966 16884 20018
rect 16828 19954 16884 19966
rect 17500 19236 17556 21196
rect 17052 19234 17556 19236
rect 17052 19182 17502 19234
rect 17554 19182 17556 19234
rect 17052 19180 17556 19182
rect 16940 18340 16996 18350
rect 16940 18246 16996 18284
rect 17052 17666 17108 19180
rect 17500 19170 17556 19180
rect 17500 18562 17556 18574
rect 17500 18510 17502 18562
rect 17554 18510 17556 18562
rect 17500 18228 17556 18510
rect 17500 18162 17556 18172
rect 17052 17614 17054 17666
rect 17106 17614 17108 17666
rect 17052 17602 17108 17614
rect 17612 17668 17668 17678
rect 17388 17554 17444 17566
rect 17388 17502 17390 17554
rect 17442 17502 17444 17554
rect 17388 17108 17444 17502
rect 17500 17556 17556 17566
rect 17500 17462 17556 17500
rect 17612 17554 17668 17612
rect 17612 17502 17614 17554
rect 17666 17502 17668 17554
rect 17612 17490 17668 17502
rect 17388 17042 17444 17052
rect 17724 15876 17780 21420
rect 17836 19348 17892 22204
rect 18060 21698 18116 23884
rect 18060 21646 18062 21698
rect 18114 21646 18116 21698
rect 18060 21252 18116 21646
rect 18060 21186 18116 21196
rect 18284 22820 18340 22830
rect 18284 20690 18340 22764
rect 18396 21364 18452 21374
rect 18396 20914 18452 21308
rect 18396 20862 18398 20914
rect 18450 20862 18452 20914
rect 18396 20850 18452 20862
rect 18284 20638 18286 20690
rect 18338 20638 18340 20690
rect 18284 20626 18340 20638
rect 18172 19348 18228 19358
rect 17836 19346 18228 19348
rect 17836 19294 18174 19346
rect 18226 19294 18228 19346
rect 17836 19292 18228 19294
rect 18172 19282 18228 19292
rect 18508 18676 18564 29484
rect 18844 29540 18900 31388
rect 19180 30100 19236 30110
rect 18956 29652 19012 29662
rect 18956 29558 19012 29596
rect 18844 28644 18900 29484
rect 19068 29314 19124 29326
rect 19068 29262 19070 29314
rect 19122 29262 19124 29314
rect 19068 28866 19124 29262
rect 19068 28814 19070 28866
rect 19122 28814 19124 28866
rect 19068 28802 19124 28814
rect 19180 28756 19236 30044
rect 19516 29652 19572 34076
rect 19628 34130 19684 34142
rect 20524 34132 20580 34142
rect 19628 34078 19630 34130
rect 19682 34078 19684 34130
rect 19628 31668 19684 34078
rect 20300 34130 20580 34132
rect 20300 34078 20526 34130
rect 20578 34078 20580 34130
rect 20300 34076 20580 34078
rect 20076 34018 20132 34030
rect 20076 33966 20078 34018
rect 20130 33966 20132 34018
rect 20076 33684 20132 33966
rect 20076 33618 20132 33628
rect 20188 33460 20244 33470
rect 20300 33460 20356 34076
rect 20524 34066 20580 34076
rect 20244 33404 20356 33460
rect 20412 33908 20468 33918
rect 20412 33458 20468 33852
rect 20412 33406 20414 33458
rect 20466 33406 20468 33458
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 20188 32676 20244 33404
rect 20412 33394 20468 33406
rect 20860 33684 20916 33694
rect 20188 32674 20692 32676
rect 20188 32622 20190 32674
rect 20242 32622 20692 32674
rect 20188 32620 20692 32622
rect 20188 32610 20244 32620
rect 20636 31780 20692 32620
rect 20636 31686 20692 31724
rect 19628 31602 19684 31612
rect 19964 31668 20020 31678
rect 19964 31666 20580 31668
rect 19964 31614 19966 31666
rect 20018 31614 20580 31666
rect 19964 31612 20580 31614
rect 19964 31602 20020 31612
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 20524 31220 20580 31612
rect 20636 31220 20692 31230
rect 20524 31218 20692 31220
rect 20524 31166 20638 31218
rect 20690 31166 20692 31218
rect 20524 31164 20692 31166
rect 20636 31154 20692 31164
rect 20748 31108 20804 31118
rect 20748 31014 20804 31052
rect 20300 30884 20356 30894
rect 20188 30882 20356 30884
rect 20188 30830 20302 30882
rect 20354 30830 20356 30882
rect 20188 30828 20356 30830
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19516 29596 19796 29652
rect 19292 28868 19348 28878
rect 19740 28868 19796 29596
rect 19292 28866 19684 28868
rect 19292 28814 19294 28866
rect 19346 28814 19684 28866
rect 19292 28812 19684 28814
rect 19292 28802 19348 28812
rect 19180 28662 19236 28700
rect 19628 28754 19684 28812
rect 19628 28702 19630 28754
rect 19682 28702 19684 28754
rect 19628 28690 19684 28702
rect 18620 28420 18676 28430
rect 18620 27858 18676 28364
rect 18844 28082 18900 28588
rect 19292 28644 19348 28654
rect 19348 28588 19460 28644
rect 19292 28578 19348 28588
rect 18844 28030 18846 28082
rect 18898 28030 18900 28082
rect 18844 28018 18900 28030
rect 19068 28532 19124 28542
rect 18620 27806 18622 27858
rect 18674 27806 18676 27858
rect 18620 26964 18676 27806
rect 19068 27858 19124 28476
rect 19404 28196 19460 28588
rect 19516 28642 19572 28654
rect 19516 28590 19518 28642
rect 19570 28590 19572 28642
rect 19516 28420 19572 28590
rect 19740 28530 19796 28812
rect 20188 28642 20244 30828
rect 20300 30818 20356 30828
rect 20748 30212 20804 30222
rect 20748 30118 20804 30156
rect 20188 28590 20190 28642
rect 20242 28590 20244 28642
rect 19740 28478 19742 28530
rect 19794 28478 19796 28530
rect 19740 28466 19796 28478
rect 19964 28532 20020 28542
rect 19964 28438 20020 28476
rect 19516 28354 19572 28364
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19404 28140 19684 28196
rect 19836 28186 20100 28196
rect 19068 27806 19070 27858
rect 19122 27806 19124 27858
rect 18956 27748 19012 27758
rect 18956 27654 19012 27692
rect 19068 27524 19124 27806
rect 18620 26628 18676 26908
rect 18732 27468 19124 27524
rect 19180 27858 19236 27870
rect 19180 27806 19182 27858
rect 19234 27806 19236 27858
rect 18732 27076 18788 27468
rect 18844 27188 18900 27198
rect 19180 27188 19236 27806
rect 18844 27186 19236 27188
rect 18844 27134 18846 27186
rect 18898 27134 19236 27186
rect 18844 27132 19236 27134
rect 18844 27122 18900 27132
rect 18732 26908 18788 27020
rect 19180 26964 19236 27132
rect 19628 27186 19684 28140
rect 20188 28084 20244 28590
rect 20076 28028 20244 28084
rect 20300 29314 20356 29326
rect 20300 29262 20302 29314
rect 20354 29262 20356 29314
rect 20300 28532 20356 29262
rect 20636 28868 20692 28878
rect 20636 28754 20692 28812
rect 20636 28702 20638 28754
rect 20690 28702 20692 28754
rect 20636 28690 20692 28702
rect 20076 27858 20132 28028
rect 20076 27806 20078 27858
rect 20130 27806 20132 27858
rect 20076 27794 20132 27806
rect 20300 27858 20356 28476
rect 20300 27806 20302 27858
rect 20354 27806 20356 27858
rect 20300 27794 20356 27806
rect 20412 27860 20468 27870
rect 19628 27134 19630 27186
rect 19682 27134 19684 27186
rect 19628 27122 19684 27134
rect 20412 27188 20468 27804
rect 20412 27094 20468 27132
rect 20636 27746 20692 27758
rect 20636 27694 20638 27746
rect 20690 27694 20692 27746
rect 19852 26964 19908 26974
rect 19180 26962 19908 26964
rect 19180 26910 19854 26962
rect 19906 26910 19908 26962
rect 19180 26908 19908 26910
rect 18732 26852 19124 26908
rect 19852 26898 19908 26908
rect 18620 26562 18676 26572
rect 19068 26516 19124 26852
rect 19964 26852 20020 26862
rect 19964 26758 20020 26796
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19068 26450 19124 26460
rect 18620 26292 18676 26302
rect 18620 26198 18676 26236
rect 19068 26290 19124 26302
rect 19068 26238 19070 26290
rect 19122 26238 19124 26290
rect 19068 26180 19124 26238
rect 19628 26290 19684 26302
rect 19628 26238 19630 26290
rect 19682 26238 19684 26290
rect 19068 26114 19124 26124
rect 19404 26178 19460 26190
rect 19404 26126 19406 26178
rect 19458 26126 19460 26178
rect 19404 23716 19460 26126
rect 19516 26066 19572 26078
rect 19516 26014 19518 26066
rect 19570 26014 19572 26066
rect 19516 24836 19572 26014
rect 19516 24770 19572 24780
rect 19516 24612 19572 24622
rect 19516 24518 19572 24556
rect 19628 24500 19684 26238
rect 20636 26290 20692 27694
rect 20636 26238 20638 26290
rect 20690 26238 20692 26290
rect 20300 25620 20356 25630
rect 20636 25620 20692 26238
rect 20748 27634 20804 27646
rect 20748 27582 20750 27634
rect 20802 27582 20804 27634
rect 20748 26292 20804 27582
rect 20860 27300 20916 33628
rect 20972 31892 21028 40124
rect 21196 40114 21252 40124
rect 21308 39618 21364 41020
rect 21308 39566 21310 39618
rect 21362 39566 21364 39618
rect 21084 39508 21140 39518
rect 21084 38500 21140 39452
rect 21308 39284 21364 39566
rect 21420 40740 21476 40750
rect 21420 39506 21476 40684
rect 21532 40628 21588 43708
rect 21644 43538 21700 43550
rect 21644 43486 21646 43538
rect 21698 43486 21700 43538
rect 21644 42980 21700 43486
rect 21980 43538 22036 45166
rect 22428 45108 22484 45118
rect 21980 43486 21982 43538
rect 22034 43486 22036 43538
rect 21980 43474 22036 43486
rect 22316 45106 22484 45108
rect 22316 45054 22430 45106
rect 22482 45054 22484 45106
rect 22316 45052 22484 45054
rect 21644 42914 21700 42924
rect 22316 43316 22372 45052
rect 22428 45042 22484 45052
rect 23212 45108 23268 45118
rect 23212 44548 23268 45052
rect 22764 44492 23268 44548
rect 22204 42868 22260 42878
rect 21644 42642 21700 42654
rect 21644 42590 21646 42642
rect 21698 42590 21700 42642
rect 21644 41300 21700 42590
rect 22092 42644 22148 42654
rect 21756 41300 21812 41310
rect 21644 41298 21812 41300
rect 21644 41246 21758 41298
rect 21810 41246 21812 41298
rect 21644 41244 21812 41246
rect 21756 41076 21812 41244
rect 21756 41010 21812 41020
rect 21532 40572 21700 40628
rect 21420 39454 21422 39506
rect 21474 39454 21476 39506
rect 21420 39442 21476 39454
rect 21532 40404 21588 40414
rect 21308 39228 21476 39284
rect 21308 38836 21364 38846
rect 21308 38742 21364 38780
rect 21196 38724 21252 38734
rect 21196 38612 21364 38668
rect 21084 38434 21140 38444
rect 21308 37940 21364 38612
rect 21420 38500 21476 39228
rect 21420 38434 21476 38444
rect 21420 38276 21476 38286
rect 21532 38276 21588 40348
rect 21644 40180 21700 40572
rect 21644 40114 21700 40124
rect 21756 40514 21812 40526
rect 21756 40462 21758 40514
rect 21810 40462 21812 40514
rect 21756 39172 21812 40462
rect 22092 39620 22148 42588
rect 22204 41970 22260 42812
rect 22316 42754 22372 43260
rect 22316 42702 22318 42754
rect 22370 42702 22372 42754
rect 22316 42690 22372 42702
rect 22540 44436 22596 44446
rect 22204 41918 22206 41970
rect 22258 41918 22260 41970
rect 22204 41906 22260 41918
rect 22540 41860 22596 44380
rect 22652 43538 22708 43550
rect 22652 43486 22654 43538
rect 22706 43486 22708 43538
rect 22652 42978 22708 43486
rect 22652 42926 22654 42978
rect 22706 42926 22708 42978
rect 22652 42914 22708 42926
rect 22764 42754 22820 44492
rect 23884 43650 23940 45948
rect 24556 46002 25172 46004
rect 24556 45950 24558 46002
rect 24610 45950 25172 46002
rect 24556 45948 25172 45950
rect 24556 45938 24612 45948
rect 24668 45780 24724 45790
rect 24668 45330 24724 45724
rect 24668 45278 24670 45330
rect 24722 45278 24724 45330
rect 24668 45266 24724 45278
rect 24556 44996 24612 45006
rect 24556 44902 24612 44940
rect 24556 44212 24612 44222
rect 23884 43598 23886 43650
rect 23938 43598 23940 43650
rect 22764 42702 22766 42754
rect 22818 42702 22820 42754
rect 22764 42690 22820 42702
rect 23212 43426 23268 43438
rect 23212 43374 23214 43426
rect 23266 43374 23268 43426
rect 22652 41860 22708 41870
rect 22540 41858 22708 41860
rect 22540 41806 22654 41858
rect 22706 41806 22708 41858
rect 22540 41804 22708 41806
rect 22652 41794 22708 41804
rect 22764 41300 22820 41310
rect 22764 40740 22820 41244
rect 22652 40516 22708 40526
rect 22428 40514 22708 40516
rect 22428 40462 22654 40514
rect 22706 40462 22708 40514
rect 22428 40460 22708 40462
rect 22204 39620 22260 39630
rect 22092 39618 22260 39620
rect 22092 39566 22206 39618
rect 22258 39566 22260 39618
rect 22092 39564 22260 39566
rect 22204 39554 22260 39564
rect 22428 39394 22484 40460
rect 22652 40450 22708 40460
rect 22428 39342 22430 39394
rect 22482 39342 22484 39394
rect 22428 39330 22484 39342
rect 22652 39396 22708 39406
rect 22764 39396 22820 40684
rect 23212 40402 23268 43374
rect 23548 43092 23604 43102
rect 23548 42754 23604 43036
rect 23884 42868 23940 43598
rect 24332 43652 24388 43662
rect 24332 43558 24388 43596
rect 23884 42802 23940 42812
rect 24108 43538 24164 43550
rect 24108 43486 24110 43538
rect 24162 43486 24164 43538
rect 24108 43204 24164 43486
rect 24444 43538 24500 43550
rect 24444 43486 24446 43538
rect 24498 43486 24500 43538
rect 24220 43428 24276 43438
rect 24444 43428 24500 43486
rect 24220 43334 24276 43372
rect 24332 43372 24500 43428
rect 24332 43316 24388 43372
rect 24556 43316 24612 44156
rect 25116 43652 25172 45948
rect 27468 45892 27524 45902
rect 28364 45892 28420 45902
rect 32172 45892 32228 45902
rect 27468 45890 28420 45892
rect 27468 45838 27470 45890
rect 27522 45838 28366 45890
rect 28418 45838 28420 45890
rect 27468 45836 28420 45838
rect 26684 45778 26740 45790
rect 26684 45726 26686 45778
rect 26738 45726 26740 45778
rect 25228 45108 25284 45118
rect 25228 45014 25284 45052
rect 25452 45106 25508 45118
rect 25452 45054 25454 45106
rect 25506 45054 25508 45106
rect 25228 43652 25284 43662
rect 24332 43250 24388 43260
rect 24444 43260 24612 43316
rect 24668 43650 25284 43652
rect 24668 43598 25230 43650
rect 25282 43598 25284 43650
rect 24668 43596 25284 43598
rect 23548 42702 23550 42754
rect 23602 42702 23604 42754
rect 23548 42644 23604 42702
rect 23996 42756 24052 42766
rect 23996 42662 24052 42700
rect 23548 42578 23604 42588
rect 24108 42420 24164 43148
rect 24108 42364 24276 42420
rect 24108 41858 24164 41870
rect 24108 41806 24110 41858
rect 24162 41806 24164 41858
rect 23996 41746 24052 41758
rect 23996 41694 23998 41746
rect 24050 41694 24052 41746
rect 23884 41300 23940 41310
rect 23996 41300 24052 41694
rect 23884 41298 24052 41300
rect 23884 41246 23886 41298
rect 23938 41246 24052 41298
rect 23884 41244 24052 41246
rect 23884 41234 23940 41244
rect 23996 41076 24052 41086
rect 23996 40514 24052 41020
rect 23996 40462 23998 40514
rect 24050 40462 24052 40514
rect 23996 40450 24052 40462
rect 23212 40350 23214 40402
rect 23266 40350 23268 40402
rect 23212 40338 23268 40350
rect 24108 40180 24164 41806
rect 24220 40404 24276 42364
rect 24444 41188 24500 43260
rect 24556 42980 24612 42990
rect 24556 42886 24612 42924
rect 24668 42756 24724 43596
rect 25228 43586 25284 43596
rect 25452 43538 25508 45054
rect 25676 45108 25732 45118
rect 25676 45014 25732 45052
rect 25788 45106 25844 45118
rect 25788 45054 25790 45106
rect 25842 45054 25844 45106
rect 25564 44996 25620 45006
rect 25564 44902 25620 44940
rect 25788 43762 25844 45054
rect 26348 45108 26404 45118
rect 26348 45014 26404 45052
rect 25788 43710 25790 43762
rect 25842 43710 25844 43762
rect 25452 43486 25454 43538
rect 25506 43486 25508 43538
rect 24668 42662 24724 42700
rect 24780 43316 24836 43326
rect 24556 42644 24612 42654
rect 24556 42550 24612 42588
rect 24668 42196 24724 42206
rect 24556 42084 24612 42094
rect 24556 41970 24612 42028
rect 24556 41918 24558 41970
rect 24610 41918 24612 41970
rect 24556 41906 24612 41918
rect 24668 41970 24724 42140
rect 24668 41918 24670 41970
rect 24722 41918 24724 41970
rect 24668 41906 24724 41918
rect 24556 41188 24612 41198
rect 24444 41186 24612 41188
rect 24444 41134 24558 41186
rect 24610 41134 24612 41186
rect 24444 41132 24612 41134
rect 24556 41122 24612 41132
rect 24444 40628 24500 40638
rect 24444 40534 24500 40572
rect 24780 40516 24836 43260
rect 25452 43204 25508 43486
rect 25676 43540 25732 43550
rect 25676 43446 25732 43484
rect 25452 43138 25508 43148
rect 25564 43426 25620 43438
rect 25564 43374 25566 43426
rect 25618 43374 25620 43426
rect 24892 42868 24948 42878
rect 25116 42868 25172 42878
rect 24948 42866 25172 42868
rect 24948 42814 25118 42866
rect 25170 42814 25172 42866
rect 24948 42812 25172 42814
rect 24892 42802 24948 42812
rect 25116 42802 25172 42812
rect 25004 42532 25060 42542
rect 25004 42438 25060 42476
rect 25564 42084 25620 43374
rect 25788 43316 25844 43710
rect 26572 44322 26628 44334
rect 26572 44270 26574 44322
rect 26626 44270 26628 44322
rect 26348 43540 26404 43550
rect 26348 43446 26404 43484
rect 25788 43250 25844 43260
rect 25564 42018 25620 42028
rect 25788 42754 25844 42766
rect 25788 42702 25790 42754
rect 25842 42702 25844 42754
rect 25788 41972 25844 42702
rect 26460 42644 26516 42654
rect 26460 42550 26516 42588
rect 25452 41858 25508 41870
rect 25452 41806 25454 41858
rect 25506 41806 25508 41858
rect 25228 40964 25284 40974
rect 25228 40962 25396 40964
rect 25228 40910 25230 40962
rect 25282 40910 25396 40962
rect 25228 40908 25396 40910
rect 25228 40898 25284 40908
rect 24220 40310 24276 40348
rect 24668 40404 24724 40414
rect 24780 40404 24836 40460
rect 24668 40402 24836 40404
rect 24668 40350 24670 40402
rect 24722 40350 24836 40402
rect 24668 40348 24836 40350
rect 25228 40402 25284 40414
rect 25228 40350 25230 40402
rect 25282 40350 25284 40402
rect 24668 40338 24724 40348
rect 24332 40290 24388 40302
rect 24332 40238 24334 40290
rect 24386 40238 24388 40290
rect 24332 40180 24388 40238
rect 24108 40124 24388 40180
rect 22652 39394 22820 39396
rect 22652 39342 22654 39394
rect 22706 39342 22820 39394
rect 22652 39340 22820 39342
rect 23100 39618 23156 39630
rect 23100 39566 23102 39618
rect 23154 39566 23156 39618
rect 22652 39330 22708 39340
rect 21756 39106 21812 39116
rect 22540 39172 22596 39182
rect 22316 39060 22372 39070
rect 22204 38836 22260 38846
rect 21756 38612 21812 38622
rect 21420 38274 21588 38276
rect 21420 38222 21422 38274
rect 21474 38222 21588 38274
rect 21420 38220 21588 38222
rect 21644 38610 21812 38612
rect 21644 38558 21758 38610
rect 21810 38558 21812 38610
rect 21644 38556 21812 38558
rect 21420 38210 21476 38220
rect 21532 38052 21588 38062
rect 21644 38052 21700 38556
rect 21756 38546 21812 38556
rect 22204 38274 22260 38780
rect 22204 38222 22206 38274
rect 22258 38222 22260 38274
rect 22204 38210 22260 38222
rect 21532 38050 21700 38052
rect 21532 37998 21534 38050
rect 21586 37998 21700 38050
rect 21532 37996 21700 37998
rect 21532 37986 21588 37996
rect 21420 37940 21476 37950
rect 20972 27636 21028 31836
rect 21196 37938 21476 37940
rect 21196 37886 21422 37938
rect 21474 37886 21476 37938
rect 21196 37884 21476 37886
rect 21196 31220 21252 37884
rect 21420 37874 21476 37884
rect 21644 37044 21700 37996
rect 22092 37940 22148 37950
rect 21644 36978 21700 36988
rect 21868 37938 22148 37940
rect 21868 37886 22094 37938
rect 22146 37886 22148 37938
rect 21868 37884 22148 37886
rect 21868 37156 21924 37884
rect 22092 37874 22148 37884
rect 22204 37940 22260 37950
rect 22316 37940 22372 39004
rect 22540 38834 22596 39116
rect 22540 38782 22542 38834
rect 22594 38782 22596 38834
rect 22540 38770 22596 38782
rect 23100 38668 23156 39566
rect 23884 39506 23940 39518
rect 23884 39454 23886 39506
rect 23938 39454 23940 39506
rect 23212 38836 23268 38846
rect 23212 38742 23268 38780
rect 23884 38668 23940 39454
rect 24444 39060 24500 39070
rect 24444 38834 24500 39004
rect 24444 38782 24446 38834
rect 24498 38782 24500 38834
rect 24444 38770 24500 38782
rect 22204 37938 22372 37940
rect 22204 37886 22206 37938
rect 22258 37886 22372 37938
rect 22204 37884 22372 37886
rect 22988 38612 23156 38668
rect 23660 38612 23940 38668
rect 23996 38724 24052 38734
rect 22988 37938 23044 38612
rect 22988 37886 22990 37938
rect 23042 37886 23044 37938
rect 22204 37874 22260 37884
rect 22988 37266 23044 37886
rect 23660 37490 23716 38612
rect 23660 37438 23662 37490
rect 23714 37438 23716 37490
rect 23660 37426 23716 37438
rect 23884 37380 23940 37390
rect 23884 37286 23940 37324
rect 23996 37378 24052 38668
rect 23996 37326 23998 37378
rect 24050 37326 24052 37378
rect 23996 37314 24052 37326
rect 24780 38052 24836 38062
rect 22988 37214 22990 37266
rect 23042 37214 23044 37266
rect 21532 36484 21588 36494
rect 21532 36390 21588 36428
rect 21644 36258 21700 36270
rect 21644 36206 21646 36258
rect 21698 36206 21700 36258
rect 21308 35812 21364 35822
rect 21644 35812 21700 36206
rect 21308 35810 21700 35812
rect 21308 35758 21310 35810
rect 21362 35758 21700 35810
rect 21308 35756 21700 35758
rect 21756 36258 21812 36270
rect 21756 36206 21758 36258
rect 21810 36206 21812 36258
rect 21308 35746 21364 35756
rect 21756 35588 21812 36206
rect 21756 35522 21812 35532
rect 21532 35252 21588 35262
rect 21308 34018 21364 34030
rect 21308 33966 21310 34018
rect 21362 33966 21364 34018
rect 21308 33460 21364 33966
rect 21308 33394 21364 33404
rect 21532 33346 21588 35196
rect 21868 34916 21924 37100
rect 22204 37156 22260 37166
rect 22204 37154 22708 37156
rect 22204 37102 22206 37154
rect 22258 37102 22708 37154
rect 22204 37100 22708 37102
rect 22204 37090 22260 37100
rect 22540 36932 22596 36942
rect 22540 36484 22596 36876
rect 22092 36482 22596 36484
rect 22092 36430 22542 36482
rect 22594 36430 22596 36482
rect 22092 36428 22596 36430
rect 21980 36258 22036 36270
rect 21980 36206 21982 36258
rect 22034 36206 22036 36258
rect 21980 35140 22036 36206
rect 22092 35698 22148 36428
rect 22540 36418 22596 36428
rect 22652 35922 22708 37100
rect 22764 37044 22820 37054
rect 22988 37044 23044 37214
rect 23548 37156 23604 37166
rect 23548 37154 24052 37156
rect 23548 37102 23550 37154
rect 23602 37102 24052 37154
rect 23548 37100 24052 37102
rect 23548 37090 23604 37100
rect 22820 36988 22932 37044
rect 22764 36978 22820 36988
rect 22652 35870 22654 35922
rect 22706 35870 22708 35922
rect 22652 35858 22708 35870
rect 22540 35700 22596 35710
rect 22092 35646 22094 35698
rect 22146 35646 22148 35698
rect 22092 35634 22148 35646
rect 22428 35698 22596 35700
rect 22428 35646 22542 35698
rect 22594 35646 22596 35698
rect 22428 35644 22596 35646
rect 21980 35074 22036 35084
rect 22316 35588 22372 35598
rect 22204 35028 22260 35038
rect 22092 34916 22148 34926
rect 21868 34914 22148 34916
rect 21868 34862 22094 34914
rect 22146 34862 22148 34914
rect 21868 34860 22148 34862
rect 22092 34850 22148 34860
rect 22204 34802 22260 34972
rect 22204 34750 22206 34802
rect 22258 34750 22260 34802
rect 22204 34738 22260 34750
rect 21868 34690 21924 34702
rect 21868 34638 21870 34690
rect 21922 34638 21924 34690
rect 21868 33572 21924 34638
rect 21868 33506 21924 33516
rect 21980 34692 22036 34702
rect 21532 33294 21534 33346
rect 21586 33294 21588 33346
rect 21532 33282 21588 33294
rect 21308 33236 21364 33246
rect 21308 33142 21364 33180
rect 21420 31892 21476 31902
rect 21308 31668 21364 31678
rect 21308 31574 21364 31612
rect 21196 31154 21252 31164
rect 21420 31332 21476 31836
rect 21644 31668 21700 31678
rect 21644 31574 21700 31612
rect 21420 31218 21476 31276
rect 21420 31166 21422 31218
rect 21474 31166 21476 31218
rect 21420 31154 21476 31166
rect 21868 31220 21924 31230
rect 21868 30994 21924 31164
rect 21868 30942 21870 30994
rect 21922 30942 21924 30994
rect 21868 30930 21924 30942
rect 21308 30212 21364 30222
rect 21308 29988 21364 30156
rect 21420 29988 21476 29998
rect 21308 29986 21476 29988
rect 21308 29934 21422 29986
rect 21474 29934 21476 29986
rect 21308 29932 21476 29934
rect 21308 28308 21364 29932
rect 21420 29922 21476 29932
rect 21532 29316 21588 29326
rect 21420 28756 21476 28766
rect 21420 28530 21476 28700
rect 21532 28754 21588 29260
rect 21532 28702 21534 28754
rect 21586 28702 21588 28754
rect 21532 28690 21588 28702
rect 21420 28478 21422 28530
rect 21474 28478 21476 28530
rect 21420 28466 21476 28478
rect 21644 28532 21700 28542
rect 21644 28438 21700 28476
rect 21308 28252 21588 28308
rect 21084 27860 21140 27870
rect 21420 27860 21476 27870
rect 21084 27858 21420 27860
rect 21084 27806 21086 27858
rect 21138 27806 21420 27858
rect 21084 27804 21420 27806
rect 21084 27794 21140 27804
rect 20972 27580 21252 27636
rect 20972 27300 21028 27310
rect 20860 27244 20972 27300
rect 20972 27234 21028 27244
rect 21084 27188 21140 27198
rect 21084 26404 21140 27132
rect 21196 26964 21252 27580
rect 21308 27186 21364 27804
rect 21420 27794 21476 27804
rect 21532 27636 21588 28252
rect 21756 27860 21812 27870
rect 21756 27766 21812 27804
rect 21532 27580 21812 27636
rect 21308 27134 21310 27186
rect 21362 27134 21364 27186
rect 21308 27122 21364 27134
rect 21532 27020 21700 27076
rect 21532 26964 21588 27020
rect 21196 26908 21588 26964
rect 21420 26404 21476 26414
rect 21084 26402 21476 26404
rect 21084 26350 21422 26402
rect 21474 26350 21476 26402
rect 21084 26348 21476 26350
rect 20748 26226 20804 26236
rect 20300 25618 20692 25620
rect 20300 25566 20302 25618
rect 20354 25566 20638 25618
rect 20690 25566 20692 25618
rect 20300 25564 20692 25566
rect 20300 25554 20356 25564
rect 20636 25554 20692 25564
rect 20188 25508 20244 25518
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20188 24722 20244 25452
rect 20748 25284 20804 25294
rect 20748 25282 21364 25284
rect 20748 25230 20750 25282
rect 20802 25230 21364 25282
rect 20748 25228 21364 25230
rect 20748 25218 20804 25228
rect 20188 24670 20190 24722
rect 20242 24670 20244 24722
rect 20188 24658 20244 24670
rect 20300 24836 20356 24846
rect 19740 24500 19796 24510
rect 19628 24444 19740 24500
rect 19740 24434 19796 24444
rect 19740 24050 19796 24062
rect 19740 23998 19742 24050
rect 19794 23998 19796 24050
rect 19740 23716 19796 23998
rect 19068 23660 19796 23716
rect 20188 23714 20244 23726
rect 20188 23662 20190 23714
rect 20242 23662 20244 23714
rect 18620 23268 18676 23278
rect 18620 23174 18676 23212
rect 18956 23156 19012 23166
rect 19068 23156 19124 23660
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 18956 23154 19124 23156
rect 18956 23102 18958 23154
rect 19010 23102 19124 23154
rect 18956 23100 19124 23102
rect 18956 20692 19012 23100
rect 19964 22260 20020 22270
rect 19964 22166 20020 22204
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20188 21812 20244 23662
rect 20300 23154 20356 24780
rect 20748 24612 20804 24622
rect 20636 24610 20804 24612
rect 20636 24558 20750 24610
rect 20802 24558 20804 24610
rect 20636 24556 20804 24558
rect 20636 24500 20692 24556
rect 20748 24546 20804 24556
rect 20300 23102 20302 23154
rect 20354 23102 20356 23154
rect 20300 23090 20356 23102
rect 20412 23826 20468 23838
rect 20412 23774 20414 23826
rect 20466 23774 20468 23826
rect 20412 23268 20468 23774
rect 20412 22484 20468 23212
rect 20412 22418 20468 22428
rect 20524 23266 20580 23278
rect 20524 23214 20526 23266
rect 20578 23214 20580 23266
rect 19852 21756 20244 21812
rect 19852 21700 19908 21756
rect 19740 21140 19796 21150
rect 19292 21028 19348 21038
rect 19292 20934 19348 20972
rect 18956 20626 19012 20636
rect 19740 20690 19796 21084
rect 19740 20638 19742 20690
rect 19794 20638 19796 20690
rect 19740 20580 19796 20638
rect 19628 20524 19740 20580
rect 19852 20690 19908 21644
rect 19964 21588 20020 21598
rect 19964 20804 20020 21532
rect 19964 20802 20356 20804
rect 19964 20750 19966 20802
rect 20018 20750 20356 20802
rect 19964 20748 20356 20750
rect 19964 20738 20020 20748
rect 19852 20638 19854 20690
rect 19906 20638 19908 20690
rect 19852 20580 19908 20638
rect 19852 20524 20244 20580
rect 18844 20020 18900 20030
rect 18844 19926 18900 19964
rect 18508 18610 18564 18620
rect 17836 18452 17892 18462
rect 18620 18452 18676 18462
rect 17836 18358 17892 18396
rect 18508 18450 18676 18452
rect 18508 18398 18622 18450
rect 18674 18398 18676 18450
rect 18508 18396 18676 18398
rect 18284 18226 18340 18238
rect 18284 18174 18286 18226
rect 18338 18174 18340 18226
rect 18172 17442 18228 17454
rect 18172 17390 18174 17442
rect 18226 17390 18228 17442
rect 18060 16884 18116 16894
rect 18172 16884 18228 17390
rect 18116 16828 18228 16884
rect 18060 16436 18116 16828
rect 18284 16548 18340 18174
rect 18396 16884 18452 16894
rect 18508 16884 18564 18396
rect 18620 18386 18676 18396
rect 18452 16828 18564 16884
rect 18620 18228 18676 18238
rect 18620 17442 18676 18172
rect 19628 17780 19684 20524
rect 19740 20514 19796 20524
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20188 20244 20244 20524
rect 20076 20188 20244 20244
rect 20076 19012 20132 20188
rect 20300 19346 20356 20748
rect 20300 19294 20302 19346
rect 20354 19294 20356 19346
rect 20300 19282 20356 19294
rect 20076 18956 20244 19012
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19964 18452 20020 18462
rect 19964 18338 20020 18396
rect 19964 18286 19966 18338
rect 20018 18286 20020 18338
rect 19964 18274 20020 18286
rect 20076 18450 20132 18462
rect 20076 18398 20078 18450
rect 20130 18398 20132 18450
rect 19292 17724 19684 17780
rect 19068 17668 19124 17678
rect 19068 17574 19124 17612
rect 18620 17390 18622 17442
rect 18674 17390 18676 17442
rect 18620 16882 18676 17390
rect 18620 16830 18622 16882
rect 18674 16830 18676 16882
rect 18396 16790 18452 16828
rect 18620 16818 18676 16830
rect 18284 16482 18340 16492
rect 19068 16660 19124 16670
rect 18060 16370 18116 16380
rect 18396 16212 18452 16222
rect 18172 16100 18228 16110
rect 18172 16006 18228 16044
rect 18396 16098 18452 16156
rect 18396 16046 18398 16098
rect 18450 16046 18452 16098
rect 18396 16034 18452 16046
rect 19068 16100 19124 16604
rect 19068 16034 19124 16044
rect 19292 16100 19348 17724
rect 19628 17666 19684 17724
rect 19628 17614 19630 17666
rect 19682 17614 19684 17666
rect 19628 17602 19684 17614
rect 19964 17556 20020 17566
rect 19964 17462 20020 17500
rect 19628 17442 19684 17454
rect 19628 17390 19630 17442
rect 19682 17390 19684 17442
rect 19628 16884 19684 17390
rect 20076 17444 20132 18398
rect 20188 17556 20244 18956
rect 20524 17668 20580 23214
rect 20636 20914 20692 24444
rect 21308 24162 21364 25228
rect 21308 24110 21310 24162
rect 21362 24110 21364 24162
rect 21308 24098 21364 24110
rect 20748 23940 20804 23950
rect 21420 23940 21476 26348
rect 21532 25732 21588 25742
rect 21532 24050 21588 25676
rect 21532 23998 21534 24050
rect 21586 23998 21588 24050
rect 21532 23986 21588 23998
rect 20748 23938 21476 23940
rect 20748 23886 20750 23938
rect 20802 23886 21476 23938
rect 20748 23884 21476 23886
rect 20748 23380 20804 23884
rect 21644 23828 21700 27020
rect 21756 25284 21812 27580
rect 21868 27634 21924 27646
rect 21868 27582 21870 27634
rect 21922 27582 21924 27634
rect 21868 26404 21924 27582
rect 21980 26908 22036 34636
rect 22316 33348 22372 35532
rect 22428 34914 22484 35644
rect 22540 35634 22596 35644
rect 22764 35698 22820 35710
rect 22764 35646 22766 35698
rect 22818 35646 22820 35698
rect 22764 35588 22820 35646
rect 22764 35522 22820 35532
rect 22428 34862 22430 34914
rect 22482 34862 22484 34914
rect 22428 34850 22484 34862
rect 22876 34244 22932 36988
rect 22988 36978 23044 36988
rect 23212 36372 23268 36382
rect 23212 36278 23268 36316
rect 23996 35924 24052 37100
rect 24668 37154 24724 37166
rect 24668 37102 24670 37154
rect 24722 37102 24724 37154
rect 23996 35830 24052 35868
rect 24556 36484 24612 36494
rect 24668 36484 24724 37102
rect 24612 36428 24724 36484
rect 24556 35922 24612 36428
rect 24780 35924 24836 37996
rect 24556 35870 24558 35922
rect 24610 35870 24612 35922
rect 24556 35858 24612 35870
rect 24668 35868 24836 35924
rect 25228 35924 25284 40350
rect 25340 39060 25396 40908
rect 25452 40628 25508 41806
rect 25788 41186 25844 41916
rect 26124 41972 26180 41982
rect 26460 41972 26516 41982
rect 26124 41970 26516 41972
rect 26124 41918 26126 41970
rect 26178 41918 26462 41970
rect 26514 41918 26516 41970
rect 26124 41916 26516 41918
rect 26124 41906 26180 41916
rect 26348 41746 26404 41758
rect 26348 41694 26350 41746
rect 26402 41694 26404 41746
rect 26348 41300 26404 41694
rect 26460 41636 26516 41916
rect 26460 41570 26516 41580
rect 26460 41300 26516 41310
rect 26348 41298 26516 41300
rect 26348 41246 26462 41298
rect 26514 41246 26516 41298
rect 26348 41244 26516 41246
rect 26460 41234 26516 41244
rect 25788 41134 25790 41186
rect 25842 41134 25844 41186
rect 25788 41122 25844 41134
rect 25452 40562 25508 40572
rect 25900 40740 25956 40750
rect 25900 40626 25956 40684
rect 25900 40574 25902 40626
rect 25954 40574 25956 40626
rect 25900 40562 25956 40574
rect 25564 40516 25620 40526
rect 25564 40422 25620 40460
rect 26012 40402 26068 40414
rect 26012 40350 26014 40402
rect 26066 40350 26068 40402
rect 26012 39956 26068 40350
rect 25340 38994 25396 39004
rect 25900 39900 26068 39956
rect 26124 40404 26180 40414
rect 25340 38724 25396 38762
rect 25340 38658 25396 38668
rect 25676 38500 25732 38510
rect 25676 37492 25732 38444
rect 25676 37490 25844 37492
rect 25676 37438 25678 37490
rect 25730 37438 25844 37490
rect 25676 37436 25844 37438
rect 25676 37426 25732 37436
rect 25564 37268 25620 37278
rect 25340 37266 25620 37268
rect 25340 37214 25566 37266
rect 25618 37214 25620 37266
rect 25340 37212 25620 37214
rect 25340 36594 25396 37212
rect 25564 37202 25620 37212
rect 25340 36542 25342 36594
rect 25394 36542 25396 36594
rect 25340 36530 25396 36542
rect 25676 36596 25732 36606
rect 25676 36502 25732 36540
rect 25564 36372 25620 36382
rect 25228 35868 25508 35924
rect 23212 35700 23268 35710
rect 23212 35606 23268 35644
rect 23772 35700 23828 35710
rect 23772 35606 23828 35644
rect 24108 35700 24164 35710
rect 24444 35700 24500 35710
rect 24108 35698 24500 35700
rect 24108 35646 24110 35698
rect 24162 35646 24446 35698
rect 24498 35646 24500 35698
rect 24108 35644 24500 35646
rect 24108 35634 24164 35644
rect 23660 35586 23716 35598
rect 23660 35534 23662 35586
rect 23714 35534 23716 35586
rect 23660 35476 23716 35534
rect 23660 35420 24164 35476
rect 23548 35252 23604 35262
rect 23548 35026 23604 35196
rect 23772 35252 23828 35262
rect 23772 35140 23828 35196
rect 23772 35138 23940 35140
rect 23772 35086 23774 35138
rect 23826 35086 23940 35138
rect 23772 35084 23940 35086
rect 23772 35074 23828 35084
rect 23548 34974 23550 35026
rect 23602 34974 23604 35026
rect 23548 34962 23604 34974
rect 23436 34914 23492 34926
rect 23436 34862 23438 34914
rect 23490 34862 23492 34914
rect 23212 34690 23268 34702
rect 23212 34638 23214 34690
rect 23266 34638 23268 34690
rect 23100 34356 23156 34366
rect 22764 34188 22932 34244
rect 22988 34300 23100 34356
rect 22540 33572 22596 33582
rect 22428 33460 22484 33470
rect 22428 33366 22484 33404
rect 22316 33254 22372 33292
rect 22540 33346 22596 33516
rect 22540 33294 22542 33346
rect 22594 33294 22596 33346
rect 22540 33282 22596 33294
rect 22652 32676 22708 32686
rect 22092 31780 22148 31790
rect 22092 31686 22148 31724
rect 22652 31332 22708 32620
rect 22540 31220 22596 31230
rect 22316 30882 22372 30894
rect 22316 30830 22318 30882
rect 22370 30830 22372 30882
rect 22316 30772 22372 30830
rect 22316 30706 22372 30716
rect 22540 30322 22596 31164
rect 22652 31218 22708 31276
rect 22652 31166 22654 31218
rect 22706 31166 22708 31218
rect 22652 31154 22708 31166
rect 22540 30270 22542 30322
rect 22594 30270 22596 30322
rect 22540 30258 22596 30270
rect 22428 29316 22484 29326
rect 22428 29222 22484 29260
rect 22428 28756 22484 28766
rect 22092 28754 22484 28756
rect 22092 28702 22430 28754
rect 22482 28702 22484 28754
rect 22092 28700 22484 28702
rect 22092 28642 22148 28700
rect 22428 28690 22484 28700
rect 22764 28756 22820 34188
rect 22876 33348 22932 33358
rect 22988 33348 23044 34300
rect 23100 34290 23156 34300
rect 23212 33796 23268 34638
rect 23436 34692 23492 34862
rect 23436 34626 23492 34636
rect 23772 34244 23828 34254
rect 23436 34188 23772 34244
rect 23436 34018 23492 34188
rect 23772 34150 23828 34188
rect 23884 34020 23940 35084
rect 23996 34356 24052 34366
rect 23996 34262 24052 34300
rect 24108 34242 24164 35420
rect 24220 35308 24276 35644
rect 24444 35634 24500 35644
rect 24220 35252 24612 35308
rect 24220 34802 24276 34814
rect 24556 34804 24612 35252
rect 24668 35028 24724 35868
rect 24780 35700 24836 35710
rect 25228 35700 25284 35710
rect 24780 35698 25284 35700
rect 24780 35646 24782 35698
rect 24834 35646 25230 35698
rect 25282 35646 25284 35698
rect 24780 35644 25284 35646
rect 24780 35634 24836 35644
rect 25228 35634 25284 35644
rect 25340 35700 25396 35710
rect 25004 35140 25060 35150
rect 25004 35046 25060 35084
rect 24668 34962 24724 34972
rect 25340 34916 25396 35644
rect 25452 35252 25508 35868
rect 25564 35810 25620 36316
rect 25564 35758 25566 35810
rect 25618 35758 25620 35810
rect 25564 35746 25620 35758
rect 25788 35698 25844 37436
rect 25788 35646 25790 35698
rect 25842 35646 25844 35698
rect 25788 35634 25844 35646
rect 25452 35186 25508 35196
rect 25116 34860 25396 34916
rect 24892 34804 24948 34814
rect 24220 34750 24222 34802
rect 24274 34750 24276 34802
rect 24220 34692 24276 34750
rect 24220 34626 24276 34636
rect 24444 34802 24948 34804
rect 24444 34750 24558 34802
rect 24610 34750 24894 34802
rect 24946 34750 24948 34802
rect 24444 34748 24948 34750
rect 24108 34190 24110 34242
rect 24162 34190 24164 34242
rect 24108 34020 24164 34190
rect 24332 34132 24388 34142
rect 24444 34132 24500 34748
rect 24556 34738 24612 34748
rect 24892 34738 24948 34748
rect 24332 34130 24500 34132
rect 24332 34078 24334 34130
rect 24386 34078 24500 34130
rect 24332 34076 24500 34078
rect 25004 34690 25060 34702
rect 25004 34638 25006 34690
rect 25058 34638 25060 34690
rect 24332 34066 24388 34076
rect 23436 33966 23438 34018
rect 23490 33966 23492 34018
rect 23436 33954 23492 33966
rect 23772 33964 23940 34020
rect 23996 33964 24164 34020
rect 23212 33730 23268 33740
rect 22876 33346 23044 33348
rect 22876 33294 22878 33346
rect 22930 33294 23044 33346
rect 22876 33292 23044 33294
rect 23548 33348 23604 33358
rect 23548 33346 23716 33348
rect 23548 33294 23550 33346
rect 23602 33294 23716 33346
rect 23548 33292 23716 33294
rect 22876 33282 22932 33292
rect 23548 33282 23604 33292
rect 23212 33234 23268 33246
rect 23212 33182 23214 33234
rect 23266 33182 23268 33234
rect 22876 33124 22932 33134
rect 22876 31890 22932 33068
rect 23212 32228 23268 33182
rect 23548 33124 23604 33134
rect 23548 33030 23604 33068
rect 22876 31838 22878 31890
rect 22930 31838 22932 31890
rect 22876 31826 22932 31838
rect 22988 32172 23268 32228
rect 23548 32564 23604 32574
rect 22988 30996 23044 32172
rect 22988 30210 23044 30940
rect 23100 31220 23156 31230
rect 23100 30882 23156 31164
rect 23100 30830 23102 30882
rect 23154 30830 23156 30882
rect 23100 30660 23156 30830
rect 23100 30594 23156 30604
rect 22988 30158 22990 30210
rect 23042 30158 23044 30210
rect 22988 30146 23044 30158
rect 23548 30100 23604 32508
rect 23660 31220 23716 33292
rect 23660 31154 23716 31164
rect 23772 31668 23828 33964
rect 23660 30996 23716 31006
rect 23772 30996 23828 31612
rect 23660 30994 23828 30996
rect 23660 30942 23662 30994
rect 23714 30942 23828 30994
rect 23660 30940 23828 30942
rect 23884 33346 23940 33358
rect 23884 33294 23886 33346
rect 23938 33294 23940 33346
rect 23660 30930 23716 30940
rect 23772 30772 23828 30782
rect 23660 30100 23716 30110
rect 23548 30044 23660 30100
rect 23660 30034 23716 30044
rect 23772 29876 23828 30716
rect 23884 30548 23940 33294
rect 23996 31108 24052 33964
rect 23996 31042 24052 31052
rect 24332 33908 24388 33918
rect 24332 33346 24388 33852
rect 24892 33796 24948 33806
rect 24332 33294 24334 33346
rect 24386 33294 24388 33346
rect 24220 30882 24276 30894
rect 24220 30830 24222 30882
rect 24274 30830 24276 30882
rect 23884 30482 23940 30492
rect 23996 30770 24052 30782
rect 23996 30718 23998 30770
rect 24050 30718 24052 30770
rect 23996 30324 24052 30718
rect 23996 30258 24052 30268
rect 24220 30324 24276 30830
rect 24108 29986 24164 29998
rect 24108 29934 24110 29986
rect 24162 29934 24164 29986
rect 24108 29876 24164 29934
rect 23772 29820 24164 29876
rect 22092 28590 22094 28642
rect 22146 28590 22148 28642
rect 22092 28578 22148 28590
rect 22540 28644 22596 28654
rect 22764 28644 22820 28700
rect 22540 28550 22596 28588
rect 22652 28588 22820 28644
rect 23212 29426 23268 29438
rect 23212 29374 23214 29426
rect 23266 29374 23268 29426
rect 23212 28654 23268 29374
rect 23772 28980 23828 29820
rect 24220 29426 24276 30268
rect 24220 29374 24222 29426
rect 24274 29374 24276 29426
rect 24220 29362 24276 29374
rect 23884 29204 23940 29214
rect 24332 29204 24388 33294
rect 24556 33348 24612 33358
rect 24556 33234 24612 33292
rect 24556 33182 24558 33234
rect 24610 33182 24612 33234
rect 24556 33170 24612 33182
rect 24892 33122 24948 33740
rect 25004 33684 25060 34638
rect 25116 34468 25172 34860
rect 25788 34804 25844 34814
rect 25788 34710 25844 34748
rect 25452 34692 25508 34702
rect 25340 34690 25508 34692
rect 25340 34638 25454 34690
rect 25506 34638 25508 34690
rect 25340 34636 25508 34638
rect 25116 34412 25284 34468
rect 25004 33618 25060 33628
rect 25228 33234 25284 34412
rect 25228 33182 25230 33234
rect 25282 33182 25284 33234
rect 25228 33170 25284 33182
rect 24892 33070 24894 33122
rect 24946 33070 24948 33122
rect 24556 32900 24612 32910
rect 24556 32674 24612 32844
rect 24556 32622 24558 32674
rect 24610 32622 24612 32674
rect 24556 32610 24612 32622
rect 24668 32564 24724 32574
rect 24668 32470 24724 32508
rect 24780 31108 24836 31118
rect 24668 30884 24724 30894
rect 24556 29988 24612 29998
rect 24668 29988 24724 30828
rect 24612 29932 24724 29988
rect 24556 29894 24612 29932
rect 24444 29316 24500 29326
rect 24444 29222 24500 29260
rect 23884 29202 24388 29204
rect 23884 29150 23886 29202
rect 23938 29150 24388 29202
rect 23884 29148 24388 29150
rect 23884 29138 23940 29148
rect 23772 28924 24164 28980
rect 23996 28756 24052 28766
rect 23996 28662 24052 28700
rect 23212 28602 23214 28654
rect 23266 28644 23268 28654
rect 23266 28602 23604 28644
rect 23212 28588 23604 28602
rect 22316 28530 22372 28542
rect 22316 28478 22318 28530
rect 22370 28478 22372 28530
rect 22316 28420 22372 28478
rect 22652 28420 22708 28588
rect 22876 28532 22932 28542
rect 22876 28530 23492 28532
rect 22876 28478 22878 28530
rect 22930 28478 23492 28530
rect 22876 28476 23492 28478
rect 22876 28466 22932 28476
rect 22316 28364 22708 28420
rect 22876 28084 22932 28094
rect 23436 28084 23492 28476
rect 22540 28082 22932 28084
rect 22540 28030 22878 28082
rect 22930 28030 22932 28082
rect 22540 28028 22932 28030
rect 22428 27748 22484 27758
rect 22540 27748 22596 28028
rect 22876 28018 22932 28028
rect 23324 28082 23492 28084
rect 23324 28030 23438 28082
rect 23490 28030 23492 28082
rect 23324 28028 23492 28030
rect 22428 27746 22596 27748
rect 22428 27694 22430 27746
rect 22482 27694 22596 27746
rect 22428 27692 22596 27694
rect 22428 27682 22484 27692
rect 21980 26852 22372 26908
rect 22316 26628 22372 26852
rect 22316 26572 22484 26628
rect 21868 26338 21924 26348
rect 22316 26402 22372 26414
rect 22316 26350 22318 26402
rect 22370 26350 22372 26402
rect 22204 26292 22260 26302
rect 22204 26198 22260 26236
rect 21980 25508 22036 25518
rect 21980 25394 22036 25452
rect 21980 25342 21982 25394
rect 22034 25342 22036 25394
rect 21980 25330 22036 25342
rect 21756 25218 21812 25228
rect 22204 24612 22260 24622
rect 22092 24556 22204 24612
rect 21980 24500 22036 24510
rect 21756 24052 21812 24062
rect 21756 23940 21812 23996
rect 21868 23940 21924 23950
rect 21756 23938 21924 23940
rect 21756 23886 21870 23938
rect 21922 23886 21924 23938
rect 21756 23884 21924 23886
rect 21868 23874 21924 23884
rect 21980 23938 22036 24444
rect 21980 23886 21982 23938
rect 22034 23886 22036 23938
rect 21980 23874 22036 23886
rect 20748 23314 20804 23324
rect 21532 23772 21700 23828
rect 21308 23156 21364 23166
rect 21308 23062 21364 23100
rect 20636 20862 20638 20914
rect 20690 20862 20692 20914
rect 20636 20850 20692 20862
rect 20748 22370 20804 22382
rect 21420 22372 21476 22382
rect 20748 22318 20750 22370
rect 20802 22318 20804 22370
rect 20748 20804 20804 22318
rect 20748 20738 20804 20748
rect 20972 22370 21476 22372
rect 20972 22318 21422 22370
rect 21474 22318 21476 22370
rect 20972 22316 21476 22318
rect 20636 20692 20692 20702
rect 20636 19346 20692 20636
rect 20748 20580 20804 20590
rect 20972 20580 21028 22316
rect 21420 22306 21476 22316
rect 20748 20578 21028 20580
rect 20748 20526 20750 20578
rect 20802 20526 21028 20578
rect 20748 20524 21028 20526
rect 21308 20690 21364 20702
rect 21308 20638 21310 20690
rect 21362 20638 21364 20690
rect 20748 20514 20804 20524
rect 20748 20356 20804 20366
rect 20748 19458 20804 20300
rect 20748 19406 20750 19458
rect 20802 19406 20804 19458
rect 20748 19394 20804 19406
rect 20636 19294 20638 19346
rect 20690 19294 20692 19346
rect 20636 19282 20692 19294
rect 21308 19348 21364 20638
rect 21420 20692 21476 20702
rect 21420 20598 21476 20636
rect 21420 19348 21476 19358
rect 21308 19346 21476 19348
rect 21308 19294 21422 19346
rect 21474 19294 21476 19346
rect 21308 19292 21476 19294
rect 21420 19282 21476 19292
rect 21532 19124 21588 23772
rect 21756 23716 21812 23726
rect 21756 23622 21812 23660
rect 21644 23604 21700 23614
rect 21644 22482 21700 23548
rect 21644 22430 21646 22482
rect 21698 22430 21700 22482
rect 21644 20802 21700 22430
rect 21868 22932 21924 22942
rect 21868 22148 21924 22876
rect 21980 22484 22036 22494
rect 22092 22484 22148 24556
rect 22204 24546 22260 24556
rect 21980 22482 22148 22484
rect 21980 22430 21982 22482
rect 22034 22430 22148 22482
rect 21980 22428 22148 22430
rect 22204 23380 22260 23390
rect 21980 22418 22036 22428
rect 21868 22054 21924 22092
rect 22092 22148 22148 22158
rect 22204 22148 22260 23324
rect 22092 22146 22260 22148
rect 22092 22094 22094 22146
rect 22146 22094 22260 22146
rect 22092 22092 22260 22094
rect 21980 21924 22036 21934
rect 21644 20750 21646 20802
rect 21698 20750 21700 20802
rect 21644 20738 21700 20750
rect 21868 21868 21980 21924
rect 21868 20690 21924 21868
rect 21980 21858 22036 21868
rect 21980 20804 22036 20814
rect 22092 20804 22148 22092
rect 21980 20802 22148 20804
rect 21980 20750 21982 20802
rect 22034 20750 22148 20802
rect 21980 20748 22148 20750
rect 21980 20738 22036 20748
rect 21868 20638 21870 20690
rect 21922 20638 21924 20690
rect 21868 20626 21924 20638
rect 21308 19068 21588 19124
rect 21308 18788 21364 19068
rect 20860 18732 21364 18788
rect 20860 18340 20916 18732
rect 20860 17892 20916 18284
rect 20860 17778 20916 17836
rect 20860 17726 20862 17778
rect 20914 17726 20916 17778
rect 20860 17714 20916 17726
rect 20972 18562 21028 18574
rect 20972 18510 20974 18562
rect 21026 18510 21028 18562
rect 20300 17556 20356 17566
rect 20188 17500 20300 17556
rect 20300 17490 20356 17500
rect 20076 17388 20244 17444
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19964 16884 20020 16894
rect 19628 16882 20132 16884
rect 19628 16830 19966 16882
rect 20018 16830 20132 16882
rect 19628 16828 20132 16830
rect 19516 16772 19572 16782
rect 19292 16034 19348 16044
rect 19404 16770 19572 16772
rect 19404 16718 19518 16770
rect 19570 16718 19572 16770
rect 19404 16716 19572 16718
rect 19404 16098 19460 16716
rect 19516 16706 19572 16716
rect 19404 16046 19406 16098
rect 19458 16046 19460 16098
rect 17724 15810 17780 15820
rect 17948 15874 18004 15886
rect 17948 15822 17950 15874
rect 18002 15822 18004 15874
rect 17948 15540 18004 15822
rect 17948 15474 18004 15484
rect 18284 15874 18340 15886
rect 18284 15822 18286 15874
rect 18338 15822 18340 15874
rect 18284 15428 18340 15822
rect 18284 15362 18340 15372
rect 18396 15876 18452 15886
rect 18396 15538 18452 15820
rect 19068 15874 19124 15886
rect 19068 15822 19070 15874
rect 19122 15822 19124 15874
rect 18396 15486 18398 15538
rect 18450 15486 18452 15538
rect 18396 15148 18452 15486
rect 18844 15540 18900 15550
rect 18844 15446 18900 15484
rect 18732 15202 18788 15214
rect 18732 15150 18734 15202
rect 18786 15150 18788 15202
rect 18396 15092 18564 15148
rect 16604 14418 16660 14430
rect 16604 14366 16606 14418
rect 16658 14366 16660 14418
rect 16604 14308 16660 14366
rect 16604 14242 16660 14252
rect 18396 14420 18452 14430
rect 18396 13972 18452 14364
rect 18284 13970 18452 13972
rect 18284 13918 18398 13970
rect 18450 13918 18452 13970
rect 18284 13916 18452 13918
rect 17948 13858 18004 13870
rect 17948 13806 17950 13858
rect 18002 13806 18004 13858
rect 17836 13746 17892 13758
rect 17836 13694 17838 13746
rect 17890 13694 17892 13746
rect 16716 13076 16772 13086
rect 16716 12402 16772 13020
rect 17724 12964 17780 12974
rect 17836 12964 17892 13694
rect 17948 13748 18004 13806
rect 17948 13682 18004 13692
rect 17948 13524 18004 13534
rect 17948 13430 18004 13468
rect 17948 12964 18004 12974
rect 17836 12962 18004 12964
rect 17836 12910 17950 12962
rect 18002 12910 18004 12962
rect 17836 12908 18004 12910
rect 17724 12870 17780 12908
rect 16716 12350 16718 12402
rect 16770 12350 16772 12402
rect 16716 12338 16772 12350
rect 17612 12738 17668 12750
rect 17612 12686 17614 12738
rect 17666 12686 17668 12738
rect 17612 12290 17668 12686
rect 17612 12238 17614 12290
rect 17666 12238 17668 12290
rect 17612 12226 17668 12238
rect 17948 12290 18004 12908
rect 18284 12962 18340 13916
rect 18396 13906 18452 13916
rect 18508 13188 18564 15092
rect 18732 14642 18788 15150
rect 18732 14590 18734 14642
rect 18786 14590 18788 14642
rect 18732 14578 18788 14590
rect 18956 14308 19012 14318
rect 18844 14306 19012 14308
rect 18844 14254 18958 14306
rect 19010 14254 19012 14306
rect 18844 14252 19012 14254
rect 18508 13122 18564 13132
rect 18732 13524 18788 13534
rect 18844 13524 18900 14252
rect 18956 14242 19012 14252
rect 18732 13522 18900 13524
rect 18732 13470 18734 13522
rect 18786 13470 18900 13522
rect 18732 13468 18900 13470
rect 18956 13860 19012 13870
rect 19068 13860 19124 15822
rect 19404 15540 19460 16046
rect 19516 16548 19572 16558
rect 19516 15540 19572 16492
rect 19628 16212 19684 16828
rect 19964 16818 20020 16828
rect 19740 16660 19796 16670
rect 19740 16566 19796 16604
rect 19628 16118 19684 16156
rect 20076 15988 20132 16828
rect 20188 16324 20244 17388
rect 20524 17108 20580 17612
rect 20636 17108 20692 17118
rect 20524 17106 20692 17108
rect 20524 17054 20638 17106
rect 20690 17054 20692 17106
rect 20524 17052 20692 17054
rect 20636 17042 20692 17052
rect 20972 16996 21028 18510
rect 21308 18450 21364 18732
rect 21868 18676 21924 18686
rect 21924 18620 22036 18676
rect 21868 18582 21924 18620
rect 21308 18398 21310 18450
rect 21362 18398 21364 18450
rect 21308 18386 21364 18398
rect 21980 18116 22036 18620
rect 22204 18564 22260 18574
rect 22204 18450 22260 18508
rect 22204 18398 22206 18450
rect 22258 18398 22260 18450
rect 22204 18386 22260 18398
rect 22316 18452 22372 26350
rect 22428 22036 22484 26572
rect 22540 24164 22596 27692
rect 22652 27858 22708 27870
rect 22652 27806 22654 27858
rect 22706 27806 22708 27858
rect 22652 25732 22708 27806
rect 22652 25666 22708 25676
rect 22988 27858 23044 27870
rect 22988 27806 22990 27858
rect 23042 27806 23044 27858
rect 22876 24612 22932 24622
rect 22876 24518 22932 24556
rect 22988 24500 23044 27806
rect 22988 24434 23044 24444
rect 22540 24108 22708 24164
rect 22428 21970 22484 21980
rect 22540 23938 22596 23950
rect 22540 23886 22542 23938
rect 22594 23886 22596 23938
rect 22428 21586 22484 21598
rect 22428 21534 22430 21586
rect 22482 21534 22484 21586
rect 22428 19908 22484 21534
rect 22540 20356 22596 23886
rect 22540 20290 22596 20300
rect 22652 21924 22708 24108
rect 22764 23938 22820 23950
rect 22764 23886 22766 23938
rect 22818 23886 22820 23938
rect 22764 23604 22820 23886
rect 22764 23538 22820 23548
rect 22988 23940 23044 23950
rect 22988 23716 23044 23884
rect 23100 23828 23156 23838
rect 23100 23734 23156 23772
rect 22764 23156 22820 23166
rect 22764 23062 22820 23100
rect 22988 22370 23044 23660
rect 23212 23714 23268 23726
rect 23212 23662 23214 23714
rect 23266 23662 23268 23714
rect 23212 23380 23268 23662
rect 23324 23492 23380 28028
rect 23436 28018 23492 28028
rect 23548 27076 23604 28588
rect 23548 27010 23604 27020
rect 23436 26962 23492 26974
rect 23436 26910 23438 26962
rect 23490 26910 23492 26962
rect 23436 26516 23492 26910
rect 23436 26450 23492 26460
rect 23996 26852 24052 26862
rect 23996 26290 24052 26796
rect 23996 26238 23998 26290
rect 24050 26238 24052 26290
rect 23996 26226 24052 26238
rect 23548 25508 23604 25518
rect 23548 24724 23604 25452
rect 23548 24722 23940 24724
rect 23548 24670 23550 24722
rect 23602 24670 23940 24722
rect 23548 24668 23940 24670
rect 23548 24658 23604 24668
rect 23884 23938 23940 24668
rect 24108 23940 24164 28924
rect 24556 28084 24612 28094
rect 24332 27746 24388 27758
rect 24332 27694 24334 27746
rect 24386 27694 24388 27746
rect 24220 27076 24276 27086
rect 24220 26982 24276 27020
rect 24332 26852 24388 27694
rect 24556 26962 24612 28028
rect 24556 26910 24558 26962
rect 24610 26910 24612 26962
rect 24556 26898 24612 26910
rect 24332 26786 24388 26796
rect 24668 26740 24724 26750
rect 24556 26402 24612 26414
rect 24556 26350 24558 26402
rect 24610 26350 24612 26402
rect 24556 26292 24612 26350
rect 24556 25844 24612 26236
rect 24556 25778 24612 25788
rect 24668 25508 24724 26684
rect 24556 25452 24724 25508
rect 24332 25060 24388 25070
rect 24332 24834 24388 25004
rect 24444 24948 24500 24958
rect 24444 24854 24500 24892
rect 24332 24782 24334 24834
rect 24386 24782 24388 24834
rect 24332 24052 24388 24782
rect 24444 24500 24500 24510
rect 24444 24406 24500 24444
rect 24332 23996 24500 24052
rect 23884 23886 23886 23938
rect 23938 23886 23940 23938
rect 23884 23828 23940 23886
rect 23660 23772 23940 23828
rect 23996 23884 24164 23940
rect 23436 23492 23492 23502
rect 23324 23436 23436 23492
rect 23436 23426 23492 23436
rect 23212 23314 23268 23324
rect 23100 23268 23156 23278
rect 23100 23174 23156 23212
rect 23212 22930 23268 22942
rect 23212 22878 23214 22930
rect 23266 22878 23268 22930
rect 22988 22318 22990 22370
rect 23042 22318 23044 22370
rect 22876 22260 22932 22270
rect 22876 22166 22932 22204
rect 22428 19814 22484 19852
rect 22652 18788 22708 21868
rect 22764 22146 22820 22158
rect 22764 22094 22766 22146
rect 22818 22094 22820 22146
rect 22764 21700 22820 22094
rect 22764 21634 22820 21644
rect 22876 22036 22932 22046
rect 22876 21140 22932 21980
rect 22764 21084 22932 21140
rect 22764 18900 22820 21084
rect 22876 20580 22932 20590
rect 22876 20486 22932 20524
rect 22988 20132 23044 22318
rect 23100 22370 23156 22382
rect 23100 22318 23102 22370
rect 23154 22318 23156 22370
rect 23100 21812 23156 22318
rect 23100 21718 23156 21756
rect 23212 22372 23268 22878
rect 23660 22484 23716 23772
rect 23996 23604 24052 23884
rect 24444 23828 24500 23996
rect 24556 24050 24612 25452
rect 24556 23998 24558 24050
rect 24610 23998 24612 24050
rect 24556 23986 24612 23998
rect 24444 23772 24724 23828
rect 24444 23716 24500 23772
rect 23772 23548 24052 23604
rect 24108 23660 24500 23716
rect 23772 22596 23828 23548
rect 23884 23380 23940 23390
rect 23884 22932 23940 23324
rect 23996 23268 24052 23278
rect 23996 23174 24052 23212
rect 24108 23266 24164 23660
rect 24556 23380 24612 23390
rect 24556 23286 24612 23324
rect 24108 23214 24110 23266
rect 24162 23214 24164 23266
rect 24108 23202 24164 23214
rect 24668 23266 24724 23772
rect 24668 23214 24670 23266
rect 24722 23214 24724 23266
rect 24668 23202 24724 23214
rect 23996 22932 24052 22942
rect 24556 22932 24612 22942
rect 23884 22930 24052 22932
rect 23884 22878 23998 22930
rect 24050 22878 24052 22930
rect 23884 22876 24052 22878
rect 23996 22866 24052 22876
rect 24444 22930 24612 22932
rect 24444 22878 24558 22930
rect 24610 22878 24612 22930
rect 24444 22876 24612 22878
rect 23772 22540 23940 22596
rect 23660 22428 23828 22484
rect 23436 22372 23492 22382
rect 23212 22370 23492 22372
rect 23212 22318 23438 22370
rect 23490 22318 23492 22370
rect 23212 22316 23492 22318
rect 23212 20802 23268 22316
rect 23436 22306 23492 22316
rect 23772 22370 23828 22428
rect 23772 22318 23774 22370
rect 23826 22318 23828 22370
rect 23772 22306 23828 22318
rect 23324 21924 23380 21934
rect 23324 21810 23380 21868
rect 23324 21758 23326 21810
rect 23378 21758 23380 21810
rect 23324 21746 23380 21758
rect 23436 21700 23492 21710
rect 23436 21606 23492 21644
rect 23212 20750 23214 20802
rect 23266 20750 23268 20802
rect 23212 20738 23268 20750
rect 23772 21362 23828 21374
rect 23772 21310 23774 21362
rect 23826 21310 23828 21362
rect 23548 20692 23604 20702
rect 23548 20598 23604 20636
rect 23772 20692 23828 21310
rect 23772 20626 23828 20636
rect 23884 20356 23940 22540
rect 23996 21812 24052 21822
rect 24332 21812 24388 21822
rect 23996 21586 24052 21756
rect 23996 21534 23998 21586
rect 24050 21534 24052 21586
rect 23996 21522 24052 21534
rect 24108 21810 24388 21812
rect 24108 21758 24334 21810
rect 24386 21758 24388 21810
rect 24108 21756 24388 21758
rect 23660 20300 23940 20356
rect 23100 20132 23156 20142
rect 22988 20130 23156 20132
rect 22988 20078 23102 20130
rect 23154 20078 23156 20130
rect 22988 20076 23156 20078
rect 23100 19796 23156 20076
rect 23548 20020 23604 20030
rect 23100 19730 23156 19740
rect 23212 20018 23604 20020
rect 23212 19966 23550 20018
rect 23602 19966 23604 20018
rect 23212 19964 23604 19966
rect 22764 18844 22932 18900
rect 22652 18732 22820 18788
rect 22316 18386 22372 18396
rect 22652 18452 22708 18462
rect 22652 18358 22708 18396
rect 21980 18060 22372 18116
rect 21420 17556 21476 17566
rect 20860 16940 21028 16996
rect 21308 17442 21364 17454
rect 21308 17390 21310 17442
rect 21362 17390 21364 17442
rect 20188 16258 20244 16268
rect 20300 16660 20356 16670
rect 20300 16212 20356 16604
rect 20412 16660 20468 16670
rect 20412 16658 20692 16660
rect 20412 16606 20414 16658
rect 20466 16606 20692 16658
rect 20412 16604 20692 16606
rect 20412 16594 20468 16604
rect 20300 16156 20580 16212
rect 20300 15988 20356 15998
rect 20076 15986 20356 15988
rect 20076 15934 20302 15986
rect 20354 15934 20356 15986
rect 20076 15932 20356 15934
rect 20300 15922 20356 15932
rect 20524 15986 20580 16156
rect 20524 15934 20526 15986
rect 20578 15934 20580 15986
rect 20524 15922 20580 15934
rect 20412 15876 20468 15886
rect 20412 15782 20468 15820
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19628 15540 19684 15550
rect 19516 15484 19628 15540
rect 19404 15474 19460 15484
rect 19628 15474 19684 15484
rect 19964 15540 20020 15550
rect 19740 15428 19796 15438
rect 19740 15334 19796 15372
rect 19964 15426 20020 15484
rect 19964 15374 19966 15426
rect 20018 15374 20020 15426
rect 19964 15362 20020 15374
rect 20188 15540 20244 15550
rect 19516 15316 19572 15326
rect 19516 15222 19572 15260
rect 20188 15314 20244 15484
rect 20188 15262 20190 15314
rect 20242 15262 20244 15314
rect 20188 15250 20244 15262
rect 20636 15316 20692 16604
rect 20860 16212 20916 16940
rect 21084 16884 21140 16894
rect 20860 16146 20916 16156
rect 20972 16772 21028 16782
rect 20972 15540 21028 16716
rect 21084 16770 21140 16828
rect 21084 16718 21086 16770
rect 21138 16718 21140 16770
rect 21084 16706 21140 16718
rect 21308 16548 21364 17390
rect 21196 16324 21252 16334
rect 21196 16098 21252 16268
rect 21196 16046 21198 16098
rect 21250 16046 21252 16098
rect 21196 16034 21252 16046
rect 20972 15446 21028 15484
rect 20748 15428 20804 15438
rect 20748 15334 20804 15372
rect 20636 15222 20692 15260
rect 21196 15316 21252 15326
rect 21308 15316 21364 16492
rect 21420 15986 21476 17500
rect 21868 17554 21924 17566
rect 21868 17502 21870 17554
rect 21922 17502 21924 17554
rect 21868 17108 21924 17502
rect 21868 17042 21924 17052
rect 21532 16772 21588 16782
rect 21532 16678 21588 16716
rect 21868 16212 21924 16222
rect 21532 16100 21588 16110
rect 21532 16006 21588 16044
rect 21420 15934 21422 15986
rect 21474 15934 21476 15986
rect 21420 15922 21476 15934
rect 21868 15538 21924 16156
rect 21868 15486 21870 15538
rect 21922 15486 21924 15538
rect 21868 15474 21924 15486
rect 21980 16210 22036 16222
rect 21980 16158 21982 16210
rect 22034 16158 22036 16210
rect 21196 15314 21364 15316
rect 21196 15262 21198 15314
rect 21250 15262 21364 15314
rect 21196 15260 21364 15262
rect 21196 15250 21252 15260
rect 19628 15204 19684 15214
rect 19180 15090 19236 15102
rect 19180 15038 19182 15090
rect 19234 15038 19236 15090
rect 19180 14418 19236 15038
rect 19628 14754 19684 15148
rect 20860 15204 20916 15242
rect 21980 15148 22036 16158
rect 22316 16100 22372 18060
rect 22764 17780 22820 18732
rect 22876 18452 22932 18844
rect 22876 18386 22932 18396
rect 23212 18564 23268 19964
rect 23548 19954 23604 19964
rect 23660 19684 23716 20300
rect 23884 20132 23940 20142
rect 23884 20038 23940 20076
rect 23548 19628 23716 19684
rect 23548 19572 23604 19628
rect 23436 19516 23604 19572
rect 23436 19124 23492 19516
rect 24108 19460 24164 21756
rect 24332 21746 24388 21756
rect 24444 21810 24500 22876
rect 24556 22866 24612 22876
rect 24556 22484 24612 22494
rect 24556 22390 24612 22428
rect 24444 21758 24446 21810
rect 24498 21758 24500 21810
rect 24444 21700 24500 21758
rect 24444 21634 24500 21644
rect 24220 21586 24276 21598
rect 24220 21534 24222 21586
rect 24274 21534 24276 21586
rect 24220 21028 24276 21534
rect 24220 20962 24276 20972
rect 24332 19906 24388 19918
rect 24332 19854 24334 19906
rect 24386 19854 24388 19906
rect 24332 19796 24388 19854
rect 24332 19730 24388 19740
rect 23548 19404 24164 19460
rect 23548 19346 23604 19404
rect 24780 19348 24836 31052
rect 24892 28084 24948 33070
rect 25228 32564 25284 32574
rect 25228 32470 25284 32508
rect 25004 31892 25060 31902
rect 25004 31798 25060 31836
rect 25340 30884 25396 34636
rect 25452 34626 25508 34636
rect 25676 34692 25732 34702
rect 25676 34598 25732 34636
rect 25900 34244 25956 39900
rect 26012 39732 26068 39742
rect 26124 39732 26180 40348
rect 26460 40292 26516 40302
rect 26012 39730 26180 39732
rect 26012 39678 26014 39730
rect 26066 39678 26180 39730
rect 26012 39676 26180 39678
rect 26236 40290 26516 40292
rect 26236 40238 26462 40290
rect 26514 40238 26516 40290
rect 26236 40236 26516 40238
rect 26012 39666 26068 39676
rect 26236 39620 26292 40236
rect 26460 40226 26516 40236
rect 26124 39564 26292 39620
rect 26012 38836 26068 38846
rect 26124 38836 26180 39564
rect 26012 38834 26180 38836
rect 26012 38782 26014 38834
rect 26066 38782 26180 38834
rect 26012 38780 26180 38782
rect 26012 38770 26068 38780
rect 26124 38724 26180 38780
rect 26236 39396 26292 39406
rect 26236 38836 26292 39340
rect 26236 38742 26292 38780
rect 26124 38658 26180 38668
rect 26572 38052 26628 44270
rect 26684 42196 26740 45726
rect 26684 42130 26740 42140
rect 27020 45108 27076 45118
rect 27468 45108 27524 45836
rect 28364 45826 28420 45836
rect 32060 45890 32228 45892
rect 32060 45838 32174 45890
rect 32226 45838 32228 45890
rect 32060 45836 32228 45838
rect 29148 45780 29204 45790
rect 29148 45686 29204 45724
rect 30604 45780 30660 45790
rect 27692 45108 27748 45118
rect 27468 45106 27748 45108
rect 27468 45054 27694 45106
rect 27746 45054 27748 45106
rect 27468 45052 27748 45054
rect 26684 41748 26740 41758
rect 26684 41654 26740 41692
rect 26796 41746 26852 41758
rect 26796 41694 26798 41746
rect 26850 41694 26852 41746
rect 26796 41076 26852 41694
rect 26796 41010 26852 41020
rect 26684 40404 26740 40414
rect 26684 40310 26740 40348
rect 26908 39844 26964 39854
rect 26908 39730 26964 39788
rect 26908 39678 26910 39730
rect 26962 39678 26964 39730
rect 26908 39666 26964 39678
rect 26684 39396 26740 39406
rect 26684 39302 26740 39340
rect 26572 37958 26628 37996
rect 26796 38722 26852 38734
rect 26796 38670 26798 38722
rect 26850 38670 26852 38722
rect 26572 37380 26628 37390
rect 26796 37380 26852 38670
rect 27020 37604 27076 45052
rect 27132 44098 27188 44110
rect 27132 44046 27134 44098
rect 27186 44046 27188 44098
rect 27132 43652 27188 44046
rect 27132 43586 27188 43596
rect 27244 43428 27300 43438
rect 27692 43428 27748 45052
rect 28476 44996 28532 45006
rect 28476 44902 28532 44940
rect 30604 44996 30660 45724
rect 31388 45666 31444 45678
rect 31612 45668 31668 45678
rect 31388 45614 31390 45666
rect 31442 45614 31444 45666
rect 31388 45332 31444 45614
rect 31388 45266 31444 45276
rect 31500 45612 31612 45668
rect 31388 45108 31444 45118
rect 31500 45108 31556 45612
rect 31612 45602 31668 45612
rect 31948 45332 32004 45342
rect 31388 45106 31556 45108
rect 31388 45054 31390 45106
rect 31442 45054 31556 45106
rect 31388 45052 31556 45054
rect 31612 45276 31948 45332
rect 31612 45106 31668 45276
rect 31948 45238 32004 45276
rect 31612 45054 31614 45106
rect 31666 45054 31668 45106
rect 31388 45042 31444 45052
rect 31612 45042 31668 45054
rect 31724 45108 31780 45118
rect 31052 44996 31108 45006
rect 30604 44994 30996 44996
rect 30604 44942 30606 44994
rect 30658 44942 30996 44994
rect 30604 44940 30996 44942
rect 30604 44930 30660 44940
rect 30940 44772 30996 44940
rect 31052 44902 31108 44940
rect 31164 44882 31220 44894
rect 31164 44830 31166 44882
rect 31218 44830 31220 44882
rect 30940 44716 31108 44772
rect 30940 44436 30996 44446
rect 30940 44342 30996 44380
rect 30268 44210 30324 44222
rect 30268 44158 30270 44210
rect 30322 44158 30324 44210
rect 27244 43426 27748 43428
rect 27244 43374 27246 43426
rect 27298 43374 27748 43426
rect 27244 43372 27748 43374
rect 28476 43652 28532 43662
rect 27244 41972 27300 43372
rect 28476 42868 28532 43596
rect 30268 43652 30324 44158
rect 31052 44210 31108 44716
rect 31164 44548 31220 44830
rect 31164 44482 31220 44492
rect 31500 44322 31556 44334
rect 31500 44270 31502 44322
rect 31554 44270 31556 44322
rect 31052 44158 31054 44210
rect 31106 44158 31108 44210
rect 31052 44146 31108 44158
rect 31276 44210 31332 44222
rect 31276 44158 31278 44210
rect 31330 44158 31332 44210
rect 29596 43428 29652 43438
rect 28476 42802 28532 42812
rect 28588 42866 28644 42878
rect 28588 42814 28590 42866
rect 28642 42814 28644 42866
rect 28588 42756 28644 42814
rect 29148 42756 29204 42766
rect 28588 42754 29204 42756
rect 28588 42702 29150 42754
rect 29202 42702 29204 42754
rect 28588 42700 29204 42702
rect 27244 41878 27300 41916
rect 29148 41972 29204 42700
rect 29148 41906 29204 41916
rect 29372 42754 29428 42766
rect 29372 42702 29374 42754
rect 29426 42702 29428 42754
rect 28028 41860 28084 41870
rect 28028 41766 28084 41804
rect 27692 41748 27748 41758
rect 27692 40626 27748 41692
rect 28588 41300 28644 41310
rect 28588 41298 28980 41300
rect 28588 41246 28590 41298
rect 28642 41246 28980 41298
rect 28588 41244 28980 41246
rect 28588 41234 28644 41244
rect 27692 40574 27694 40626
rect 27746 40574 27748 40626
rect 27692 40562 27748 40574
rect 28924 40626 28980 41244
rect 28924 40574 28926 40626
rect 28978 40574 28980 40626
rect 28028 40516 28084 40526
rect 27244 40404 27300 40414
rect 27468 40404 27524 40414
rect 27244 40402 27524 40404
rect 27244 40350 27246 40402
rect 27298 40350 27470 40402
rect 27522 40350 27524 40402
rect 27244 40348 27524 40350
rect 27244 40338 27300 40348
rect 27244 39618 27300 39630
rect 27244 39566 27246 39618
rect 27298 39566 27300 39618
rect 27020 37538 27076 37548
rect 27132 38836 27188 38846
rect 27244 38836 27300 39566
rect 27132 38834 27300 38836
rect 27132 38782 27134 38834
rect 27186 38782 27300 38834
rect 27132 38780 27300 38782
rect 27356 39508 27412 40348
rect 27468 40338 27524 40348
rect 27804 40404 27860 40414
rect 27804 40310 27860 40348
rect 28028 40402 28084 40460
rect 28028 40350 28030 40402
rect 28082 40350 28084 40402
rect 28028 40338 28084 40350
rect 28364 40516 28420 40526
rect 28252 39844 28308 39854
rect 26572 37378 26852 37380
rect 26572 37326 26574 37378
rect 26626 37326 26852 37378
rect 26572 37324 26852 37326
rect 26572 37044 26628 37324
rect 26572 36978 26628 36988
rect 26348 35924 26404 35934
rect 26012 35588 26068 35598
rect 26012 35494 26068 35532
rect 26348 35476 26404 35868
rect 26908 35924 26964 35934
rect 27132 35924 27188 38780
rect 26908 35922 27188 35924
rect 26908 35870 26910 35922
rect 26962 35870 27188 35922
rect 26908 35868 27188 35870
rect 27244 37716 27300 37726
rect 26908 35858 26964 35868
rect 27244 35812 27300 37660
rect 27356 36036 27412 39452
rect 27692 39618 27748 39630
rect 27692 39566 27694 39618
rect 27746 39566 27748 39618
rect 27692 38946 27748 39566
rect 27692 38894 27694 38946
rect 27746 38894 27748 38946
rect 27692 38668 27748 38894
rect 27580 38612 27748 38668
rect 28252 38668 28308 39788
rect 28364 39620 28420 40460
rect 28924 40516 28980 40574
rect 28924 40450 28980 40460
rect 29372 41076 29428 42702
rect 29484 42756 29540 42766
rect 29484 41298 29540 42700
rect 29484 41246 29486 41298
rect 29538 41246 29540 41298
rect 29484 41234 29540 41246
rect 28476 40404 28532 40414
rect 28476 40310 28532 40348
rect 28700 40402 28756 40414
rect 28700 40350 28702 40402
rect 28754 40350 28756 40402
rect 28700 39956 28756 40350
rect 29148 40402 29204 40414
rect 29148 40350 29150 40402
rect 29202 40350 29204 40402
rect 28924 40292 28980 40302
rect 28924 40198 28980 40236
rect 29148 40180 29204 40350
rect 29148 40114 29204 40124
rect 28700 39900 29204 39956
rect 29148 39842 29204 39900
rect 29148 39790 29150 39842
rect 29202 39790 29204 39842
rect 29148 39778 29204 39790
rect 28476 39620 28532 39630
rect 28364 39618 28532 39620
rect 28364 39566 28478 39618
rect 28530 39566 28532 39618
rect 28364 39564 28532 39566
rect 28476 39554 28532 39564
rect 29260 39620 29316 39630
rect 29148 39508 29204 39518
rect 28588 39394 28644 39406
rect 28588 39342 28590 39394
rect 28642 39342 28644 39394
rect 28252 38612 28420 38668
rect 27580 37490 27636 38612
rect 27580 37438 27582 37490
rect 27634 37438 27636 37490
rect 27580 37426 27636 37438
rect 27804 37716 27860 37726
rect 27580 37266 27636 37278
rect 27580 37214 27582 37266
rect 27634 37214 27636 37266
rect 27580 36148 27636 37214
rect 27804 37266 27860 37660
rect 27804 37214 27806 37266
rect 27858 37214 27860 37266
rect 27804 37202 27860 37214
rect 27804 36372 27860 36382
rect 27804 36370 28196 36372
rect 27804 36318 27806 36370
rect 27858 36318 28196 36370
rect 27804 36316 28196 36318
rect 27804 36306 27860 36316
rect 27580 36092 27972 36148
rect 27356 35980 27860 36036
rect 27356 35812 27412 35822
rect 27244 35810 27412 35812
rect 27244 35758 27358 35810
rect 27410 35758 27412 35810
rect 27244 35756 27412 35758
rect 27356 35746 27412 35756
rect 26348 35028 26404 35420
rect 26684 35698 26740 35710
rect 26684 35646 26686 35698
rect 26738 35646 26740 35698
rect 26684 35364 26740 35646
rect 27692 35700 27748 35710
rect 27692 35606 27748 35644
rect 26684 35298 26740 35308
rect 25900 34178 25956 34188
rect 26012 35026 26404 35028
rect 26012 34974 26350 35026
rect 26402 34974 26404 35026
rect 26012 34972 26404 34974
rect 25788 34130 25844 34142
rect 25788 34078 25790 34130
rect 25842 34078 25844 34130
rect 25452 34018 25508 34030
rect 25452 33966 25454 34018
rect 25506 33966 25508 34018
rect 25452 31556 25508 33966
rect 25788 33012 25844 34078
rect 26012 34020 26068 34972
rect 26348 34962 26404 34972
rect 27020 34802 27076 34814
rect 27020 34750 27022 34802
rect 27074 34750 27076 34802
rect 26908 34692 26964 34702
rect 26460 34690 26964 34692
rect 26460 34638 26910 34690
rect 26962 34638 26964 34690
rect 26460 34636 26964 34638
rect 26460 34242 26516 34636
rect 26908 34626 26964 34636
rect 26460 34190 26462 34242
rect 26514 34190 26516 34242
rect 26460 34178 26516 34190
rect 25788 32946 25844 32956
rect 25900 33964 26068 34020
rect 25676 31892 25732 31902
rect 25732 31836 25844 31892
rect 25676 31826 25732 31836
rect 25676 31556 25732 31566
rect 25452 31500 25676 31556
rect 25564 31220 25620 31230
rect 25564 31126 25620 31164
rect 25676 30996 25732 31500
rect 25676 30930 25732 30940
rect 25340 30828 25620 30884
rect 25340 30548 25396 30558
rect 25396 30492 25508 30548
rect 25340 30482 25396 30492
rect 25452 30434 25508 30492
rect 25452 30382 25454 30434
rect 25506 30382 25508 30434
rect 25452 30370 25508 30382
rect 25564 30210 25620 30828
rect 25564 30158 25566 30210
rect 25618 30158 25620 30210
rect 25564 30146 25620 30158
rect 25004 30100 25060 30110
rect 25004 29986 25060 30044
rect 25004 29934 25006 29986
rect 25058 29934 25060 29986
rect 25004 29428 25060 29934
rect 25452 29988 25508 29998
rect 25788 29988 25844 31836
rect 25900 31778 25956 33964
rect 26796 33684 26852 33694
rect 26012 33348 26068 33358
rect 26068 33292 26180 33348
rect 26012 33254 26068 33292
rect 26012 32564 26068 32574
rect 26012 31890 26068 32508
rect 26012 31838 26014 31890
rect 26066 31838 26068 31890
rect 26012 31826 26068 31838
rect 25900 31726 25902 31778
rect 25954 31726 25956 31778
rect 25900 31714 25956 31726
rect 26124 31778 26180 33292
rect 26236 33122 26292 33134
rect 26236 33070 26238 33122
rect 26290 33070 26292 33122
rect 26236 32452 26292 33070
rect 26236 32386 26292 32396
rect 26684 32674 26740 32686
rect 26684 32622 26686 32674
rect 26738 32622 26740 32674
rect 26684 31892 26740 32622
rect 26684 31826 26740 31836
rect 26124 31726 26126 31778
rect 26178 31726 26180 31778
rect 26124 31444 26180 31726
rect 26796 31778 26852 33628
rect 26908 33458 26964 33470
rect 26908 33406 26910 33458
rect 26962 33406 26964 33458
rect 26908 32004 26964 33406
rect 27020 33460 27076 34750
rect 27020 33394 27076 33404
rect 27468 34692 27524 34702
rect 27356 33122 27412 33134
rect 27356 33070 27358 33122
rect 27410 33070 27412 33122
rect 27356 32900 27412 33070
rect 26908 31938 26964 31948
rect 27244 32844 27356 32900
rect 26796 31726 26798 31778
rect 26850 31726 26852 31778
rect 26572 31556 26628 31594
rect 26572 31490 26628 31500
rect 26012 31388 26180 31444
rect 26796 31444 26852 31726
rect 26908 31780 26964 31790
rect 27132 31780 27188 31790
rect 26908 31778 27132 31780
rect 26908 31726 26910 31778
rect 26962 31726 27132 31778
rect 26908 31724 27132 31726
rect 26908 31714 26964 31724
rect 27132 31714 27188 31724
rect 27020 31556 27076 31566
rect 27020 31554 27188 31556
rect 27020 31502 27022 31554
rect 27074 31502 27188 31554
rect 27020 31500 27188 31502
rect 27020 31490 27076 31500
rect 25900 31220 25956 31230
rect 26012 31220 26068 31388
rect 26796 31378 26852 31388
rect 25900 31218 26068 31220
rect 25900 31166 25902 31218
rect 25954 31166 26068 31218
rect 25900 31164 26068 31166
rect 26572 31332 26628 31342
rect 26572 31218 26628 31276
rect 26572 31166 26574 31218
rect 26626 31166 26628 31218
rect 25900 31154 25956 31164
rect 26572 31154 26628 31166
rect 26796 31220 26852 31230
rect 26796 31126 26852 31164
rect 27020 31220 27076 31230
rect 27132 31220 27188 31500
rect 27076 31218 27188 31220
rect 27076 31166 27134 31218
rect 27186 31166 27188 31218
rect 27076 31164 27188 31166
rect 27244 31220 27300 32844
rect 27356 32834 27412 32844
rect 27468 33124 27524 34636
rect 27580 33348 27636 33358
rect 27580 33254 27636 33292
rect 27692 33124 27748 33134
rect 27468 33068 27692 33124
rect 27468 32788 27524 33068
rect 27692 33030 27748 33068
rect 27468 32722 27524 32732
rect 27468 32228 27524 32238
rect 27356 31780 27412 31790
rect 27356 31686 27412 31724
rect 27356 31220 27412 31230
rect 27244 31218 27412 31220
rect 27244 31166 27358 31218
rect 27410 31166 27412 31218
rect 27244 31164 27412 31166
rect 27020 31154 27076 31164
rect 27132 31126 27188 31164
rect 27356 31154 27412 31164
rect 26124 30994 26180 31006
rect 26124 30942 26126 30994
rect 26178 30942 26180 30994
rect 26124 30884 26180 30942
rect 26124 30818 26180 30828
rect 26684 30882 26740 30894
rect 26684 30830 26686 30882
rect 26738 30830 26740 30882
rect 26460 30212 26516 30222
rect 26684 30212 26740 30830
rect 27244 30882 27300 30894
rect 27244 30830 27246 30882
rect 27298 30830 27300 30882
rect 26796 30212 26852 30222
rect 26684 30210 26852 30212
rect 26684 30158 26798 30210
rect 26850 30158 26852 30210
rect 26684 30156 26852 30158
rect 26460 30118 26516 30156
rect 26796 30146 26852 30156
rect 27132 30210 27188 30222
rect 27132 30158 27134 30210
rect 27186 30158 27188 30210
rect 25900 30100 25956 30110
rect 25900 30006 25956 30044
rect 26236 30100 26292 30110
rect 25452 29986 25844 29988
rect 25452 29934 25454 29986
rect 25506 29934 25844 29986
rect 25452 29932 25844 29934
rect 26012 29986 26068 29998
rect 26012 29934 26014 29986
rect 26066 29934 26068 29986
rect 25452 29922 25508 29932
rect 25340 29428 25396 29438
rect 25004 29426 25396 29428
rect 25004 29374 25342 29426
rect 25394 29374 25396 29426
rect 25004 29372 25396 29374
rect 24892 28018 24948 28028
rect 24892 26962 24948 26974
rect 24892 26910 24894 26962
rect 24946 26910 24948 26962
rect 24892 26852 24948 26910
rect 24892 25620 24948 26796
rect 24892 25554 24948 25564
rect 25116 25506 25172 29372
rect 25340 29362 25396 29372
rect 26012 28756 26068 29934
rect 26236 29652 26292 30044
rect 26236 29596 26628 29652
rect 26012 28690 26068 28700
rect 26124 28754 26180 28766
rect 26124 28702 26126 28754
rect 26178 28702 26180 28754
rect 26124 28644 26180 28702
rect 26124 28578 26180 28588
rect 26236 28084 26292 28094
rect 26124 27860 26180 27870
rect 25340 27748 25396 27758
rect 25340 27746 25732 27748
rect 25340 27694 25342 27746
rect 25394 27694 25732 27746
rect 25340 27692 25732 27694
rect 25340 27682 25396 27692
rect 25228 27634 25284 27646
rect 25228 27582 25230 27634
rect 25282 27582 25284 27634
rect 25228 26740 25284 27582
rect 25228 26674 25284 26684
rect 25452 27524 25508 27534
rect 25228 26404 25284 26414
rect 25452 26404 25508 27468
rect 25676 27186 25732 27692
rect 25676 27134 25678 27186
rect 25730 27134 25732 27186
rect 25676 27122 25732 27134
rect 25788 27300 25844 27310
rect 25676 26964 25732 27002
rect 25676 26898 25732 26908
rect 25788 26850 25844 27244
rect 26012 27188 26068 27198
rect 26012 27074 26068 27132
rect 26012 27022 26014 27074
rect 26066 27022 26068 27074
rect 26012 27010 26068 27022
rect 25788 26798 25790 26850
rect 25842 26798 25844 26850
rect 25788 26786 25844 26798
rect 25788 26516 25844 26526
rect 25788 26422 25844 26460
rect 25452 26348 25620 26404
rect 25228 26290 25284 26348
rect 25228 26238 25230 26290
rect 25282 26238 25284 26290
rect 25228 26226 25284 26238
rect 25564 26292 25620 26348
rect 25676 26292 25732 26302
rect 25564 26290 25732 26292
rect 25564 26238 25678 26290
rect 25730 26238 25732 26290
rect 25564 26236 25732 26238
rect 25452 26178 25508 26190
rect 25452 26126 25454 26178
rect 25506 26126 25508 26178
rect 25452 25732 25508 26126
rect 25452 25666 25508 25676
rect 25116 25454 25118 25506
rect 25170 25454 25172 25506
rect 25116 25442 25172 25454
rect 25116 25284 25172 25294
rect 25004 25228 25116 25284
rect 23548 19294 23550 19346
rect 23602 19294 23604 19346
rect 23548 19282 23604 19294
rect 23772 19292 24836 19348
rect 24892 20804 24948 20814
rect 23436 19068 23604 19124
rect 23212 18452 23268 18508
rect 23548 18452 23604 19068
rect 23212 18450 23380 18452
rect 23212 18398 23214 18450
rect 23266 18398 23380 18450
rect 23212 18396 23380 18398
rect 23212 18386 23268 18396
rect 23324 17890 23380 18396
rect 23548 18450 23716 18452
rect 23548 18398 23550 18450
rect 23602 18398 23716 18450
rect 23548 18396 23716 18398
rect 23548 18386 23604 18396
rect 23324 17838 23326 17890
rect 23378 17838 23380 17890
rect 23324 17826 23380 17838
rect 23436 17892 23492 17902
rect 22540 17724 22764 17780
rect 22428 17554 22484 17566
rect 22428 17502 22430 17554
rect 22482 17502 22484 17554
rect 22428 17108 22484 17502
rect 22428 17042 22484 17052
rect 22316 16006 22372 16044
rect 22428 15316 22484 15326
rect 22540 15316 22596 17724
rect 22764 17714 22820 17724
rect 23436 17778 23492 17836
rect 23660 17890 23716 18396
rect 23660 17838 23662 17890
rect 23714 17838 23716 17890
rect 23660 17826 23716 17838
rect 23436 17726 23438 17778
rect 23490 17726 23492 17778
rect 23436 17714 23492 17726
rect 22764 17554 22820 17566
rect 22764 17502 22766 17554
rect 22818 17502 22820 17554
rect 22652 17444 22708 17454
rect 22652 17350 22708 17388
rect 22764 16772 22820 17502
rect 22988 17556 23044 17566
rect 22988 17554 23268 17556
rect 22988 17502 22990 17554
rect 23042 17502 23268 17554
rect 22988 17500 23268 17502
rect 22988 17490 23044 17500
rect 22764 16706 22820 16716
rect 23100 17108 23156 17118
rect 23100 16100 23156 17052
rect 23212 16210 23268 17500
rect 23660 17444 23716 17454
rect 23660 16994 23716 17388
rect 23660 16942 23662 16994
rect 23714 16942 23716 16994
rect 23660 16930 23716 16942
rect 23212 16158 23214 16210
rect 23266 16158 23268 16210
rect 23212 16146 23268 16158
rect 23324 16772 23380 16782
rect 22876 16098 23156 16100
rect 22876 16046 23102 16098
rect 23154 16046 23156 16098
rect 22876 16044 23156 16046
rect 22876 15538 22932 16044
rect 23100 16034 23156 16044
rect 23324 16098 23380 16716
rect 23324 16046 23326 16098
rect 23378 16046 23380 16098
rect 23324 16034 23380 16046
rect 23772 16100 23828 19292
rect 24892 19236 24948 20748
rect 25004 20132 25060 25228
rect 25116 25218 25172 25228
rect 25452 25284 25508 25294
rect 25452 24836 25508 25228
rect 25452 24770 25508 24780
rect 25340 24724 25396 24734
rect 25340 24630 25396 24668
rect 25228 23828 25284 23838
rect 25228 23266 25284 23772
rect 25228 23214 25230 23266
rect 25282 23214 25284 23266
rect 25228 23202 25284 23214
rect 25116 23044 25172 23054
rect 25116 20802 25172 22988
rect 25340 22930 25396 22942
rect 25340 22878 25342 22930
rect 25394 22878 25396 22930
rect 25228 21476 25284 21486
rect 25228 21382 25284 21420
rect 25116 20750 25118 20802
rect 25170 20750 25172 20802
rect 25116 20738 25172 20750
rect 25340 20692 25396 22878
rect 25564 22932 25620 26236
rect 25676 26226 25732 26236
rect 25900 26290 25956 26302
rect 25900 26238 25902 26290
rect 25954 26238 25956 26290
rect 25788 24724 25844 24734
rect 25788 24630 25844 24668
rect 25900 24500 25956 26238
rect 25900 24434 25956 24444
rect 26012 26292 26068 26302
rect 25788 23716 25844 23726
rect 25788 23266 25844 23660
rect 25788 23214 25790 23266
rect 25842 23214 25844 23266
rect 25788 23202 25844 23214
rect 25564 22866 25620 22876
rect 25676 22930 25732 22942
rect 25676 22878 25678 22930
rect 25730 22878 25732 22930
rect 25676 22484 25732 22878
rect 25676 22418 25732 22428
rect 26012 20804 26068 26236
rect 26124 23940 26180 27804
rect 26236 27524 26292 28028
rect 26572 28082 26628 29596
rect 26796 29540 26852 29550
rect 26572 28030 26574 28082
rect 26626 28030 26628 28082
rect 26572 28018 26628 28030
rect 26684 28644 26740 28654
rect 26684 27970 26740 28588
rect 26684 27918 26686 27970
rect 26738 27918 26740 27970
rect 26684 27906 26740 27918
rect 26236 27458 26292 27468
rect 26796 27076 26852 29484
rect 27132 28642 27188 30158
rect 27244 30212 27300 30830
rect 27244 30146 27300 30156
rect 27468 30210 27524 32172
rect 27692 31778 27748 31790
rect 27692 31726 27694 31778
rect 27746 31726 27748 31778
rect 27692 31668 27748 31726
rect 27804 31780 27860 35980
rect 27916 35700 27972 36092
rect 28140 35922 28196 36316
rect 28140 35870 28142 35922
rect 28194 35870 28196 35922
rect 28140 35858 28196 35870
rect 28252 36260 28308 36270
rect 28252 35810 28308 36204
rect 28252 35758 28254 35810
rect 28306 35758 28308 35810
rect 28252 35746 28308 35758
rect 27916 35634 27972 35644
rect 27916 34692 27972 34702
rect 27916 33124 27972 34636
rect 28252 33346 28308 33358
rect 28252 33294 28254 33346
rect 28306 33294 28308 33346
rect 28252 33236 28308 33294
rect 28364 33348 28420 38612
rect 28588 38612 28644 39342
rect 28588 38546 28644 38556
rect 29148 38836 29204 39452
rect 29148 38274 29204 38780
rect 29260 38668 29316 39564
rect 29372 39058 29428 41020
rect 29596 39508 29652 43372
rect 29708 43316 29764 43326
rect 29708 42978 29764 43260
rect 29708 42926 29710 42978
rect 29762 42926 29764 42978
rect 29708 42914 29764 42926
rect 30156 42868 30212 42878
rect 29932 42866 30212 42868
rect 29932 42814 30158 42866
rect 30210 42814 30212 42866
rect 29932 42812 30212 42814
rect 29932 41636 29988 42812
rect 30156 42802 30212 42812
rect 30044 42644 30100 42654
rect 30044 42550 30100 42588
rect 30268 42532 30324 43596
rect 30604 44098 30660 44110
rect 30604 44046 30606 44098
rect 30658 44046 30660 44098
rect 30604 43540 30660 44046
rect 31276 43652 31332 44158
rect 31276 43586 31332 43596
rect 30604 43474 30660 43484
rect 31164 43540 31220 43550
rect 30604 43316 30660 43326
rect 30380 42756 30436 42766
rect 30380 42662 30436 42700
rect 30604 42754 30660 43260
rect 30604 42702 30606 42754
rect 30658 42702 30660 42754
rect 30604 42690 30660 42702
rect 31164 42866 31220 43484
rect 31388 43316 31444 43326
rect 31500 43316 31556 44270
rect 31444 43260 31556 43316
rect 31388 42978 31444 43260
rect 31388 42926 31390 42978
rect 31442 42926 31444 42978
rect 31388 42914 31444 42926
rect 31724 42978 31780 45052
rect 31948 44324 32004 44334
rect 31948 44230 32004 44268
rect 32060 43876 32116 45836
rect 32172 45826 32228 45836
rect 32620 45890 32676 46398
rect 32620 45838 32622 45890
rect 32674 45838 32676 45890
rect 32620 45826 32676 45838
rect 33180 46450 33236 46462
rect 33180 46398 33182 46450
rect 33234 46398 33236 46450
rect 33068 45780 33124 45790
rect 33068 45686 33124 45724
rect 32508 45444 32564 45454
rect 32284 45108 32340 45118
rect 32284 45014 32340 45052
rect 32508 44996 32564 45388
rect 32396 44994 32564 44996
rect 32396 44942 32510 44994
rect 32562 44942 32564 44994
rect 32396 44940 32564 44942
rect 32284 44548 32340 44558
rect 32284 44454 32340 44492
rect 32060 43820 32228 43876
rect 31724 42926 31726 42978
rect 31778 42926 31780 42978
rect 31724 42914 31780 42926
rect 31948 43538 32004 43550
rect 31948 43486 31950 43538
rect 32002 43486 32004 43538
rect 31164 42814 31166 42866
rect 31218 42814 31220 42866
rect 30156 42476 30324 42532
rect 30156 41858 30212 42476
rect 30828 42082 30884 42094
rect 30828 42030 30830 42082
rect 30882 42030 30884 42082
rect 30492 41972 30548 41982
rect 30492 41878 30548 41916
rect 30156 41806 30158 41858
rect 30210 41806 30212 41858
rect 30156 41794 30212 41806
rect 29932 41570 29988 41580
rect 30716 41412 30772 41422
rect 30828 41412 30884 42030
rect 31164 41412 31220 42814
rect 31948 42084 32004 43486
rect 32172 42644 32228 43820
rect 32396 43764 32452 44940
rect 32508 44930 32564 44940
rect 32620 45108 32676 45118
rect 32620 44546 32676 45052
rect 32620 44494 32622 44546
rect 32674 44494 32676 44546
rect 32620 44482 32676 44494
rect 33180 44434 33236 46398
rect 40348 46450 40404 46462
rect 40348 46398 40350 46450
rect 40402 46398 40404 46450
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 38220 45890 38276 45902
rect 38220 45838 38222 45890
rect 38274 45838 38276 45890
rect 33740 45778 33796 45790
rect 33740 45726 33742 45778
rect 33794 45726 33796 45778
rect 33404 45666 33460 45678
rect 33404 45614 33406 45666
rect 33458 45614 33460 45666
rect 33404 45444 33460 45614
rect 33404 45378 33460 45388
rect 33740 45108 33796 45726
rect 34412 45778 34468 45790
rect 34412 45726 34414 45778
rect 34466 45726 34468 45778
rect 33852 45668 33908 45678
rect 33852 45574 33908 45612
rect 33964 45666 34020 45678
rect 33964 45614 33966 45666
rect 34018 45614 34020 45666
rect 33964 45444 34020 45614
rect 33964 45378 34020 45388
rect 34412 45332 34468 45726
rect 37884 45778 37940 45790
rect 37884 45726 37886 45778
rect 37938 45726 37940 45778
rect 34412 45266 34468 45276
rect 34524 45666 34580 45678
rect 34524 45614 34526 45666
rect 34578 45614 34580 45666
rect 33740 45042 33796 45052
rect 33404 44996 33460 45006
rect 34524 44996 34580 45614
rect 33180 44382 33182 44434
rect 33234 44382 33236 44434
rect 33180 44370 33236 44382
rect 33292 44940 33404 44996
rect 33292 44436 33348 44940
rect 33404 44902 33460 44940
rect 33852 44940 34580 44996
rect 34636 45666 34692 45678
rect 34636 45614 34638 45666
rect 34690 45614 34692 45666
rect 34636 44996 34692 45614
rect 36316 45108 36372 45118
rect 36316 45106 36596 45108
rect 36316 45054 36318 45106
rect 36370 45054 36596 45106
rect 36316 45052 36596 45054
rect 36316 45042 36372 45052
rect 33852 44546 33908 44940
rect 34636 44930 34692 44940
rect 35532 44994 35588 45006
rect 35532 44942 35534 44994
rect 35586 44942 35588 44994
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 33852 44494 33854 44546
rect 33906 44494 33908 44546
rect 33852 44482 33908 44494
rect 33964 44548 34020 44558
rect 32508 44324 32564 44334
rect 32508 44322 33124 44324
rect 32508 44270 32510 44322
rect 32562 44270 33124 44322
rect 32508 44268 33124 44270
rect 32508 44258 32564 44268
rect 32620 44098 32676 44110
rect 32620 44046 32622 44098
rect 32674 44046 32676 44098
rect 32396 43708 32564 43764
rect 31948 42018 32004 42028
rect 32060 42588 32228 42644
rect 31276 41858 31332 41870
rect 31276 41806 31278 41858
rect 31330 41806 31332 41858
rect 31276 41636 31332 41806
rect 31276 41570 31332 41580
rect 30604 41410 31108 41412
rect 30604 41358 30718 41410
rect 30770 41358 31108 41410
rect 30604 41356 31108 41358
rect 29708 41186 29764 41198
rect 29708 41134 29710 41186
rect 29762 41134 29764 41186
rect 29708 40964 29764 41134
rect 29708 40898 29764 40908
rect 30604 40964 30660 41356
rect 30716 41346 30772 41356
rect 30492 40740 30548 40750
rect 30492 40626 30548 40684
rect 30492 40574 30494 40626
rect 30546 40574 30548 40626
rect 30492 40562 30548 40574
rect 30604 40626 30660 40908
rect 30604 40574 30606 40626
rect 30658 40574 30660 40626
rect 30604 40562 30660 40574
rect 30940 41186 30996 41198
rect 30940 41134 30942 41186
rect 30994 41134 30996 41186
rect 30156 40402 30212 40414
rect 30156 40350 30158 40402
rect 30210 40350 30212 40402
rect 29372 39006 29374 39058
rect 29426 39006 29428 39058
rect 29372 38994 29428 39006
rect 29484 39452 29652 39508
rect 29708 39618 29764 39630
rect 29708 39566 29710 39618
rect 29762 39566 29764 39618
rect 29708 39508 29764 39566
rect 30044 39620 30100 39630
rect 30044 39526 30100 39564
rect 29260 38612 29428 38668
rect 29148 38222 29150 38274
rect 29202 38222 29204 38274
rect 29148 38210 29204 38222
rect 29372 38162 29428 38612
rect 29372 38110 29374 38162
rect 29426 38110 29428 38162
rect 28588 37826 28644 37838
rect 28588 37774 28590 37826
rect 28642 37774 28644 37826
rect 28588 37716 28644 37774
rect 28644 37660 28868 37716
rect 28588 37650 28644 37660
rect 28588 37266 28644 37278
rect 28588 37214 28590 37266
rect 28642 37214 28644 37266
rect 28588 36482 28644 37214
rect 28588 36430 28590 36482
rect 28642 36430 28644 36482
rect 28588 34804 28644 36430
rect 28812 35922 28868 37660
rect 28924 37268 28980 37278
rect 29148 37268 29204 37278
rect 28924 37266 29204 37268
rect 28924 37214 28926 37266
rect 28978 37214 29150 37266
rect 29202 37214 29204 37266
rect 28924 37212 29204 37214
rect 28924 37202 28980 37212
rect 29148 37202 29204 37212
rect 29260 36596 29316 36606
rect 29260 36482 29316 36540
rect 29260 36430 29262 36482
rect 29314 36430 29316 36482
rect 29260 36418 29316 36430
rect 29372 36260 29428 38110
rect 29484 37492 29540 39452
rect 29708 39442 29764 39452
rect 29708 38948 29764 38958
rect 29596 38946 29764 38948
rect 29596 38894 29710 38946
rect 29762 38894 29764 38946
rect 29596 38892 29764 38894
rect 29596 38612 29652 38892
rect 29708 38882 29764 38892
rect 30156 38668 30212 40350
rect 30380 40402 30436 40414
rect 30380 40350 30382 40402
rect 30434 40350 30436 40402
rect 30268 39844 30324 39854
rect 30268 39750 30324 39788
rect 29596 38052 29652 38556
rect 29708 38612 30212 38668
rect 30380 38836 30436 40350
rect 30716 40404 30772 40414
rect 30940 40404 30996 41134
rect 30772 40348 30996 40404
rect 30716 40310 30772 40348
rect 31052 40068 31108 41356
rect 31164 41356 31892 41412
rect 31164 41186 31220 41356
rect 31164 41134 31166 41186
rect 31218 41134 31220 41186
rect 31164 41122 31220 41134
rect 31836 41186 31892 41356
rect 32060 41188 32116 42588
rect 32396 42530 32452 42542
rect 32396 42478 32398 42530
rect 32450 42478 32452 42530
rect 32396 42084 32452 42478
rect 32396 42018 32452 42028
rect 32508 41860 32564 43708
rect 32620 42532 32676 44046
rect 33068 43764 33124 44268
rect 33180 43764 33236 43774
rect 33068 43762 33236 43764
rect 33068 43710 33182 43762
rect 33234 43710 33236 43762
rect 33068 43708 33236 43710
rect 33180 43698 33236 43708
rect 33068 43316 33124 43326
rect 33068 43222 33124 43260
rect 33292 43092 33348 44380
rect 33964 44436 34020 44492
rect 34188 44548 34244 44558
rect 34188 44454 34244 44492
rect 35532 44548 35588 44942
rect 35532 44482 35588 44492
rect 34076 44436 34132 44446
rect 33964 44434 34132 44436
rect 33964 44382 34078 44434
rect 34130 44382 34132 44434
rect 33964 44380 34132 44382
rect 33628 44324 33684 44334
rect 33628 43764 33684 44268
rect 33628 43698 33684 43708
rect 33740 43764 33796 43774
rect 33964 43764 34020 44380
rect 34076 44370 34132 44380
rect 35868 44100 35924 44110
rect 35420 44098 35924 44100
rect 35420 44046 35870 44098
rect 35922 44046 35924 44098
rect 35420 44044 35924 44046
rect 33740 43762 34580 43764
rect 33740 43710 33742 43762
rect 33794 43710 34580 43762
rect 33740 43708 34580 43710
rect 33740 43698 33796 43708
rect 33404 43540 33460 43550
rect 33404 43446 33460 43484
rect 33964 43538 34020 43550
rect 33964 43486 33966 43538
rect 34018 43486 34020 43538
rect 33068 43036 33348 43092
rect 33068 42866 33124 43036
rect 33068 42814 33070 42866
rect 33122 42814 33124 42866
rect 33068 42802 33124 42814
rect 33628 42756 33684 42766
rect 33628 42662 33684 42700
rect 33180 42532 33236 42542
rect 32620 42476 32788 42532
rect 32396 41804 32564 41860
rect 32732 41860 32788 42476
rect 33180 42530 33572 42532
rect 33180 42478 33182 42530
rect 33234 42478 33572 42530
rect 33180 42476 33572 42478
rect 33180 42466 33236 42476
rect 33404 42308 33460 42318
rect 32396 41524 32452 41804
rect 32732 41794 32788 41804
rect 33068 41858 33124 41870
rect 33068 41806 33070 41858
rect 33122 41806 33124 41858
rect 33068 41524 33124 41806
rect 33180 41748 33236 41758
rect 33180 41746 33348 41748
rect 33180 41694 33182 41746
rect 33234 41694 33348 41746
rect 33180 41692 33348 41694
rect 33180 41682 33236 41692
rect 32396 41468 33124 41524
rect 31836 41134 31838 41186
rect 31890 41134 31892 41186
rect 31836 41122 31892 41134
rect 31948 41132 32116 41188
rect 32284 41188 32340 41198
rect 32396 41188 32452 41468
rect 32284 41186 32452 41188
rect 32284 41134 32286 41186
rect 32338 41134 32452 41186
rect 32284 41132 32452 41134
rect 32508 41188 32564 41198
rect 32844 41188 32900 41198
rect 32508 41186 32900 41188
rect 32508 41134 32510 41186
rect 32562 41134 32846 41186
rect 32898 41134 32900 41186
rect 32508 41132 32900 41134
rect 31276 40962 31332 40974
rect 31276 40910 31278 40962
rect 31330 40910 31332 40962
rect 31276 40740 31332 40910
rect 31388 40964 31444 40974
rect 31388 40870 31444 40908
rect 31276 40684 31668 40740
rect 31612 40626 31668 40684
rect 31612 40574 31614 40626
rect 31666 40574 31668 40626
rect 31388 40516 31444 40526
rect 31388 40422 31444 40460
rect 30716 40012 31108 40068
rect 31164 40404 31220 40414
rect 29708 38162 29764 38612
rect 30380 38274 30436 38780
rect 30380 38222 30382 38274
rect 30434 38222 30436 38274
rect 30380 38210 30436 38222
rect 30492 39620 30548 39630
rect 30492 38276 30548 39564
rect 30716 39618 30772 40012
rect 31052 39620 31108 39630
rect 30716 39566 30718 39618
rect 30770 39566 30772 39618
rect 30716 39554 30772 39566
rect 30940 39564 31052 39620
rect 30828 39396 30884 39406
rect 30940 39396 30996 39564
rect 31052 39554 31108 39564
rect 30828 39394 30996 39396
rect 30828 39342 30830 39394
rect 30882 39342 30996 39394
rect 30828 39340 30996 39342
rect 30828 39330 30884 39340
rect 31164 38668 31220 40348
rect 31500 40404 31556 40414
rect 31500 40310 31556 40348
rect 31276 40180 31332 40190
rect 31276 39058 31332 40124
rect 31276 39006 31278 39058
rect 31330 39006 31332 39058
rect 31276 38994 31332 39006
rect 31500 40180 31556 40190
rect 31388 38722 31444 38734
rect 31388 38670 31390 38722
rect 31442 38670 31444 38722
rect 31164 38612 31332 38668
rect 30828 38276 30884 38286
rect 30492 38274 30884 38276
rect 30492 38222 30830 38274
rect 30882 38222 30884 38274
rect 30492 38220 30884 38222
rect 30828 38210 30884 38220
rect 29708 38110 29710 38162
rect 29762 38110 29764 38162
rect 29708 38098 29764 38110
rect 29596 37958 29652 37996
rect 30380 38052 30436 38062
rect 30268 37940 30324 37950
rect 29484 37426 29540 37436
rect 29820 37828 29876 37838
rect 30268 37828 30324 37884
rect 30380 37938 30436 37996
rect 30380 37886 30382 37938
rect 30434 37886 30436 37938
rect 30380 37874 30436 37886
rect 30940 37938 30996 37950
rect 30940 37886 30942 37938
rect 30994 37886 30996 37938
rect 29820 37826 30324 37828
rect 29820 37774 29822 37826
rect 29874 37774 30324 37826
rect 29820 37772 30324 37774
rect 29820 36596 29876 37772
rect 29820 36530 29876 36540
rect 29932 37154 29988 37166
rect 29932 37102 29934 37154
rect 29986 37102 29988 37154
rect 29708 36372 29764 36382
rect 29708 36278 29764 36316
rect 28812 35870 28814 35922
rect 28866 35870 28868 35922
rect 28812 35858 28868 35870
rect 28924 36204 29428 36260
rect 29484 36258 29540 36270
rect 29484 36206 29486 36258
rect 29538 36206 29540 36258
rect 28588 34738 28644 34748
rect 28924 34468 28980 36204
rect 29148 36036 29204 36046
rect 29148 35922 29204 35980
rect 29148 35870 29150 35922
rect 29202 35870 29204 35922
rect 29148 35700 29204 35870
rect 29484 35812 29540 36206
rect 29596 36260 29652 36270
rect 29596 36166 29652 36204
rect 29820 36258 29876 36270
rect 29820 36206 29822 36258
rect 29874 36206 29876 36258
rect 29596 36036 29652 36046
rect 29596 35922 29652 35980
rect 29596 35870 29598 35922
rect 29650 35870 29652 35922
rect 29596 35858 29652 35870
rect 29372 35700 29428 35710
rect 29148 35634 29204 35644
rect 29260 35644 29372 35700
rect 29260 35026 29316 35644
rect 29372 35634 29428 35644
rect 29260 34974 29262 35026
rect 29314 34974 29316 35026
rect 29260 34962 29316 34974
rect 29484 34916 29540 35756
rect 29484 34850 29540 34860
rect 29820 35588 29876 36206
rect 29932 35922 29988 37102
rect 30940 37156 30996 37886
rect 30604 36596 30660 36606
rect 29932 35870 29934 35922
rect 29986 35870 29988 35922
rect 29932 35858 29988 35870
rect 30044 36594 30660 36596
rect 30044 36542 30606 36594
rect 30658 36542 30660 36594
rect 30044 36540 30660 36542
rect 30044 35810 30100 36540
rect 30604 36530 30660 36540
rect 30940 36484 30996 37100
rect 31164 37268 31220 37278
rect 31052 36484 31108 36494
rect 30940 36482 31108 36484
rect 30940 36430 31054 36482
rect 31106 36430 31108 36482
rect 30940 36428 31108 36430
rect 31052 36418 31108 36428
rect 30604 36260 30660 36270
rect 30044 35758 30046 35810
rect 30098 35758 30100 35810
rect 30044 35746 30100 35758
rect 30492 36258 30660 36260
rect 30492 36206 30606 36258
rect 30658 36206 30660 36258
rect 30492 36204 30660 36206
rect 30380 35700 30436 35710
rect 30492 35700 30548 36204
rect 30604 36194 30660 36204
rect 30716 36258 30772 36270
rect 30716 36206 30718 36258
rect 30770 36206 30772 36258
rect 30716 36148 30772 36206
rect 30716 36082 30772 36092
rect 30940 36258 30996 36270
rect 30940 36206 30942 36258
rect 30994 36206 30996 36258
rect 30828 35922 30884 35934
rect 30828 35870 30830 35922
rect 30882 35870 30884 35922
rect 30828 35812 30884 35870
rect 30940 35812 30996 36206
rect 30828 35756 30940 35812
rect 30940 35746 30996 35756
rect 30380 35698 30548 35700
rect 30380 35646 30382 35698
rect 30434 35646 30548 35698
rect 30380 35644 30548 35646
rect 30380 35588 30436 35644
rect 29820 35532 30436 35588
rect 29372 34692 29428 34730
rect 29372 34626 29428 34636
rect 29708 34692 29764 34702
rect 28588 34412 29316 34468
rect 28588 34018 28644 34412
rect 28588 33966 28590 34018
rect 28642 33966 28644 34018
rect 28588 33954 28644 33966
rect 29036 34132 29092 34142
rect 29036 33908 29092 34076
rect 29036 33852 29204 33908
rect 28364 33292 28756 33348
rect 28252 33170 28308 33180
rect 28588 33124 28644 33134
rect 27916 33122 28084 33124
rect 27916 33070 27918 33122
rect 27970 33070 28084 33122
rect 27916 33068 28084 33070
rect 27916 33058 27972 33068
rect 28028 32788 28084 33068
rect 28588 33030 28644 33068
rect 28028 32722 28084 32732
rect 28140 33012 28196 33022
rect 27916 32676 27972 32686
rect 27916 32582 27972 32620
rect 28028 32450 28084 32462
rect 28028 32398 28030 32450
rect 28082 32398 28084 32450
rect 27804 31714 27860 31724
rect 27916 32228 27972 32238
rect 27916 31778 27972 32172
rect 27916 31726 27918 31778
rect 27970 31726 27972 31778
rect 27916 31714 27972 31726
rect 27692 31602 27748 31612
rect 27804 31556 27860 31566
rect 27804 31462 27860 31500
rect 27916 31332 27972 31342
rect 27580 31108 27636 31118
rect 27580 31014 27636 31052
rect 27916 31108 27972 31276
rect 27916 31042 27972 31052
rect 28028 30994 28084 32398
rect 28028 30942 28030 30994
rect 28082 30942 28084 30994
rect 28028 30930 28084 30942
rect 28140 30996 28196 32956
rect 28476 33012 28532 33022
rect 28476 32788 28532 32956
rect 28476 32562 28532 32732
rect 28476 32510 28478 32562
rect 28530 32510 28532 32562
rect 28476 32498 28532 32510
rect 28588 31780 28644 31790
rect 28364 31556 28420 31566
rect 28364 31554 28532 31556
rect 28364 31502 28366 31554
rect 28418 31502 28532 31554
rect 28364 31500 28532 31502
rect 28364 31490 28420 31500
rect 28476 31332 28532 31500
rect 28476 31266 28532 31276
rect 28252 30996 28308 31006
rect 28140 30994 28532 30996
rect 28140 30942 28254 30994
rect 28306 30942 28532 30994
rect 28140 30940 28532 30942
rect 28252 30930 28308 30940
rect 27692 30882 27748 30894
rect 27692 30830 27694 30882
rect 27746 30830 27748 30882
rect 27692 30548 27748 30830
rect 27468 30158 27470 30210
rect 27522 30158 27524 30210
rect 27132 28590 27134 28642
rect 27186 28590 27188 28642
rect 27132 28084 27188 28590
rect 27244 29986 27300 29998
rect 27244 29934 27246 29986
rect 27298 29934 27300 29986
rect 27244 28420 27300 29934
rect 27468 29988 27524 30158
rect 27468 29922 27524 29932
rect 27580 30492 27972 30548
rect 27580 29764 27636 30492
rect 27916 30434 27972 30492
rect 27916 30382 27918 30434
rect 27970 30382 27972 30434
rect 27916 30370 27972 30382
rect 27692 30100 27748 30110
rect 27692 30006 27748 30044
rect 28252 29986 28308 29998
rect 28252 29934 28254 29986
rect 28306 29934 28308 29986
rect 27468 29708 27636 29764
rect 28028 29764 28084 29774
rect 27356 29540 27412 29550
rect 27356 29446 27412 29484
rect 27468 28868 27524 29708
rect 27468 28812 27748 28868
rect 27468 28754 27524 28812
rect 27468 28702 27470 28754
rect 27522 28702 27524 28754
rect 27468 28690 27524 28702
rect 27580 28644 27636 28654
rect 27244 28364 27524 28420
rect 27356 28196 27412 28206
rect 27132 28018 27188 28028
rect 27244 28140 27356 28196
rect 26236 26962 26292 26974
rect 26236 26910 26238 26962
rect 26290 26910 26292 26962
rect 26236 26908 26292 26910
rect 26572 26964 26628 27002
rect 26236 26852 26516 26908
rect 26572 26898 26628 26908
rect 26460 24612 26516 26852
rect 26684 26292 26740 26302
rect 26796 26292 26852 27020
rect 27020 27188 27076 27198
rect 26908 26852 26964 26862
rect 26908 26758 26964 26796
rect 26684 26290 26852 26292
rect 26684 26238 26686 26290
rect 26738 26238 26852 26290
rect 26684 26236 26852 26238
rect 26684 26226 26740 26236
rect 27020 25394 27076 27132
rect 27244 26908 27300 28140
rect 27356 28130 27412 28140
rect 27356 27300 27412 27310
rect 27356 27186 27412 27244
rect 27356 27134 27358 27186
rect 27410 27134 27412 27186
rect 27356 27122 27412 27134
rect 27020 25342 27022 25394
rect 27074 25342 27076 25394
rect 27020 25330 27076 25342
rect 27132 26852 27300 26908
rect 26796 25172 26852 25182
rect 26124 23874 26180 23884
rect 26236 24556 26740 24612
rect 26236 23266 26292 24556
rect 26684 24050 26740 24556
rect 26684 23998 26686 24050
rect 26738 23998 26740 24050
rect 26684 23986 26740 23998
rect 26684 23828 26740 23838
rect 26236 23214 26238 23266
rect 26290 23214 26292 23266
rect 26236 23202 26292 23214
rect 26460 23266 26516 23278
rect 26460 23214 26462 23266
rect 26514 23214 26516 23266
rect 26348 23044 26404 23054
rect 26348 22950 26404 22988
rect 26460 21476 26516 23214
rect 26684 22482 26740 23772
rect 26684 22430 26686 22482
rect 26738 22430 26740 22482
rect 26684 22418 26740 22430
rect 26460 21410 26516 21420
rect 26460 20804 26516 20814
rect 26012 20802 26516 20804
rect 26012 20750 26462 20802
rect 26514 20750 26516 20802
rect 26012 20748 26516 20750
rect 26460 20738 26516 20748
rect 25900 20692 25956 20702
rect 25340 20690 25956 20692
rect 25340 20638 25902 20690
rect 25954 20638 25956 20690
rect 25340 20636 25956 20638
rect 25900 20626 25956 20636
rect 25900 20132 25956 20142
rect 25004 20066 25060 20076
rect 25676 20130 25956 20132
rect 25676 20078 25902 20130
rect 25954 20078 25956 20130
rect 25676 20076 25956 20078
rect 25564 20018 25620 20030
rect 25564 19966 25566 20018
rect 25618 19966 25620 20018
rect 24332 19234 24948 19236
rect 24332 19222 24894 19234
rect 24332 19170 24334 19222
rect 24386 19182 24894 19222
rect 24946 19182 24948 19234
rect 24386 19180 24948 19182
rect 24386 19170 24388 19180
rect 24332 19158 24388 19170
rect 24108 18340 24164 18350
rect 24108 18246 24164 18284
rect 24220 17890 24276 17902
rect 24220 17838 24222 17890
rect 24274 17838 24276 17890
rect 23884 17780 23940 17790
rect 23884 17686 23940 17724
rect 23772 16098 24164 16100
rect 23772 16046 23774 16098
rect 23826 16046 24164 16098
rect 23772 16044 24164 16046
rect 23772 16034 23828 16044
rect 23996 15876 24052 15886
rect 23996 15782 24052 15820
rect 22876 15486 22878 15538
rect 22930 15486 22932 15538
rect 22876 15474 22932 15486
rect 23436 15540 23492 15550
rect 23436 15446 23492 15484
rect 24108 15538 24164 16044
rect 24108 15486 24110 15538
rect 24162 15486 24164 15538
rect 24108 15474 24164 15486
rect 22428 15314 22540 15316
rect 22428 15262 22430 15314
rect 22482 15262 22540 15314
rect 22428 15260 22540 15262
rect 22428 15250 22484 15260
rect 22540 15222 22596 15260
rect 23548 15314 23604 15326
rect 23548 15262 23550 15314
rect 23602 15262 23604 15314
rect 20860 15138 20916 15148
rect 19628 14702 19630 14754
rect 19682 14702 19684 14754
rect 19628 14690 19684 14702
rect 21868 15092 22036 15148
rect 23548 15148 23604 15262
rect 21308 14642 21364 14654
rect 21308 14590 21310 14642
rect 21362 14590 21364 14642
rect 19180 14366 19182 14418
rect 19234 14366 19236 14418
rect 19180 14354 19236 14366
rect 19404 14530 19460 14542
rect 19404 14478 19406 14530
rect 19458 14478 19460 14530
rect 19404 14418 19460 14478
rect 19404 14366 19406 14418
rect 19458 14366 19460 14418
rect 19404 14354 19460 14366
rect 19852 14530 19908 14542
rect 19852 14478 19854 14530
rect 19906 14478 19908 14530
rect 19516 14308 19572 14318
rect 19852 14308 19908 14478
rect 20300 14420 20356 14430
rect 20300 14326 20356 14364
rect 19516 14214 19572 14252
rect 19628 14252 19908 14308
rect 20412 14306 20468 14318
rect 20412 14254 20414 14306
rect 20466 14254 20468 14306
rect 18956 13858 19124 13860
rect 18956 13806 18958 13858
rect 19010 13806 19124 13858
rect 18956 13804 19124 13806
rect 18732 13074 18788 13468
rect 18732 13022 18734 13074
rect 18786 13022 18788 13074
rect 18732 13010 18788 13022
rect 18284 12910 18286 12962
rect 18338 12910 18340 12962
rect 18284 12898 18340 12910
rect 18844 12964 18900 12974
rect 18172 12852 18228 12862
rect 18172 12758 18228 12796
rect 18508 12852 18564 12862
rect 17948 12238 17950 12290
rect 18002 12238 18004 12290
rect 17948 12226 18004 12238
rect 16604 12178 16660 12190
rect 16604 12126 16606 12178
rect 16658 12126 16660 12178
rect 16604 11284 16660 12126
rect 16940 12180 16996 12190
rect 17388 12180 17444 12190
rect 16940 12178 17444 12180
rect 16940 12126 16942 12178
rect 16994 12126 17390 12178
rect 17442 12126 17444 12178
rect 16940 12124 17444 12126
rect 16940 12114 16996 12124
rect 17388 12114 17444 12124
rect 16716 12068 16772 12078
rect 16716 11506 16772 12012
rect 17836 12068 17892 12078
rect 17836 11974 17892 12012
rect 18508 12066 18564 12796
rect 18508 12014 18510 12066
rect 18562 12014 18564 12066
rect 18508 12002 18564 12014
rect 16716 11454 16718 11506
rect 16770 11454 16772 11506
rect 16716 11442 16772 11454
rect 18172 11732 18228 11742
rect 16604 11218 16660 11228
rect 18172 10610 18228 11676
rect 18844 11506 18900 12908
rect 18956 12962 19012 13804
rect 19516 13188 19572 13198
rect 19628 13188 19684 14252
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19572 13132 19684 13188
rect 19516 13122 19572 13132
rect 18956 12910 18958 12962
rect 19010 12910 19012 12962
rect 18956 12898 19012 12910
rect 19852 12964 19908 12974
rect 19852 12870 19908 12908
rect 20300 12964 20356 12974
rect 20300 12870 20356 12908
rect 18844 11454 18846 11506
rect 18898 11454 18900 11506
rect 18844 11442 18900 11454
rect 19068 12850 19124 12862
rect 19068 12798 19070 12850
rect 19122 12798 19124 12850
rect 19068 11396 19124 12798
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19068 11330 19124 11340
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 20412 10836 20468 14254
rect 20524 14306 20580 14318
rect 20524 14254 20526 14306
rect 20578 14254 20580 14306
rect 20524 12964 20580 14254
rect 21308 13860 21364 14590
rect 21308 13794 21364 13804
rect 21756 14532 21812 14542
rect 21756 13858 21812 14476
rect 21756 13806 21758 13858
rect 21810 13806 21812 13858
rect 21084 13524 21140 13534
rect 21140 13468 21252 13524
rect 21084 13458 21140 13468
rect 20524 12898 20580 12908
rect 20860 12740 20916 12750
rect 20860 12646 20916 12684
rect 20636 12068 20692 12078
rect 20636 12066 21140 12068
rect 20636 12014 20638 12066
rect 20690 12014 21140 12066
rect 20636 12012 21140 12014
rect 20636 12002 20692 12012
rect 20412 10770 20468 10780
rect 18172 10558 18174 10610
rect 18226 10558 18228 10610
rect 18172 10546 18228 10558
rect 16268 10444 16548 10500
rect 18844 10498 18900 10510
rect 18844 10446 18846 10498
rect 18898 10446 18900 10498
rect 16268 9268 16324 10444
rect 18844 10050 18900 10446
rect 18844 9998 18846 10050
rect 18898 9998 18900 10050
rect 18844 9986 18900 9998
rect 20972 10498 21028 10510
rect 20972 10446 20974 10498
rect 21026 10446 21028 10498
rect 16940 9938 16996 9950
rect 16940 9886 16942 9938
rect 16994 9886 16996 9938
rect 16828 9268 16884 9278
rect 16268 9266 16828 9268
rect 16268 9214 16270 9266
rect 16322 9214 16828 9266
rect 16268 9212 16828 9214
rect 16268 9202 16324 9212
rect 16828 9174 16884 9212
rect 16044 8484 16100 9100
rect 16044 8418 16100 8428
rect 16604 8484 16660 8494
rect 16268 8260 16324 8270
rect 16268 8166 16324 8204
rect 16044 8034 16100 8046
rect 16044 7982 16046 8034
rect 16098 7982 16100 8034
rect 16044 7924 16100 7982
rect 16156 8036 16212 8046
rect 16156 7942 16212 7980
rect 16044 7858 16100 7868
rect 16380 6804 16436 6814
rect 15932 5954 15988 5964
rect 16044 6802 16436 6804
rect 16044 6750 16382 6802
rect 16434 6750 16436 6802
rect 16044 6748 16436 6750
rect 16044 6468 16100 6748
rect 16380 6738 16436 6748
rect 16492 6804 16548 6814
rect 15148 5854 15150 5906
rect 15202 5854 15204 5906
rect 15148 5842 15204 5854
rect 15036 4958 15038 5010
rect 15090 4958 15092 5010
rect 15036 4946 15092 4958
rect 15148 5572 15204 5582
rect 14252 4398 14254 4450
rect 14306 4398 14308 4450
rect 14252 4386 14308 4398
rect 13580 4286 13582 4338
rect 13634 4286 13636 4338
rect 13580 4274 13636 4286
rect 7084 4174 7086 4226
rect 7138 4174 7140 4226
rect 7084 4162 7140 4174
rect 7532 4228 7588 4238
rect 4476 3948 4740 3958
rect 6972 3948 7476 4004
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 7420 3778 7476 3948
rect 7420 3726 7422 3778
rect 7474 3726 7476 3778
rect 7420 3714 7476 3726
rect 7532 3666 7588 4172
rect 7532 3614 7534 3666
rect 7586 3614 7588 3666
rect 7532 3602 7588 3614
rect 13132 4226 13188 4238
rect 13132 4174 13134 4226
rect 13186 4174 13188 4226
rect 7756 3554 7812 3566
rect 7756 3502 7758 3554
rect 7810 3502 7812 3554
rect 7756 3444 7812 3502
rect 13132 3556 13188 4174
rect 13132 3490 13188 3500
rect 7756 3378 7812 3388
rect 8204 3444 8260 3454
rect 8204 3350 8260 3388
rect 15148 3444 15204 5516
rect 15260 5236 15316 5246
rect 15708 5236 15764 5246
rect 15260 5234 15764 5236
rect 15260 5182 15262 5234
rect 15314 5182 15710 5234
rect 15762 5182 15764 5234
rect 15260 5180 15764 5182
rect 15260 5170 15316 5180
rect 15708 5170 15764 5180
rect 16044 5124 16100 6412
rect 16268 6580 16324 6590
rect 16268 6130 16324 6524
rect 16268 6078 16270 6130
rect 16322 6078 16324 6130
rect 16268 6066 16324 6078
rect 16156 6020 16212 6030
rect 16156 5926 16212 5964
rect 16380 6020 16436 6030
rect 16492 6020 16548 6748
rect 16380 6018 16548 6020
rect 16380 5966 16382 6018
rect 16434 5966 16548 6018
rect 16380 5964 16548 5966
rect 16380 5954 16436 5964
rect 16156 5124 16212 5134
rect 16044 5122 16212 5124
rect 16044 5070 16158 5122
rect 16210 5070 16212 5122
rect 16044 5068 16212 5070
rect 16156 5058 16212 5068
rect 16604 5124 16660 8428
rect 16716 8370 16772 8382
rect 16716 8318 16718 8370
rect 16770 8318 16772 8370
rect 16716 8260 16772 8318
rect 16716 8194 16772 8204
rect 16716 8036 16772 8046
rect 16716 7942 16772 7980
rect 16828 8034 16884 8046
rect 16828 7982 16830 8034
rect 16882 7982 16884 8034
rect 16716 7364 16772 7374
rect 16828 7364 16884 7982
rect 16716 7362 16884 7364
rect 16716 7310 16718 7362
rect 16770 7310 16884 7362
rect 16716 7308 16884 7310
rect 16716 6690 16772 7308
rect 16940 6692 16996 9886
rect 17500 9828 17556 9838
rect 18060 9828 18116 9838
rect 17500 9826 18116 9828
rect 17500 9774 17502 9826
rect 17554 9774 18062 9826
rect 18114 9774 18116 9826
rect 17500 9772 18116 9774
rect 17276 9716 17332 9726
rect 17276 9604 17332 9660
rect 17164 9602 17332 9604
rect 17164 9550 17278 9602
rect 17330 9550 17332 9602
rect 17164 9548 17332 9550
rect 17052 8034 17108 8046
rect 17052 7982 17054 8034
rect 17106 7982 17108 8034
rect 17052 7028 17108 7982
rect 17164 7924 17220 9548
rect 17276 9538 17332 9548
rect 17500 9268 17556 9772
rect 18060 9762 18116 9772
rect 18844 9826 18900 9838
rect 18844 9774 18846 9826
rect 18898 9774 18900 9826
rect 18844 9716 18900 9774
rect 20972 9828 21028 10446
rect 21084 10500 21140 12012
rect 21196 10612 21252 13468
rect 21308 13188 21364 13198
rect 21308 13074 21364 13132
rect 21308 13022 21310 13074
rect 21362 13022 21364 13074
rect 21308 13010 21364 13022
rect 21420 12180 21476 12190
rect 21756 12180 21812 13806
rect 21420 12178 21812 12180
rect 21420 12126 21422 12178
rect 21474 12126 21758 12178
rect 21810 12126 21812 12178
rect 21420 12124 21812 12126
rect 21420 11844 21476 12124
rect 21756 12114 21812 12124
rect 21868 12740 21924 15092
rect 23436 15090 23492 15102
rect 23548 15092 23828 15148
rect 23436 15038 23438 15090
rect 23490 15038 23492 15090
rect 23436 14642 23492 15038
rect 23436 14590 23438 14642
rect 23490 14590 23492 14642
rect 23436 14578 23492 14590
rect 22428 13860 22484 13870
rect 22428 13076 22484 13804
rect 23212 13748 23268 13758
rect 22428 13074 23156 13076
rect 22428 13022 22430 13074
rect 22482 13022 23156 13074
rect 22428 13020 23156 13022
rect 22428 13010 22484 13020
rect 23100 12962 23156 13020
rect 23100 12910 23102 12962
rect 23154 12910 23156 12962
rect 23100 12898 23156 12910
rect 21420 11778 21476 11788
rect 21868 11394 21924 12684
rect 22540 12740 22596 12750
rect 22540 12290 22596 12684
rect 22540 12238 22542 12290
rect 22594 12238 22596 12290
rect 22540 12226 22596 12238
rect 21868 11342 21870 11394
rect 21922 11342 21924 11394
rect 21868 11060 21924 11342
rect 21868 10994 21924 11004
rect 22204 11956 22260 11966
rect 22204 11506 22260 11900
rect 22204 11454 22206 11506
rect 22258 11454 22260 11506
rect 21532 10836 21588 10846
rect 21532 10742 21588 10780
rect 21308 10612 21364 10622
rect 21196 10610 21364 10612
rect 21196 10558 21310 10610
rect 21362 10558 21364 10610
rect 21196 10556 21364 10558
rect 21308 10546 21364 10556
rect 21084 10444 21252 10500
rect 21196 10388 21252 10444
rect 21420 10498 21476 10510
rect 21420 10446 21422 10498
rect 21474 10446 21476 10498
rect 21420 10388 21476 10446
rect 21196 10332 21476 10388
rect 20972 9762 21028 9772
rect 21308 9826 21364 9838
rect 21532 9828 21588 9838
rect 21308 9774 21310 9826
rect 21362 9774 21364 9826
rect 18844 9650 18900 9660
rect 19180 9714 19236 9726
rect 19180 9662 19182 9714
rect 19234 9662 19236 9714
rect 17500 9202 17556 9212
rect 18732 9604 18788 9614
rect 17388 9156 17444 9166
rect 17388 9044 17444 9100
rect 17388 9042 17668 9044
rect 17388 8990 17390 9042
rect 17442 8990 17668 9042
rect 17388 8988 17668 8990
rect 17388 8978 17444 8988
rect 17276 8148 17332 8158
rect 17276 8054 17332 8092
rect 17388 8036 17444 8046
rect 17276 7924 17332 7934
rect 17164 7868 17276 7924
rect 17276 7858 17332 7868
rect 17052 6972 17332 7028
rect 17052 6804 17108 6814
rect 17052 6710 17108 6748
rect 16716 6638 16718 6690
rect 16770 6638 16772 6690
rect 16716 6626 16772 6638
rect 16828 6636 16996 6692
rect 16604 5030 16660 5068
rect 15708 5012 15764 5022
rect 15708 4918 15764 4956
rect 15820 5012 15876 5022
rect 15820 5010 15988 5012
rect 15820 4958 15822 5010
rect 15874 4958 15988 5010
rect 15820 4956 15988 4958
rect 15820 4946 15876 4956
rect 15932 4452 15988 4956
rect 16044 4900 16100 4910
rect 16044 4806 16100 4844
rect 16380 4452 16436 4462
rect 15932 4396 16380 4452
rect 16380 4226 16436 4396
rect 16380 4174 16382 4226
rect 16434 4174 16436 4226
rect 16380 4162 16436 4174
rect 16828 4004 16884 6636
rect 16940 6466 16996 6478
rect 16940 6414 16942 6466
rect 16994 6414 16996 6466
rect 16940 6132 16996 6414
rect 17164 6468 17220 6478
rect 17164 6374 17220 6412
rect 17276 6132 17332 6972
rect 17388 6692 17444 7980
rect 17612 7586 17668 8988
rect 18172 8932 18228 8942
rect 18172 8930 18452 8932
rect 18172 8878 18174 8930
rect 18226 8878 18452 8930
rect 18172 8876 18452 8878
rect 18172 8866 18228 8876
rect 18396 8482 18452 8876
rect 18396 8430 18398 8482
rect 18450 8430 18452 8482
rect 18396 8418 18452 8430
rect 18732 8370 18788 9548
rect 18732 8318 18734 8370
rect 18786 8318 18788 8370
rect 18732 8306 18788 8318
rect 19180 8372 19236 9662
rect 20524 9492 20580 9502
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 20300 9436 20524 9492
rect 20580 9436 20692 9492
rect 20300 8930 20356 9436
rect 20524 9426 20580 9436
rect 20300 8878 20302 8930
rect 20354 8878 20356 8930
rect 20300 8866 20356 8878
rect 19180 8306 19236 8316
rect 20188 8370 20244 8382
rect 20188 8318 20190 8370
rect 20242 8318 20244 8370
rect 18060 8260 18116 8270
rect 18060 8166 18116 8204
rect 18396 8258 18452 8270
rect 18396 8206 18398 8258
rect 18450 8206 18452 8258
rect 17612 7534 17614 7586
rect 17666 7534 17668 7586
rect 17612 7522 17668 7534
rect 17724 8148 17780 8158
rect 17724 6804 17780 8092
rect 17836 8034 17892 8046
rect 17836 7982 17838 8034
rect 17890 7982 17892 8034
rect 17836 7924 17892 7982
rect 17836 7858 17892 7868
rect 17948 8034 18004 8046
rect 17948 7982 17950 8034
rect 18002 7982 18004 8034
rect 17836 6804 17892 6814
rect 17724 6802 17892 6804
rect 17724 6750 17838 6802
rect 17890 6750 17892 6802
rect 17724 6748 17892 6750
rect 17836 6738 17892 6748
rect 17388 6690 17780 6692
rect 17388 6638 17390 6690
rect 17442 6638 17780 6690
rect 17388 6636 17780 6638
rect 17388 6626 17444 6636
rect 17612 6132 17668 6142
rect 17276 6076 17612 6132
rect 16940 6066 16996 6076
rect 16380 3948 16884 4004
rect 17052 6020 17108 6030
rect 16380 3554 16436 3948
rect 16380 3502 16382 3554
rect 16434 3502 16436 3554
rect 16380 3490 16436 3502
rect 15148 3378 15204 3388
rect 17052 3442 17108 5964
rect 17388 5012 17444 5022
rect 17164 5010 17444 5012
rect 17164 4958 17390 5010
rect 17442 4958 17444 5010
rect 17164 4956 17444 4958
rect 17164 3666 17220 4956
rect 17388 4946 17444 4956
rect 17500 4900 17556 6076
rect 17612 6066 17668 6076
rect 17612 5796 17668 5806
rect 17612 5702 17668 5740
rect 17724 5684 17780 6636
rect 17948 6580 18004 7982
rect 18396 7924 18452 8206
rect 19628 8258 19684 8270
rect 19628 8206 19630 8258
rect 19682 8206 19684 8258
rect 19404 8036 19460 8046
rect 19404 7942 19460 7980
rect 18396 7858 18452 7868
rect 19628 7700 19684 8206
rect 20188 8260 20244 8318
rect 20188 8194 20244 8204
rect 20636 8258 20692 9436
rect 20860 8930 20916 8942
rect 20860 8878 20862 8930
rect 20914 8878 20916 8930
rect 20860 8484 20916 8878
rect 21196 8932 21252 8942
rect 21196 8838 21252 8876
rect 20860 8418 20916 8428
rect 20636 8206 20638 8258
rect 20690 8206 20692 8258
rect 20636 8194 20692 8206
rect 20300 8148 20356 8158
rect 21308 8148 21364 9774
rect 21420 9772 21532 9828
rect 21420 9268 21476 9772
rect 21532 9762 21588 9772
rect 21868 9828 21924 9838
rect 21868 9734 21924 9772
rect 21532 9602 21588 9614
rect 21532 9550 21534 9602
rect 21586 9550 21588 9602
rect 21532 9492 21588 9550
rect 21644 9604 21700 9614
rect 21644 9510 21700 9548
rect 21756 9602 21812 9614
rect 21756 9550 21758 9602
rect 21810 9550 21812 9602
rect 21532 9426 21588 9436
rect 21420 9212 21588 9268
rect 21420 8372 21476 8382
rect 21420 8278 21476 8316
rect 21532 8258 21588 9212
rect 21532 8206 21534 8258
rect 21586 8206 21588 8258
rect 21532 8194 21588 8206
rect 21420 8148 21476 8158
rect 21308 8092 21420 8148
rect 20300 8054 20356 8092
rect 21420 8054 21476 8092
rect 20188 8036 20244 8046
rect 20188 7942 20244 7980
rect 20524 8034 20580 8046
rect 20524 7982 20526 8034
rect 20578 7982 20580 8034
rect 20524 7924 20580 7982
rect 21756 8034 21812 9550
rect 21980 8932 22036 8942
rect 21980 8258 22036 8876
rect 21980 8206 21982 8258
rect 22034 8206 22036 8258
rect 21980 8194 22036 8206
rect 21756 7982 21758 8034
rect 21810 7982 21812 8034
rect 21756 7924 21812 7982
rect 19836 7868 20100 7878
rect 20524 7868 21812 7924
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19740 7700 19796 7710
rect 19628 7644 19740 7700
rect 19740 7634 19796 7644
rect 20300 7700 20356 7710
rect 17948 6514 18004 6524
rect 19964 6580 20020 6590
rect 19964 6486 20020 6524
rect 19292 6468 19348 6478
rect 17948 5908 18004 5918
rect 17948 5814 18004 5852
rect 18172 5684 18228 5694
rect 17724 5628 18004 5684
rect 17948 5348 18004 5628
rect 17500 4564 17556 4844
rect 17836 5236 17892 5246
rect 17612 4564 17668 4574
rect 17500 4562 17668 4564
rect 17500 4510 17614 4562
rect 17666 4510 17668 4562
rect 17500 4508 17668 4510
rect 17612 4498 17668 4508
rect 17836 4562 17892 5180
rect 17836 4510 17838 4562
rect 17890 4510 17892 4562
rect 17836 4498 17892 4510
rect 17948 4562 18004 5292
rect 17948 4510 17950 4562
rect 18002 4510 18004 4562
rect 17948 4498 18004 4510
rect 17388 4452 17444 4462
rect 17388 4358 17444 4396
rect 17724 4226 17780 4238
rect 17724 4174 17726 4226
rect 17778 4174 17780 4226
rect 17724 3892 17780 4174
rect 17276 3836 17780 3892
rect 17276 3778 17332 3836
rect 17276 3726 17278 3778
rect 17330 3726 17332 3778
rect 17276 3714 17332 3726
rect 17164 3614 17166 3666
rect 17218 3614 17220 3666
rect 17164 3602 17220 3614
rect 17612 3556 17668 3566
rect 17612 3462 17668 3500
rect 17052 3390 17054 3442
rect 17106 3390 17108 3442
rect 17052 3378 17108 3390
rect 18172 3388 18228 5628
rect 18956 5684 19012 5694
rect 18956 5590 19012 5628
rect 18508 5124 18564 5134
rect 18508 4338 18564 5068
rect 19292 4450 19348 6412
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 20076 5908 20132 5918
rect 19516 5236 19572 5246
rect 19572 5180 19908 5236
rect 19516 5142 19572 5180
rect 19852 5122 19908 5180
rect 19852 5070 19854 5122
rect 19906 5070 19908 5122
rect 19852 5058 19908 5070
rect 20076 5010 20132 5852
rect 20300 5348 20356 7644
rect 21756 6804 21812 7868
rect 21756 6748 21924 6804
rect 20748 6690 20804 6702
rect 20748 6638 20750 6690
rect 20802 6638 20804 6690
rect 20748 6580 20804 6638
rect 21308 6580 21364 6590
rect 20748 6514 20804 6524
rect 20972 6578 21364 6580
rect 20972 6526 21310 6578
rect 21362 6526 21364 6578
rect 20972 6524 21364 6526
rect 20860 6132 20916 6142
rect 20860 6038 20916 6076
rect 20972 5684 21028 6524
rect 21308 6514 21364 6524
rect 21756 6580 21812 6590
rect 21420 6468 21476 6478
rect 21420 6374 21476 6412
rect 21532 6466 21588 6478
rect 21532 6414 21534 6466
rect 21586 6414 21588 6466
rect 21532 6020 21588 6414
rect 21532 5954 21588 5964
rect 21196 5908 21252 5918
rect 21196 5814 21252 5852
rect 21756 5908 21812 6524
rect 21868 6020 21924 6748
rect 21980 6020 22036 6030
rect 21868 5964 21980 6020
rect 21756 5906 21924 5908
rect 21756 5854 21758 5906
rect 21810 5854 21924 5906
rect 21756 5852 21924 5854
rect 21756 5842 21812 5852
rect 20300 5282 20356 5292
rect 20412 5628 21028 5684
rect 21308 5796 21364 5806
rect 20412 5234 20468 5628
rect 20412 5182 20414 5234
rect 20466 5182 20468 5234
rect 20412 5170 20468 5182
rect 20524 5348 20580 5358
rect 20524 5122 20580 5292
rect 20524 5070 20526 5122
rect 20578 5070 20580 5122
rect 20524 5058 20580 5070
rect 21308 5122 21364 5740
rect 21532 5796 21588 5806
rect 21532 5234 21588 5740
rect 21532 5182 21534 5234
rect 21586 5182 21588 5234
rect 21532 5170 21588 5182
rect 21308 5070 21310 5122
rect 21362 5070 21364 5122
rect 21308 5058 21364 5070
rect 21644 5124 21700 5134
rect 21644 5030 21700 5068
rect 20076 4958 20078 5010
rect 20130 4958 20132 5010
rect 20076 4946 20132 4958
rect 20300 4898 20356 4910
rect 20300 4846 20302 4898
rect 20354 4846 20356 4898
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19292 4398 19294 4450
rect 19346 4398 19348 4450
rect 19292 4386 19348 4398
rect 18508 4286 18510 4338
rect 18562 4286 18564 4338
rect 18508 4274 18564 4286
rect 20300 4228 20356 4846
rect 20300 4162 20356 4172
rect 21084 4340 21140 4350
rect 20860 3668 20916 3678
rect 3836 3332 3892 3342
rect 5516 3332 5572 3342
rect 6972 3332 7028 3342
rect 8540 3332 8596 3342
rect 10108 3332 10164 3342
rect 11676 3332 11732 3342
rect 3612 3330 3892 3332
rect 3612 3278 3838 3330
rect 3890 3278 3892 3330
rect 3612 3276 3892 3278
rect 3612 800 3668 3276
rect 3836 3266 3892 3276
rect 5180 3330 5572 3332
rect 5180 3278 5518 3330
rect 5570 3278 5572 3330
rect 5180 3276 5572 3278
rect 5180 800 5236 3276
rect 5516 3266 5572 3276
rect 6748 3330 7028 3332
rect 6748 3278 6974 3330
rect 7026 3278 7028 3330
rect 6748 3276 7028 3278
rect 6748 800 6804 3276
rect 6972 3266 7028 3276
rect 8316 3330 8596 3332
rect 8316 3278 8542 3330
rect 8594 3278 8596 3330
rect 8316 3276 8596 3278
rect 8316 800 8372 3276
rect 8540 3266 8596 3276
rect 9884 3330 10164 3332
rect 9884 3278 10110 3330
rect 10162 3278 10164 3330
rect 9884 3276 10164 3278
rect 9884 800 9940 3276
rect 10108 3266 10164 3276
rect 11452 3330 11732 3332
rect 11452 3278 11678 3330
rect 11730 3278 11732 3330
rect 11452 3276 11732 3278
rect 11452 800 11508 3276
rect 11676 3266 11732 3276
rect 12572 3332 12628 3342
rect 12572 3330 13076 3332
rect 12572 3278 12574 3330
rect 12626 3278 13076 3330
rect 12572 3276 13076 3278
rect 12572 3266 12628 3276
rect 13020 800 13076 3276
rect 13468 3330 13524 3342
rect 13468 3278 13470 3330
rect 13522 3278 13524 3330
rect 13468 1762 13524 3278
rect 15372 3330 15428 3342
rect 15372 3278 15374 3330
rect 15426 3278 15428 3330
rect 13468 1710 13470 1762
rect 13522 1710 13524 1762
rect 13468 1698 13524 1710
rect 14588 1762 14644 1774
rect 14588 1710 14590 1762
rect 14642 1710 14644 1762
rect 14588 800 14644 1710
rect 3584 0 3696 800
rect 5152 0 5264 800
rect 6720 0 6832 800
rect 8288 0 8400 800
rect 9856 0 9968 800
rect 11424 0 11536 800
rect 12992 0 13104 800
rect 14560 0 14672 800
rect 15372 756 15428 3278
rect 17948 3332 18228 3388
rect 19292 3442 19348 3454
rect 19292 3390 19294 3442
rect 19346 3390 19348 3442
rect 17948 2884 18004 3332
rect 17724 2828 18004 2884
rect 15820 924 16212 980
rect 15820 756 15876 924
rect 16156 800 16212 924
rect 17724 800 17780 2828
rect 19292 800 19348 3390
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20860 800 20916 3612
rect 21084 3554 21140 4284
rect 21868 4338 21924 5852
rect 21980 5010 22036 5964
rect 22204 5572 22260 11454
rect 23212 11394 23268 13692
rect 23212 11342 23214 11394
rect 23266 11342 23268 11394
rect 23212 11330 23268 11342
rect 23324 13074 23380 13086
rect 23324 13022 23326 13074
rect 23378 13022 23380 13074
rect 23324 12964 23380 13022
rect 23772 13074 23828 15092
rect 24220 14644 24276 17838
rect 24332 17780 24388 17790
rect 24332 17686 24388 17724
rect 24444 16884 24500 19180
rect 24892 19170 24948 19180
rect 25004 19796 25060 19806
rect 25004 19012 25060 19740
rect 24668 18956 25060 19012
rect 24668 18674 24724 18956
rect 24668 18622 24670 18674
rect 24722 18622 24724 18674
rect 24668 18610 24724 18622
rect 25228 18452 25284 18462
rect 24444 16790 24500 16828
rect 24556 18340 24612 18350
rect 24556 16436 24612 18284
rect 24220 14578 24276 14588
rect 24444 16380 24612 16436
rect 24892 17444 24948 17454
rect 25228 17444 25284 18396
rect 25340 17890 25396 17902
rect 25340 17838 25342 17890
rect 25394 17838 25396 17890
rect 25340 17778 25396 17838
rect 25340 17726 25342 17778
rect 25394 17726 25396 17778
rect 25340 17714 25396 17726
rect 24892 17442 25284 17444
rect 24892 17390 24894 17442
rect 24946 17390 25284 17442
rect 24892 17388 25284 17390
rect 25452 17444 25508 17454
rect 24444 15540 24500 16380
rect 24108 14532 24164 14542
rect 24108 14438 24164 14476
rect 23772 13022 23774 13074
rect 23826 13022 23828 13074
rect 23772 13010 23828 13022
rect 23884 13746 23940 13758
rect 23884 13694 23886 13746
rect 23938 13694 23940 13746
rect 23884 13636 23940 13694
rect 24444 13748 24500 15484
rect 24444 13682 24500 13692
rect 24556 16098 24612 16110
rect 24556 16046 24558 16098
rect 24610 16046 24612 16098
rect 23324 11394 23380 12908
rect 23324 11342 23326 11394
rect 23378 11342 23380 11394
rect 23324 11330 23380 11342
rect 23436 12068 23492 12078
rect 23436 11394 23492 12012
rect 23436 11342 23438 11394
rect 23490 11342 23492 11394
rect 23436 11330 23492 11342
rect 23772 11956 23828 11966
rect 23772 11394 23828 11900
rect 23772 11342 23774 11394
rect 23826 11342 23828 11394
rect 23772 11330 23828 11342
rect 22764 11170 22820 11182
rect 22764 11118 22766 11170
rect 22818 11118 22820 11170
rect 22764 11060 22820 11118
rect 22764 10994 22820 11004
rect 23436 10052 23492 10062
rect 23436 9940 23492 9996
rect 23436 9938 23716 9940
rect 23436 9886 23438 9938
rect 23490 9886 23716 9938
rect 23436 9884 23716 9886
rect 23436 9874 23492 9884
rect 22652 9714 22708 9726
rect 22652 9662 22654 9714
rect 22706 9662 22708 9714
rect 22652 8932 22708 9662
rect 22652 8866 22708 8876
rect 22764 9602 22820 9614
rect 22764 9550 22766 9602
rect 22818 9550 22820 9602
rect 22428 8484 22484 8494
rect 22428 7476 22484 8428
rect 22764 8258 22820 9550
rect 23324 8930 23380 8942
rect 23324 8878 23326 8930
rect 23378 8878 23380 8930
rect 22764 8206 22766 8258
rect 22818 8206 22820 8258
rect 22764 8194 22820 8206
rect 22988 8260 23044 8270
rect 22988 8166 23044 8204
rect 23212 8258 23268 8270
rect 23212 8206 23214 8258
rect 23266 8206 23268 8258
rect 22540 8148 22596 8158
rect 22540 7700 22596 8092
rect 22988 7700 23044 7710
rect 22540 7698 23044 7700
rect 22540 7646 22990 7698
rect 23042 7646 23044 7698
rect 22540 7644 23044 7646
rect 22988 7634 23044 7644
rect 23212 7588 23268 8206
rect 23324 8034 23380 8878
rect 23324 7982 23326 8034
rect 23378 7982 23380 8034
rect 23324 7970 23380 7982
rect 23660 8148 23716 9884
rect 23884 9938 23940 13580
rect 24332 12964 24388 12974
rect 24220 12962 24388 12964
rect 24220 12910 24334 12962
rect 24386 12910 24388 12962
rect 24220 12908 24388 12910
rect 24108 12740 24164 12750
rect 24108 12646 24164 12684
rect 24108 11620 24164 11630
rect 24220 11620 24276 12908
rect 24332 12898 24388 12908
rect 24108 11618 24276 11620
rect 24108 11566 24110 11618
rect 24162 11566 24276 11618
rect 24108 11564 24276 11566
rect 24108 11554 24164 11564
rect 23884 9886 23886 9938
rect 23938 9886 23940 9938
rect 23884 9874 23940 9886
rect 24220 9828 24276 9838
rect 24108 9826 24276 9828
rect 24108 9774 24222 9826
rect 24274 9774 24276 9826
rect 24108 9772 24276 9774
rect 24108 9044 24164 9772
rect 24220 9762 24276 9772
rect 24108 9042 24276 9044
rect 24108 8990 24110 9042
rect 24162 8990 24276 9042
rect 24108 8988 24276 8990
rect 24108 8978 24164 8988
rect 23772 8370 23828 8382
rect 23772 8318 23774 8370
rect 23826 8318 23828 8370
rect 23772 8260 23828 8318
rect 23772 8194 23828 8204
rect 23884 8372 23940 8382
rect 23660 7588 23716 8092
rect 23884 8146 23940 8316
rect 23884 8094 23886 8146
rect 23938 8094 23940 8146
rect 23884 8082 23940 8094
rect 24108 8370 24164 8382
rect 24108 8318 24110 8370
rect 24162 8318 24164 8370
rect 24108 8036 24164 8318
rect 24108 7970 24164 7980
rect 23772 7588 23828 7598
rect 23660 7586 23828 7588
rect 23660 7534 23774 7586
rect 23826 7534 23828 7586
rect 23660 7532 23828 7534
rect 23212 7522 23268 7532
rect 23772 7522 23828 7532
rect 24108 7588 24164 7598
rect 24108 7494 24164 7532
rect 22652 7476 22708 7486
rect 22428 7420 22652 7476
rect 22428 6916 22484 7420
rect 22652 7382 22708 7420
rect 23324 7474 23380 7486
rect 23324 7422 23326 7474
rect 23378 7422 23380 7474
rect 22428 6850 22484 6860
rect 23324 6804 23380 7422
rect 23996 7474 24052 7486
rect 23996 7422 23998 7474
rect 24050 7422 24052 7474
rect 23324 6748 23604 6804
rect 23548 6692 23604 6748
rect 23548 6636 23716 6692
rect 22428 5796 22484 5806
rect 22428 5702 22484 5740
rect 22204 5506 22260 5516
rect 22316 5684 22372 5694
rect 22316 5122 22372 5628
rect 22764 5572 22820 5582
rect 22540 5348 22596 5358
rect 22540 5346 22708 5348
rect 22540 5294 22542 5346
rect 22594 5294 22708 5346
rect 22540 5292 22708 5294
rect 22540 5282 22596 5292
rect 22316 5070 22318 5122
rect 22370 5070 22372 5122
rect 22316 5058 22372 5070
rect 21980 4958 21982 5010
rect 22034 4958 22036 5010
rect 21980 4946 22036 4958
rect 22428 4900 22484 4910
rect 22428 4898 22596 4900
rect 22428 4846 22430 4898
rect 22482 4846 22596 4898
rect 22428 4844 22596 4846
rect 22428 4834 22484 4844
rect 21868 4286 21870 4338
rect 21922 4286 21924 4338
rect 21868 4274 21924 4286
rect 22428 4452 22484 4462
rect 21420 4228 21476 4238
rect 21420 4134 21476 4172
rect 22092 3668 22148 3678
rect 22092 3574 22148 3612
rect 21084 3502 21086 3554
rect 21138 3502 21140 3554
rect 21084 3490 21140 3502
rect 22428 800 22484 4396
rect 22540 4450 22596 4844
rect 22540 4398 22542 4450
rect 22594 4398 22596 4450
rect 22540 4386 22596 4398
rect 22652 3780 22708 5292
rect 22764 5122 22820 5516
rect 23660 5348 23716 6636
rect 22764 5070 22766 5122
rect 22818 5070 22820 5122
rect 22764 5058 22820 5070
rect 23436 5236 23492 5246
rect 23436 5122 23492 5180
rect 23436 5070 23438 5122
rect 23490 5070 23492 5122
rect 23436 5058 23492 5070
rect 23548 5234 23604 5246
rect 23548 5182 23550 5234
rect 23602 5182 23604 5234
rect 23548 5124 23604 5182
rect 23660 5124 23716 5292
rect 23996 6132 24052 7422
rect 24220 6580 24276 8988
rect 24556 8372 24612 16046
rect 24668 16100 24724 16110
rect 24668 14642 24724 16044
rect 24668 14590 24670 14642
rect 24722 14590 24724 14642
rect 24668 14578 24724 14590
rect 24780 15316 24836 15326
rect 24668 12292 24724 12302
rect 24668 12066 24724 12236
rect 24668 12014 24670 12066
rect 24722 12014 24724 12066
rect 24668 12002 24724 12014
rect 24780 9268 24836 15260
rect 24892 13636 24948 17388
rect 25340 17108 25396 17118
rect 25228 16884 25284 16894
rect 25228 16098 25284 16828
rect 25228 16046 25230 16098
rect 25282 16046 25284 16098
rect 25228 16034 25284 16046
rect 25340 16882 25396 17052
rect 25340 16830 25342 16882
rect 25394 16830 25396 16882
rect 25340 15148 25396 16830
rect 25452 15316 25508 17388
rect 25564 16660 25620 19966
rect 25676 19346 25732 20076
rect 25900 20066 25956 20076
rect 26796 20020 26852 25116
rect 27020 23828 27076 23838
rect 27020 23734 27076 23772
rect 27132 23380 27188 26852
rect 27356 26404 27412 26414
rect 27468 26404 27524 28364
rect 27580 27858 27636 28588
rect 27580 27806 27582 27858
rect 27634 27806 27636 27858
rect 27580 27794 27636 27806
rect 27692 27746 27748 28812
rect 27804 28420 27860 28430
rect 27804 27858 27860 28364
rect 27916 28418 27972 28430
rect 27916 28366 27918 28418
rect 27970 28366 27972 28418
rect 27916 28196 27972 28366
rect 27916 28130 27972 28140
rect 28028 28082 28084 29708
rect 28252 28532 28308 29934
rect 28476 29540 28532 30940
rect 28476 29474 28532 29484
rect 28588 29316 28644 31724
rect 28252 28466 28308 28476
rect 28364 29260 28644 29316
rect 28028 28030 28030 28082
rect 28082 28030 28084 28082
rect 28028 28018 28084 28030
rect 27804 27806 27806 27858
rect 27858 27806 27860 27858
rect 27804 27794 27860 27806
rect 27692 27694 27694 27746
rect 27746 27694 27748 27746
rect 27692 27682 27748 27694
rect 27356 26402 27524 26404
rect 27356 26350 27358 26402
rect 27410 26350 27524 26402
rect 27356 26348 27524 26350
rect 28028 26852 28084 26862
rect 27356 26338 27412 26348
rect 28028 25732 28084 26796
rect 27692 25730 28084 25732
rect 27692 25678 28030 25730
rect 28082 25678 28084 25730
rect 27692 25676 28084 25678
rect 27244 25506 27300 25518
rect 27244 25454 27246 25506
rect 27298 25454 27300 25506
rect 27244 24052 27300 25454
rect 27244 23938 27300 23996
rect 27244 23886 27246 23938
rect 27298 23886 27300 23938
rect 27244 23874 27300 23886
rect 27580 23940 27636 23950
rect 27356 23716 27412 23726
rect 27356 23622 27412 23660
rect 27468 23714 27524 23726
rect 27468 23662 27470 23714
rect 27522 23662 27524 23714
rect 27468 23604 27524 23662
rect 27468 23380 27524 23548
rect 27132 23314 27188 23324
rect 27244 23324 27524 23380
rect 27132 23156 27188 23166
rect 27244 23156 27300 23324
rect 27132 23154 27300 23156
rect 27132 23102 27134 23154
rect 27186 23102 27300 23154
rect 27132 23100 27300 23102
rect 27132 23090 27188 23100
rect 27468 23044 27524 23054
rect 27580 23044 27636 23884
rect 27692 23938 27748 25676
rect 28028 25666 28084 25676
rect 27804 25396 27860 25406
rect 27804 25302 27860 25340
rect 27916 25282 27972 25294
rect 27916 25230 27918 25282
rect 27970 25230 27972 25282
rect 27916 24052 27972 25230
rect 27916 23986 27972 23996
rect 27692 23886 27694 23938
rect 27746 23886 27748 23938
rect 27692 23874 27748 23886
rect 28140 23940 28196 23950
rect 28140 23846 28196 23884
rect 28028 23714 28084 23726
rect 28028 23662 28030 23714
rect 28082 23662 28084 23714
rect 28028 23156 28084 23662
rect 28028 23090 28084 23100
rect 27468 23042 27636 23044
rect 27468 22990 27470 23042
rect 27522 22990 27636 23042
rect 27468 22988 27636 22990
rect 27468 22978 27524 22988
rect 27356 22148 27412 22158
rect 27132 22146 27412 22148
rect 27132 22094 27358 22146
rect 27410 22094 27412 22146
rect 27132 22092 27412 22094
rect 27132 21026 27188 22092
rect 27356 22082 27412 22092
rect 27468 22146 27524 22158
rect 27468 22094 27470 22146
rect 27522 22094 27524 22146
rect 27356 21700 27412 21710
rect 27468 21700 27524 22094
rect 27580 22146 27636 22158
rect 27804 22148 27860 22158
rect 27580 22094 27582 22146
rect 27634 22094 27636 22146
rect 27580 21812 27636 22094
rect 27580 21746 27636 21756
rect 27692 22092 27804 22148
rect 27356 21698 27524 21700
rect 27356 21646 27358 21698
rect 27410 21646 27524 21698
rect 27356 21644 27524 21646
rect 27356 21634 27412 21644
rect 27692 21588 27748 22092
rect 27804 22054 27860 22092
rect 27132 20974 27134 21026
rect 27186 20974 27188 21026
rect 27132 20962 27188 20974
rect 27468 21532 27748 21588
rect 28028 21586 28084 21598
rect 28028 21534 28030 21586
rect 28082 21534 28084 21586
rect 26796 19926 26852 19964
rect 25676 19294 25678 19346
rect 25730 19294 25732 19346
rect 25676 19282 25732 19294
rect 26348 19908 26404 19918
rect 26348 18452 26404 19852
rect 26348 18386 26404 18396
rect 27468 18340 27524 21532
rect 27804 21476 27860 21486
rect 27804 20802 27860 21420
rect 27804 20750 27806 20802
rect 27858 20750 27860 20802
rect 27804 20738 27860 20750
rect 27580 20690 27636 20702
rect 27580 20638 27582 20690
rect 27634 20638 27636 20690
rect 27580 20244 27636 20638
rect 27580 20178 27636 20188
rect 27692 20690 27748 20702
rect 27692 20638 27694 20690
rect 27746 20638 27748 20690
rect 27692 20020 27748 20638
rect 27692 19954 27748 19964
rect 27468 18274 27524 18284
rect 27804 19346 27860 19358
rect 27804 19294 27806 19346
rect 27858 19294 27860 19346
rect 25788 17780 25844 17790
rect 25788 17666 25844 17724
rect 27692 17780 27748 17790
rect 25788 17614 25790 17666
rect 25842 17614 25844 17666
rect 25788 17602 25844 17614
rect 26348 17666 26404 17678
rect 26348 17614 26350 17666
rect 26402 17614 26404 17666
rect 25676 17554 25732 17566
rect 25676 17502 25678 17554
rect 25730 17502 25732 17554
rect 25676 16884 25732 17502
rect 26348 17556 26404 17614
rect 26348 17490 26404 17500
rect 26908 17668 26964 17678
rect 26908 17106 26964 17612
rect 26908 17054 26910 17106
rect 26962 17054 26964 17106
rect 26908 17042 26964 17054
rect 27132 17666 27188 17678
rect 27132 17614 27134 17666
rect 27186 17614 27188 17666
rect 26012 16884 26068 16894
rect 25676 16882 26068 16884
rect 25676 16830 26014 16882
rect 26066 16830 26068 16882
rect 25676 16828 26068 16830
rect 26012 16818 26068 16828
rect 26236 16772 26292 16782
rect 26124 16770 26292 16772
rect 26124 16718 26238 16770
rect 26290 16718 26292 16770
rect 26124 16716 26292 16718
rect 25676 16660 25732 16670
rect 25564 16658 25732 16660
rect 25564 16606 25678 16658
rect 25730 16606 25732 16658
rect 25564 16604 25732 16606
rect 25676 16594 25732 16604
rect 26124 16212 26180 16716
rect 26236 16706 26292 16716
rect 25900 16156 26180 16212
rect 26908 16548 26964 16558
rect 25900 15652 25956 16156
rect 26012 15988 26068 15998
rect 26012 15986 26180 15988
rect 26012 15934 26014 15986
rect 26066 15934 26180 15986
rect 26012 15932 26180 15934
rect 26012 15922 26068 15932
rect 25900 15596 26068 15652
rect 26012 15540 26068 15596
rect 25564 15316 25620 15326
rect 25452 15314 25620 15316
rect 25452 15262 25566 15314
rect 25618 15262 25620 15314
rect 25452 15260 25620 15262
rect 25564 15250 25620 15260
rect 25900 15316 25956 15326
rect 25228 15092 25396 15148
rect 25788 15204 25844 15242
rect 25788 15138 25844 15148
rect 25004 14644 25060 14654
rect 25004 14550 25060 14588
rect 24892 13570 24948 13580
rect 25228 12516 25284 15092
rect 25900 13972 25956 15260
rect 26012 15314 26068 15484
rect 26124 15426 26180 15932
rect 26124 15374 26126 15426
rect 26178 15374 26180 15426
rect 26124 15362 26180 15374
rect 26908 15426 26964 16492
rect 27132 16212 27188 17614
rect 27692 17666 27748 17724
rect 27692 17614 27694 17666
rect 27746 17614 27748 17666
rect 27692 17602 27748 17614
rect 26908 15374 26910 15426
rect 26962 15374 26964 15426
rect 26012 15262 26014 15314
rect 26066 15262 26068 15314
rect 26012 15148 26068 15262
rect 26236 15204 26292 15214
rect 26460 15204 26516 15214
rect 26292 15202 26516 15204
rect 26292 15150 26462 15202
rect 26514 15150 26516 15202
rect 26292 15148 26516 15150
rect 26012 15092 26180 15148
rect 25900 13970 26068 13972
rect 25900 13918 25902 13970
rect 25954 13918 26068 13970
rect 25900 13916 26068 13918
rect 25900 13906 25956 13916
rect 25340 13636 25396 13646
rect 25340 13542 25396 13580
rect 26012 12964 26068 13916
rect 25564 12962 26068 12964
rect 25564 12910 26014 12962
rect 26066 12910 26068 12962
rect 25564 12908 26068 12910
rect 26124 12964 26180 15092
rect 26236 13746 26292 15148
rect 26460 15138 26516 15148
rect 26908 15148 26964 15374
rect 27020 15876 27076 15886
rect 27020 15426 27076 15820
rect 27020 15374 27022 15426
rect 27074 15374 27076 15426
rect 27020 15362 27076 15374
rect 27132 15426 27188 16156
rect 27244 17556 27300 17566
rect 27244 15876 27300 17500
rect 27804 17556 27860 19294
rect 28028 18564 28084 21534
rect 28364 20804 28420 29260
rect 28476 28642 28532 28654
rect 28476 28590 28478 28642
rect 28530 28590 28532 28642
rect 28476 28084 28532 28590
rect 28588 28530 28644 28542
rect 28588 28478 28590 28530
rect 28642 28478 28644 28530
rect 28588 28420 28644 28478
rect 28588 28354 28644 28364
rect 28476 28018 28532 28028
rect 28700 26908 28756 33292
rect 28812 32564 28868 32574
rect 29036 32564 29092 32574
rect 28812 32470 28868 32508
rect 28924 32562 29092 32564
rect 28924 32510 29038 32562
rect 29090 32510 29092 32562
rect 28924 32508 29092 32510
rect 28924 30100 28980 32508
rect 29036 32498 29092 32508
rect 29148 31778 29204 33852
rect 29260 33346 29316 34412
rect 29708 34242 29764 34636
rect 29708 34190 29710 34242
rect 29762 34190 29764 34242
rect 29708 34178 29764 34190
rect 29484 33460 29540 33470
rect 29484 33366 29540 33404
rect 29260 33294 29262 33346
rect 29314 33294 29316 33346
rect 29260 33282 29316 33294
rect 29372 33348 29428 33358
rect 29372 33254 29428 33292
rect 29820 33346 29876 35532
rect 30492 35476 30548 35644
rect 30492 35410 30548 35420
rect 30604 35698 30660 35710
rect 30604 35646 30606 35698
rect 30658 35646 30660 35698
rect 30604 35364 30660 35646
rect 30716 35700 30772 35710
rect 30716 35606 30772 35644
rect 31052 35700 31108 35710
rect 31052 35606 31108 35644
rect 31164 35476 31220 37212
rect 30604 35298 30660 35308
rect 31052 35420 31220 35476
rect 29932 34804 29988 34814
rect 29932 34132 29988 34748
rect 29932 34066 29988 34076
rect 29820 33294 29822 33346
rect 29874 33294 29876 33346
rect 29820 33282 29876 33294
rect 30268 33570 30324 33582
rect 30268 33518 30270 33570
rect 30322 33518 30324 33570
rect 29596 33122 29652 33134
rect 29596 33070 29598 33122
rect 29650 33070 29652 33122
rect 29596 32900 29652 33070
rect 29372 32562 29428 32574
rect 29372 32510 29374 32562
rect 29426 32510 29428 32562
rect 29260 32450 29316 32462
rect 29260 32398 29262 32450
rect 29314 32398 29316 32450
rect 29260 32004 29316 32398
rect 29372 32228 29428 32510
rect 29372 32162 29428 32172
rect 29596 32116 29652 32844
rect 30268 33012 30324 33518
rect 30716 33570 30772 33582
rect 30716 33518 30718 33570
rect 30770 33518 30772 33570
rect 30716 33458 30772 33518
rect 30716 33406 30718 33458
rect 30770 33406 30772 33458
rect 30716 33394 30772 33406
rect 30268 32786 30324 32956
rect 30268 32734 30270 32786
rect 30322 32734 30324 32786
rect 30268 32722 30324 32734
rect 30380 33236 30436 33246
rect 30380 33122 30436 33180
rect 30380 33070 30382 33122
rect 30434 33070 30436 33122
rect 30380 32788 30436 33070
rect 30380 32722 30436 32732
rect 29820 32676 29876 32686
rect 29820 32582 29876 32620
rect 29596 32060 30100 32116
rect 29260 31948 29988 32004
rect 29932 31890 29988 31948
rect 29932 31838 29934 31890
rect 29986 31838 29988 31890
rect 29932 31826 29988 31838
rect 29148 31726 29150 31778
rect 29202 31726 29204 31778
rect 29148 31714 29204 31726
rect 29036 31556 29092 31566
rect 29036 31106 29092 31500
rect 30044 31220 30100 32060
rect 29036 31054 29038 31106
rect 29090 31054 29092 31106
rect 29036 31042 29092 31054
rect 29932 31164 30100 31220
rect 30268 31668 30324 31678
rect 28924 30034 28980 30044
rect 29372 29316 29428 29326
rect 29148 28642 29204 28654
rect 29148 28590 29150 28642
rect 29202 28590 29204 28642
rect 29148 28420 29204 28590
rect 29260 28532 29316 28542
rect 29260 28438 29316 28476
rect 29148 27858 29204 28364
rect 29372 28084 29428 29260
rect 29148 27806 29150 27858
rect 29202 27806 29204 27858
rect 29148 27748 29204 27806
rect 29148 27682 29204 27692
rect 29260 28082 29428 28084
rect 29260 28030 29374 28082
rect 29426 28030 29428 28082
rect 29260 28028 29428 28030
rect 28700 26852 28868 26908
rect 28812 26740 28868 26852
rect 28812 26674 28868 26684
rect 28924 26180 28980 26190
rect 28476 25396 28532 25406
rect 28476 25302 28532 25340
rect 28588 25172 28644 25182
rect 28588 24834 28644 25116
rect 28588 24782 28590 24834
rect 28642 24782 28644 24834
rect 28588 24770 28644 24782
rect 28476 23828 28532 23838
rect 28476 23734 28532 23772
rect 28588 23716 28644 23726
rect 28588 23622 28644 23660
rect 28924 22932 28980 26124
rect 29148 23940 29204 23950
rect 29148 23846 29204 23884
rect 29260 23268 29316 28028
rect 29372 28018 29428 28028
rect 29484 28532 29540 28542
rect 29484 27972 29540 28476
rect 29820 27972 29876 27982
rect 29484 27970 29876 27972
rect 29484 27918 29486 27970
rect 29538 27918 29822 27970
rect 29874 27918 29876 27970
rect 29484 27916 29876 27918
rect 29484 27906 29540 27916
rect 29820 27906 29876 27916
rect 29596 27748 29652 27758
rect 29596 26514 29652 27692
rect 29596 26462 29598 26514
rect 29650 26462 29652 26514
rect 29596 26450 29652 26462
rect 29708 27636 29764 27646
rect 29708 25284 29764 27580
rect 29596 25282 29764 25284
rect 29596 25230 29710 25282
rect 29762 25230 29764 25282
rect 29596 25228 29764 25230
rect 29372 24052 29428 24062
rect 29372 23938 29428 23996
rect 29372 23886 29374 23938
rect 29426 23886 29428 23938
rect 29372 23874 29428 23886
rect 29596 23938 29652 25228
rect 29708 25218 29764 25228
rect 29820 26964 29876 27002
rect 29596 23886 29598 23938
rect 29650 23886 29652 23938
rect 29596 23874 29652 23886
rect 29820 23938 29876 26908
rect 29932 26908 29988 31164
rect 30268 30324 30324 31612
rect 31052 31444 31108 35420
rect 31164 34580 31220 34590
rect 31164 33458 31220 34524
rect 31164 33406 31166 33458
rect 31218 33406 31220 33458
rect 31164 33124 31220 33406
rect 31276 33460 31332 38612
rect 31388 37940 31444 38670
rect 31500 38668 31556 40124
rect 31612 39732 31668 40574
rect 31948 40516 32004 41132
rect 32284 41122 32340 41132
rect 32508 41122 32564 41132
rect 32844 41122 32900 41132
rect 33292 41186 33348 41692
rect 33292 41134 33294 41186
rect 33346 41134 33348 41186
rect 33292 41122 33348 41134
rect 32956 41074 33012 41086
rect 32956 41022 32958 41074
rect 33010 41022 33012 41074
rect 32060 40964 32116 40974
rect 32060 40870 32116 40908
rect 32172 40962 32228 40974
rect 32172 40910 32174 40962
rect 32226 40910 32228 40962
rect 31836 40460 32004 40516
rect 32172 40516 32228 40910
rect 32508 40964 32564 40974
rect 32732 40964 32788 40974
rect 32396 40628 32452 40638
rect 32396 40534 32452 40572
rect 32284 40516 32340 40526
rect 32172 40514 32340 40516
rect 32172 40462 32286 40514
rect 32338 40462 32340 40514
rect 32172 40460 32340 40462
rect 31836 40180 31892 40460
rect 32060 40404 32116 40414
rect 32172 40404 32228 40460
rect 32284 40450 32340 40460
rect 32060 40402 32228 40404
rect 32060 40350 32062 40402
rect 32114 40350 32228 40402
rect 32060 40348 32228 40350
rect 32060 40338 32116 40348
rect 31836 40114 31892 40124
rect 31948 40292 32004 40302
rect 31836 39732 31892 39742
rect 31612 39730 31892 39732
rect 31612 39678 31838 39730
rect 31890 39678 31892 39730
rect 31612 39676 31892 39678
rect 31836 39666 31892 39676
rect 31948 39058 32004 40236
rect 32396 40180 32452 40190
rect 32060 40178 32452 40180
rect 32060 40126 32398 40178
rect 32450 40126 32452 40178
rect 32060 40124 32452 40126
rect 32060 39842 32116 40124
rect 32396 40114 32452 40124
rect 32060 39790 32062 39842
rect 32114 39790 32116 39842
rect 32060 39778 32116 39790
rect 31948 39006 31950 39058
rect 32002 39006 32004 39058
rect 31948 38994 32004 39006
rect 32284 39618 32340 39630
rect 32284 39566 32286 39618
rect 32338 39566 32340 39618
rect 31724 38946 31780 38958
rect 31724 38894 31726 38946
rect 31778 38894 31780 38946
rect 31612 38836 31668 38846
rect 31724 38836 31780 38894
rect 32172 38948 32228 38958
rect 32172 38854 32228 38892
rect 31668 38780 31780 38836
rect 31948 38836 32004 38846
rect 31612 38770 31668 38780
rect 31948 38668 32004 38780
rect 31500 38612 31668 38668
rect 31948 38612 32116 38668
rect 31388 37874 31444 37884
rect 31500 37826 31556 37838
rect 31500 37774 31502 37826
rect 31554 37774 31556 37826
rect 31500 36260 31556 37774
rect 31500 36194 31556 36204
rect 31388 35812 31444 35822
rect 31388 35718 31444 35756
rect 31500 35588 31556 35598
rect 31500 35364 31556 35532
rect 31500 35298 31556 35308
rect 31612 33570 31668 38612
rect 32060 38050 32116 38612
rect 32284 38610 32340 39566
rect 32396 39396 32452 39406
rect 32396 38946 32452 39340
rect 32396 38894 32398 38946
rect 32450 38894 32452 38946
rect 32396 38882 32452 38894
rect 32508 38668 32564 40908
rect 32620 40908 32732 40964
rect 32620 39284 32676 40908
rect 32732 40898 32788 40908
rect 32956 40740 33012 41022
rect 33404 41076 33460 42252
rect 33516 41524 33572 42476
rect 33964 42308 34020 43486
rect 34524 43538 34580 43708
rect 35420 43762 35476 44044
rect 35868 44034 35924 44044
rect 36204 44100 36260 44110
rect 36204 44098 36484 44100
rect 36204 44046 36206 44098
rect 36258 44046 36484 44098
rect 36204 44044 36484 44046
rect 36204 44034 36260 44044
rect 35420 43710 35422 43762
rect 35474 43710 35476 43762
rect 34524 43486 34526 43538
rect 34578 43486 34580 43538
rect 34524 43474 34580 43486
rect 34748 43540 34804 43550
rect 34748 43446 34804 43484
rect 34972 43538 35028 43550
rect 34972 43486 34974 43538
rect 35026 43486 35028 43538
rect 34972 43428 35028 43486
rect 35308 43428 35364 43438
rect 34972 43426 35364 43428
rect 34972 43374 35310 43426
rect 35362 43374 35364 43426
rect 34972 43372 35364 43374
rect 35308 43362 35364 43372
rect 34412 43316 34468 43326
rect 34300 43314 34468 43316
rect 34300 43262 34414 43314
rect 34466 43262 34468 43314
rect 34300 43260 34468 43262
rect 34300 42866 34356 43260
rect 34412 43250 34468 43260
rect 34524 43316 34580 43326
rect 34300 42814 34302 42866
rect 34354 42814 34356 42866
rect 34300 42802 34356 42814
rect 33964 42242 34020 42252
rect 33964 42084 34020 42094
rect 33516 41468 33796 41524
rect 33740 41188 33796 41468
rect 33740 41094 33796 41132
rect 33404 41010 33460 41020
rect 33852 41076 33908 41086
rect 33852 40982 33908 41020
rect 33516 40962 33572 40974
rect 33516 40910 33518 40962
rect 33570 40910 33572 40962
rect 33516 40740 33572 40910
rect 33628 40964 33684 40974
rect 33628 40962 33796 40964
rect 33628 40910 33630 40962
rect 33682 40910 33796 40962
rect 33628 40908 33796 40910
rect 33628 40898 33684 40908
rect 32956 40684 33572 40740
rect 32732 39508 32788 39518
rect 32956 39508 33012 39518
rect 32732 39506 33012 39508
rect 32732 39454 32734 39506
rect 32786 39454 32958 39506
rect 33010 39454 33012 39506
rect 32732 39452 33012 39454
rect 32732 39442 32788 39452
rect 32956 39442 33012 39452
rect 33068 39394 33124 39406
rect 33068 39342 33070 39394
rect 33122 39342 33124 39394
rect 32620 39228 32788 39284
rect 32284 38558 32286 38610
rect 32338 38558 32340 38610
rect 32284 38546 32340 38558
rect 32396 38612 32564 38668
rect 32620 39060 32676 39070
rect 32396 38388 32452 38612
rect 32284 38332 32452 38388
rect 32060 37998 32062 38050
rect 32114 37998 32116 38050
rect 32060 37986 32116 37998
rect 32172 38164 32228 38174
rect 32172 37938 32228 38108
rect 32172 37886 32174 37938
rect 32226 37886 32228 37938
rect 32172 37874 32228 37886
rect 32060 37156 32116 37166
rect 32060 37062 32116 37100
rect 31948 36482 32004 36494
rect 31948 36430 31950 36482
rect 32002 36430 32004 36482
rect 31724 35698 31780 35710
rect 31724 35646 31726 35698
rect 31778 35646 31780 35698
rect 31724 35364 31780 35646
rect 31724 35298 31780 35308
rect 31836 35700 31892 35710
rect 31836 35028 31892 35644
rect 31724 34972 31892 35028
rect 31724 34020 31780 34972
rect 31836 34804 31892 34814
rect 31948 34804 32004 36430
rect 32060 35924 32116 35934
rect 32284 35924 32340 38332
rect 32508 38274 32564 38286
rect 32508 38222 32510 38274
rect 32562 38222 32564 38274
rect 32396 38052 32452 38062
rect 32508 38052 32564 38222
rect 32396 38050 32564 38052
rect 32396 37998 32398 38050
rect 32450 37998 32564 38050
rect 32396 37996 32564 37998
rect 32396 37986 32452 37996
rect 32620 37156 32676 39004
rect 32732 38668 32788 39228
rect 33068 38836 33124 39342
rect 33292 38946 33348 38958
rect 33292 38894 33294 38946
rect 33346 38894 33348 38946
rect 33180 38836 33236 38846
rect 33068 38834 33236 38836
rect 33068 38782 33182 38834
rect 33234 38782 33236 38834
rect 33068 38780 33236 38782
rect 33180 38770 33236 38780
rect 33292 38836 33348 38894
rect 32732 38612 33012 38668
rect 32956 38274 33012 38612
rect 32956 38222 32958 38274
rect 33010 38222 33012 38274
rect 32956 38210 33012 38222
rect 32732 38164 32788 38174
rect 32732 38070 32788 38108
rect 33180 38164 33236 38174
rect 33292 38164 33348 38780
rect 33180 38162 33348 38164
rect 33180 38110 33182 38162
rect 33234 38110 33348 38162
rect 33180 38108 33348 38110
rect 33180 38098 33236 38108
rect 32060 35922 32340 35924
rect 32060 35870 32062 35922
rect 32114 35870 32340 35922
rect 32060 35868 32340 35870
rect 32508 37100 32676 37156
rect 33180 37156 33236 37166
rect 32060 35858 32116 35868
rect 32172 35700 32228 35710
rect 32172 35606 32228 35644
rect 32172 35476 32228 35486
rect 31892 34748 32004 34804
rect 32060 35364 32116 35374
rect 31836 34738 31892 34748
rect 31836 34020 31892 34030
rect 31724 34018 31892 34020
rect 31724 33966 31838 34018
rect 31890 33966 31892 34018
rect 31724 33964 31892 33966
rect 31836 33954 31892 33964
rect 31612 33518 31614 33570
rect 31666 33518 31668 33570
rect 31612 33506 31668 33518
rect 31276 33394 31332 33404
rect 32060 33458 32116 35308
rect 32172 34354 32228 35420
rect 32172 34302 32174 34354
rect 32226 34302 32228 34354
rect 32172 34290 32228 34302
rect 32396 34130 32452 34142
rect 32396 34078 32398 34130
rect 32450 34078 32452 34130
rect 32060 33406 32062 33458
rect 32114 33406 32116 33458
rect 32060 33394 32116 33406
rect 32172 33908 32228 33918
rect 31164 33058 31220 33068
rect 31612 33124 31668 33134
rect 32060 33124 32116 33134
rect 31612 33122 32116 33124
rect 31612 33070 31614 33122
rect 31666 33070 32062 33122
rect 32114 33070 32116 33122
rect 31612 33068 32116 33070
rect 31612 33058 31668 33068
rect 32060 32116 32116 33068
rect 32060 32050 32116 32060
rect 32060 31892 32116 31902
rect 31612 31890 32116 31892
rect 31612 31838 32062 31890
rect 32114 31838 32116 31890
rect 31612 31836 32116 31838
rect 31164 31444 31220 31454
rect 31052 31388 31164 31444
rect 31164 31378 31220 31388
rect 31612 31106 31668 31836
rect 31612 31054 31614 31106
rect 31666 31054 31668 31106
rect 31612 31042 31668 31054
rect 31724 30994 31780 31006
rect 31724 30942 31726 30994
rect 31778 30942 31780 30994
rect 31164 30882 31220 30894
rect 31164 30830 31166 30882
rect 31218 30830 31220 30882
rect 31052 30324 31108 30334
rect 30268 30322 30548 30324
rect 30268 30270 30270 30322
rect 30322 30270 30548 30322
rect 30268 30268 30548 30270
rect 30268 30258 30324 30268
rect 30492 30212 30548 30268
rect 30716 30212 30772 30222
rect 30492 30210 30996 30212
rect 30492 30158 30718 30210
rect 30770 30158 30996 30210
rect 30492 30156 30996 30158
rect 30716 30146 30772 30156
rect 30380 30098 30436 30110
rect 30380 30046 30382 30098
rect 30434 30046 30436 30098
rect 30380 29988 30436 30046
rect 30268 29932 30380 29988
rect 30268 28420 30324 29932
rect 30380 29894 30436 29932
rect 30828 29986 30884 29998
rect 30828 29934 30830 29986
rect 30882 29934 30884 29986
rect 30604 28420 30660 28430
rect 30268 28354 30324 28364
rect 30492 28418 30660 28420
rect 30492 28366 30606 28418
rect 30658 28366 30660 28418
rect 30492 28364 30660 28366
rect 30044 28084 30100 28094
rect 30044 27990 30100 28028
rect 30156 27860 30212 27870
rect 30156 27746 30212 27804
rect 30156 27694 30158 27746
rect 30210 27694 30212 27746
rect 30156 27298 30212 27694
rect 30492 27524 30548 28364
rect 30604 28354 30660 28364
rect 30716 28420 30772 28430
rect 30716 27858 30772 28364
rect 30716 27806 30718 27858
rect 30770 27806 30772 27858
rect 30716 27794 30772 27806
rect 30492 27458 30548 27468
rect 30828 27300 30884 29934
rect 30940 28644 30996 30156
rect 31052 30210 31108 30268
rect 31052 30158 31054 30210
rect 31106 30158 31108 30210
rect 31052 30146 31108 30158
rect 31164 29988 31220 30830
rect 31388 30492 31668 30548
rect 31388 30436 31444 30492
rect 31388 30342 31444 30380
rect 31500 30324 31556 30334
rect 31500 30098 31556 30268
rect 31500 30046 31502 30098
rect 31554 30046 31556 30098
rect 31500 30034 31556 30046
rect 31164 29922 31220 29932
rect 31612 28868 31668 30492
rect 31724 30098 31780 30942
rect 31724 30046 31726 30098
rect 31778 30046 31780 30098
rect 31724 29988 31780 30046
rect 31724 29922 31780 29932
rect 31836 30994 31892 31006
rect 31836 30942 31838 30994
rect 31890 30942 31892 30994
rect 31836 29764 31892 30942
rect 32060 30324 32116 31836
rect 32172 31220 32228 33852
rect 32284 33236 32340 33246
rect 32396 33236 32452 34078
rect 32284 33234 32452 33236
rect 32284 33182 32286 33234
rect 32338 33182 32452 33234
rect 32284 33180 32452 33182
rect 32284 33170 32340 33180
rect 32396 32564 32452 33180
rect 32508 32788 32564 37100
rect 33180 37062 33236 37100
rect 33068 37044 33124 37054
rect 32620 37042 33124 37044
rect 32620 36990 33070 37042
rect 33122 36990 33124 37042
rect 32620 36988 33124 36990
rect 32620 36594 32676 36988
rect 33068 36978 33124 36988
rect 32620 36542 32622 36594
rect 32674 36542 32676 36594
rect 32620 36530 32676 36542
rect 33180 36932 33236 36942
rect 33068 36372 33124 36382
rect 32956 36316 33068 36372
rect 32956 33460 33012 36316
rect 33068 36306 33124 36316
rect 33068 35698 33124 35710
rect 33068 35646 33070 35698
rect 33122 35646 33124 35698
rect 33068 35364 33124 35646
rect 33068 35298 33124 35308
rect 33068 34804 33124 34814
rect 33068 34130 33124 34748
rect 33068 34078 33070 34130
rect 33122 34078 33124 34130
rect 33068 34066 33124 34078
rect 33068 33460 33124 33470
rect 32956 33458 33124 33460
rect 32956 33406 33070 33458
rect 33122 33406 33124 33458
rect 32956 33404 33124 33406
rect 33068 33348 33124 33404
rect 33068 33282 33124 33292
rect 32508 32732 33012 32788
rect 32284 31220 32340 31230
rect 32172 31218 32340 31220
rect 32172 31166 32286 31218
rect 32338 31166 32340 31218
rect 32172 31164 32340 31166
rect 32284 31154 32340 31164
rect 32060 30230 32116 30268
rect 31836 29698 31892 29708
rect 32172 30100 32228 30110
rect 32172 29986 32228 30044
rect 32172 29934 32174 29986
rect 32226 29934 32228 29986
rect 31724 29316 31780 29326
rect 31724 29314 31892 29316
rect 31724 29262 31726 29314
rect 31778 29262 31892 29314
rect 31724 29260 31892 29262
rect 31724 29250 31780 29260
rect 31164 28644 31220 28654
rect 30940 28642 31220 28644
rect 30940 28590 31166 28642
rect 31218 28590 31220 28642
rect 30940 28588 31220 28590
rect 31164 28578 31220 28588
rect 31164 28420 31220 28430
rect 31164 27858 31220 28364
rect 31164 27806 31166 27858
rect 31218 27806 31220 27858
rect 31164 27794 31220 27806
rect 31276 28084 31332 28094
rect 31276 27524 31332 28028
rect 31612 27860 31668 28812
rect 31724 27860 31780 27870
rect 31612 27858 31780 27860
rect 31612 27806 31726 27858
rect 31778 27806 31780 27858
rect 31612 27804 31780 27806
rect 31724 27794 31780 27804
rect 31836 27860 31892 29260
rect 31948 29202 32004 29214
rect 31948 29150 31950 29202
rect 32002 29150 32004 29202
rect 31948 28084 32004 29150
rect 32172 28532 32228 29934
rect 32284 29652 32340 29662
rect 32396 29652 32452 32508
rect 32284 29650 32452 29652
rect 32284 29598 32286 29650
rect 32338 29598 32452 29650
rect 32284 29596 32452 29598
rect 32284 29586 32340 29596
rect 32284 28532 32340 28542
rect 32172 28530 32340 28532
rect 32172 28478 32286 28530
rect 32338 28478 32340 28530
rect 32172 28476 32340 28478
rect 32172 28420 32228 28476
rect 32284 28466 32340 28476
rect 32172 28354 32228 28364
rect 31948 28018 32004 28028
rect 32060 28196 32116 28206
rect 31948 27860 32004 27870
rect 31892 27858 32004 27860
rect 31892 27806 31950 27858
rect 32002 27806 32004 27858
rect 31892 27804 32004 27806
rect 31836 27766 31892 27804
rect 31948 27794 32004 27804
rect 31276 27468 31668 27524
rect 30156 27246 30158 27298
rect 30210 27246 30212 27298
rect 30156 27234 30212 27246
rect 30380 27244 30884 27300
rect 30380 27186 30436 27244
rect 30380 27134 30382 27186
rect 30434 27134 30436 27186
rect 30380 27122 30436 27134
rect 29932 26852 30100 26908
rect 29820 23886 29822 23938
rect 29874 23886 29876 23938
rect 29820 23874 29876 23886
rect 29484 23828 29540 23838
rect 29484 23734 29540 23772
rect 29372 23716 29428 23726
rect 29372 23268 29428 23660
rect 29596 23268 29652 23278
rect 29372 23266 29652 23268
rect 29372 23214 29598 23266
rect 29650 23214 29652 23266
rect 29372 23212 29652 23214
rect 29260 23202 29316 23212
rect 29596 23202 29652 23212
rect 28924 22876 29204 22932
rect 29148 22484 29204 22876
rect 29148 22390 29204 22428
rect 29596 22372 29652 22382
rect 28476 22148 28532 22158
rect 28476 22054 28532 22092
rect 28812 21812 28868 21822
rect 29484 21812 29540 21822
rect 29596 21812 29652 22316
rect 28812 21718 28868 21756
rect 28924 21810 29652 21812
rect 28924 21758 29486 21810
rect 29538 21758 29652 21810
rect 28924 21756 29652 21758
rect 30044 21812 30100 26852
rect 30156 25506 30212 25518
rect 30156 25454 30158 25506
rect 30210 25454 30212 25506
rect 30156 23828 30212 25454
rect 30716 25396 30772 27244
rect 31500 27188 31556 27198
rect 31500 27094 31556 27132
rect 31500 26964 31556 26974
rect 31388 26850 31444 26862
rect 31388 26798 31390 26850
rect 31442 26798 31444 26850
rect 30828 25620 30884 25630
rect 31388 25620 31444 26798
rect 30828 25618 31444 25620
rect 30828 25566 30830 25618
rect 30882 25566 31444 25618
rect 30828 25564 31444 25566
rect 30828 25554 30884 25564
rect 30268 25340 31332 25396
rect 30268 24050 30324 25340
rect 31276 24724 31332 25340
rect 31276 24722 31444 24724
rect 31276 24670 31278 24722
rect 31330 24670 31444 24722
rect 31276 24668 31444 24670
rect 31276 24658 31332 24668
rect 31388 24500 31444 24668
rect 31500 24722 31556 26908
rect 31612 25060 31668 27468
rect 32060 26964 32116 28140
rect 32284 27636 32340 27646
rect 32284 27634 32452 27636
rect 32284 27582 32286 27634
rect 32338 27582 32452 27634
rect 32284 27580 32452 27582
rect 32284 27570 32340 27580
rect 32284 27412 32340 27422
rect 32284 27186 32340 27356
rect 32284 27134 32286 27186
rect 32338 27134 32340 27186
rect 32284 27122 32340 27134
rect 32396 27076 32452 27580
rect 32844 27412 32900 27422
rect 32508 27244 32788 27300
rect 32508 27188 32564 27244
rect 32508 27122 32564 27132
rect 32732 27186 32788 27244
rect 32732 27134 32734 27186
rect 32786 27134 32788 27186
rect 32732 27122 32788 27134
rect 32396 27010 32452 27020
rect 32620 27076 32676 27114
rect 32620 27010 32676 27020
rect 32844 27074 32900 27356
rect 32844 27022 32846 27074
rect 32898 27022 32900 27074
rect 32844 27010 32900 27022
rect 32060 26898 32116 26908
rect 32844 26908 32900 26918
rect 32732 26740 32788 26750
rect 31612 24994 31668 25004
rect 32508 25284 32564 25294
rect 31500 24670 31502 24722
rect 31554 24670 31556 24722
rect 31500 24658 31556 24670
rect 32508 24946 32564 25228
rect 32508 24894 32510 24946
rect 32562 24894 32564 24946
rect 31836 24500 31892 24510
rect 31388 24444 31668 24500
rect 31164 24276 31220 24286
rect 30492 24164 30548 24174
rect 30492 24070 30548 24108
rect 30268 23998 30270 24050
rect 30322 23998 30324 24050
rect 30268 23986 30324 23998
rect 30156 23492 30212 23772
rect 30828 23716 30884 23726
rect 30828 23714 30996 23716
rect 30828 23662 30830 23714
rect 30882 23662 30996 23714
rect 30828 23660 30996 23662
rect 30828 23650 30884 23660
rect 30156 23436 30324 23492
rect 30268 23154 30324 23436
rect 30268 23102 30270 23154
rect 30322 23102 30324 23154
rect 30268 23090 30324 23102
rect 30716 23154 30772 23166
rect 30716 23102 30718 23154
rect 30770 23102 30772 23154
rect 30156 21812 30212 21822
rect 30044 21810 30212 21812
rect 30044 21758 30158 21810
rect 30210 21758 30212 21810
rect 30044 21756 30212 21758
rect 28476 21586 28532 21598
rect 28476 21534 28478 21586
rect 28530 21534 28532 21586
rect 28476 21476 28532 21534
rect 28476 21410 28532 21420
rect 28812 21588 28868 21598
rect 28924 21588 28980 21756
rect 29484 21746 29540 21756
rect 28812 21586 28980 21588
rect 28812 21534 28814 21586
rect 28866 21534 28980 21586
rect 28812 21532 28980 21534
rect 29036 21586 29092 21598
rect 29036 21534 29038 21586
rect 29090 21534 29092 21586
rect 28364 20748 28532 20804
rect 28364 20578 28420 20590
rect 28364 20526 28366 20578
rect 28418 20526 28420 20578
rect 28364 20244 28420 20526
rect 28364 20178 28420 20188
rect 28364 20020 28420 20030
rect 28476 20020 28532 20748
rect 28420 19964 28532 20020
rect 28364 19926 28420 19964
rect 28476 18900 28532 19964
rect 28476 18834 28532 18844
rect 27804 17490 27860 17500
rect 27916 18562 28084 18564
rect 27916 18510 28030 18562
rect 28082 18510 28084 18562
rect 27916 18508 28084 18510
rect 27356 17444 27412 17454
rect 27356 17350 27412 17388
rect 27356 16996 27412 17006
rect 27356 16770 27412 16940
rect 27916 16884 27972 18508
rect 28028 18498 28084 18508
rect 28028 17780 28084 17790
rect 28028 17686 28084 17724
rect 28812 17780 28868 21532
rect 29036 20244 29092 21534
rect 29484 21028 29540 21038
rect 29484 20934 29540 20972
rect 29596 20690 29652 20702
rect 29596 20638 29598 20690
rect 29650 20638 29652 20690
rect 29596 20580 29652 20638
rect 29932 20692 29988 20702
rect 30044 20692 30100 21756
rect 30156 21746 30212 21756
rect 29932 20690 30100 20692
rect 29932 20638 29934 20690
rect 29986 20638 30100 20690
rect 29932 20636 30100 20638
rect 30492 21700 30548 21710
rect 29932 20626 29988 20636
rect 29596 20514 29652 20524
rect 30268 20580 30324 20590
rect 30268 20486 30324 20524
rect 29036 20178 29092 20188
rect 29484 20244 29540 20254
rect 29484 19908 29540 20188
rect 30380 20132 30436 20142
rect 29484 19906 29652 19908
rect 29484 19854 29486 19906
rect 29538 19854 29652 19906
rect 29484 19852 29652 19854
rect 29484 19842 29540 19852
rect 29260 19236 29316 19246
rect 29148 19180 29260 19236
rect 29148 19122 29204 19180
rect 29260 19170 29316 19180
rect 29148 19070 29150 19122
rect 29202 19070 29204 19122
rect 29148 19058 29204 19070
rect 29260 19012 29316 19022
rect 29260 19010 29540 19012
rect 29260 18958 29262 19010
rect 29314 18958 29540 19010
rect 29260 18956 29540 18958
rect 29260 18946 29316 18956
rect 28812 17714 28868 17724
rect 29148 17780 29204 17790
rect 29148 17686 29204 17724
rect 28588 17554 28644 17566
rect 28588 17502 28590 17554
rect 28642 17502 28644 17554
rect 28252 17442 28308 17454
rect 28252 17390 28254 17442
rect 28306 17390 28308 17442
rect 27356 16718 27358 16770
rect 27410 16718 27412 16770
rect 27356 16706 27412 16718
rect 27804 16828 27916 16884
rect 27356 15876 27412 15886
rect 27244 15820 27356 15876
rect 27356 15810 27412 15820
rect 27132 15374 27134 15426
rect 27186 15374 27188 15426
rect 27132 15362 27188 15374
rect 27692 15540 27748 15550
rect 27692 15314 27748 15484
rect 27692 15262 27694 15314
rect 27746 15262 27748 15314
rect 27692 15250 27748 15262
rect 26908 15092 27076 15148
rect 26236 13694 26238 13746
rect 26290 13694 26292 13746
rect 26236 13682 26292 13694
rect 26460 14644 26516 14654
rect 26460 13972 26516 14588
rect 27020 14420 27076 15092
rect 27580 15090 27636 15102
rect 27580 15038 27582 15090
rect 27634 15038 27636 15090
rect 27132 14644 27188 14654
rect 27580 14644 27636 15038
rect 27132 14642 27636 14644
rect 27132 14590 27134 14642
rect 27186 14590 27636 14642
rect 27132 14588 27636 14590
rect 27132 14578 27188 14588
rect 27804 14530 27860 16828
rect 27916 16818 27972 16828
rect 28028 16996 28084 17006
rect 27916 15316 27972 15326
rect 27916 15222 27972 15260
rect 28028 15148 28084 16940
rect 28140 16212 28196 16222
rect 28140 16118 28196 16156
rect 28140 15316 28196 15326
rect 28140 15222 28196 15260
rect 27804 14478 27806 14530
rect 27858 14478 27860 14530
rect 27804 14466 27860 14478
rect 27916 15092 28084 15148
rect 27020 14364 27524 14420
rect 26460 13746 26516 13916
rect 27468 13970 27524 14364
rect 27916 14084 27972 15092
rect 28252 14754 28308 17390
rect 28476 17442 28532 17454
rect 28476 17390 28478 17442
rect 28530 17390 28532 17442
rect 28476 16324 28532 17390
rect 28588 16660 28644 17502
rect 29484 16994 29540 18956
rect 29484 16942 29486 16994
rect 29538 16942 29540 16994
rect 29484 16930 29540 16942
rect 28588 16594 28644 16604
rect 29596 16548 29652 19852
rect 30380 19684 30436 20076
rect 30492 19796 30548 21644
rect 30716 21028 30772 23102
rect 30828 22484 30884 22494
rect 30828 21812 30884 22428
rect 30828 21586 30884 21756
rect 30828 21534 30830 21586
rect 30882 21534 30884 21586
rect 30828 21522 30884 21534
rect 30716 20962 30772 20972
rect 30716 20580 30772 20590
rect 30716 20486 30772 20524
rect 30940 20020 30996 23660
rect 31052 21476 31108 21486
rect 31052 21382 31108 21420
rect 31164 21364 31220 24220
rect 31276 23492 31332 23502
rect 31276 23154 31332 23436
rect 31276 23102 31278 23154
rect 31330 23102 31332 23154
rect 31276 22932 31332 23102
rect 31612 23154 31668 24444
rect 31612 23102 31614 23154
rect 31666 23102 31668 23154
rect 31612 23090 31668 23102
rect 31724 24498 31892 24500
rect 31724 24446 31838 24498
rect 31890 24446 31892 24498
rect 31724 24444 31892 24446
rect 31276 22866 31332 22876
rect 31724 22372 31780 24444
rect 31836 24434 31892 24444
rect 31948 23828 32004 23838
rect 31836 23156 31892 23166
rect 31836 23062 31892 23100
rect 31388 22316 31780 22372
rect 31948 22370 32004 23772
rect 32508 23156 32564 24894
rect 32508 23090 32564 23100
rect 31948 22318 31950 22370
rect 32002 22318 32004 22370
rect 31276 22260 31332 22270
rect 31276 22166 31332 22204
rect 31276 21588 31332 21598
rect 31276 21494 31332 21532
rect 31164 21298 31220 21308
rect 31388 20804 31444 22316
rect 31724 22148 31780 22158
rect 31724 21810 31780 22092
rect 31724 21758 31726 21810
rect 31778 21758 31780 21810
rect 31724 21746 31780 21758
rect 31836 21812 31892 21822
rect 31836 21586 31892 21756
rect 31836 21534 31838 21586
rect 31890 21534 31892 21586
rect 31836 21522 31892 21534
rect 30940 19954 30996 19964
rect 31052 20748 31780 20804
rect 30492 19730 30548 19740
rect 30380 19618 30436 19628
rect 31052 19460 31108 20748
rect 30604 19458 31108 19460
rect 30604 19406 31054 19458
rect 31106 19406 31108 19458
rect 30604 19404 31108 19406
rect 30044 19236 30100 19246
rect 30044 19142 30100 19180
rect 30380 19236 30436 19246
rect 30604 19236 30660 19404
rect 31052 19394 31108 19404
rect 31164 20580 31220 20590
rect 30380 19234 30660 19236
rect 30380 19182 30382 19234
rect 30434 19182 30660 19234
rect 30380 19180 30660 19182
rect 30716 19236 30772 19246
rect 31164 19236 31220 20524
rect 31500 19908 31556 19918
rect 31500 19814 31556 19852
rect 30380 19170 30436 19180
rect 29708 19122 29764 19134
rect 29708 19070 29710 19122
rect 29762 19070 29764 19122
rect 29708 16996 29764 19070
rect 30156 19124 30212 19134
rect 30156 19030 30212 19068
rect 29932 19012 29988 19022
rect 29932 18918 29988 18956
rect 29708 16930 29764 16940
rect 30044 18900 30100 18910
rect 29484 16492 29652 16548
rect 29708 16660 29764 16670
rect 28476 16268 29092 16324
rect 28588 16100 28644 16110
rect 28588 16006 28644 16044
rect 28476 15988 28532 15998
rect 28476 15894 28532 15932
rect 29036 15538 29092 16268
rect 29036 15486 29038 15538
rect 29090 15486 29092 15538
rect 29036 15474 29092 15486
rect 29148 16212 29204 16222
rect 29148 15540 29204 16156
rect 29372 16210 29428 16222
rect 29372 16158 29374 16210
rect 29426 16158 29428 16210
rect 29260 16100 29316 16110
rect 29372 16100 29428 16158
rect 29316 16044 29428 16100
rect 29260 16034 29316 16044
rect 29260 15540 29316 15550
rect 29148 15538 29316 15540
rect 29148 15486 29262 15538
rect 29314 15486 29316 15538
rect 29148 15484 29316 15486
rect 29260 15474 29316 15484
rect 28700 15426 28756 15438
rect 28700 15374 28702 15426
rect 28754 15374 28756 15426
rect 28588 15316 28644 15326
rect 28476 15204 28532 15242
rect 28588 15222 28644 15260
rect 28476 15138 28532 15148
rect 28252 14702 28254 14754
rect 28306 14702 28308 14754
rect 27468 13918 27470 13970
rect 27522 13918 27524 13970
rect 27468 13906 27524 13918
rect 27692 14028 27972 14084
rect 28028 14420 28084 14430
rect 26460 13694 26462 13746
rect 26514 13694 26516 13746
rect 26460 13682 26516 13694
rect 27356 13748 27412 13758
rect 26236 12964 26292 12974
rect 26572 12964 26628 12974
rect 26124 12962 26404 12964
rect 26124 12910 26238 12962
rect 26290 12910 26404 12962
rect 26124 12908 26404 12910
rect 25228 12450 25284 12460
rect 25452 12738 25508 12750
rect 25452 12686 25454 12738
rect 25506 12686 25508 12738
rect 25452 12628 25508 12686
rect 25228 11956 25284 11966
rect 25228 11862 25284 11900
rect 25452 10836 25508 12572
rect 25564 12178 25620 12908
rect 26012 12898 26068 12908
rect 26236 12898 26292 12908
rect 25564 12126 25566 12178
rect 25618 12126 25620 12178
rect 25564 12114 25620 12126
rect 25676 12738 25732 12750
rect 25900 12740 25956 12750
rect 25676 12686 25678 12738
rect 25730 12686 25732 12738
rect 25676 12068 25732 12686
rect 25788 12684 25900 12740
rect 25788 12292 25844 12684
rect 25900 12646 25956 12684
rect 26124 12516 26180 12526
rect 26348 12516 26404 12908
rect 26572 12870 26628 12908
rect 26908 12852 26964 12862
rect 26908 12758 26964 12796
rect 27020 12852 27076 12862
rect 27244 12852 27300 12862
rect 27020 12850 27244 12852
rect 27020 12798 27022 12850
rect 27074 12798 27244 12850
rect 27020 12796 27244 12798
rect 27020 12786 27076 12796
rect 27244 12786 27300 12796
rect 26460 12740 26516 12750
rect 26460 12646 26516 12684
rect 26180 12460 26292 12516
rect 26348 12460 26852 12516
rect 26124 12450 26180 12460
rect 26236 12404 26292 12460
rect 26236 12348 26404 12404
rect 25788 12198 25844 12236
rect 25676 12002 25732 12012
rect 26236 12178 26292 12190
rect 26236 12126 26238 12178
rect 26290 12126 26292 12178
rect 26236 12068 26292 12126
rect 26236 12002 26292 12012
rect 25788 11396 25844 11406
rect 25788 11394 26180 11396
rect 25788 11342 25790 11394
rect 25842 11342 26180 11394
rect 25788 11340 26180 11342
rect 25788 11330 25844 11340
rect 25228 10780 25508 10836
rect 25004 10500 25060 10510
rect 25004 9938 25060 10444
rect 25116 10052 25172 10062
rect 25228 10052 25284 10780
rect 25172 9996 25284 10052
rect 25340 10610 25396 10622
rect 25340 10558 25342 10610
rect 25394 10558 25396 10610
rect 25116 9986 25172 9996
rect 25004 9886 25006 9938
rect 25058 9886 25060 9938
rect 25004 9874 25060 9886
rect 24780 9266 25284 9268
rect 24780 9214 24782 9266
rect 24834 9214 25284 9266
rect 24780 9212 25284 9214
rect 24780 9202 24836 9212
rect 25228 9042 25284 9212
rect 25340 9156 25396 10558
rect 25564 10610 25620 10622
rect 25564 10558 25566 10610
rect 25618 10558 25620 10610
rect 25564 9380 25620 10558
rect 25788 10612 25844 10622
rect 25788 10610 26068 10612
rect 25788 10558 25790 10610
rect 25842 10558 26068 10610
rect 25788 10556 26068 10558
rect 25788 10546 25844 10556
rect 25676 10500 25732 10510
rect 25676 10406 25732 10444
rect 25564 9324 25844 9380
rect 25788 9266 25844 9324
rect 25788 9214 25790 9266
rect 25842 9214 25844 9266
rect 25452 9156 25508 9166
rect 25340 9100 25452 9156
rect 25452 9090 25508 9100
rect 25676 9098 25732 9110
rect 25228 8990 25230 9042
rect 25282 8990 25284 9042
rect 25228 8978 25284 8990
rect 25676 9046 25678 9098
rect 25730 9046 25732 9098
rect 25676 8484 25732 9046
rect 24556 7924 24612 8316
rect 25564 8428 25732 8484
rect 25228 8148 25284 8158
rect 25228 8054 25284 8092
rect 25452 8148 25508 8158
rect 24556 7858 24612 7868
rect 24332 7250 24388 7262
rect 24332 7198 24334 7250
rect 24386 7198 24388 7250
rect 24332 6692 24388 7198
rect 24556 7250 24612 7262
rect 24556 7198 24558 7250
rect 24610 7198 24612 7250
rect 24556 6916 24612 7198
rect 25452 7252 25508 8092
rect 25564 8146 25620 8428
rect 25564 8094 25566 8146
rect 25618 8094 25620 8146
rect 25564 8036 25620 8094
rect 25676 8260 25732 8270
rect 25676 8146 25732 8204
rect 25676 8094 25678 8146
rect 25730 8094 25732 8146
rect 25676 8082 25732 8094
rect 25788 8148 25844 9214
rect 26012 9266 26068 10556
rect 26124 9604 26180 11340
rect 26124 9538 26180 9548
rect 26236 9828 26292 9838
rect 26012 9214 26014 9266
rect 26066 9214 26068 9266
rect 25900 9156 25956 9166
rect 25900 9062 25956 9100
rect 26012 8932 26068 9214
rect 26012 8866 26068 8876
rect 25900 8260 25956 8270
rect 26236 8260 26292 9772
rect 25900 8258 26292 8260
rect 25900 8206 25902 8258
rect 25954 8206 26238 8258
rect 26290 8206 26292 8258
rect 25900 8204 26292 8206
rect 25900 8194 25956 8204
rect 26236 8194 26292 8204
rect 25788 8082 25844 8092
rect 25564 7970 25620 7980
rect 25564 7476 25620 7486
rect 26012 7476 26068 7486
rect 25564 7474 25844 7476
rect 25564 7422 25566 7474
rect 25618 7422 25844 7474
rect 25564 7420 25844 7422
rect 25564 7410 25620 7420
rect 25452 7196 25620 7252
rect 24612 6860 24724 6916
rect 24556 6850 24612 6860
rect 24332 6626 24388 6636
rect 24220 6486 24276 6524
rect 23996 6076 24612 6132
rect 23772 5124 23828 5134
rect 23660 5068 23772 5124
rect 23548 5058 23604 5068
rect 23772 5010 23828 5068
rect 23996 5122 24052 6076
rect 24556 5794 24612 6076
rect 24556 5742 24558 5794
rect 24610 5742 24612 5794
rect 24556 5730 24612 5742
rect 24668 5236 24724 6860
rect 24668 5142 24724 5180
rect 24780 6692 24836 6702
rect 23996 5070 23998 5122
rect 24050 5070 24052 5122
rect 23996 5058 24052 5070
rect 24780 5122 24836 6636
rect 25228 6020 25284 6030
rect 25228 5926 25284 5964
rect 25340 5908 25396 5918
rect 25452 5908 25508 5918
rect 25396 5906 25508 5908
rect 25396 5854 25454 5906
rect 25506 5854 25508 5906
rect 25396 5852 25508 5854
rect 25116 5236 25172 5246
rect 25340 5236 25396 5852
rect 25452 5842 25508 5852
rect 24780 5070 24782 5122
rect 24834 5070 24836 5122
rect 24780 5058 24836 5070
rect 24892 5234 25396 5236
rect 24892 5182 25118 5234
rect 25170 5182 25396 5234
rect 24892 5180 25396 5182
rect 23772 4958 23774 5010
rect 23826 4958 23828 5010
rect 23772 4946 23828 4958
rect 23548 4900 23604 4910
rect 23548 4806 23604 4844
rect 24668 4226 24724 4238
rect 24668 4174 24670 4226
rect 24722 4174 24724 4226
rect 22652 3714 22708 3724
rect 24556 3780 24612 3790
rect 24556 3686 24612 3724
rect 24668 3556 24724 4174
rect 24892 3778 24948 5180
rect 25116 5170 25172 5180
rect 25564 4900 25620 7196
rect 25788 5012 25844 7420
rect 26012 6690 26068 7420
rect 26236 7364 26292 7374
rect 26236 7270 26292 7308
rect 26012 6638 26014 6690
rect 26066 6638 26068 6690
rect 26012 6626 26068 6638
rect 26124 6692 26180 6702
rect 26012 5794 26068 5806
rect 26012 5742 26014 5794
rect 26066 5742 26068 5794
rect 25900 5684 25956 5694
rect 25900 5590 25956 5628
rect 26012 5124 26068 5742
rect 25676 4900 25732 4910
rect 25564 4898 25732 4900
rect 25564 4846 25678 4898
rect 25730 4846 25732 4898
rect 25564 4844 25732 4846
rect 25228 4452 25284 4462
rect 25228 4358 25284 4396
rect 24892 3726 24894 3778
rect 24946 3726 24948 3778
rect 24892 3714 24948 3726
rect 25676 3556 25732 4844
rect 25788 4338 25844 4956
rect 25788 4286 25790 4338
rect 25842 4286 25844 4338
rect 25788 4274 25844 4286
rect 25900 5068 26068 5124
rect 26124 5124 26180 6636
rect 25900 4228 25956 5068
rect 26012 4900 26068 4910
rect 26124 4900 26180 5068
rect 26012 4898 26180 4900
rect 26012 4846 26014 4898
rect 26066 4846 26180 4898
rect 26012 4844 26180 4846
rect 26348 5460 26404 12348
rect 26684 12292 26740 12302
rect 26684 12198 26740 12236
rect 26796 12178 26852 12460
rect 26796 12126 26798 12178
rect 26850 12126 26852 12178
rect 26796 12114 26852 12126
rect 26460 12066 26516 12078
rect 26460 12014 26462 12066
rect 26514 12014 26516 12066
rect 26460 11506 26516 12014
rect 26460 11454 26462 11506
rect 26514 11454 26516 11506
rect 26460 11442 26516 11454
rect 27132 9940 27188 9950
rect 27020 9938 27188 9940
rect 27020 9886 27134 9938
rect 27186 9886 27188 9938
rect 27020 9884 27188 9886
rect 26796 9044 26852 9054
rect 26684 9042 26852 9044
rect 26684 8990 26798 9042
rect 26850 8990 26852 9042
rect 26684 8988 26852 8990
rect 26460 8034 26516 8046
rect 26460 7982 26462 8034
rect 26514 7982 26516 8034
rect 26460 6804 26516 7982
rect 26460 6018 26516 6748
rect 26572 7364 26628 7374
rect 26572 6130 26628 7308
rect 26684 6692 26740 8988
rect 26796 8978 26852 8988
rect 27020 9042 27076 9884
rect 27132 9874 27188 9884
rect 27020 8990 27022 9042
rect 27074 8990 27076 9042
rect 27020 8932 27076 8990
rect 27132 9044 27188 9054
rect 27132 8950 27188 8988
rect 27020 8866 27076 8876
rect 26684 6626 26740 6636
rect 26796 8146 26852 8158
rect 26796 8094 26798 8146
rect 26850 8094 26852 8146
rect 26572 6078 26574 6130
rect 26626 6078 26628 6130
rect 26572 6066 26628 6078
rect 26460 5966 26462 6018
rect 26514 5966 26516 6018
rect 26460 5796 26516 5966
rect 26684 6020 26740 6030
rect 26796 6020 26852 8094
rect 27356 6356 27412 13692
rect 27692 13746 27748 14028
rect 28028 13970 28084 14364
rect 28028 13918 28030 13970
rect 28082 13918 28084 13970
rect 28028 13906 28084 13918
rect 27692 13694 27694 13746
rect 27746 13694 27748 13746
rect 27692 13076 27748 13694
rect 27692 13010 27748 13020
rect 27804 13858 27860 13870
rect 27804 13806 27806 13858
rect 27858 13806 27860 13858
rect 27804 12292 27860 13806
rect 28252 13858 28308 14702
rect 28364 14308 28420 14318
rect 28364 14214 28420 14252
rect 28476 14308 28532 14318
rect 28700 14308 28756 15374
rect 29372 15426 29428 16044
rect 29484 15652 29540 16492
rect 29708 16210 29764 16604
rect 29708 16158 29710 16210
rect 29762 16158 29764 16210
rect 29708 16146 29764 16158
rect 29596 15876 29652 15886
rect 29596 15782 29652 15820
rect 29820 15876 29876 15886
rect 29820 15782 29876 15820
rect 29484 15596 29652 15652
rect 29372 15374 29374 15426
rect 29426 15374 29428 15426
rect 29372 15362 29428 15374
rect 28476 14306 28756 14308
rect 28476 14254 28478 14306
rect 28530 14254 28756 14306
rect 28476 14252 28756 14254
rect 29372 14530 29428 14542
rect 29372 14478 29374 14530
rect 29426 14478 29428 14530
rect 28364 13972 28420 13982
rect 28476 13972 28532 14252
rect 28420 13916 28532 13972
rect 28700 13972 28756 13982
rect 29372 13972 29428 14478
rect 28700 13970 29428 13972
rect 28700 13918 28702 13970
rect 28754 13918 29428 13970
rect 28700 13916 29428 13918
rect 29484 14418 29540 14430
rect 29484 14366 29486 14418
rect 29538 14366 29540 14418
rect 28364 13878 28420 13916
rect 28700 13906 28756 13916
rect 28252 13806 28254 13858
rect 28306 13806 28308 13858
rect 28252 13794 28308 13806
rect 28588 13748 28644 13758
rect 28812 13748 28868 13758
rect 28588 13746 28868 13748
rect 28588 13694 28590 13746
rect 28642 13694 28814 13746
rect 28866 13694 28868 13746
rect 28588 13692 28868 13694
rect 28588 13682 28644 13692
rect 28812 13682 28868 13692
rect 29484 13188 29540 14366
rect 29484 13122 29540 13132
rect 29372 13076 29428 13086
rect 29372 12982 29428 13020
rect 29148 12964 29204 12974
rect 29596 12964 29652 15596
rect 30044 15314 30100 18844
rect 30716 18676 30772 19180
rect 31052 19180 31220 19236
rect 31388 19796 31444 19806
rect 30716 18610 30772 18620
rect 30940 19012 30996 19022
rect 30940 18450 30996 18956
rect 30940 18398 30942 18450
rect 30994 18398 30996 18450
rect 30940 18386 30996 18398
rect 31052 18228 31108 19180
rect 30940 18172 31108 18228
rect 31164 18562 31220 18574
rect 31164 18510 31166 18562
rect 31218 18510 31220 18562
rect 30828 17780 30884 17790
rect 30828 16996 30884 17724
rect 30380 16994 30884 16996
rect 30380 16942 30830 16994
rect 30882 16942 30884 16994
rect 30380 16940 30884 16942
rect 30268 16884 30324 16894
rect 30268 16790 30324 16828
rect 30380 16210 30436 16940
rect 30828 16930 30884 16940
rect 30380 16158 30382 16210
rect 30434 16158 30436 16210
rect 30380 16146 30436 16158
rect 30716 16210 30772 16222
rect 30716 16158 30718 16210
rect 30770 16158 30772 16210
rect 30716 15988 30772 16158
rect 30716 15922 30772 15932
rect 30268 15876 30324 15886
rect 30268 15782 30324 15820
rect 30044 15262 30046 15314
rect 30098 15262 30100 15314
rect 30044 15148 30100 15262
rect 29820 15092 30100 15148
rect 30604 15316 30660 15326
rect 29708 14642 29764 14654
rect 29708 14590 29710 14642
rect 29762 14590 29764 14642
rect 29708 13074 29764 14590
rect 29708 13022 29710 13074
rect 29762 13022 29764 13074
rect 29708 13010 29764 13022
rect 27804 12226 27860 12236
rect 29036 12962 29204 12964
rect 29036 12910 29150 12962
rect 29202 12910 29204 12962
rect 29036 12908 29204 12910
rect 29036 12292 29092 12908
rect 29148 12898 29204 12908
rect 29484 12908 29652 12964
rect 29820 12964 29876 15092
rect 30604 14530 30660 15260
rect 30604 14478 30606 14530
rect 30658 14478 30660 14530
rect 30604 14466 30660 14478
rect 30156 14420 30212 14430
rect 30156 14326 30212 14364
rect 29932 14308 29988 14318
rect 29932 13858 29988 14252
rect 29932 13806 29934 13858
rect 29986 13806 29988 13858
rect 29932 13794 29988 13806
rect 30604 13858 30660 13870
rect 30604 13806 30606 13858
rect 30658 13806 30660 13858
rect 30156 13748 30212 13758
rect 30156 13654 30212 13692
rect 29820 12908 30212 12964
rect 29036 12198 29092 12236
rect 29148 12740 29204 12750
rect 28924 12068 28980 12078
rect 28588 12066 28980 12068
rect 28588 12014 28926 12066
rect 28978 12014 28980 12066
rect 28588 12012 28980 12014
rect 28588 11506 28644 12012
rect 28924 12002 28980 12012
rect 28588 11454 28590 11506
rect 28642 11454 28644 11506
rect 28588 11442 28644 11454
rect 29148 10498 29204 12684
rect 29484 11284 29540 12908
rect 29708 12852 29764 12862
rect 29596 12796 29708 12852
rect 29596 12738 29652 12796
rect 29708 12786 29764 12796
rect 29596 12686 29598 12738
rect 29650 12686 29652 12738
rect 29596 12674 29652 12686
rect 29820 12740 29876 12750
rect 29820 12180 29876 12684
rect 29820 12114 29876 12124
rect 29596 11508 29652 11518
rect 30156 11508 30212 12908
rect 30604 12740 30660 13806
rect 30716 13746 30772 13758
rect 30716 13694 30718 13746
rect 30770 13694 30772 13746
rect 30716 12852 30772 13694
rect 30716 12786 30772 12796
rect 30604 12674 30660 12684
rect 30940 12404 30996 18172
rect 31164 17220 31220 18510
rect 31276 17554 31332 17566
rect 31276 17502 31278 17554
rect 31330 17502 31332 17554
rect 31276 17332 31332 17502
rect 31276 17266 31332 17276
rect 31052 17164 31220 17220
rect 31052 17106 31108 17164
rect 31052 17054 31054 17106
rect 31106 17054 31108 17106
rect 31052 15204 31108 17054
rect 31164 16996 31220 17006
rect 31164 16902 31220 16940
rect 31276 16884 31332 16894
rect 31388 16884 31444 19740
rect 31500 19012 31556 19022
rect 31500 18918 31556 18956
rect 31500 18564 31556 18574
rect 31500 18470 31556 18508
rect 31724 18450 31780 20748
rect 31836 20132 31892 20142
rect 31836 19908 31892 20076
rect 31948 20020 32004 22318
rect 32172 22930 32228 22942
rect 32172 22878 32174 22930
rect 32226 22878 32228 22930
rect 32060 22036 32116 22046
rect 32060 20914 32116 21980
rect 32060 20862 32062 20914
rect 32114 20862 32116 20914
rect 32060 20850 32116 20862
rect 31948 19964 32116 20020
rect 31836 19842 31892 19852
rect 31948 19796 32004 19806
rect 31948 19702 32004 19740
rect 31948 19236 32004 19246
rect 32060 19236 32116 19964
rect 31948 19234 32116 19236
rect 31948 19182 31950 19234
rect 32002 19182 32116 19234
rect 31948 19180 32116 19182
rect 31948 19170 32004 19180
rect 31724 18398 31726 18450
rect 31778 18398 31780 18450
rect 31724 18386 31780 18398
rect 32060 17666 32116 17678
rect 32060 17614 32062 17666
rect 32114 17614 32116 17666
rect 31836 17332 31892 17342
rect 31276 16882 31444 16884
rect 31276 16830 31278 16882
rect 31330 16830 31444 16882
rect 31276 16828 31444 16830
rect 31500 17108 31556 17118
rect 31724 17108 31780 17118
rect 31500 16882 31556 17052
rect 31500 16830 31502 16882
rect 31554 16830 31556 16882
rect 31276 16772 31332 16828
rect 31276 16706 31332 16716
rect 31276 15988 31332 15998
rect 31276 15426 31332 15932
rect 31500 15540 31556 16830
rect 31500 15474 31556 15484
rect 31612 17052 31724 17108
rect 31612 15538 31668 17052
rect 31724 17042 31780 17052
rect 31836 17106 31892 17276
rect 31836 17054 31838 17106
rect 31890 17054 31892 17106
rect 31836 17042 31892 17054
rect 31948 16996 32004 17006
rect 31948 16902 32004 16940
rect 32060 16884 32116 17614
rect 32060 16818 32116 16828
rect 31612 15486 31614 15538
rect 31666 15486 31668 15538
rect 31612 15474 31668 15486
rect 31836 15540 31892 15550
rect 31276 15374 31278 15426
rect 31330 15374 31332 15426
rect 31276 15362 31332 15374
rect 31724 15428 31780 15438
rect 31724 15334 31780 15372
rect 31500 15314 31556 15326
rect 31500 15262 31502 15314
rect 31554 15262 31556 15314
rect 31500 15204 31556 15262
rect 31052 15148 31556 15204
rect 31500 15092 31668 15148
rect 31052 13748 31108 13758
rect 31052 13074 31108 13692
rect 31388 13748 31444 13758
rect 31388 13654 31444 13692
rect 31612 13746 31668 15092
rect 31836 13972 31892 15484
rect 31948 13972 32004 13982
rect 31836 13970 32004 13972
rect 31836 13918 31950 13970
rect 32002 13918 32004 13970
rect 31836 13916 32004 13918
rect 31612 13694 31614 13746
rect 31666 13694 31668 13746
rect 31052 13022 31054 13074
rect 31106 13022 31108 13074
rect 31052 13010 31108 13022
rect 31612 12852 31668 13694
rect 31836 13748 31892 13758
rect 31836 13654 31892 13692
rect 31724 13636 31780 13646
rect 31724 13542 31780 13580
rect 31052 12796 31668 12852
rect 31052 12516 31108 12796
rect 31948 12740 32004 13916
rect 31612 12684 32004 12740
rect 32060 13300 32116 13310
rect 31052 12460 31220 12516
rect 30940 12348 31108 12404
rect 30492 12292 30548 12302
rect 30380 12236 30492 12292
rect 30380 12178 30436 12236
rect 30492 12226 30548 12236
rect 30380 12126 30382 12178
rect 30434 12126 30436 12178
rect 30380 12114 30436 12126
rect 30940 12180 30996 12190
rect 30940 12086 30996 12124
rect 31052 12068 31108 12348
rect 31164 12402 31220 12460
rect 31164 12350 31166 12402
rect 31218 12350 31220 12402
rect 31164 12338 31220 12350
rect 31388 12404 31444 12414
rect 31388 12310 31444 12348
rect 31276 12292 31332 12302
rect 31276 12198 31332 12236
rect 31612 12178 31668 12684
rect 32060 12404 32116 13244
rect 32060 12310 32116 12348
rect 31612 12126 31614 12178
rect 31666 12126 31668 12178
rect 31612 12114 31668 12126
rect 31052 12012 31444 12068
rect 30492 11956 30548 11966
rect 30492 11954 31332 11956
rect 30492 11902 30494 11954
rect 30546 11902 31332 11954
rect 30492 11900 31332 11902
rect 30492 11890 30548 11900
rect 30268 11508 30324 11518
rect 29596 11506 30324 11508
rect 29596 11454 29598 11506
rect 29650 11454 30270 11506
rect 30322 11454 30324 11506
rect 29596 11452 30324 11454
rect 29596 11442 29652 11452
rect 30268 11442 30324 11452
rect 30492 11394 30548 11406
rect 30492 11342 30494 11394
rect 30546 11342 30548 11394
rect 29932 11284 29988 11294
rect 30492 11284 30548 11342
rect 29484 11282 30548 11284
rect 29484 11230 29934 11282
rect 29986 11230 30548 11282
rect 29484 11228 30548 11230
rect 29932 11218 29988 11228
rect 30492 10724 30548 11228
rect 30828 11172 30884 11182
rect 30828 11078 30884 11116
rect 30492 10658 30548 10668
rect 31276 10722 31332 11900
rect 31276 10670 31278 10722
rect 31330 10670 31332 10722
rect 31276 10658 31332 10670
rect 29148 10446 29150 10498
rect 29202 10446 29204 10498
rect 29148 10434 29204 10446
rect 27916 10052 27972 10062
rect 27692 10050 27972 10052
rect 27692 9998 27918 10050
rect 27970 9998 27972 10050
rect 27692 9996 27972 9998
rect 27580 9828 27636 9838
rect 27580 9734 27636 9772
rect 27468 9716 27524 9726
rect 27468 9622 27524 9660
rect 27580 8820 27636 8830
rect 27692 8820 27748 9996
rect 27916 9986 27972 9996
rect 27580 8818 27748 8820
rect 27580 8766 27582 8818
rect 27634 8766 27748 8818
rect 27580 8764 27748 8766
rect 27804 9826 27860 9838
rect 27804 9774 27806 9826
rect 27858 9774 27860 9826
rect 27468 8372 27524 8382
rect 27580 8372 27636 8764
rect 27468 8370 27636 8372
rect 27468 8318 27470 8370
rect 27522 8318 27636 8370
rect 27468 8316 27636 8318
rect 27804 8372 27860 9774
rect 30716 9826 30772 9838
rect 30716 9774 30718 9826
rect 30770 9774 30772 9826
rect 28700 9716 28756 9726
rect 27916 9604 27972 9614
rect 27916 9042 27972 9548
rect 28700 9154 28756 9660
rect 30716 9604 30772 9774
rect 30716 9538 30772 9548
rect 28700 9102 28702 9154
rect 28754 9102 28756 9154
rect 28700 9090 28756 9102
rect 27916 8990 27918 9042
rect 27970 8990 27972 9042
rect 27916 8978 27972 8990
rect 29596 9044 29652 9054
rect 27468 6580 27524 8316
rect 27804 8306 27860 8316
rect 29148 8932 29204 8942
rect 27692 8258 27748 8270
rect 27692 8206 27694 8258
rect 27746 8206 27748 8258
rect 27692 8148 27748 8206
rect 28140 8204 28532 8260
rect 28140 8148 28196 8204
rect 27692 8092 28196 8148
rect 28252 8036 28308 8046
rect 28252 7942 28308 7980
rect 28364 7362 28420 8204
rect 28476 8146 28532 8204
rect 29148 8258 29204 8876
rect 29260 8372 29316 8382
rect 29260 8278 29316 8316
rect 29148 8206 29150 8258
rect 29202 8206 29204 8258
rect 29148 8194 29204 8206
rect 29596 8258 29652 8988
rect 30828 9044 30884 9054
rect 30828 8930 30884 8988
rect 30828 8878 30830 8930
rect 30882 8878 30884 8930
rect 30828 8866 30884 8878
rect 30380 8372 30436 8382
rect 30380 8370 31220 8372
rect 30380 8318 30382 8370
rect 30434 8318 31220 8370
rect 30380 8316 31220 8318
rect 30380 8306 30436 8316
rect 29596 8206 29598 8258
rect 29650 8206 29652 8258
rect 29596 8194 29652 8206
rect 28476 8094 28478 8146
rect 28530 8094 28532 8146
rect 28476 8082 28532 8094
rect 28588 8148 28644 8158
rect 29484 8148 29540 8158
rect 30044 8148 30100 8158
rect 28588 8146 29092 8148
rect 28588 8094 28590 8146
rect 28642 8094 29092 8146
rect 28588 8092 29092 8094
rect 28588 8082 28644 8092
rect 28364 7310 28366 7362
rect 28418 7310 28420 7362
rect 27468 6514 27524 6524
rect 28252 6916 28308 6926
rect 28252 6578 28308 6860
rect 28364 6692 28420 7310
rect 29036 7362 29092 8092
rect 29484 8054 29540 8092
rect 29820 8146 30100 8148
rect 29820 8094 30046 8146
rect 30098 8094 30100 8146
rect 29820 8092 30100 8094
rect 29820 7364 29876 8092
rect 30044 8082 30100 8092
rect 30268 8036 30324 8046
rect 30268 8034 30436 8036
rect 30268 7982 30270 8034
rect 30322 7982 30436 8034
rect 30268 7980 30436 7982
rect 30268 7970 30324 7980
rect 29036 7310 29038 7362
rect 29090 7310 29092 7362
rect 29036 7140 29092 7310
rect 29036 7074 29092 7084
rect 29260 7308 29876 7364
rect 29260 6802 29316 7308
rect 29260 6750 29262 6802
rect 29314 6750 29316 6802
rect 29260 6738 29316 6750
rect 29596 7140 29652 7150
rect 28364 6626 28420 6636
rect 29372 6692 29428 6702
rect 29372 6598 29428 6636
rect 29596 6690 29652 7084
rect 30268 7140 30324 7150
rect 30268 6914 30324 7084
rect 30268 6862 30270 6914
rect 30322 6862 30324 6914
rect 30268 6850 30324 6862
rect 30380 6804 30436 7980
rect 31164 7586 31220 8316
rect 31164 7534 31166 7586
rect 31218 7534 31220 7586
rect 31164 7522 31220 7534
rect 29596 6638 29598 6690
rect 29650 6638 29652 6690
rect 29596 6626 29652 6638
rect 30044 6692 30100 6702
rect 30044 6598 30100 6636
rect 28252 6526 28254 6578
rect 28306 6526 28308 6578
rect 28252 6514 28308 6526
rect 29148 6580 29204 6590
rect 29148 6486 29204 6524
rect 28588 6468 28644 6478
rect 28588 6374 28644 6412
rect 29596 6468 29652 6478
rect 27356 6290 27412 6300
rect 26684 6018 26852 6020
rect 26684 5966 26686 6018
rect 26738 5966 26852 6018
rect 26684 5964 26852 5966
rect 26684 5954 26740 5964
rect 26460 5740 26740 5796
rect 26348 5236 26404 5404
rect 26460 5236 26516 5246
rect 26348 5234 26516 5236
rect 26348 5182 26462 5234
rect 26514 5182 26516 5234
rect 26348 5180 26516 5182
rect 26348 4900 26404 5180
rect 26460 5170 26516 5180
rect 26012 4834 26068 4844
rect 26348 4834 26404 4844
rect 25900 4162 25956 4172
rect 26572 4226 26628 4238
rect 26572 4174 26574 4226
rect 26626 4174 26628 4226
rect 26572 3778 26628 4174
rect 26572 3726 26574 3778
rect 26626 3726 26628 3778
rect 26572 3714 26628 3726
rect 26684 3780 26740 5740
rect 29260 5794 29316 5806
rect 29260 5742 29262 5794
rect 29314 5742 29316 5794
rect 26908 5572 26964 5582
rect 26908 5234 26964 5516
rect 26908 5182 26910 5234
rect 26962 5182 26964 5234
rect 26908 5170 26964 5182
rect 29148 5236 29204 5246
rect 29148 5142 29204 5180
rect 27804 5124 27860 5134
rect 27804 5010 27860 5068
rect 27804 4958 27806 5010
rect 27858 4958 27860 5010
rect 27804 4946 27860 4958
rect 29260 5012 29316 5742
rect 29596 5234 29652 6412
rect 29596 5182 29598 5234
rect 29650 5182 29652 5234
rect 29596 5170 29652 5182
rect 30044 5348 30100 5358
rect 28140 4900 28196 4910
rect 28588 4900 28644 4910
rect 28140 4898 28532 4900
rect 28140 4846 28142 4898
rect 28194 4846 28532 4898
rect 28140 4844 28532 4846
rect 28140 4834 28196 4844
rect 28476 4228 28532 4844
rect 28588 4898 28868 4900
rect 28588 4846 28590 4898
rect 28642 4846 28868 4898
rect 28588 4844 28868 4846
rect 28588 4834 28644 4844
rect 28700 4228 28756 4238
rect 28476 4226 28756 4228
rect 28476 4174 28702 4226
rect 28754 4174 28756 4226
rect 28476 4172 28756 4174
rect 26908 3780 26964 3790
rect 26684 3778 26964 3780
rect 26684 3726 26910 3778
rect 26962 3726 26964 3778
rect 26684 3724 26964 3726
rect 26908 3714 26964 3724
rect 28588 3666 28644 4172
rect 28700 4162 28756 4172
rect 28700 3780 28756 3790
rect 28700 3686 28756 3724
rect 28588 3614 28590 3666
rect 28642 3614 28644 3666
rect 28588 3602 28644 3614
rect 26572 3556 26628 3566
rect 25676 3554 26628 3556
rect 25676 3502 26574 3554
rect 26626 3502 26628 3554
rect 25676 3500 26628 3502
rect 24668 3442 24724 3500
rect 26572 3490 26628 3500
rect 24668 3390 24670 3442
rect 24722 3390 24724 3442
rect 24668 3378 24724 3390
rect 23996 3332 24052 3342
rect 23996 800 24052 3276
rect 25228 3332 25284 3342
rect 25788 3332 25844 3342
rect 27356 3332 27412 3342
rect 25228 3238 25284 3276
rect 25564 3330 25844 3332
rect 25564 3278 25790 3330
rect 25842 3278 25844 3330
rect 25564 3276 25844 3278
rect 25564 800 25620 3276
rect 25788 3266 25844 3276
rect 27132 3330 27412 3332
rect 27132 3278 27358 3330
rect 27410 3278 27412 3330
rect 27132 3276 27412 3278
rect 27132 800 27188 3276
rect 27356 3266 27412 3276
rect 28812 2436 28868 4844
rect 29260 4338 29316 4956
rect 29260 4286 29262 4338
rect 29314 4286 29316 4338
rect 29260 4274 29316 4286
rect 29484 5124 29540 5134
rect 29260 3780 29316 3790
rect 29484 3780 29540 5068
rect 30044 4450 30100 5292
rect 30268 5348 30324 5358
rect 30380 5348 30436 6748
rect 30940 6916 30996 6926
rect 30940 6690 30996 6860
rect 30940 6638 30942 6690
rect 30994 6638 30996 6690
rect 30940 6626 30996 6638
rect 30604 6468 30660 6478
rect 30604 6374 30660 6412
rect 31052 6466 31108 6478
rect 31052 6414 31054 6466
rect 31106 6414 31108 6466
rect 31052 6356 31108 6414
rect 31052 6290 31108 6300
rect 31276 6466 31332 6478
rect 31276 6414 31278 6466
rect 31330 6414 31332 6466
rect 30268 5346 30436 5348
rect 30268 5294 30270 5346
rect 30322 5294 30436 5346
rect 30268 5292 30436 5294
rect 31052 5684 31108 5694
rect 30268 5282 30324 5292
rect 31052 5234 31108 5628
rect 31276 5348 31332 6414
rect 31276 5282 31332 5292
rect 31052 5182 31054 5234
rect 31106 5182 31108 5234
rect 31052 5170 31108 5182
rect 30492 5124 30548 5134
rect 30492 5010 30548 5068
rect 30492 4958 30494 5010
rect 30546 4958 30548 5010
rect 30492 4946 30548 4958
rect 30380 4900 30436 4910
rect 30380 4806 30436 4844
rect 30044 4398 30046 4450
rect 30098 4398 30100 4450
rect 30044 4386 30100 4398
rect 29316 3724 29540 3780
rect 29260 3714 29316 3724
rect 30268 3666 30324 3678
rect 30268 3614 30270 3666
rect 30322 3614 30324 3666
rect 29036 3556 29092 3566
rect 29036 3462 29092 3500
rect 28700 2380 28868 2436
rect 28700 800 28756 2380
rect 30268 800 30324 3614
rect 31388 3444 31444 12012
rect 31948 11844 32004 11854
rect 31948 11282 32004 11788
rect 31948 11230 31950 11282
rect 32002 11230 32004 11282
rect 31948 10610 32004 11230
rect 31948 10558 31950 10610
rect 32002 10558 32004 10610
rect 31500 10388 31556 10398
rect 31500 9938 31556 10332
rect 31500 9886 31502 9938
rect 31554 9886 31556 9938
rect 31500 9874 31556 9886
rect 31948 9604 32004 10558
rect 31948 9538 32004 9548
rect 32172 9044 32228 22878
rect 32732 22484 32788 26684
rect 32844 23156 32900 26852
rect 32956 25844 33012 32732
rect 33180 32676 33236 36876
rect 33516 36372 33572 40684
rect 33740 40628 33796 40908
rect 33740 40516 33796 40572
rect 33852 40516 33908 40526
rect 33740 40514 33908 40516
rect 33740 40462 33854 40514
rect 33906 40462 33908 40514
rect 33740 40460 33908 40462
rect 33852 40450 33908 40460
rect 33628 40404 33684 40414
rect 33628 40310 33684 40348
rect 33740 38836 33796 38846
rect 33740 38742 33796 38780
rect 33964 38668 34020 42028
rect 34300 41412 34356 41422
rect 34188 41410 34356 41412
rect 34188 41358 34302 41410
rect 34354 41358 34356 41410
rect 34188 41356 34356 41358
rect 34076 40180 34132 40190
rect 34188 40180 34244 41356
rect 34300 41346 34356 41356
rect 34300 41188 34356 41198
rect 34300 41094 34356 41132
rect 34524 40740 34580 43260
rect 35420 43316 35476 43710
rect 35644 43764 35700 43774
rect 35644 43650 35700 43708
rect 35644 43598 35646 43650
rect 35698 43598 35700 43650
rect 35644 43586 35700 43598
rect 35420 43250 35476 43260
rect 36428 43538 36484 44044
rect 36428 43486 36430 43538
rect 36482 43486 36484 43538
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 36428 42866 36484 43486
rect 36428 42814 36430 42866
rect 36482 42814 36484 42866
rect 36428 42802 36484 42814
rect 36540 42756 36596 45052
rect 36988 44996 37044 45006
rect 37212 44996 37268 45006
rect 36988 44994 37212 44996
rect 36988 44942 36990 44994
rect 37042 44942 37212 44994
rect 36988 44940 37212 44942
rect 36988 44930 37044 44940
rect 36988 44324 37044 44334
rect 36652 43764 36708 43774
rect 36652 43538 36708 43708
rect 36988 43762 37044 44268
rect 36988 43710 36990 43762
rect 37042 43710 37044 43762
rect 36988 43698 37044 43710
rect 37100 44322 37156 44334
rect 37100 44270 37102 44322
rect 37154 44270 37156 44322
rect 36652 43486 36654 43538
rect 36706 43486 36708 43538
rect 36652 43474 36708 43486
rect 37100 43540 37156 44270
rect 37212 43764 37268 44940
rect 37884 44436 37940 45726
rect 38220 45780 38276 45838
rect 38556 45780 38612 45790
rect 38220 45724 38500 45780
rect 37996 45668 38052 45678
rect 37996 45574 38052 45612
rect 38444 45556 38500 45724
rect 37996 44436 38052 44446
rect 37884 44434 38052 44436
rect 37884 44382 37998 44434
rect 38050 44382 38052 44434
rect 37884 44380 38052 44382
rect 37996 44370 38052 44380
rect 37212 43698 37268 43708
rect 37436 44322 37492 44334
rect 37436 44270 37438 44322
rect 37490 44270 37492 44322
rect 37436 43988 37492 44270
rect 38332 44100 38388 44110
rect 37100 43474 37156 43484
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 36540 41188 36596 42700
rect 36652 42308 36708 42318
rect 36652 41970 36708 42252
rect 36652 41918 36654 41970
rect 36706 41918 36708 41970
rect 36652 41906 36708 41918
rect 36988 42082 37044 42094
rect 36988 42030 36990 42082
rect 37042 42030 37044 42082
rect 36988 41748 37044 42030
rect 37436 41972 37492 43932
rect 38108 44098 38388 44100
rect 38108 44046 38334 44098
rect 38386 44046 38388 44098
rect 38108 44044 38388 44046
rect 38108 43540 38164 44044
rect 38332 44034 38388 44044
rect 38444 43876 38500 45500
rect 38556 44324 38612 45724
rect 39116 45668 39172 45678
rect 39340 45668 39396 45678
rect 39116 45218 39172 45612
rect 39116 45166 39118 45218
rect 39170 45166 39172 45218
rect 39116 45154 39172 45166
rect 39228 45612 39340 45668
rect 38556 44230 38612 44268
rect 39228 43988 39284 45612
rect 39340 45602 39396 45612
rect 39900 45106 39956 45118
rect 39900 45054 39902 45106
rect 39954 45054 39956 45106
rect 39676 44884 39732 44894
rect 39340 44212 39396 44222
rect 39340 44210 39508 44212
rect 39340 44158 39342 44210
rect 39394 44158 39508 44210
rect 39340 44156 39508 44158
rect 39340 44146 39396 44156
rect 39228 43932 39396 43988
rect 38332 43820 38500 43876
rect 38220 43764 38276 43774
rect 38220 43670 38276 43708
rect 38108 43446 38164 43484
rect 37884 42980 37940 42990
rect 37884 42642 37940 42924
rect 37884 42590 37886 42642
rect 37938 42590 37940 42642
rect 37884 42578 37940 42590
rect 37548 42530 37604 42542
rect 37548 42478 37550 42530
rect 37602 42478 37604 42530
rect 37548 42308 37604 42478
rect 37548 42242 37604 42252
rect 37884 41972 37940 41982
rect 37436 41970 37940 41972
rect 37436 41918 37886 41970
rect 37938 41918 37940 41970
rect 37436 41916 37940 41918
rect 38332 41972 38388 43820
rect 39228 43764 39284 43774
rect 38556 43652 38612 43662
rect 38444 43540 38500 43550
rect 38444 43446 38500 43484
rect 38556 43538 38612 43596
rect 39004 43652 39060 43662
rect 39004 43558 39060 43596
rect 38556 43486 38558 43538
rect 38610 43486 38612 43538
rect 38556 43474 38612 43486
rect 39228 43538 39284 43708
rect 39228 43486 39230 43538
rect 39282 43486 39284 43538
rect 39228 43474 39284 43486
rect 38780 43428 38836 43438
rect 38780 43426 39172 43428
rect 38780 43374 38782 43426
rect 38834 43374 39172 43426
rect 38780 43372 39172 43374
rect 38780 43362 38836 43372
rect 39116 43092 39172 43372
rect 39340 43204 39396 43932
rect 39452 43708 39508 44156
rect 39676 43988 39732 44828
rect 39452 43652 39620 43708
rect 39340 43148 39508 43204
rect 39116 43036 39396 43092
rect 39004 42868 39060 42878
rect 38444 41972 38500 41982
rect 38332 41970 38500 41972
rect 38332 41918 38446 41970
rect 38498 41918 38500 41970
rect 38332 41916 38500 41918
rect 37324 41748 37380 41758
rect 36988 41682 37044 41692
rect 37100 41746 37380 41748
rect 37100 41694 37326 41746
rect 37378 41694 37380 41746
rect 37100 41692 37380 41694
rect 34636 41076 34692 41086
rect 34636 40982 34692 41020
rect 35084 41074 35140 41086
rect 35084 41022 35086 41074
rect 35138 41022 35140 41074
rect 34972 40962 35028 40974
rect 34972 40910 34974 40962
rect 35026 40910 35028 40962
rect 34524 40684 34692 40740
rect 34412 40516 34468 40526
rect 34076 40178 34244 40180
rect 34076 40126 34078 40178
rect 34130 40126 34244 40178
rect 34076 40124 34244 40126
rect 34300 40460 34412 40516
rect 34300 40402 34356 40460
rect 34412 40450 34468 40460
rect 34524 40516 34580 40526
rect 34636 40516 34692 40684
rect 34524 40514 34692 40516
rect 34524 40462 34526 40514
rect 34578 40462 34692 40514
rect 34524 40460 34692 40462
rect 34524 40450 34580 40460
rect 34300 40350 34302 40402
rect 34354 40350 34356 40402
rect 34076 39844 34132 40124
rect 34076 39778 34132 39788
rect 34300 39508 34356 40350
rect 34412 40290 34468 40302
rect 34412 40238 34414 40290
rect 34466 40238 34468 40290
rect 34412 39844 34468 40238
rect 34412 39778 34468 39788
rect 34636 39844 34692 40460
rect 34972 40516 35028 40910
rect 34972 40450 35028 40460
rect 34524 39508 34580 39518
rect 34300 39506 34580 39508
rect 34300 39454 34526 39506
rect 34578 39454 34580 39506
rect 34300 39452 34580 39454
rect 34524 39442 34580 39452
rect 34636 39506 34692 39788
rect 34636 39454 34638 39506
rect 34690 39454 34692 39506
rect 34636 39442 34692 39454
rect 34860 39508 34916 39518
rect 34860 39414 34916 39452
rect 34188 39396 34244 39406
rect 34076 39394 34244 39396
rect 34076 39342 34190 39394
rect 34242 39342 34244 39394
rect 34076 39340 34244 39342
rect 34076 39060 34132 39340
rect 34188 39330 34244 39340
rect 34972 39396 35028 39406
rect 34972 39302 35028 39340
rect 34076 38834 34132 39004
rect 34076 38782 34078 38834
rect 34130 38782 34132 38834
rect 34076 38770 34132 38782
rect 34188 39172 34244 39182
rect 33964 38612 34132 38668
rect 33628 38052 33684 38062
rect 33628 37958 33684 37996
rect 33740 37604 33796 37614
rect 33740 37490 33796 37548
rect 33740 37438 33742 37490
rect 33794 37438 33796 37490
rect 33740 37426 33796 37438
rect 33628 37268 33684 37278
rect 33628 37044 33684 37212
rect 33964 37266 34020 37278
rect 33964 37214 33966 37266
rect 34018 37214 34020 37266
rect 33852 37156 33908 37166
rect 33852 37062 33908 37100
rect 33628 36978 33684 36988
rect 33516 36306 33572 36316
rect 33964 36932 34020 37214
rect 33404 35924 33460 35934
rect 33964 35924 34020 36876
rect 34076 36036 34132 38612
rect 34188 37380 34244 39116
rect 35084 39172 35140 41022
rect 35532 41076 35588 41086
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35420 39732 35476 39742
rect 35308 39620 35364 39630
rect 35308 39526 35364 39564
rect 35420 39396 35476 39676
rect 35420 39330 35476 39340
rect 35084 39106 35140 39116
rect 35196 38836 35252 38846
rect 34748 38834 35252 38836
rect 34748 38782 35198 38834
rect 35250 38782 35252 38834
rect 34748 38780 35252 38782
rect 34300 38612 34356 38622
rect 34300 38162 34356 38556
rect 34300 38110 34302 38162
rect 34354 38110 34356 38162
rect 34300 38098 34356 38110
rect 34748 37940 34804 38780
rect 35196 38770 35252 38780
rect 35532 38668 35588 41020
rect 36092 41074 36148 41086
rect 36092 41022 36094 41074
rect 36146 41022 36148 41074
rect 35980 40964 36036 40974
rect 35868 40962 36036 40964
rect 35868 40910 35982 40962
rect 36034 40910 36036 40962
rect 35868 40908 36036 40910
rect 35644 39620 35700 39630
rect 35644 39526 35700 39564
rect 35756 39508 35812 39518
rect 35756 39414 35812 39452
rect 35868 38946 35924 40908
rect 35980 40898 36036 40908
rect 35980 39732 36036 39742
rect 36092 39732 36148 41022
rect 36540 40516 36596 41132
rect 35980 39730 36092 39732
rect 35980 39678 35982 39730
rect 36034 39678 36092 39730
rect 35980 39676 36092 39678
rect 35980 39666 36036 39676
rect 36092 39638 36148 39676
rect 36204 40514 36596 40516
rect 36204 40462 36542 40514
rect 36594 40462 36596 40514
rect 36204 40460 36596 40462
rect 35868 38894 35870 38946
rect 35922 38894 35924 38946
rect 35868 38882 35924 38894
rect 36092 39396 36148 39406
rect 36092 38834 36148 39340
rect 36092 38782 36094 38834
rect 36146 38782 36148 38834
rect 36092 38770 36148 38782
rect 35084 38612 35140 38622
rect 35532 38612 35924 38668
rect 35084 38518 35140 38556
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 34748 37884 34916 37940
rect 34748 37492 34804 37502
rect 34748 37398 34804 37436
rect 34860 37490 34916 37884
rect 34860 37438 34862 37490
rect 34914 37438 34916 37490
rect 34860 37426 34916 37438
rect 35644 37604 35700 37614
rect 35644 37490 35700 37548
rect 35644 37438 35646 37490
rect 35698 37438 35700 37490
rect 35196 37380 35252 37390
rect 34188 37378 34580 37380
rect 34188 37326 34190 37378
rect 34242 37326 34580 37378
rect 34188 37324 34580 37326
rect 34188 37314 34244 37324
rect 34524 37044 34580 37324
rect 35196 37286 35252 37324
rect 34636 37268 34692 37278
rect 34636 37174 34692 37212
rect 34972 37266 35028 37278
rect 34972 37214 34974 37266
rect 35026 37214 35028 37266
rect 34524 36988 34804 37044
rect 34748 36594 34804 36988
rect 34972 36932 35028 37214
rect 35644 37156 35700 37438
rect 35644 37090 35700 37100
rect 34972 36866 35028 36876
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 34748 36542 34750 36594
rect 34802 36542 34804 36594
rect 34748 36530 34804 36542
rect 34076 35980 34244 36036
rect 33404 35922 34020 35924
rect 33404 35870 33406 35922
rect 33458 35870 34020 35922
rect 33404 35868 34020 35870
rect 33404 35858 33460 35868
rect 33628 34020 33684 35868
rect 34076 35586 34132 35598
rect 34076 35534 34078 35586
rect 34130 35534 34132 35586
rect 33964 35474 34020 35486
rect 33964 35422 33966 35474
rect 34018 35422 34020 35474
rect 33852 34244 33908 34254
rect 33964 34244 34020 35422
rect 34076 34356 34132 35534
rect 34188 35028 34244 35980
rect 34188 34914 34244 34972
rect 34188 34862 34190 34914
rect 34242 34862 34244 34914
rect 34188 34850 34244 34862
rect 34524 35588 34580 35598
rect 34524 34804 34580 35532
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35420 35028 35476 35038
rect 35420 34934 35476 34972
rect 34524 34738 34580 34748
rect 34076 34290 34132 34300
rect 33852 34242 34020 34244
rect 33852 34190 33854 34242
rect 33906 34190 34020 34242
rect 33852 34188 34020 34190
rect 33852 34178 33908 34188
rect 33852 34020 33908 34030
rect 33628 33964 33852 34020
rect 35868 34020 35924 38612
rect 36204 38052 36260 40460
rect 36540 40450 36596 40460
rect 36316 39844 36372 39854
rect 36316 39730 36372 39788
rect 36316 39678 36318 39730
rect 36370 39678 36372 39730
rect 36316 39666 36372 39678
rect 37100 39620 37156 41692
rect 37324 41682 37380 41692
rect 37324 41188 37380 41198
rect 37324 41094 37380 41132
rect 37324 39732 37380 39742
rect 37324 39638 37380 39676
rect 36428 39508 36484 39518
rect 36988 39508 37044 39518
rect 36428 39506 37044 39508
rect 36428 39454 36430 39506
rect 36482 39454 36990 39506
rect 37042 39454 37044 39506
rect 36428 39452 37044 39454
rect 36428 39442 36484 39452
rect 36988 39442 37044 39452
rect 36988 38948 37044 38958
rect 36988 38834 37044 38892
rect 36988 38782 36990 38834
rect 37042 38782 37044 38834
rect 36988 38770 37044 38782
rect 37100 38836 37156 39564
rect 37436 39618 37492 41916
rect 37884 41906 37940 41916
rect 38444 41906 38500 41916
rect 38892 41972 38948 41982
rect 37660 41746 37716 41758
rect 38444 41748 38500 41758
rect 37660 41694 37662 41746
rect 37714 41694 37716 41746
rect 37660 39620 37716 41694
rect 38108 41746 38500 41748
rect 38108 41694 38446 41746
rect 38498 41694 38500 41746
rect 38108 41692 38500 41694
rect 38108 41298 38164 41692
rect 38444 41682 38500 41692
rect 38780 41746 38836 41758
rect 38780 41694 38782 41746
rect 38834 41694 38836 41746
rect 38108 41246 38110 41298
rect 38162 41246 38164 41298
rect 38108 41234 38164 41246
rect 37436 39566 37438 39618
rect 37490 39566 37492 39618
rect 37436 39554 37492 39566
rect 37548 39618 37716 39620
rect 37548 39566 37662 39618
rect 37714 39566 37716 39618
rect 37548 39564 37716 39566
rect 37212 39394 37268 39406
rect 37212 39342 37214 39394
rect 37266 39342 37268 39394
rect 37212 39172 37268 39342
rect 37548 39172 37604 39564
rect 37660 39554 37716 39564
rect 38668 40852 38724 40862
rect 37212 39106 37268 39116
rect 37436 39116 37604 39172
rect 38444 39284 38500 39294
rect 37212 38836 37268 38846
rect 37100 38834 37268 38836
rect 37100 38782 37214 38834
rect 37266 38782 37268 38834
rect 37100 38780 37268 38782
rect 37212 38770 37268 38780
rect 36428 38724 36484 38762
rect 36428 38658 36484 38668
rect 36204 37986 36260 37996
rect 36428 38164 36484 38174
rect 36092 37492 36148 37502
rect 36092 37398 36148 37436
rect 36428 37380 36484 38108
rect 37436 38164 37492 39116
rect 38444 38946 38500 39228
rect 38444 38894 38446 38946
rect 38498 38894 38500 38946
rect 38444 38882 38500 38894
rect 37548 38836 37604 38846
rect 37772 38836 37828 38846
rect 37548 38834 37828 38836
rect 37548 38782 37550 38834
rect 37602 38782 37774 38834
rect 37826 38782 37828 38834
rect 37548 38780 37828 38782
rect 37548 38770 37604 38780
rect 37772 38770 37828 38780
rect 37996 38836 38052 38846
rect 37996 38742 38052 38780
rect 38108 38834 38164 38846
rect 38108 38782 38110 38834
rect 38162 38782 38164 38834
rect 38108 38724 38164 38782
rect 38108 38658 38164 38668
rect 38668 38668 38724 40796
rect 38780 39730 38836 41694
rect 38892 40404 38948 41916
rect 38892 40310 38948 40348
rect 38780 39678 38782 39730
rect 38834 39678 38836 39730
rect 38780 39666 38836 39678
rect 38668 38612 38836 38668
rect 37436 38098 37492 38108
rect 36428 37314 36484 37324
rect 36540 38052 36596 38062
rect 36428 36260 36484 36270
rect 36092 36148 36148 36158
rect 36092 35922 36148 36092
rect 36092 35870 36094 35922
rect 36146 35870 36148 35922
rect 36092 35858 36148 35870
rect 35980 35700 36036 35710
rect 35980 34692 36036 35644
rect 36316 35698 36372 35710
rect 36316 35646 36318 35698
rect 36370 35646 36372 35698
rect 36316 35140 36372 35646
rect 36316 35074 36372 35084
rect 36428 34916 36484 36204
rect 36540 35698 36596 37996
rect 37100 38052 37156 38062
rect 37100 37266 37156 37996
rect 37100 37214 37102 37266
rect 37154 37214 37156 37266
rect 37100 37202 37156 37214
rect 38108 38052 38164 38062
rect 37884 37154 37940 37166
rect 37884 37102 37886 37154
rect 37938 37102 37940 37154
rect 37884 36594 37940 37102
rect 38108 36706 38164 37996
rect 38780 37716 38836 38612
rect 38780 37650 38836 37660
rect 38108 36654 38110 36706
rect 38162 36654 38164 36706
rect 38108 36642 38164 36654
rect 38780 37156 38836 37166
rect 37884 36542 37886 36594
rect 37938 36542 37940 36594
rect 37884 36530 37940 36542
rect 37660 36482 37716 36494
rect 38332 36484 38388 36494
rect 37660 36430 37662 36482
rect 37714 36430 37716 36482
rect 36540 35646 36542 35698
rect 36594 35646 36596 35698
rect 36540 35634 36596 35646
rect 36988 36370 37044 36382
rect 36988 36318 36990 36370
rect 37042 36318 37044 36370
rect 36988 35700 37044 36318
rect 37324 36372 37380 36382
rect 37548 36372 37604 36382
rect 37324 36370 37604 36372
rect 37324 36318 37326 36370
rect 37378 36318 37550 36370
rect 37602 36318 37604 36370
rect 37324 36316 37604 36318
rect 37324 36306 37380 36316
rect 37548 36306 37604 36316
rect 37100 36260 37156 36270
rect 37100 36166 37156 36204
rect 36988 35634 37044 35644
rect 37100 35924 37156 35934
rect 36988 35140 37044 35150
rect 36988 35046 37044 35084
rect 36428 34860 36932 34916
rect 36092 34692 36148 34702
rect 35980 34690 36148 34692
rect 35980 34638 36094 34690
rect 36146 34638 36148 34690
rect 35980 34636 36148 34638
rect 36092 34468 36148 34636
rect 36092 34402 36148 34412
rect 36428 34690 36484 34702
rect 36428 34638 36430 34690
rect 36482 34638 36484 34690
rect 36316 34130 36372 34142
rect 36316 34078 36318 34130
rect 36370 34078 36372 34130
rect 35980 34020 36036 34030
rect 36316 34020 36372 34078
rect 35868 34018 36372 34020
rect 35868 33966 35982 34018
rect 36034 33966 36372 34018
rect 35868 33964 36372 33966
rect 33740 33348 33796 33358
rect 33180 32610 33236 32620
rect 33404 32676 33460 32686
rect 33404 32582 33460 32620
rect 33740 32674 33796 33292
rect 33852 32788 33908 33964
rect 35980 33954 36036 33964
rect 36428 33908 36484 34638
rect 36652 34356 36708 34366
rect 36652 34262 36708 34300
rect 36540 34130 36596 34142
rect 36540 34078 36542 34130
rect 36594 34078 36596 34130
rect 36540 34020 36596 34078
rect 36764 34132 36820 34142
rect 36764 34038 36820 34076
rect 36540 33954 36596 33964
rect 36428 33842 36484 33852
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35868 33460 35924 33470
rect 35196 33236 35252 33246
rect 34860 33234 35252 33236
rect 34860 33182 35198 33234
rect 35250 33182 35252 33234
rect 34860 33180 35252 33182
rect 33964 32788 34020 32798
rect 33852 32786 34020 32788
rect 33852 32734 33966 32786
rect 34018 32734 34020 32786
rect 33852 32732 34020 32734
rect 33964 32722 34020 32732
rect 34076 32788 34132 32798
rect 34076 32786 34804 32788
rect 34076 32734 34078 32786
rect 34130 32734 34804 32786
rect 34076 32732 34804 32734
rect 34076 32722 34132 32732
rect 33740 32622 33742 32674
rect 33794 32622 33796 32674
rect 33740 32610 33796 32622
rect 34748 32674 34804 32732
rect 34860 32786 34916 33180
rect 35196 33170 35252 33180
rect 34860 32734 34862 32786
rect 34914 32734 34916 32786
rect 34860 32722 34916 32734
rect 35420 33124 35476 33134
rect 34748 32622 34750 32674
rect 34802 32622 34804 32674
rect 34748 32610 34804 32622
rect 33068 32564 33124 32574
rect 33068 32470 33124 32508
rect 34188 32562 34244 32574
rect 34188 32510 34190 32562
rect 34242 32510 34244 32562
rect 34188 32452 34244 32510
rect 34300 32564 34356 32574
rect 34300 32470 34356 32508
rect 35420 32562 35476 33068
rect 35420 32510 35422 32562
rect 35474 32510 35476 32562
rect 33404 32116 33460 32126
rect 33180 31556 33236 31566
rect 33180 30660 33236 31500
rect 33404 30884 33460 32060
rect 33964 31890 34020 31902
rect 33964 31838 33966 31890
rect 34018 31838 34020 31890
rect 33964 31668 34020 31838
rect 33516 31556 33572 31566
rect 33516 31462 33572 31500
rect 33964 31220 34020 31612
rect 34188 31556 34244 32396
rect 35420 32452 35476 32510
rect 35868 32452 35924 33404
rect 35980 33348 36036 33358
rect 35980 33346 36148 33348
rect 35980 33294 35982 33346
rect 36034 33294 36148 33346
rect 35980 33292 36148 33294
rect 35980 33282 36036 33292
rect 36092 32564 36148 33292
rect 36428 33124 36484 33134
rect 36428 33030 36484 33068
rect 36540 32564 36596 32574
rect 36092 32562 36596 32564
rect 36092 32510 36542 32562
rect 36594 32510 36596 32562
rect 36092 32508 36596 32510
rect 35980 32452 36036 32462
rect 35868 32450 36148 32452
rect 35868 32398 35982 32450
rect 36034 32398 36148 32450
rect 35868 32396 36148 32398
rect 35420 32386 35476 32396
rect 35980 32386 36036 32396
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 34636 31556 34692 31566
rect 34188 31554 34692 31556
rect 34188 31502 34638 31554
rect 34690 31502 34692 31554
rect 34188 31500 34692 31502
rect 33964 31154 34020 31164
rect 33404 30882 33572 30884
rect 33404 30830 33406 30882
rect 33458 30830 33572 30882
rect 33404 30828 33572 30830
rect 33404 30818 33460 30828
rect 33180 30594 33236 30604
rect 33516 30324 33572 30828
rect 34300 30882 34356 30894
rect 34300 30830 34302 30882
rect 34354 30830 34356 30882
rect 34076 30436 34132 30446
rect 34076 30342 34132 30380
rect 33516 30258 33572 30268
rect 34188 30324 34244 30334
rect 34076 30212 34132 30222
rect 34188 30212 34244 30268
rect 34076 30210 34244 30212
rect 34076 30158 34078 30210
rect 34130 30158 34244 30210
rect 34076 30156 34244 30158
rect 34300 30212 34356 30830
rect 34636 30548 34692 31500
rect 34636 30482 34692 30492
rect 34748 31556 34804 31566
rect 35196 31556 35252 31566
rect 34748 30436 34804 31500
rect 35084 31554 35252 31556
rect 35084 31502 35198 31554
rect 35250 31502 35252 31554
rect 35084 31500 35252 31502
rect 34076 30146 34132 30156
rect 34300 30146 34356 30156
rect 34636 30324 34692 30334
rect 33404 30100 33460 30110
rect 33740 30100 33796 30110
rect 33404 30098 33740 30100
rect 33404 30046 33406 30098
rect 33458 30046 33740 30098
rect 33404 30044 33740 30046
rect 33404 30034 33460 30044
rect 33740 30006 33796 30044
rect 33068 29988 33124 29998
rect 34412 29988 34468 29998
rect 33068 29986 33348 29988
rect 33068 29934 33070 29986
rect 33122 29934 33348 29986
rect 33068 29932 33348 29934
rect 33068 29922 33124 29932
rect 33292 29428 33348 29932
rect 33852 29986 34468 29988
rect 33852 29934 34414 29986
rect 34466 29934 34468 29986
rect 33852 29932 34468 29934
rect 33628 29652 33684 29690
rect 33628 29586 33684 29596
rect 33852 29650 33908 29932
rect 33852 29598 33854 29650
rect 33906 29598 33908 29650
rect 33852 29586 33908 29598
rect 33740 29540 33796 29550
rect 33740 29446 33796 29484
rect 33404 29428 33460 29438
rect 33292 29426 33460 29428
rect 33292 29374 33406 29426
rect 33458 29374 33460 29426
rect 33292 29372 33460 29374
rect 33292 28642 33348 28654
rect 33292 28590 33294 28642
rect 33346 28590 33348 28642
rect 33292 28196 33348 28590
rect 33292 28130 33348 28140
rect 33180 27746 33236 27758
rect 33180 27694 33182 27746
rect 33234 27694 33236 27746
rect 33180 27300 33236 27694
rect 33292 27748 33348 27758
rect 33292 27654 33348 27692
rect 33180 27234 33236 27244
rect 33180 27074 33236 27086
rect 33180 27022 33182 27074
rect 33234 27022 33236 27074
rect 33068 26852 33124 26862
rect 33068 26758 33124 26796
rect 32956 25788 33124 25844
rect 32956 25620 33012 25630
rect 32956 25526 33012 25564
rect 33068 24948 33124 25788
rect 33180 25620 33236 27022
rect 33404 27076 33460 29372
rect 33516 28868 33572 28878
rect 33516 28774 33572 28812
rect 33852 28868 33908 28878
rect 33852 28774 33908 28812
rect 33964 28756 34020 29932
rect 34412 29922 34468 29932
rect 34076 29428 34132 29438
rect 34076 29334 34132 29372
rect 34524 29426 34580 29438
rect 34524 29374 34526 29426
rect 34578 29374 34580 29426
rect 33964 28700 34132 28756
rect 33852 28420 33908 28430
rect 33740 27860 33796 27870
rect 33852 27860 33908 28364
rect 34076 27972 34132 28700
rect 34188 28644 34244 28654
rect 34188 28642 34356 28644
rect 34188 28590 34190 28642
rect 34242 28590 34356 28642
rect 34188 28588 34356 28590
rect 34188 28578 34244 28588
rect 34076 27916 34244 27972
rect 33852 27804 34132 27860
rect 33740 27766 33796 27804
rect 33964 27300 34020 27310
rect 33964 27186 34020 27244
rect 33964 27134 33966 27186
rect 34018 27134 34020 27186
rect 33964 27122 34020 27134
rect 34076 27188 34132 27804
rect 33404 26290 33460 27020
rect 33852 27076 33908 27114
rect 33852 27010 33908 27020
rect 34076 27074 34132 27132
rect 34076 27022 34078 27074
rect 34130 27022 34132 27074
rect 34076 27010 34132 27022
rect 34188 27076 34244 27916
rect 34300 27524 34356 28588
rect 34524 27860 34580 29374
rect 34636 27972 34692 30268
rect 34748 30210 34804 30380
rect 34748 30158 34750 30210
rect 34802 30158 34804 30210
rect 34748 30146 34804 30158
rect 34860 30996 34916 31006
rect 35084 30996 35140 31500
rect 35196 31490 35252 31500
rect 35980 31554 36036 31566
rect 35980 31502 35982 31554
rect 36034 31502 36036 31554
rect 35980 31444 36036 31502
rect 35980 31108 36036 31388
rect 35644 31052 36036 31108
rect 34860 30994 35084 30996
rect 34860 30942 34862 30994
rect 34914 30942 35084 30994
rect 34860 30940 35084 30942
rect 34748 28644 34804 28654
rect 34748 28084 34804 28588
rect 34860 28420 34916 30940
rect 35084 30902 35140 30940
rect 35308 30994 35364 31006
rect 35308 30942 35310 30994
rect 35362 30942 35364 30994
rect 35308 30772 35364 30942
rect 35644 30772 35700 31052
rect 35756 30884 35812 30894
rect 35980 30884 36036 30894
rect 35756 30882 35924 30884
rect 35756 30830 35758 30882
rect 35810 30830 35924 30882
rect 35756 30828 35924 30830
rect 35756 30818 35812 30828
rect 35308 30716 35700 30772
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35420 30436 35476 30446
rect 35084 30100 35140 30110
rect 35084 30006 35140 30044
rect 35420 30098 35476 30380
rect 35420 30046 35422 30098
rect 35474 30046 35476 30098
rect 35420 30034 35476 30046
rect 34972 29540 35028 29550
rect 34972 28644 35028 29484
rect 35196 29316 35252 29326
rect 35084 29314 35252 29316
rect 35084 29262 35198 29314
rect 35250 29262 35252 29314
rect 35084 29260 35252 29262
rect 35084 28868 35140 29260
rect 35196 29250 35252 29260
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 28868 35252 28878
rect 35084 28866 35252 28868
rect 35084 28814 35198 28866
rect 35250 28814 35252 28866
rect 35084 28812 35252 28814
rect 35196 28802 35252 28812
rect 35084 28644 35140 28654
rect 34972 28642 35140 28644
rect 34972 28590 35086 28642
rect 35138 28590 35140 28642
rect 34972 28588 35140 28590
rect 35084 28578 35140 28588
rect 34860 28364 35140 28420
rect 34748 28028 35028 28084
rect 34636 27916 34804 27972
rect 34524 27794 34580 27804
rect 34412 27748 34468 27758
rect 34412 27654 34468 27692
rect 34300 27468 34692 27524
rect 34300 27076 34356 27086
rect 34188 27074 34356 27076
rect 34188 27022 34302 27074
rect 34354 27022 34356 27074
rect 34188 27020 34356 27022
rect 34188 26908 34244 27020
rect 34300 27010 34356 27020
rect 34524 27076 34580 27086
rect 34524 26982 34580 27020
rect 33852 26852 34244 26908
rect 33740 26628 33796 26638
rect 33404 26238 33406 26290
rect 33458 26238 33460 26290
rect 33404 26226 33460 26238
rect 33628 26292 33684 26302
rect 33740 26292 33796 26572
rect 33852 26514 33908 26796
rect 33852 26462 33854 26514
rect 33906 26462 33908 26514
rect 33852 26450 33908 26462
rect 34636 26628 34692 27468
rect 34636 26514 34692 26572
rect 34636 26462 34638 26514
rect 34690 26462 34692 26514
rect 34636 26450 34692 26462
rect 33628 26290 33796 26292
rect 33628 26238 33630 26290
rect 33682 26238 33796 26290
rect 33628 26236 33796 26238
rect 34076 26290 34132 26302
rect 34076 26238 34078 26290
rect 34130 26238 34132 26290
rect 33628 26226 33684 26236
rect 33516 26178 33572 26190
rect 33516 26126 33518 26178
rect 33570 26126 33572 26178
rect 33180 25554 33236 25564
rect 33292 25620 33348 25630
rect 33516 25620 33572 26126
rect 33292 25618 33572 25620
rect 33292 25566 33294 25618
rect 33346 25566 33572 25618
rect 33292 25564 33572 25566
rect 33740 25620 33796 25630
rect 33292 25554 33348 25564
rect 33740 25526 33796 25564
rect 33404 25284 33460 25294
rect 33852 25284 33908 25294
rect 33404 25282 33572 25284
rect 33404 25230 33406 25282
rect 33458 25230 33572 25282
rect 33404 25228 33572 25230
rect 33404 25218 33460 25228
rect 33516 24948 33572 25228
rect 33852 25190 33908 25228
rect 33068 24892 33460 24948
rect 33516 24892 33908 24948
rect 33068 24722 33124 24734
rect 33068 24670 33070 24722
rect 33122 24670 33124 24722
rect 33068 23828 33124 24670
rect 33124 23772 33236 23828
rect 33068 23762 33124 23772
rect 33068 23156 33124 23166
rect 32844 23154 33124 23156
rect 32844 23102 33070 23154
rect 33122 23102 33124 23154
rect 32844 23100 33124 23102
rect 32732 22428 33012 22484
rect 32284 22260 32340 22270
rect 32844 22260 32900 22270
rect 32284 22166 32340 22204
rect 32732 22258 32900 22260
rect 32732 22206 32846 22258
rect 32898 22206 32900 22258
rect 32732 22204 32900 22206
rect 32396 22146 32452 22158
rect 32396 22094 32398 22146
rect 32450 22094 32452 22146
rect 32284 22036 32340 22046
rect 32396 22036 32452 22094
rect 32620 22148 32676 22158
rect 32620 22054 32676 22092
rect 32340 21980 32452 22036
rect 32284 21970 32340 21980
rect 32396 21812 32452 21822
rect 32732 21812 32788 22204
rect 32844 22194 32900 22204
rect 32396 21810 32788 21812
rect 32396 21758 32398 21810
rect 32450 21758 32788 21810
rect 32396 21756 32788 21758
rect 32844 22036 32900 22046
rect 32396 21746 32452 21756
rect 32284 21586 32340 21598
rect 32284 21534 32286 21586
rect 32338 21534 32340 21586
rect 32284 21476 32340 21534
rect 32508 21588 32564 21598
rect 32844 21588 32900 21980
rect 32564 21532 32900 21588
rect 32508 21494 32564 21532
rect 32284 19796 32340 21420
rect 32956 20020 33012 22428
rect 33068 21810 33124 23100
rect 33180 22370 33236 23772
rect 33292 23156 33348 23166
rect 33292 23062 33348 23100
rect 33180 22318 33182 22370
rect 33234 22318 33236 22370
rect 33180 22306 33236 22318
rect 33404 21924 33460 24892
rect 33852 24834 33908 24892
rect 33852 24782 33854 24834
rect 33906 24782 33908 24834
rect 33852 24770 33908 24782
rect 34076 24612 34132 26238
rect 34076 24546 34132 24556
rect 34636 23716 34692 23726
rect 34412 23660 34636 23716
rect 34300 23156 34356 23166
rect 34300 23062 34356 23100
rect 33852 23044 33908 23054
rect 33068 21758 33070 21810
rect 33122 21758 33124 21810
rect 33068 21746 33124 21758
rect 33180 21868 33460 21924
rect 33628 23042 33908 23044
rect 33628 22990 33854 23042
rect 33906 22990 33908 23042
rect 33628 22988 33908 22990
rect 32732 19964 33012 20020
rect 33180 20132 33236 21868
rect 33404 21698 33460 21710
rect 33404 21646 33406 21698
rect 33458 21646 33460 21698
rect 33292 20244 33348 20254
rect 33404 20244 33460 21646
rect 33348 20188 33460 20244
rect 33628 21588 33684 22988
rect 33852 22978 33908 22988
rect 33628 20242 33684 21532
rect 33740 22820 33796 22830
rect 33740 20804 33796 22764
rect 33964 22260 34020 22270
rect 33964 22166 34020 22204
rect 34412 21924 34468 23660
rect 34636 23650 34692 23660
rect 34748 23380 34804 27916
rect 34860 27748 34916 27758
rect 34860 23492 34916 27692
rect 34972 27186 35028 28028
rect 34972 27134 34974 27186
rect 35026 27134 35028 27186
rect 34972 23716 35028 27134
rect 34972 23650 35028 23660
rect 34860 23436 35028 23492
rect 34748 23314 34804 23324
rect 34972 23154 35028 23436
rect 34972 23102 34974 23154
rect 35026 23102 35028 23154
rect 34748 23044 34804 23054
rect 34748 22036 34804 22988
rect 34972 22932 35028 23102
rect 34972 22866 35028 22876
rect 34748 21970 34804 21980
rect 35084 21924 35140 28364
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35420 27188 35476 27198
rect 35420 27094 35476 27132
rect 35532 26908 35588 30716
rect 35868 29986 35924 30828
rect 35868 29934 35870 29986
rect 35922 29934 35924 29986
rect 35868 29652 35924 29934
rect 35868 29586 35924 29596
rect 35980 28754 36036 30828
rect 36092 30772 36148 32396
rect 36540 31780 36596 32508
rect 36540 31714 36596 31724
rect 36540 31554 36596 31566
rect 36540 31502 36542 31554
rect 36594 31502 36596 31554
rect 36204 31332 36260 31342
rect 36204 30882 36260 31276
rect 36540 30996 36596 31502
rect 36540 30902 36596 30940
rect 36204 30830 36206 30882
rect 36258 30830 36260 30882
rect 36204 30818 36260 30830
rect 36764 30884 36820 30894
rect 36876 30884 36932 34860
rect 37100 34914 37156 35868
rect 37660 35924 37716 36430
rect 37660 35858 37716 35868
rect 37996 36482 38388 36484
rect 37996 36430 38334 36482
rect 38386 36430 38388 36482
rect 37996 36428 38388 36430
rect 37324 35586 37380 35598
rect 37324 35534 37326 35586
rect 37378 35534 37380 35586
rect 37324 35026 37380 35534
rect 37548 35476 37604 35486
rect 37548 35138 37604 35420
rect 37996 35252 38052 36428
rect 38332 36418 38388 36428
rect 37548 35086 37550 35138
rect 37602 35086 37604 35138
rect 37548 35074 37604 35086
rect 37772 35196 38052 35252
rect 37772 35138 37828 35196
rect 37772 35086 37774 35138
rect 37826 35086 37828 35138
rect 37772 35074 37828 35086
rect 37324 34974 37326 35026
rect 37378 34974 37380 35026
rect 37324 34962 37380 34974
rect 37100 34862 37102 34914
rect 37154 34862 37156 34914
rect 37100 34850 37156 34862
rect 36988 34130 37044 34142
rect 36988 34078 36990 34130
rect 37042 34078 37044 34130
rect 36988 32564 37044 34078
rect 37436 34020 37492 34030
rect 37436 34018 37604 34020
rect 37436 33966 37438 34018
rect 37490 33966 37604 34018
rect 37436 33964 37604 33966
rect 37436 33954 37492 33964
rect 37324 33348 37380 33358
rect 37324 33254 37380 33292
rect 37548 33346 37604 33964
rect 37548 33294 37550 33346
rect 37602 33294 37604 33346
rect 37548 33236 37604 33294
rect 37996 33348 38052 35196
rect 38556 36372 38612 36382
rect 38556 34914 38612 36316
rect 38556 34862 38558 34914
rect 38610 34862 38612 34914
rect 38556 34850 38612 34862
rect 38220 34802 38276 34814
rect 38220 34750 38222 34802
rect 38274 34750 38276 34802
rect 38220 34468 38276 34750
rect 38220 34402 38276 34412
rect 38332 34804 38388 34814
rect 37996 33282 38052 33292
rect 38220 34244 38276 34254
rect 38220 33908 38276 34188
rect 38220 33346 38276 33852
rect 38220 33294 38222 33346
rect 38274 33294 38276 33346
rect 38220 33282 38276 33294
rect 37548 33170 37604 33180
rect 37884 33236 37940 33246
rect 37884 33142 37940 33180
rect 37436 33122 37492 33134
rect 37436 33070 37438 33122
rect 37490 33070 37492 33122
rect 37436 32788 37492 33070
rect 37212 32732 37492 32788
rect 37212 32674 37268 32732
rect 37212 32622 37214 32674
rect 37266 32622 37268 32674
rect 37212 32610 37268 32622
rect 36988 32498 37044 32508
rect 37772 31892 37828 31902
rect 37548 31780 37604 31790
rect 37100 31556 37156 31566
rect 37100 31462 37156 31500
rect 37436 31556 37492 31566
rect 37436 31462 37492 31500
rect 37436 30996 37492 31006
rect 37548 30996 37604 31724
rect 37772 31554 37828 31836
rect 38332 31890 38388 34748
rect 38668 34018 38724 34030
rect 38668 33966 38670 34018
rect 38722 33966 38724 34018
rect 38556 33348 38612 33358
rect 38556 33234 38612 33292
rect 38556 33182 38558 33234
rect 38610 33182 38612 33234
rect 38556 33170 38612 33182
rect 38668 32004 38724 33966
rect 38780 33572 38836 37100
rect 38892 34692 38948 34702
rect 38892 34598 38948 34636
rect 39004 34356 39060 42812
rect 39340 42754 39396 43036
rect 39340 42702 39342 42754
rect 39394 42702 39396 42754
rect 39340 42690 39396 42702
rect 39452 41860 39508 43148
rect 39228 41804 39508 41860
rect 39564 42754 39620 43652
rect 39676 43538 39732 43932
rect 39676 43486 39678 43538
rect 39730 43486 39732 43538
rect 39676 43474 39732 43486
rect 39788 44322 39844 44334
rect 39788 44270 39790 44322
rect 39842 44270 39844 44322
rect 39788 43876 39844 44270
rect 39900 44324 39956 45054
rect 39900 44258 39956 44268
rect 40124 44322 40180 44334
rect 40124 44270 40126 44322
rect 40178 44270 40180 44322
rect 39788 43538 39844 43820
rect 40124 43652 40180 44270
rect 40348 44212 40404 46398
rect 41804 46450 41860 46462
rect 41804 46398 41806 46450
rect 41858 46398 41860 46450
rect 41580 45778 41636 45790
rect 41580 45726 41582 45778
rect 41634 45726 41636 45778
rect 40684 45444 40740 45454
rect 40236 44156 40404 44212
rect 40572 44210 40628 44222
rect 40572 44158 40574 44210
rect 40626 44158 40628 44210
rect 40236 43708 40292 44156
rect 40460 44100 40516 44110
rect 40348 44098 40516 44100
rect 40348 44046 40462 44098
rect 40514 44046 40516 44098
rect 40348 44044 40516 44046
rect 40348 43876 40404 44044
rect 40460 44034 40516 44044
rect 40348 43810 40404 43820
rect 40460 43764 40516 43774
rect 40572 43708 40628 44158
rect 40236 43652 40404 43708
rect 40124 43586 40180 43596
rect 40348 43650 40404 43652
rect 40348 43598 40350 43650
rect 40402 43598 40404 43650
rect 40348 43586 40404 43598
rect 40460 43652 40628 43708
rect 39788 43486 39790 43538
rect 39842 43486 39844 43538
rect 39788 43474 39844 43486
rect 40012 43316 40068 43326
rect 39788 42980 39844 42990
rect 39788 42886 39844 42924
rect 39564 42702 39566 42754
rect 39618 42702 39620 42754
rect 39228 34580 39284 41804
rect 39452 41636 39508 41646
rect 39452 39618 39508 41580
rect 39564 40964 39620 42702
rect 39900 42644 39956 42654
rect 39900 42550 39956 42588
rect 39900 41860 39956 41870
rect 39900 41766 39956 41804
rect 40012 41636 40068 43260
rect 40236 43316 40292 43326
rect 40236 43314 40404 43316
rect 40236 43262 40238 43314
rect 40290 43262 40404 43314
rect 40236 43260 40404 43262
rect 40236 43250 40292 43260
rect 40236 43092 40292 43102
rect 40236 42756 40292 43036
rect 40124 42754 40292 42756
rect 40124 42702 40238 42754
rect 40290 42702 40292 42754
rect 40124 42700 40292 42702
rect 40124 41860 40180 42700
rect 40236 42690 40292 42700
rect 40236 42532 40292 42542
rect 40348 42532 40404 43260
rect 40292 42476 40404 42532
rect 40236 42194 40292 42476
rect 40236 42142 40238 42194
rect 40290 42142 40292 42194
rect 40236 42130 40292 42142
rect 40124 41794 40180 41804
rect 40348 41858 40404 41870
rect 40348 41806 40350 41858
rect 40402 41806 40404 41858
rect 40348 41748 40404 41806
rect 40348 41682 40404 41692
rect 40012 41570 40068 41580
rect 40236 41300 40292 41310
rect 40236 41206 40292 41244
rect 39676 40964 39732 40974
rect 39564 40908 39676 40964
rect 39676 39730 39732 40908
rect 40348 40628 40404 40638
rect 40460 40628 40516 43652
rect 40572 43092 40628 43102
rect 40684 43092 40740 45388
rect 41020 45108 41076 45118
rect 41020 45014 41076 45052
rect 40908 44884 40964 44894
rect 40908 44790 40964 44828
rect 41580 44548 41636 45726
rect 41692 45780 41748 45790
rect 41692 45686 41748 45724
rect 41804 45778 41860 46398
rect 43148 46004 43204 46014
rect 43260 46004 43316 49200
rect 45276 47124 45332 47134
rect 43148 46002 43260 46004
rect 43148 45950 43150 46002
rect 43202 45950 43260 46002
rect 43148 45948 43260 45950
rect 43148 45938 43204 45948
rect 43260 45910 43316 45948
rect 44940 46004 44996 46014
rect 45276 46004 45332 47068
rect 44940 46002 45332 46004
rect 44940 45950 44942 46002
rect 44994 45950 45332 46002
rect 44940 45948 45332 45950
rect 44940 45938 44996 45948
rect 43820 45892 43876 45902
rect 43820 45798 43876 45836
rect 45276 45890 45332 45948
rect 45276 45838 45278 45890
rect 45330 45838 45332 45890
rect 45276 45826 45332 45838
rect 41804 45726 41806 45778
rect 41858 45726 41860 45778
rect 41804 45714 41860 45726
rect 45500 45780 45556 45790
rect 45836 45780 45892 45790
rect 45500 45778 45892 45780
rect 45500 45726 45502 45778
rect 45554 45726 45838 45778
rect 45890 45726 45892 45778
rect 45500 45724 45892 45726
rect 45500 45714 45556 45724
rect 45836 45714 45892 45724
rect 46620 45780 46676 45790
rect 42252 45666 42308 45678
rect 42252 45614 42254 45666
rect 42306 45614 42308 45666
rect 41692 44996 41748 45006
rect 41692 44902 41748 44940
rect 41020 44324 41076 44334
rect 41020 44230 41076 44268
rect 41468 44324 41524 44334
rect 41132 43762 41188 43774
rect 41132 43710 41134 43762
rect 41186 43710 41188 43762
rect 41132 43708 41188 43710
rect 41020 43650 41076 43662
rect 41132 43652 41412 43708
rect 41020 43598 41022 43650
rect 41074 43598 41076 43650
rect 40908 43538 40964 43550
rect 40908 43486 40910 43538
rect 40962 43486 40964 43538
rect 40908 43316 40964 43486
rect 40908 43250 40964 43260
rect 40628 43036 40740 43092
rect 40572 43026 40628 43036
rect 41020 42868 41076 43598
rect 40908 42812 41076 42868
rect 40572 42756 40628 42794
rect 40572 42690 40628 42700
rect 40684 42756 40740 42766
rect 40908 42756 40964 42812
rect 40684 42754 40964 42756
rect 40684 42702 40686 42754
rect 40738 42702 40964 42754
rect 40684 42700 40964 42702
rect 41356 42756 41412 43652
rect 40684 42532 40740 42700
rect 41020 42644 41076 42654
rect 40908 42642 41076 42644
rect 40908 42590 41022 42642
rect 41074 42590 41076 42642
rect 40908 42588 41076 42590
rect 40684 42466 40740 42476
rect 40796 42530 40852 42542
rect 40796 42478 40798 42530
rect 40850 42478 40852 42530
rect 40796 42084 40852 42478
rect 40572 42028 40852 42084
rect 40572 41860 40628 42028
rect 40908 41972 40964 42588
rect 41020 42578 41076 42588
rect 41356 42082 41412 42700
rect 41468 42754 41524 44268
rect 41468 42702 41470 42754
rect 41522 42702 41524 42754
rect 41468 42690 41524 42702
rect 41580 42196 41636 44492
rect 41692 44210 41748 44222
rect 41692 44158 41694 44210
rect 41746 44158 41748 44210
rect 41692 43708 41748 44158
rect 42028 43876 42084 43886
rect 41692 43652 41972 43708
rect 41580 42194 41860 42196
rect 41580 42142 41582 42194
rect 41634 42142 41860 42194
rect 41580 42140 41860 42142
rect 41580 42130 41636 42140
rect 41356 42030 41358 42082
rect 41410 42030 41412 42082
rect 41356 42018 41412 42030
rect 40572 41794 40628 41804
rect 40684 41916 40964 41972
rect 41020 41972 41076 41982
rect 41020 41970 41188 41972
rect 41020 41918 41022 41970
rect 41074 41918 41188 41970
rect 41020 41916 41188 41918
rect 40684 41410 40740 41916
rect 41020 41906 41076 41916
rect 41132 41860 41188 41916
rect 41132 41804 41524 41860
rect 40908 41746 40964 41758
rect 40908 41694 40910 41746
rect 40962 41694 40964 41746
rect 40908 41636 40964 41694
rect 41020 41748 41076 41758
rect 41076 41692 41412 41748
rect 41020 41682 41076 41692
rect 40908 41570 40964 41580
rect 40684 41358 40686 41410
rect 40738 41358 40740 41410
rect 40684 41346 40740 41358
rect 40908 41300 40964 41310
rect 40572 41074 40628 41086
rect 40572 41022 40574 41074
rect 40626 41022 40628 41074
rect 40572 40964 40628 41022
rect 40572 40898 40628 40908
rect 40684 40962 40740 40974
rect 40684 40910 40686 40962
rect 40738 40910 40740 40962
rect 40404 40572 40516 40628
rect 39676 39678 39678 39730
rect 39730 39678 39732 39730
rect 39676 39666 39732 39678
rect 39900 40516 39956 40526
rect 39452 39566 39454 39618
rect 39506 39566 39508 39618
rect 39452 39554 39508 39566
rect 39788 39508 39844 39518
rect 39788 39058 39844 39452
rect 39788 39006 39790 39058
rect 39842 39006 39844 39058
rect 39788 38994 39844 39006
rect 39676 38836 39732 38846
rect 39788 38836 39844 38846
rect 39676 38834 39788 38836
rect 39676 38782 39678 38834
rect 39730 38782 39788 38834
rect 39676 38780 39788 38782
rect 39676 38770 39732 38780
rect 39788 38500 39844 38780
rect 39788 38434 39844 38444
rect 39900 38834 39956 40460
rect 39900 38782 39902 38834
rect 39954 38782 39956 38834
rect 39900 38276 39956 38782
rect 40124 38722 40180 38734
rect 40124 38670 40126 38722
rect 40178 38670 40180 38722
rect 40124 38668 40180 38670
rect 40348 38722 40404 40572
rect 40684 40516 40740 40910
rect 40684 40450 40740 40460
rect 40908 40402 40964 41244
rect 40908 40350 40910 40402
rect 40962 40350 40964 40402
rect 40908 39618 40964 40350
rect 41356 41298 41412 41692
rect 41356 41246 41358 41298
rect 41410 41246 41412 41298
rect 40908 39566 40910 39618
rect 40962 39566 40964 39618
rect 40908 39554 40964 39566
rect 41244 39618 41300 39630
rect 41244 39566 41246 39618
rect 41298 39566 41300 39618
rect 40460 39394 40516 39406
rect 40460 39342 40462 39394
rect 40514 39342 40516 39394
rect 40460 38836 40516 39342
rect 40460 38770 40516 38780
rect 41132 38836 41188 38846
rect 41244 38836 41300 39566
rect 41132 38834 41300 38836
rect 41132 38782 41134 38834
rect 41186 38782 41300 38834
rect 41132 38780 41300 38782
rect 41356 39506 41412 41246
rect 41468 40516 41524 41804
rect 41692 41748 41748 41758
rect 41692 41654 41748 41692
rect 41468 40402 41524 40460
rect 41468 40350 41470 40402
rect 41522 40350 41524 40402
rect 41468 40338 41524 40350
rect 41804 40180 41860 42140
rect 41916 42084 41972 43652
rect 42028 43538 42084 43820
rect 42028 43486 42030 43538
rect 42082 43486 42084 43538
rect 42028 43474 42084 43486
rect 42252 43428 42308 45614
rect 43596 45668 43652 45678
rect 43596 45574 43652 45612
rect 45948 45666 46004 45678
rect 45948 45614 45950 45666
rect 46002 45614 46004 45666
rect 42924 45106 42980 45118
rect 42924 45054 42926 45106
rect 42978 45054 42980 45106
rect 42924 44996 42980 45054
rect 42924 43708 42980 44940
rect 43708 44996 43764 45006
rect 42476 43652 42532 43662
rect 42924 43652 43092 43708
rect 42476 43558 42532 43596
rect 42588 43428 42644 43438
rect 42252 43372 42588 43428
rect 42252 42980 42308 42990
rect 42140 42644 42196 42654
rect 42140 42550 42196 42588
rect 42028 42084 42084 42094
rect 41916 42082 42084 42084
rect 41916 42030 42030 42082
rect 42082 42030 42084 42082
rect 41916 42028 42084 42030
rect 42028 42018 42084 42028
rect 42140 41972 42196 41982
rect 42252 41972 42308 42924
rect 42140 41970 42308 41972
rect 42140 41918 42142 41970
rect 42194 41918 42308 41970
rect 42140 41916 42308 41918
rect 42588 41970 42644 43372
rect 42588 41918 42590 41970
rect 42642 41918 42644 41970
rect 42140 41906 42196 41916
rect 42588 41906 42644 41918
rect 43036 41970 43092 43652
rect 43372 43428 43428 43438
rect 43372 43334 43428 43372
rect 43036 41918 43038 41970
rect 43090 41918 43092 41970
rect 42364 41748 42420 41758
rect 42364 41654 42420 41692
rect 41916 40404 41972 40414
rect 41916 40310 41972 40348
rect 42588 40404 42644 40414
rect 43036 40404 43092 41918
rect 43484 41860 43540 41870
rect 43484 41298 43540 41804
rect 43484 41246 43486 41298
rect 43538 41246 43540 41298
rect 43484 41234 43540 41246
rect 42588 40310 42644 40348
rect 42924 40348 43036 40404
rect 41804 40124 42196 40180
rect 41692 39730 41748 39742
rect 41692 39678 41694 39730
rect 41746 39678 41748 39730
rect 41692 39620 41748 39678
rect 42028 39620 42084 39630
rect 41356 39454 41358 39506
rect 41410 39454 41412 39506
rect 40348 38670 40350 38722
rect 40402 38670 40404 38722
rect 40124 38612 40292 38668
rect 39676 38220 39956 38276
rect 40124 38500 40180 38510
rect 39676 38162 39732 38220
rect 39676 38110 39678 38162
rect 39730 38110 39732 38162
rect 39676 38098 39732 38110
rect 40124 38052 40180 38444
rect 40236 38388 40292 38612
rect 40236 38322 40292 38332
rect 40124 37492 40180 37996
rect 40348 38052 40404 38670
rect 40348 37986 40404 37996
rect 40124 37426 40180 37436
rect 41020 37492 41076 37502
rect 41020 37398 41076 37436
rect 40012 37156 40068 37166
rect 40012 37062 40068 37100
rect 40908 37156 40964 37166
rect 40908 37062 40964 37100
rect 40348 37044 40404 37054
rect 40348 36706 40404 36988
rect 40348 36654 40350 36706
rect 40402 36654 40404 36706
rect 40348 36642 40404 36654
rect 39900 36484 39956 36494
rect 39788 36372 39844 36382
rect 39788 36278 39844 36316
rect 39900 35922 39956 36428
rect 40572 36482 40628 36494
rect 40572 36430 40574 36482
rect 40626 36430 40628 36482
rect 39900 35870 39902 35922
rect 39954 35870 39956 35922
rect 39788 35700 39844 35710
rect 39452 35698 39844 35700
rect 39452 35646 39790 35698
rect 39842 35646 39844 35698
rect 39452 35644 39844 35646
rect 39452 35586 39508 35644
rect 39788 35634 39844 35644
rect 39452 35534 39454 35586
rect 39506 35534 39508 35586
rect 39452 35522 39508 35534
rect 39900 35476 39956 35870
rect 40012 36370 40068 36382
rect 40012 36318 40014 36370
rect 40066 36318 40068 36370
rect 40012 35924 40068 36318
rect 40124 36372 40180 36382
rect 40124 36370 40292 36372
rect 40124 36318 40126 36370
rect 40178 36318 40292 36370
rect 40124 36316 40292 36318
rect 40124 36306 40180 36316
rect 40012 35858 40068 35868
rect 39900 35410 39956 35420
rect 40236 35028 40292 36316
rect 40572 35476 40628 36430
rect 41132 36484 41188 38780
rect 41356 38722 41412 39454
rect 41356 38670 41358 38722
rect 41410 38670 41412 38722
rect 41356 38658 41412 38670
rect 41468 39618 42084 39620
rect 41468 39566 42030 39618
rect 42082 39566 42084 39618
rect 41468 39564 42084 39566
rect 41468 38388 41524 39564
rect 42028 39554 42084 39564
rect 42140 39060 42196 40124
rect 42588 39618 42644 39630
rect 42588 39566 42590 39618
rect 42642 39566 42644 39618
rect 42476 39508 42532 39518
rect 42476 39414 42532 39452
rect 42364 39396 42420 39406
rect 42364 39302 42420 39340
rect 42140 38834 42196 39004
rect 42140 38782 42142 38834
rect 42194 38782 42196 38834
rect 42140 38770 42196 38782
rect 41916 38722 41972 38734
rect 41916 38670 41918 38722
rect 41970 38670 41972 38722
rect 41916 38612 41972 38670
rect 42588 38668 42644 39566
rect 41804 38556 41916 38612
rect 41244 38332 41524 38388
rect 41580 38388 41636 38398
rect 41244 38050 41300 38332
rect 41244 37998 41246 38050
rect 41298 37998 41300 38050
rect 41244 37986 41300 37998
rect 41580 37940 41636 38332
rect 41356 37884 41636 37940
rect 41356 36594 41412 37884
rect 41356 36542 41358 36594
rect 41410 36542 41412 36594
rect 41356 36530 41412 36542
rect 41580 37268 41636 37278
rect 41132 36418 41188 36428
rect 40572 35410 40628 35420
rect 41020 36370 41076 36382
rect 41020 36318 41022 36370
rect 41074 36318 41076 36370
rect 40460 35028 40516 35038
rect 40236 35026 40516 35028
rect 40236 34974 40462 35026
rect 40514 34974 40516 35026
rect 40236 34972 40516 34974
rect 40460 34962 40516 34972
rect 39788 34916 39844 34926
rect 39788 34822 39844 34860
rect 39228 34514 39284 34524
rect 39340 34690 39396 34702
rect 39340 34638 39342 34690
rect 39394 34638 39396 34690
rect 39004 34290 39060 34300
rect 39340 34244 39396 34638
rect 39676 34244 39732 34254
rect 40012 34244 40068 34254
rect 39340 34242 39956 34244
rect 39340 34190 39678 34242
rect 39730 34190 39956 34242
rect 39340 34188 39956 34190
rect 39676 34178 39732 34188
rect 39340 34018 39396 34030
rect 39340 33966 39342 34018
rect 39394 33966 39396 34018
rect 39340 33572 39396 33966
rect 38780 33506 38836 33516
rect 39004 33516 39396 33572
rect 39788 34020 39844 34030
rect 38780 33348 38836 33358
rect 38780 33254 38836 33292
rect 38668 31938 38724 31948
rect 38780 33124 38836 33134
rect 39004 33124 39060 33516
rect 39788 33460 39844 33964
rect 39900 33908 39956 34188
rect 40012 34150 40068 34188
rect 40348 34242 40404 34254
rect 40348 34190 40350 34242
rect 40402 34190 40404 34242
rect 39900 33852 40068 33908
rect 39340 33404 39844 33460
rect 38836 33068 39060 33124
rect 39116 33348 39172 33358
rect 39116 33122 39172 33292
rect 39116 33070 39118 33122
rect 39170 33070 39172 33122
rect 38332 31838 38334 31890
rect 38386 31838 38388 31890
rect 38332 31826 38388 31838
rect 38780 31780 38836 33068
rect 39116 33058 39172 33070
rect 39228 33234 39284 33246
rect 39228 33182 39230 33234
rect 39282 33182 39284 33234
rect 39228 33124 39284 33182
rect 37772 31502 37774 31554
rect 37826 31502 37828 31554
rect 37772 31444 37828 31502
rect 37772 31378 37828 31388
rect 38668 31724 38836 31780
rect 38668 31666 38724 31724
rect 38668 31614 38670 31666
rect 38722 31614 38724 31666
rect 38668 31444 38724 31614
rect 38668 31378 38724 31388
rect 38780 31556 38836 31566
rect 39228 31556 39284 33068
rect 39340 32450 39396 33404
rect 39788 33346 39844 33404
rect 39788 33294 39790 33346
rect 39842 33294 39844 33346
rect 39788 33282 39844 33294
rect 40012 33346 40068 33852
rect 40012 33294 40014 33346
rect 40066 33294 40068 33346
rect 39452 33236 39508 33246
rect 39900 33236 39956 33246
rect 39452 33234 39732 33236
rect 39452 33182 39454 33234
rect 39506 33182 39732 33234
rect 39452 33180 39732 33182
rect 39452 33170 39508 33180
rect 39676 32788 39732 33180
rect 39900 33142 39956 33180
rect 39788 32788 39844 32798
rect 39676 32786 39844 32788
rect 39676 32734 39790 32786
rect 39842 32734 39844 32786
rect 39676 32732 39844 32734
rect 39788 32722 39844 32732
rect 39676 32564 39732 32574
rect 39676 32470 39732 32508
rect 39900 32564 39956 32574
rect 40012 32564 40068 33294
rect 40348 33234 40404 34190
rect 40908 34244 40964 34254
rect 40908 34150 40964 34188
rect 41020 34020 41076 36318
rect 41244 35700 41300 35710
rect 41020 33954 41076 33964
rect 41132 35644 41244 35700
rect 41132 34916 41188 35644
rect 41244 35634 41300 35644
rect 40908 33348 40964 33358
rect 41132 33348 41188 34860
rect 41244 35476 41300 35486
rect 41244 34354 41300 35420
rect 41244 34302 41246 34354
rect 41298 34302 41300 34354
rect 41244 34290 41300 34302
rect 41580 33684 41636 37212
rect 41804 37044 41860 38556
rect 41916 38546 41972 38556
rect 42028 38612 42644 38668
rect 42700 38948 42756 38958
rect 42028 38610 42084 38612
rect 42028 38558 42030 38610
rect 42082 38558 42084 38610
rect 41916 38052 41972 38062
rect 41916 37958 41972 37996
rect 41916 37268 41972 37278
rect 42028 37268 42084 38558
rect 42588 37492 42644 37502
rect 42700 37492 42756 38892
rect 42588 37490 42756 37492
rect 42588 37438 42590 37490
rect 42642 37438 42756 37490
rect 42588 37436 42756 37438
rect 42588 37426 42644 37436
rect 41916 37266 42084 37268
rect 41916 37214 41918 37266
rect 41970 37214 42084 37266
rect 41916 37212 42084 37214
rect 41916 37202 41972 37212
rect 41692 35924 41748 35934
rect 41804 35924 41860 36988
rect 42252 36260 42308 36270
rect 42700 36260 42756 36270
rect 42252 36258 42756 36260
rect 42252 36206 42254 36258
rect 42306 36206 42702 36258
rect 42754 36206 42756 36258
rect 42252 36204 42756 36206
rect 42252 36194 42308 36204
rect 41916 35924 41972 35934
rect 41804 35922 41972 35924
rect 41804 35870 41918 35922
rect 41970 35870 41972 35922
rect 41804 35868 41972 35870
rect 41692 35830 41748 35868
rect 41916 35858 41972 35868
rect 42028 35700 42084 35710
rect 42476 35700 42532 35710
rect 42028 35698 42420 35700
rect 42028 35646 42030 35698
rect 42082 35646 42420 35698
rect 42028 35644 42420 35646
rect 42028 35634 42084 35644
rect 42364 35364 42420 35644
rect 42476 35606 42532 35644
rect 42700 35588 42756 36204
rect 42700 35522 42756 35532
rect 42812 35476 42868 35486
rect 42364 35308 42644 35364
rect 42588 35026 42644 35308
rect 42588 34974 42590 35026
rect 42642 34974 42644 35026
rect 42588 34962 42644 34974
rect 42812 35028 42868 35420
rect 42924 35140 42980 40348
rect 43036 40338 43092 40348
rect 43708 39732 43764 44940
rect 44828 44994 44884 45006
rect 44828 44942 44830 44994
rect 44882 44942 44884 44994
rect 43820 44548 43876 44558
rect 43820 44434 43876 44492
rect 43820 44382 43822 44434
rect 43874 44382 43876 44434
rect 43820 44370 43876 44382
rect 44828 44324 44884 44942
rect 44828 44230 44884 44268
rect 45612 44210 45668 44222
rect 45612 44158 45614 44210
rect 45666 44158 45668 44210
rect 45612 43708 45668 44158
rect 44828 43652 44884 43662
rect 44828 43558 44884 43596
rect 44940 43652 45668 43708
rect 43820 43538 43876 43550
rect 43820 43486 43822 43538
rect 43874 43486 43876 43538
rect 43820 42532 43876 43486
rect 44268 43428 44324 43438
rect 44604 43428 44660 43438
rect 44268 43426 44660 43428
rect 44268 43374 44270 43426
rect 44322 43374 44606 43426
rect 44658 43374 44660 43426
rect 44268 43372 44660 43374
rect 44268 43362 44324 43372
rect 44604 43362 44660 43372
rect 44940 43426 44996 43652
rect 45724 43540 45780 43550
rect 44940 43374 44942 43426
rect 44994 43374 44996 43426
rect 44940 43362 44996 43374
rect 45276 43426 45332 43438
rect 45276 43374 45278 43426
rect 45330 43374 45332 43426
rect 44268 42868 44324 42878
rect 44268 42866 45108 42868
rect 44268 42814 44270 42866
rect 44322 42814 45108 42866
rect 44268 42812 45108 42814
rect 44268 42802 44324 42812
rect 44940 42644 44996 42654
rect 44940 42550 44996 42588
rect 44828 42532 44884 42542
rect 43820 42530 44884 42532
rect 43820 42478 44830 42530
rect 44882 42478 44884 42530
rect 43820 42476 44884 42478
rect 44268 41188 44324 41198
rect 44268 41094 44324 41132
rect 44604 40404 44660 40414
rect 44604 40310 44660 40348
rect 43708 39676 44324 39732
rect 44044 39508 44100 39518
rect 43932 39506 44100 39508
rect 43932 39454 44046 39506
rect 44098 39454 44100 39506
rect 43932 39452 44100 39454
rect 43484 39396 43540 39406
rect 43148 39060 43204 39070
rect 43148 38966 43204 39004
rect 43036 38834 43092 38846
rect 43036 38782 43038 38834
rect 43090 38782 43092 38834
rect 43036 38612 43092 38782
rect 43036 38546 43092 38556
rect 43372 38834 43428 38846
rect 43372 38782 43374 38834
rect 43426 38782 43428 38834
rect 43148 38388 43204 38398
rect 43036 38332 43148 38388
rect 43036 38050 43092 38332
rect 43148 38322 43204 38332
rect 43148 38164 43204 38174
rect 43148 38070 43204 38108
rect 43036 37998 43038 38050
rect 43090 37998 43092 38050
rect 43036 37986 43092 37998
rect 43036 37380 43092 37390
rect 43036 36706 43092 37324
rect 43036 36654 43038 36706
rect 43090 36654 43092 36706
rect 43036 36642 43092 36654
rect 43260 36484 43316 36494
rect 43372 36484 43428 38782
rect 43484 38050 43540 39340
rect 43820 39394 43876 39406
rect 43820 39342 43822 39394
rect 43874 39342 43876 39394
rect 43820 39172 43876 39342
rect 43820 39106 43876 39116
rect 43708 38836 43764 38846
rect 43708 38742 43764 38780
rect 43932 38668 43988 39452
rect 44044 39442 44100 39452
rect 43708 38612 43988 38668
rect 44156 39394 44212 39406
rect 44156 39342 44158 39394
rect 44210 39342 44212 39394
rect 44156 38834 44212 39342
rect 44156 38782 44158 38834
rect 44210 38782 44212 38834
rect 43596 38164 43652 38174
rect 43708 38164 43764 38612
rect 44156 38276 44212 38782
rect 44156 38210 44212 38220
rect 43596 38162 43764 38164
rect 43596 38110 43598 38162
rect 43650 38110 43764 38162
rect 43596 38108 43764 38110
rect 43932 38164 43988 38174
rect 43596 38098 43652 38108
rect 43484 37998 43486 38050
rect 43538 37998 43540 38050
rect 43484 37986 43540 37998
rect 43708 37826 43764 37838
rect 43708 37774 43710 37826
rect 43762 37774 43764 37826
rect 43708 37380 43764 37774
rect 43708 37314 43764 37324
rect 43820 37828 43876 37838
rect 43260 36482 43428 36484
rect 43260 36430 43262 36482
rect 43314 36430 43428 36482
rect 43260 36428 43428 36430
rect 43820 36594 43876 37772
rect 43932 37266 43988 38108
rect 44156 38050 44212 38062
rect 44156 37998 44158 38050
rect 44210 37998 44212 38050
rect 44156 37940 44212 37998
rect 44156 37874 44212 37884
rect 43932 37214 43934 37266
rect 43986 37214 43988 37266
rect 43932 37202 43988 37214
rect 44268 36708 44324 39676
rect 44380 39396 44436 39406
rect 44380 39302 44436 39340
rect 44716 38668 44772 42476
rect 44828 42466 44884 42476
rect 45052 40404 45108 42812
rect 45276 42644 45332 43374
rect 45612 43092 45668 43102
rect 45612 42754 45668 43036
rect 45612 42702 45614 42754
rect 45666 42702 45668 42754
rect 45500 42644 45556 42654
rect 45276 42642 45556 42644
rect 45276 42590 45502 42642
rect 45554 42590 45556 42642
rect 45276 42588 45556 42590
rect 45500 42084 45556 42588
rect 45612 42644 45668 42702
rect 45724 42756 45780 43484
rect 45724 42662 45780 42700
rect 45612 42578 45668 42588
rect 45500 42018 45556 42028
rect 45276 41300 45332 41310
rect 45276 41298 45444 41300
rect 45276 41246 45278 41298
rect 45330 41246 45444 41298
rect 45276 41244 45444 41246
rect 45276 41234 45332 41244
rect 45388 40404 45444 41244
rect 45948 40852 46004 45614
rect 46508 45666 46564 45678
rect 46508 45614 46510 45666
rect 46562 45614 46564 45666
rect 46508 45556 46564 45614
rect 46508 43652 46564 45500
rect 46396 42756 46452 42766
rect 46396 42662 46452 42700
rect 46172 42532 46228 42542
rect 46284 42532 46340 42542
rect 46172 42530 46284 42532
rect 46172 42478 46174 42530
rect 46226 42478 46284 42530
rect 46172 42476 46284 42478
rect 46172 42466 46228 42476
rect 45948 40786 46004 40796
rect 45612 40404 45668 40414
rect 45052 40402 45332 40404
rect 45052 40350 45054 40402
rect 45106 40350 45332 40402
rect 45052 40348 45332 40350
rect 45388 40402 45668 40404
rect 45388 40350 45614 40402
rect 45666 40350 45668 40402
rect 45388 40348 45668 40350
rect 45052 40338 45108 40348
rect 45276 40292 45332 40348
rect 45276 40236 45444 40292
rect 44940 39844 44996 39854
rect 44940 39750 44996 39788
rect 45276 39730 45332 39742
rect 45276 39678 45278 39730
rect 45330 39678 45332 39730
rect 44828 39620 44884 39630
rect 45276 39620 45332 39678
rect 44828 39618 45332 39620
rect 44828 39566 44830 39618
rect 44882 39566 45332 39618
rect 44828 39564 45332 39566
rect 44828 39554 44884 39564
rect 45276 39060 45332 39564
rect 45276 38994 45332 39004
rect 44940 38948 44996 38958
rect 44940 38834 44996 38892
rect 45052 38948 45108 38958
rect 45052 38946 45220 38948
rect 45052 38894 45054 38946
rect 45106 38894 45220 38946
rect 45052 38892 45220 38894
rect 45052 38882 45108 38892
rect 44940 38782 44942 38834
rect 44994 38782 44996 38834
rect 44940 38770 44996 38782
rect 44380 38612 44436 38622
rect 44716 38612 44884 38668
rect 44380 38610 44548 38612
rect 44380 38558 44382 38610
rect 44434 38558 44548 38610
rect 44380 38556 44548 38558
rect 44380 38546 44436 38556
rect 44492 37378 44548 38556
rect 44492 37326 44494 37378
rect 44546 37326 44548 37378
rect 44492 37314 44548 37326
rect 44828 38050 44884 38612
rect 44828 37998 44830 38050
rect 44882 37998 44884 38050
rect 44268 36642 44324 36652
rect 43820 36542 43822 36594
rect 43874 36542 43876 36594
rect 43260 36418 43316 36428
rect 43148 35588 43204 35598
rect 43596 35588 43652 35598
rect 43148 35586 43540 35588
rect 43148 35534 43150 35586
rect 43202 35534 43540 35586
rect 43148 35532 43540 35534
rect 43148 35522 43204 35532
rect 43260 35364 43316 35374
rect 42924 35084 43204 35140
rect 42812 34972 43092 35028
rect 43036 34914 43092 34972
rect 43036 34862 43038 34914
rect 43090 34862 43092 34914
rect 43036 34850 43092 34862
rect 43148 34692 43204 35084
rect 43260 35138 43316 35308
rect 43260 35086 43262 35138
rect 43314 35086 43316 35138
rect 43260 35074 43316 35086
rect 43484 35026 43540 35532
rect 43484 34974 43486 35026
rect 43538 34974 43540 35026
rect 43484 34962 43540 34974
rect 43596 34804 43652 35532
rect 43820 35140 43876 36542
rect 43932 36484 43988 36494
rect 44828 36484 44884 37998
rect 44940 38052 44996 38062
rect 44940 36596 44996 37996
rect 45164 37940 45220 38892
rect 45388 38946 45444 40236
rect 45388 38894 45390 38946
rect 45442 38894 45444 38946
rect 45388 38882 45444 38894
rect 45052 37828 45108 37838
rect 45052 37734 45108 37772
rect 45164 37826 45220 37884
rect 45164 37774 45166 37826
rect 45218 37774 45220 37826
rect 45164 37762 45220 37774
rect 45500 37492 45556 40348
rect 45612 40338 45668 40348
rect 45724 40402 45780 40414
rect 45724 40350 45726 40402
rect 45778 40350 45780 40402
rect 45724 40180 45780 40350
rect 45724 40114 45780 40124
rect 46284 40290 46340 42476
rect 46284 40238 46286 40290
rect 46338 40238 46340 40290
rect 45836 39060 45892 39070
rect 45836 38966 45892 39004
rect 45612 38834 45668 38846
rect 45612 38782 45614 38834
rect 45666 38782 45668 38834
rect 45612 38388 45668 38782
rect 45724 38836 45780 38846
rect 45724 38742 45780 38780
rect 45948 38836 46004 38846
rect 45612 38322 45668 38332
rect 45724 38052 45780 38062
rect 45724 37958 45780 37996
rect 45836 37940 45892 37950
rect 45836 37846 45892 37884
rect 45500 37426 45556 37436
rect 44940 36594 45332 36596
rect 44940 36542 44942 36594
rect 44994 36542 45332 36594
rect 44940 36540 45332 36542
rect 44940 36530 44996 36540
rect 43932 36482 44884 36484
rect 43932 36430 43934 36482
rect 43986 36430 44884 36482
rect 43932 36428 44884 36430
rect 43932 36418 43988 36428
rect 44828 36260 44884 36270
rect 44828 35364 44884 36204
rect 44828 35298 44884 35308
rect 44940 35588 44996 35598
rect 43820 35084 44436 35140
rect 43596 34710 43652 34748
rect 43820 34804 43876 34814
rect 43820 34802 44212 34804
rect 43820 34750 43822 34802
rect 43874 34750 44212 34802
rect 43820 34748 44212 34750
rect 43820 34738 43876 34748
rect 42476 34356 42532 34366
rect 42140 34132 42196 34142
rect 42140 34038 42196 34076
rect 41580 33618 41636 33628
rect 41692 34018 41748 34030
rect 41692 33966 41694 34018
rect 41746 33966 41748 34018
rect 40908 33346 41188 33348
rect 40908 33294 40910 33346
rect 40962 33294 41188 33346
rect 40908 33292 41188 33294
rect 40908 33282 40964 33292
rect 40348 33182 40350 33234
rect 40402 33182 40404 33234
rect 40348 33012 40404 33182
rect 40236 32956 40348 33012
rect 40236 32674 40292 32956
rect 40348 32946 40404 32956
rect 40236 32622 40238 32674
rect 40290 32622 40292 32674
rect 40236 32610 40292 32622
rect 39900 32562 40068 32564
rect 39900 32510 39902 32562
rect 39954 32510 40068 32562
rect 39900 32508 40068 32510
rect 41132 32562 41188 33292
rect 41580 33348 41636 33358
rect 41580 33254 41636 33292
rect 41692 33124 41748 33966
rect 41692 33058 41748 33068
rect 42476 34018 42532 34300
rect 43148 34130 43204 34636
rect 43148 34078 43150 34130
rect 43202 34078 43204 34130
rect 43148 34066 43204 34078
rect 43708 34692 43764 34702
rect 42476 33966 42478 34018
rect 42530 33966 42532 34018
rect 41132 32510 41134 32562
rect 41186 32510 41188 32562
rect 39340 32398 39342 32450
rect 39394 32398 39396 32450
rect 39340 32386 39396 32398
rect 38780 31554 39284 31556
rect 38780 31502 38782 31554
rect 38834 31502 39284 31554
rect 38780 31500 39284 31502
rect 39564 31780 39620 31790
rect 38780 31220 38836 31500
rect 37436 30994 37604 30996
rect 37436 30942 37438 30994
rect 37490 30942 37604 30994
rect 37436 30940 37604 30942
rect 38668 31164 38836 31220
rect 37436 30930 37492 30940
rect 36820 30828 36932 30884
rect 38108 30882 38164 30894
rect 38108 30830 38110 30882
rect 38162 30830 38164 30882
rect 36764 30818 36820 30828
rect 36092 30706 36148 30716
rect 36428 30212 36484 30222
rect 36988 30212 37044 30222
rect 35980 28702 35982 28754
rect 36034 28702 36036 28754
rect 35980 28690 36036 28702
rect 36204 30210 37044 30212
rect 36204 30158 36430 30210
rect 36482 30158 36990 30210
rect 37042 30158 37044 30210
rect 36204 30156 37044 30158
rect 35532 26852 35812 26908
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35420 23154 35476 23166
rect 35420 23102 35422 23154
rect 35474 23102 35476 23154
rect 35420 23044 35476 23102
rect 35532 23156 35588 23166
rect 35532 23062 35588 23100
rect 35644 23154 35700 23166
rect 35644 23102 35646 23154
rect 35698 23102 35700 23154
rect 35420 22978 35476 22988
rect 35532 22932 35588 22942
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35084 21868 35252 21924
rect 34412 21858 34468 21868
rect 34188 21700 34244 21710
rect 34188 21606 34244 21644
rect 34636 21700 34692 21710
rect 34636 21606 34692 21644
rect 33964 21588 34020 21598
rect 34412 21588 34468 21598
rect 35084 21588 35140 21598
rect 33964 21586 34132 21588
rect 33964 21534 33966 21586
rect 34018 21534 34132 21586
rect 33964 21532 34132 21534
rect 33964 21522 34020 21532
rect 34076 21140 34132 21532
rect 34412 21494 34468 21532
rect 34860 21586 35140 21588
rect 34860 21534 35086 21586
rect 35138 21534 35140 21586
rect 34860 21532 35140 21534
rect 34300 21474 34356 21486
rect 34300 21422 34302 21474
rect 34354 21422 34356 21474
rect 34300 21364 34356 21422
rect 34860 21364 34916 21532
rect 35084 21522 35140 21532
rect 34300 21308 34916 21364
rect 34972 21362 35028 21374
rect 35196 21364 35252 21868
rect 35532 21810 35588 22876
rect 35644 22148 35700 23102
rect 35644 22082 35700 22092
rect 35532 21758 35534 21810
rect 35586 21758 35588 21810
rect 35532 21746 35588 21758
rect 34972 21310 34974 21362
rect 35026 21310 35028 21362
rect 34972 21252 35028 21310
rect 34972 21186 35028 21196
rect 35084 21308 35252 21364
rect 34076 21084 34244 21140
rect 33964 20804 34020 20814
rect 33740 20802 34020 20804
rect 33740 20750 33966 20802
rect 34018 20750 34020 20802
rect 33740 20748 34020 20750
rect 33964 20738 34020 20748
rect 33628 20190 33630 20242
rect 33682 20190 33684 20242
rect 33292 20150 33348 20188
rect 32396 19908 32452 19918
rect 32396 19814 32452 19852
rect 32284 19730 32340 19740
rect 32508 19794 32564 19806
rect 32508 19742 32510 19794
rect 32562 19742 32564 19794
rect 32508 19348 32564 19742
rect 32620 19348 32676 19358
rect 32508 19346 32676 19348
rect 32508 19294 32622 19346
rect 32674 19294 32676 19346
rect 32508 19292 32676 19294
rect 32620 19282 32676 19292
rect 32732 19124 32788 19964
rect 32844 19796 32900 19806
rect 32900 19740 33012 19796
rect 32844 19730 32900 19740
rect 32284 19068 32788 19124
rect 32284 18452 32340 19068
rect 32284 18450 32452 18452
rect 32284 18398 32286 18450
rect 32338 18398 32452 18450
rect 32284 18396 32452 18398
rect 32284 18386 32340 18396
rect 32396 17666 32452 18396
rect 32396 17614 32398 17666
rect 32450 17614 32452 17666
rect 32396 17602 32452 17614
rect 32732 17444 32788 17454
rect 32732 17350 32788 17388
rect 32284 17108 32340 17118
rect 32284 16994 32340 17052
rect 32284 16942 32286 16994
rect 32338 16942 32340 16994
rect 32284 16930 32340 16942
rect 32396 16660 32452 16670
rect 32396 16658 32900 16660
rect 32396 16606 32398 16658
rect 32450 16606 32900 16658
rect 32396 16604 32900 16606
rect 32396 16594 32452 16604
rect 32844 16210 32900 16604
rect 32844 16158 32846 16210
rect 32898 16158 32900 16210
rect 32844 16146 32900 16158
rect 32956 14532 33012 19740
rect 33180 19236 33236 20076
rect 33180 19170 33236 19180
rect 33404 20018 33460 20030
rect 33404 19966 33406 20018
rect 33458 19966 33460 20018
rect 33180 18338 33236 18350
rect 33180 18286 33182 18338
rect 33234 18286 33236 18338
rect 33180 18228 33236 18286
rect 33180 18162 33236 18172
rect 33180 17666 33236 17678
rect 33180 17614 33182 17666
rect 33234 17614 33236 17666
rect 33180 17444 33236 17614
rect 33180 17378 33236 17388
rect 32956 14466 33012 14476
rect 33292 16772 33348 16782
rect 33180 13748 33236 13758
rect 33180 13654 33236 13692
rect 32396 13636 32452 13646
rect 32396 13542 32452 13580
rect 32508 13524 32564 13534
rect 32508 13522 33124 13524
rect 32508 13470 32510 13522
rect 32562 13470 33124 13522
rect 32508 13468 33124 13470
rect 32508 13458 32564 13468
rect 33068 13076 33124 13468
rect 33180 13076 33236 13086
rect 33068 13074 33236 13076
rect 33068 13022 33182 13074
rect 33234 13022 33236 13074
rect 33068 13020 33236 13022
rect 33180 13010 33236 13020
rect 33292 12852 33348 16716
rect 33404 15428 33460 19966
rect 33516 19908 33572 19918
rect 33516 19814 33572 19852
rect 33516 19236 33572 19246
rect 33516 17778 33572 19180
rect 33628 19124 33684 20190
rect 34188 20244 34244 21084
rect 35084 20468 35140 21308
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35756 20804 35812 26852
rect 36204 25172 36260 30156
rect 36428 30146 36484 30156
rect 36988 30146 37044 30156
rect 38108 29652 38164 30830
rect 38108 29586 38164 29596
rect 37324 29428 37380 29438
rect 36428 29316 36484 29326
rect 36428 28644 36484 29260
rect 37324 29314 37380 29372
rect 37324 29262 37326 29314
rect 37378 29262 37380 29314
rect 37324 29250 37380 29262
rect 37884 29316 37940 29326
rect 37884 29222 37940 29260
rect 38332 29314 38388 29326
rect 38332 29262 38334 29314
rect 38386 29262 38388 29314
rect 36428 28550 36484 28588
rect 36988 28532 37044 28542
rect 36988 27860 37044 28476
rect 36540 27746 36596 27758
rect 36540 27694 36542 27746
rect 36594 27694 36596 27746
rect 36540 27076 36596 27694
rect 36540 27010 36596 27020
rect 36988 26908 37044 27804
rect 37772 28308 37828 28318
rect 37660 27748 37716 27758
rect 37436 27746 37716 27748
rect 37436 27694 37662 27746
rect 37714 27694 37716 27746
rect 37436 27692 37716 27694
rect 37436 27298 37492 27692
rect 37660 27682 37716 27692
rect 37436 27246 37438 27298
rect 37490 27246 37492 27298
rect 37436 27234 37492 27246
rect 37772 27298 37828 28252
rect 38332 28308 38388 29262
rect 38668 29204 38724 31164
rect 39564 29540 39620 31724
rect 39900 31668 39956 32508
rect 41132 32498 41188 32510
rect 41916 32450 41972 32462
rect 41916 32398 41918 32450
rect 41970 32398 41972 32450
rect 41916 31892 41972 32398
rect 41916 31826 41972 31836
rect 42364 31890 42420 31902
rect 42364 31838 42366 31890
rect 42418 31838 42420 31890
rect 39900 31602 39956 31612
rect 40236 31668 40292 31678
rect 40236 31574 40292 31612
rect 41916 31668 41972 31678
rect 41356 31556 41412 31566
rect 41356 31218 41412 31500
rect 41356 31166 41358 31218
rect 41410 31166 41412 31218
rect 41356 31154 41412 31166
rect 41916 31218 41972 31612
rect 41916 31166 41918 31218
rect 41970 31166 41972 31218
rect 41916 31154 41972 31166
rect 40908 30994 40964 31006
rect 40908 30942 40910 30994
rect 40962 30942 40964 30994
rect 40236 30882 40292 30894
rect 40236 30830 40238 30882
rect 40290 30830 40292 30882
rect 39900 29652 39956 29662
rect 39564 29484 39732 29540
rect 38780 29426 38836 29438
rect 38780 29374 38782 29426
rect 38834 29374 38836 29426
rect 38780 29316 38836 29374
rect 39116 29316 39172 29326
rect 38780 29260 39116 29316
rect 39116 29250 39172 29260
rect 39228 29316 39284 29326
rect 39564 29316 39620 29326
rect 39228 29314 39620 29316
rect 39228 29262 39230 29314
rect 39282 29262 39566 29314
rect 39618 29262 39620 29314
rect 39228 29260 39620 29262
rect 39228 29250 39284 29260
rect 39564 29250 39620 29260
rect 38668 29148 38836 29204
rect 38668 28532 38724 28542
rect 38668 28438 38724 28476
rect 38332 28242 38388 28252
rect 38668 27860 38724 27870
rect 38780 27860 38836 29148
rect 39676 28532 39732 29484
rect 39788 29538 39844 29550
rect 39788 29486 39790 29538
rect 39842 29486 39844 29538
rect 39788 28756 39844 29486
rect 39900 29314 39956 29596
rect 40236 29540 40292 30830
rect 40908 30436 40964 30942
rect 40908 30370 40964 30380
rect 41132 30994 41188 31006
rect 41132 30942 41134 30994
rect 41186 30942 41188 30994
rect 41132 30772 41188 30942
rect 41580 30996 41636 31006
rect 41692 30996 41748 31006
rect 41580 30994 41692 30996
rect 41580 30942 41582 30994
rect 41634 30942 41692 30994
rect 41580 30940 41692 30942
rect 41580 30930 41636 30940
rect 41244 30884 41300 30894
rect 41244 30790 41300 30828
rect 40348 29540 40404 29550
rect 40908 29540 40964 29550
rect 40236 29538 40964 29540
rect 40236 29486 40350 29538
rect 40402 29486 40910 29538
rect 40962 29486 40964 29538
rect 40236 29484 40964 29486
rect 40348 29474 40404 29484
rect 40908 29474 40964 29484
rect 40012 29428 40068 29438
rect 40068 29372 40180 29428
rect 40012 29362 40068 29372
rect 39900 29262 39902 29314
rect 39954 29262 39956 29314
rect 39900 29250 39956 29262
rect 39788 28690 39844 28700
rect 40012 29204 40068 29214
rect 39676 28466 39732 28476
rect 40012 28084 40068 29148
rect 38724 27804 38836 27860
rect 39900 28028 40068 28084
rect 38668 27794 38724 27804
rect 39788 27748 39844 27758
rect 37772 27246 37774 27298
rect 37826 27246 37828 27298
rect 37772 27234 37828 27246
rect 38780 27746 39844 27748
rect 38780 27694 39790 27746
rect 39842 27694 39844 27746
rect 38780 27692 39844 27694
rect 38444 27188 38500 27198
rect 38220 27186 38500 27188
rect 38220 27134 38446 27186
rect 38498 27134 38500 27186
rect 38220 27132 38500 27134
rect 37548 27074 37604 27086
rect 37548 27022 37550 27074
rect 37602 27022 37604 27074
rect 37548 26908 37604 27022
rect 37996 27076 38052 27086
rect 38220 27076 38276 27132
rect 38444 27122 38500 27132
rect 37996 27074 38276 27076
rect 37996 27022 37998 27074
rect 38050 27022 38276 27074
rect 37996 27020 38276 27022
rect 38668 27076 38724 27086
rect 38780 27076 38836 27692
rect 39788 27682 39844 27692
rect 38668 27074 38836 27076
rect 38668 27022 38670 27074
rect 38722 27022 38836 27074
rect 38668 27020 38836 27022
rect 37996 27010 38052 27020
rect 38668 27010 38724 27020
rect 38332 26962 38388 26974
rect 38332 26910 38334 26962
rect 38386 26910 38388 26962
rect 38332 26908 38388 26910
rect 38556 26964 38612 26974
rect 36204 25106 36260 25116
rect 36316 26852 37044 26908
rect 37436 26852 37604 26908
rect 37772 26852 38388 26908
rect 38444 26852 38612 26908
rect 36316 24722 36372 26852
rect 36428 25508 36484 25518
rect 36988 25508 37044 25518
rect 37212 25508 37268 25518
rect 36428 25414 36484 25452
rect 36764 25506 37044 25508
rect 36764 25454 36990 25506
rect 37042 25454 37044 25506
rect 36764 25452 37044 25454
rect 36316 24670 36318 24722
rect 36370 24670 36372 24722
rect 36316 24658 36372 24670
rect 35980 24612 36036 24622
rect 35980 24518 36036 24556
rect 36428 23938 36484 23950
rect 36428 23886 36430 23938
rect 36482 23886 36484 23938
rect 36428 23828 36484 23886
rect 36428 23762 36484 23772
rect 36316 23268 36372 23278
rect 35980 23154 36036 23166
rect 35980 23102 35982 23154
rect 36034 23102 36036 23154
rect 35980 22932 36036 23102
rect 36316 23154 36372 23212
rect 36540 23268 36596 23278
rect 36764 23268 36820 25452
rect 36988 25396 37044 25452
rect 36988 25330 37044 25340
rect 37100 25506 37268 25508
rect 37100 25454 37214 25506
rect 37266 25454 37268 25506
rect 37100 25452 37268 25454
rect 37100 24836 37156 25452
rect 37212 25442 37268 25452
rect 37324 25508 37380 25518
rect 37324 25414 37380 25452
rect 36876 24780 37156 24836
rect 37212 25172 37268 25182
rect 36876 23380 36932 24780
rect 37100 24610 37156 24622
rect 37100 24558 37102 24610
rect 37154 24558 37156 24610
rect 36876 23314 36932 23324
rect 36988 23380 37044 23390
rect 37100 23380 37156 24558
rect 36988 23378 37156 23380
rect 36988 23326 36990 23378
rect 37042 23326 37156 23378
rect 36988 23324 37156 23326
rect 36988 23314 37044 23324
rect 36540 23266 36820 23268
rect 36540 23214 36542 23266
rect 36594 23214 36820 23266
rect 36540 23212 36820 23214
rect 36540 23202 36596 23212
rect 36316 23102 36318 23154
rect 36370 23102 36372 23154
rect 36092 23044 36148 23054
rect 36092 22950 36148 22988
rect 35980 22372 36036 22876
rect 35980 22306 36036 22316
rect 36092 22482 36148 22494
rect 36092 22430 36094 22482
rect 36146 22430 36148 22482
rect 36092 21924 36148 22430
rect 36092 21858 36148 21868
rect 36316 21586 36372 23102
rect 36876 23154 36932 23166
rect 36876 23102 36878 23154
rect 36930 23102 36932 23154
rect 36876 23044 36932 23102
rect 36876 22978 36932 22988
rect 37100 23044 37156 23054
rect 37100 22950 37156 22988
rect 37212 22708 37268 25116
rect 37324 25060 37380 25070
rect 37324 23492 37380 25004
rect 37324 23426 37380 23436
rect 37436 23380 37492 26852
rect 37548 26740 37604 26750
rect 37548 26514 37604 26684
rect 37548 26462 37550 26514
rect 37602 26462 37604 26514
rect 37548 26292 37604 26462
rect 37548 26226 37604 26236
rect 37324 23156 37380 23166
rect 37436 23156 37492 23324
rect 37324 23154 37492 23156
rect 37324 23102 37326 23154
rect 37378 23102 37492 23154
rect 37324 23100 37492 23102
rect 37660 25508 37716 25518
rect 37324 23090 37380 23100
rect 37212 22652 37380 22708
rect 36316 21534 36318 21586
rect 36370 21534 36372 21586
rect 36316 21522 36372 21534
rect 36988 22370 37044 22382
rect 36988 22318 36990 22370
rect 37042 22318 37044 22370
rect 34860 20412 35140 20468
rect 35308 20748 35812 20804
rect 35980 21474 36036 21486
rect 35980 21422 35982 21474
rect 36034 21422 36036 21474
rect 35980 21364 36036 21422
rect 36876 21476 36932 21486
rect 36876 21382 36932 21420
rect 34188 20178 34244 20188
rect 34524 20356 34580 20366
rect 33852 20132 33908 20142
rect 33852 20038 33908 20076
rect 33628 19058 33684 19068
rect 33740 20020 33796 20030
rect 33628 18564 33684 18574
rect 33740 18564 33796 19964
rect 34300 20020 34356 20030
rect 34300 19926 34356 19964
rect 33628 18562 33796 18564
rect 33628 18510 33630 18562
rect 33682 18510 33796 18562
rect 33628 18508 33796 18510
rect 33628 18498 33684 18508
rect 33516 17726 33518 17778
rect 33570 17726 33572 17778
rect 33516 16548 33572 17726
rect 33516 16482 33572 16492
rect 33628 16884 33684 16894
rect 33628 16098 33684 16828
rect 33628 16046 33630 16098
rect 33682 16046 33684 16098
rect 33628 16034 33684 16046
rect 33404 15148 33460 15372
rect 33516 15426 33572 15438
rect 33516 15374 33518 15426
rect 33570 15374 33572 15426
rect 33516 15316 33572 15374
rect 33516 15250 33572 15260
rect 33404 15092 33684 15148
rect 33180 12796 33348 12852
rect 33180 11284 33236 12796
rect 33628 12740 33684 15092
rect 33740 14644 33796 18508
rect 33852 18562 33908 18574
rect 33852 18510 33854 18562
rect 33906 18510 33908 18562
rect 33852 18228 33908 18510
rect 34300 18564 34356 18574
rect 34300 18338 34356 18508
rect 34300 18286 34302 18338
rect 34354 18286 34356 18338
rect 33852 18162 33908 18172
rect 33964 18226 34020 18238
rect 33964 18174 33966 18226
rect 34018 18174 34020 18226
rect 33964 17668 34020 18174
rect 33964 17602 34020 17612
rect 34188 17892 34244 17902
rect 33964 17444 34020 17454
rect 33964 15876 34020 17388
rect 33852 15874 34020 15876
rect 33852 15822 33966 15874
rect 34018 15822 34020 15874
rect 33852 15820 34020 15822
rect 33852 15538 33908 15820
rect 33964 15810 34020 15820
rect 33852 15486 33854 15538
rect 33906 15486 33908 15538
rect 33852 15474 33908 15486
rect 34188 15652 34244 17836
rect 34188 15314 34244 15596
rect 34188 15262 34190 15314
rect 34242 15262 34244 15314
rect 34188 15250 34244 15262
rect 34300 15148 34356 18286
rect 34524 17780 34580 20300
rect 34748 20132 34804 20142
rect 34636 19794 34692 19806
rect 34636 19742 34638 19794
rect 34690 19742 34692 19794
rect 34636 18452 34692 19742
rect 34748 19346 34804 20076
rect 34748 19294 34750 19346
rect 34802 19294 34804 19346
rect 34748 19282 34804 19294
rect 34860 18676 34916 20412
rect 35084 20244 35140 20254
rect 34636 18386 34692 18396
rect 34748 18620 34916 18676
rect 34972 19906 35028 19918
rect 34972 19854 34974 19906
rect 35026 19854 35028 19906
rect 34524 17686 34580 17724
rect 34748 17668 34804 18620
rect 34972 18564 35028 19854
rect 35084 19012 35140 20188
rect 35308 20130 35364 20748
rect 35980 20692 36036 21308
rect 35532 20636 36036 20692
rect 35532 20578 35588 20636
rect 36092 20580 36148 20590
rect 35532 20526 35534 20578
rect 35586 20526 35588 20578
rect 35532 20356 35588 20526
rect 35532 20290 35588 20300
rect 35868 20578 36148 20580
rect 35868 20526 36094 20578
rect 36146 20526 36148 20578
rect 35868 20524 36148 20526
rect 35308 20078 35310 20130
rect 35362 20078 35364 20130
rect 35308 19794 35364 20078
rect 35308 19742 35310 19794
rect 35362 19742 35364 19794
rect 35308 19730 35364 19742
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35868 19460 35924 20524
rect 36092 20514 36148 20524
rect 36540 20244 36596 20254
rect 36428 20188 36540 20244
rect 35308 19404 35924 19460
rect 35980 19906 36036 19918
rect 35980 19854 35982 19906
rect 36034 19854 36036 19906
rect 35196 19012 35252 19022
rect 35084 19010 35252 19012
rect 35084 18958 35198 19010
rect 35250 18958 35252 19010
rect 35084 18956 35252 18958
rect 34972 18498 35028 18508
rect 35084 18676 35140 18686
rect 34860 18452 34916 18462
rect 34860 18358 34916 18396
rect 35084 18228 35140 18620
rect 35196 18450 35252 18956
rect 35196 18398 35198 18450
rect 35250 18398 35252 18450
rect 35196 18386 35252 18398
rect 35308 19010 35364 19404
rect 35420 19236 35476 19246
rect 35420 19142 35476 19180
rect 35308 18958 35310 19010
rect 35362 18958 35364 19010
rect 34972 18172 35140 18228
rect 35308 18228 35364 18958
rect 35532 19124 35588 19134
rect 35532 18676 35588 19068
rect 35756 19124 35812 19134
rect 35756 19030 35812 19068
rect 35644 18676 35700 18686
rect 35532 18674 35700 18676
rect 35532 18622 35646 18674
rect 35698 18622 35700 18674
rect 35532 18620 35700 18622
rect 35644 18610 35700 18620
rect 35420 18564 35476 18574
rect 35420 18470 35476 18508
rect 35868 18564 35924 18574
rect 35868 18470 35924 18508
rect 35532 18450 35588 18462
rect 35532 18398 35534 18450
rect 35586 18398 35588 18450
rect 35532 18340 35588 18398
rect 35980 18340 36036 19854
rect 36092 19908 36148 19918
rect 36092 19814 36148 19852
rect 36092 19236 36148 19246
rect 36148 19180 36260 19236
rect 36092 19170 36148 19180
rect 36204 19122 36260 19180
rect 36204 19070 36206 19122
rect 36258 19070 36260 19122
rect 36204 19058 36260 19070
rect 35532 18284 36036 18340
rect 36316 19010 36372 19022
rect 36316 18958 36318 19010
rect 36370 18958 36372 19010
rect 36316 18340 36372 18958
rect 36316 18274 36372 18284
rect 36428 18562 36484 20188
rect 36540 20178 36596 20188
rect 36540 20020 36596 20030
rect 36988 20020 37044 22318
rect 37212 21476 37268 21486
rect 37212 21382 37268 21420
rect 37212 20578 37268 20590
rect 37212 20526 37214 20578
rect 37266 20526 37268 20578
rect 37212 20244 37268 20526
rect 37212 20178 37268 20188
rect 36540 20018 37156 20020
rect 36540 19966 36542 20018
rect 36594 19966 37156 20018
rect 36540 19964 37156 19966
rect 36540 19954 36596 19964
rect 36540 18676 36596 18686
rect 36540 18674 36932 18676
rect 36540 18622 36542 18674
rect 36594 18622 36932 18674
rect 36540 18620 36932 18622
rect 36540 18610 36596 18620
rect 36428 18510 36430 18562
rect 36482 18510 36484 18562
rect 35308 18172 35588 18228
rect 34860 17668 34916 17678
rect 34748 17666 34916 17668
rect 34748 17614 34862 17666
rect 34914 17614 34916 17666
rect 34748 17612 34916 17614
rect 34524 17556 34580 17566
rect 34524 15986 34580 17500
rect 34860 17332 34916 17612
rect 34860 17266 34916 17276
rect 34972 16322 35028 18172
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35420 17668 35476 17678
rect 35532 17668 35588 18172
rect 35420 17666 35588 17668
rect 35420 17614 35422 17666
rect 35474 17614 35588 17666
rect 35420 17612 35588 17614
rect 35644 17780 35700 17790
rect 35420 17556 35476 17612
rect 35420 17490 35476 17500
rect 34972 16270 34974 16322
rect 35026 16270 35028 16322
rect 34972 16210 35028 16270
rect 35084 16884 35140 16894
rect 35084 16770 35140 16828
rect 35084 16718 35086 16770
rect 35138 16718 35140 16770
rect 35084 16324 35140 16718
rect 35644 16884 35700 17724
rect 36428 17556 36484 18510
rect 36764 18450 36820 18462
rect 36764 18398 36766 18450
rect 36818 18398 36820 18450
rect 36428 17554 36708 17556
rect 36428 17502 36430 17554
rect 36482 17502 36708 17554
rect 36428 17500 36708 17502
rect 36428 17490 36484 17500
rect 36092 17444 36148 17454
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35308 16324 35364 16334
rect 35084 16268 35252 16324
rect 34972 16158 34974 16210
rect 35026 16158 35028 16210
rect 34972 16146 35028 16158
rect 34524 15934 34526 15986
rect 34578 15934 34580 15986
rect 34524 15876 34580 15934
rect 34524 15810 34580 15820
rect 35084 15426 35140 15438
rect 35084 15374 35086 15426
rect 35138 15374 35140 15426
rect 34748 15314 34804 15326
rect 34748 15262 34750 15314
rect 34802 15262 34804 15314
rect 34748 15204 34804 15262
rect 35084 15148 35140 15374
rect 34300 15092 34468 15148
rect 34748 15138 34804 15148
rect 33740 14578 33796 14588
rect 34300 13634 34356 13646
rect 34300 13582 34302 13634
rect 34354 13582 34356 13634
rect 34188 13522 34244 13534
rect 34188 13470 34190 13522
rect 34242 13470 34244 13522
rect 33628 12674 33684 12684
rect 33852 12962 33908 12974
rect 33852 12910 33854 12962
rect 33906 12910 33908 12962
rect 33292 12180 33348 12190
rect 33852 12180 33908 12910
rect 34188 12852 34244 13470
rect 34300 13076 34356 13582
rect 34412 13300 34468 15092
rect 34860 15092 35140 15148
rect 35196 15148 35252 16268
rect 35308 16322 35476 16324
rect 35308 16270 35310 16322
rect 35362 16270 35476 16322
rect 35308 16268 35476 16270
rect 35308 16258 35364 16268
rect 35420 16098 35476 16268
rect 35420 16046 35422 16098
rect 35474 16046 35476 16098
rect 35420 16034 35476 16046
rect 35644 16098 35700 16828
rect 35644 16046 35646 16098
rect 35698 16046 35700 16098
rect 35644 16034 35700 16046
rect 35868 17442 36148 17444
rect 35868 17390 36094 17442
rect 36146 17390 36148 17442
rect 35868 17388 36148 17390
rect 35868 16210 35924 17388
rect 36092 17378 36148 17388
rect 35868 16158 35870 16210
rect 35922 16158 35924 16210
rect 35420 15764 35476 15774
rect 35420 15538 35476 15708
rect 35420 15486 35422 15538
rect 35474 15486 35476 15538
rect 35420 15474 35476 15486
rect 35756 15540 35812 15550
rect 35196 15092 35588 15148
rect 34748 14644 34804 14654
rect 34748 14550 34804 14588
rect 34860 13412 34916 15092
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35308 14644 35364 14654
rect 35308 14530 35364 14588
rect 35308 14478 35310 14530
rect 35362 14478 35364 14530
rect 35308 14466 35364 14478
rect 34748 13356 34916 13412
rect 35084 14306 35140 14318
rect 35084 14254 35086 14306
rect 35138 14254 35140 14306
rect 34468 13244 34692 13300
rect 34412 13234 34468 13244
rect 34412 13076 34468 13086
rect 34300 13074 34468 13076
rect 34300 13022 34414 13074
rect 34466 13022 34468 13074
rect 34300 13020 34468 13022
rect 34412 13010 34468 13020
rect 34188 12786 34244 12796
rect 33292 12178 33908 12180
rect 33292 12126 33294 12178
rect 33346 12126 33908 12178
rect 33292 12124 33908 12126
rect 33964 12740 34020 12750
rect 33292 11844 33348 12124
rect 33292 11778 33348 11788
rect 33964 11620 34020 12684
rect 34412 12738 34468 12750
rect 34412 12686 34414 12738
rect 34466 12686 34468 12738
rect 34412 12628 34468 12686
rect 34524 12740 34580 12778
rect 34524 12674 34580 12684
rect 34300 12516 34356 12526
rect 34188 12292 34244 12302
rect 34076 12180 34132 12190
rect 34188 12180 34244 12236
rect 34076 12178 34244 12180
rect 34076 12126 34078 12178
rect 34130 12126 34244 12178
rect 34076 12124 34244 12126
rect 34076 12114 34132 12124
rect 33964 11564 34132 11620
rect 33852 11508 33908 11518
rect 33740 11452 33852 11508
rect 33180 11228 33572 11284
rect 33404 11060 33460 11070
rect 32284 10836 32340 10846
rect 32620 10836 32676 10846
rect 32284 10164 32340 10780
rect 32508 10780 32620 10836
rect 32508 10722 32564 10780
rect 32620 10770 32676 10780
rect 33404 10834 33460 11004
rect 33404 10782 33406 10834
rect 33458 10782 33460 10834
rect 33404 10770 33460 10782
rect 32508 10670 32510 10722
rect 32562 10670 32564 10722
rect 32508 10658 32564 10670
rect 33516 10610 33572 11228
rect 33628 10836 33684 10846
rect 33628 10742 33684 10780
rect 33740 10834 33796 11452
rect 33852 11442 33908 11452
rect 33740 10782 33742 10834
rect 33794 10782 33796 10834
rect 33740 10770 33796 10782
rect 33964 11396 34020 11406
rect 33964 10724 34020 11340
rect 33516 10558 33518 10610
rect 33570 10558 33572 10610
rect 32396 10388 32452 10398
rect 32396 10294 32452 10332
rect 32284 9828 32340 10108
rect 32284 9772 32564 9828
rect 32508 9268 32564 9772
rect 33516 9716 33572 10558
rect 33852 10722 34020 10724
rect 33852 10670 33966 10722
rect 34018 10670 34020 10722
rect 33852 10668 34020 10670
rect 33852 10388 33908 10668
rect 33964 10658 34020 10668
rect 33628 10332 33908 10388
rect 33628 9938 33684 10332
rect 33628 9886 33630 9938
rect 33682 9886 33684 9938
rect 33628 9874 33684 9886
rect 33516 9660 33684 9716
rect 32508 9174 32564 9212
rect 33516 9268 33572 9278
rect 32172 8978 32228 8988
rect 33292 9044 33348 9054
rect 31500 8258 31556 8270
rect 31500 8206 31502 8258
rect 31554 8206 31556 8258
rect 31500 7476 31556 8206
rect 32172 8148 32228 8158
rect 32172 8146 32452 8148
rect 32172 8094 32174 8146
rect 32226 8094 32452 8146
rect 32172 8092 32452 8094
rect 32172 8082 32228 8092
rect 32396 7698 32452 8092
rect 32396 7646 32398 7698
rect 32450 7646 32452 7698
rect 32396 7634 32452 7646
rect 32508 8036 32564 8046
rect 32508 7586 32564 7980
rect 32508 7534 32510 7586
rect 32562 7534 32564 7586
rect 32508 7522 32564 7534
rect 32732 7924 32788 7934
rect 31948 7476 32004 7486
rect 31500 7420 31948 7476
rect 31500 5122 31556 7420
rect 31948 7382 32004 7420
rect 32508 6804 32564 6814
rect 32172 6692 32228 6702
rect 32172 6598 32228 6636
rect 31612 6466 31668 6478
rect 31612 6414 31614 6466
rect 31666 6414 31668 6466
rect 31612 6356 31668 6414
rect 31612 6290 31668 6300
rect 32508 6466 32564 6748
rect 32508 6414 32510 6466
rect 32562 6414 32564 6466
rect 32284 5908 32340 5918
rect 32508 5908 32564 6414
rect 32732 6356 32788 7868
rect 33292 7474 33348 8988
rect 33516 9042 33572 9212
rect 33516 8990 33518 9042
rect 33570 8990 33572 9042
rect 33516 8978 33572 8990
rect 33628 7924 33684 9660
rect 34076 9156 34132 11564
rect 34300 10724 34356 12460
rect 34412 11060 34468 12572
rect 34412 10994 34468 11004
rect 33628 7858 33684 7868
rect 33740 9100 34132 9156
rect 34188 10668 34356 10724
rect 33516 7588 33572 7598
rect 33628 7588 33684 7598
rect 33516 7586 33628 7588
rect 33516 7534 33518 7586
rect 33570 7534 33628 7586
rect 33516 7532 33628 7534
rect 33516 7522 33572 7532
rect 33292 7422 33294 7474
rect 33346 7422 33348 7474
rect 33292 7410 33348 7422
rect 32956 6916 33012 6926
rect 32956 6578 33012 6860
rect 33292 6692 33348 6702
rect 33292 6598 33348 6636
rect 32956 6526 32958 6578
rect 33010 6526 33012 6578
rect 32956 6514 33012 6526
rect 32732 6290 32788 6300
rect 32284 5906 32564 5908
rect 32284 5854 32286 5906
rect 32338 5854 32564 5906
rect 32284 5852 32564 5854
rect 33404 6020 33460 6030
rect 32284 5842 32340 5852
rect 33180 5796 33236 5806
rect 33180 5702 33236 5740
rect 33068 5684 33124 5694
rect 32172 5682 33124 5684
rect 32172 5630 33070 5682
rect 33122 5630 33124 5682
rect 32172 5628 33124 5630
rect 32172 5234 32228 5628
rect 33068 5618 33124 5628
rect 32172 5182 32174 5234
rect 32226 5182 32228 5234
rect 32172 5170 32228 5182
rect 31500 5070 31502 5122
rect 31554 5070 31556 5122
rect 31500 5058 31556 5070
rect 32956 4900 33012 4910
rect 32284 4340 32340 4350
rect 32172 4226 32228 4238
rect 32172 4174 32174 4226
rect 32226 4174 32228 4226
rect 31836 3668 31892 3678
rect 31500 3444 31556 3454
rect 31388 3388 31500 3444
rect 31500 3378 31556 3388
rect 31836 800 31892 3612
rect 32172 3556 32228 4174
rect 32172 3490 32228 3500
rect 32284 3554 32340 4284
rect 32956 3666 33012 4844
rect 33292 4564 33348 4574
rect 33292 4470 33348 4508
rect 32956 3614 32958 3666
rect 33010 3614 33012 3666
rect 32956 3602 33012 3614
rect 32284 3502 32286 3554
rect 32338 3502 32340 3554
rect 32284 3490 32340 3502
rect 33404 800 33460 5964
rect 33628 5906 33684 7532
rect 33740 6916 33796 9100
rect 33740 6130 33796 6860
rect 34076 8932 34132 8942
rect 33740 6078 33742 6130
rect 33794 6078 33796 6130
rect 33740 6066 33796 6078
rect 33852 6802 33908 6814
rect 33852 6750 33854 6802
rect 33906 6750 33908 6802
rect 33852 6020 33908 6750
rect 33852 5954 33908 5964
rect 33964 6132 34020 6142
rect 34076 6132 34132 8876
rect 34188 6916 34244 10668
rect 34300 10500 34356 10510
rect 34300 10406 34356 10444
rect 34636 9940 34692 13244
rect 34748 12962 34804 13356
rect 34972 13300 35028 13310
rect 34748 12910 34750 12962
rect 34802 12910 34804 12962
rect 34748 11508 34804 12910
rect 34748 11442 34804 11452
rect 34860 13244 34972 13300
rect 34860 10724 34916 13244
rect 34972 13234 35028 13244
rect 34972 12852 35028 12862
rect 34972 12758 35028 12796
rect 35084 12628 35140 14254
rect 35532 13746 35588 15092
rect 35756 14644 35812 15484
rect 35868 15314 35924 16158
rect 36428 17332 36484 17342
rect 36428 16210 36484 17276
rect 36428 16158 36430 16210
rect 36482 16158 36484 16210
rect 36428 16100 36484 16158
rect 36428 16034 36484 16044
rect 36540 16884 36596 16894
rect 35868 15262 35870 15314
rect 35922 15262 35924 15314
rect 35868 15250 35924 15262
rect 35980 15986 36036 15998
rect 35980 15934 35982 15986
rect 36034 15934 36036 15986
rect 35980 15148 36036 15934
rect 36540 15538 36596 16828
rect 36540 15486 36542 15538
rect 36594 15486 36596 15538
rect 36540 15474 36596 15486
rect 36092 15428 36148 15438
rect 36092 15334 36148 15372
rect 36428 15316 36484 15326
rect 35980 15092 36260 15148
rect 35756 14578 35812 14588
rect 35868 14532 35924 14542
rect 35868 14438 35924 14476
rect 35980 14420 36036 14430
rect 35980 14326 36036 14364
rect 36092 14308 36148 14318
rect 36092 14214 36148 14252
rect 35532 13694 35534 13746
rect 35586 13694 35588 13746
rect 35532 13682 35588 13694
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 36204 13076 36260 15092
rect 36316 13860 36372 13870
rect 36428 13860 36484 15260
rect 36316 13858 36484 13860
rect 36316 13806 36318 13858
rect 36370 13806 36484 13858
rect 36316 13804 36484 13806
rect 36540 14530 36596 14542
rect 36540 14478 36542 14530
rect 36594 14478 36596 14530
rect 36316 13794 36372 13804
rect 36540 13188 36596 14478
rect 36652 14084 36708 17500
rect 36764 16212 36820 18398
rect 36876 16884 36932 18620
rect 37100 18452 37156 19964
rect 37212 19908 37268 19918
rect 37212 19814 37268 19852
rect 36876 16828 37044 16884
rect 36764 16146 36820 16156
rect 36652 14018 36708 14028
rect 36876 16100 36932 16110
rect 36540 13122 36596 13132
rect 36204 13020 36372 13076
rect 35084 12562 35140 12572
rect 36204 12852 36260 12862
rect 36204 12068 36260 12796
rect 36204 11974 36260 12012
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 34636 9874 34692 9884
rect 34748 10668 34916 10724
rect 34972 11508 35028 11518
rect 34412 9604 34468 9614
rect 34748 9604 34804 10668
rect 34860 10500 34916 10510
rect 34860 9826 34916 10444
rect 34860 9774 34862 9826
rect 34914 9774 34916 9826
rect 34860 9762 34916 9774
rect 34972 9828 35028 11452
rect 35196 11172 35252 11182
rect 35084 11116 35196 11172
rect 35084 9938 35140 11116
rect 35196 11106 35252 11116
rect 35532 11060 35588 11070
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35532 10052 35588 11004
rect 35756 10612 35812 10622
rect 35084 9886 35086 9938
rect 35138 9886 35140 9938
rect 35084 9874 35140 9886
rect 35420 9996 35588 10052
rect 35644 10556 35756 10612
rect 34972 9734 35028 9772
rect 35420 9826 35476 9996
rect 35420 9774 35422 9826
rect 35474 9774 35476 9826
rect 35420 9716 35476 9774
rect 35420 9650 35476 9660
rect 35196 9604 35252 9614
rect 34748 9548 35196 9604
rect 34412 9510 34468 9548
rect 35196 9510 35252 9548
rect 35196 9268 35252 9278
rect 35196 9154 35252 9212
rect 35196 9102 35198 9154
rect 35250 9102 35252 9154
rect 35196 9090 35252 9102
rect 35308 9156 35364 9166
rect 35308 9062 35364 9100
rect 35644 9044 35700 10556
rect 35756 10546 35812 10556
rect 35980 9940 36036 9950
rect 35756 9826 35812 9838
rect 35756 9774 35758 9826
rect 35810 9774 35812 9826
rect 35756 9716 35812 9774
rect 35980 9826 36036 9884
rect 35980 9774 35982 9826
rect 36034 9774 36036 9826
rect 35980 9762 36036 9774
rect 36204 9828 36260 9838
rect 36204 9734 36260 9772
rect 35756 9650 35812 9660
rect 35868 9604 35924 9614
rect 35924 9548 36036 9604
rect 35868 9538 35924 9548
rect 35532 9042 35700 9044
rect 35532 8990 35646 9042
rect 35698 8990 35700 9042
rect 35532 8988 35700 8990
rect 34748 8932 34804 8942
rect 34524 8930 34804 8932
rect 34524 8878 34750 8930
rect 34802 8878 34804 8930
rect 34524 8876 34804 8878
rect 34300 8372 34356 8382
rect 34300 8278 34356 8316
rect 34188 6692 34244 6860
rect 34188 6626 34244 6636
rect 34524 6468 34580 8876
rect 34748 8866 34804 8876
rect 34972 8932 35028 8942
rect 35028 8876 35140 8932
rect 34972 8866 35028 8876
rect 34860 8818 34916 8830
rect 34860 8766 34862 8818
rect 34914 8766 34916 8818
rect 34860 8260 34916 8766
rect 34636 8204 34916 8260
rect 35084 8258 35140 8876
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35084 8206 35086 8258
rect 35138 8206 35140 8258
rect 34636 6580 34692 8204
rect 34748 8034 34804 8046
rect 34748 7982 34750 8034
rect 34802 7982 34804 8034
rect 34748 7588 34804 7982
rect 34860 8034 34916 8046
rect 34860 7982 34862 8034
rect 34914 7982 34916 8034
rect 34860 7924 34916 7982
rect 34972 8036 35028 8046
rect 34972 7942 35028 7980
rect 34860 7858 34916 7868
rect 34748 7522 34804 7532
rect 34636 6514 34692 6524
rect 34524 6402 34580 6412
rect 33964 6130 34132 6132
rect 33964 6078 33966 6130
rect 34018 6078 34132 6130
rect 33964 6076 34132 6078
rect 33628 5854 33630 5906
rect 33682 5854 33684 5906
rect 33516 5236 33572 5246
rect 33516 4450 33572 5180
rect 33628 5124 33684 5854
rect 33852 5796 33908 5806
rect 33852 5702 33908 5740
rect 33628 5058 33684 5068
rect 33964 4788 34020 6076
rect 34972 6020 35028 6030
rect 34972 5926 35028 5964
rect 34188 5908 34244 5918
rect 34860 5908 34916 5918
rect 34244 5852 34356 5908
rect 34188 5814 34244 5852
rect 34300 5234 34356 5852
rect 34860 5814 34916 5852
rect 34300 5182 34302 5234
rect 34354 5182 34356 5234
rect 34300 5170 34356 5182
rect 34748 5236 34804 5246
rect 34748 5142 34804 5180
rect 34636 5124 34692 5134
rect 34636 5030 34692 5068
rect 35084 5122 35140 8206
rect 35196 8372 35252 8382
rect 35196 8258 35252 8316
rect 35196 8206 35198 8258
rect 35250 8206 35252 8258
rect 35196 8194 35252 8206
rect 35532 7586 35588 8988
rect 35644 8978 35700 8988
rect 35644 8372 35700 8382
rect 35644 8278 35700 8316
rect 35756 8034 35812 8046
rect 35756 7982 35758 8034
rect 35810 7982 35812 8034
rect 35756 7700 35812 7982
rect 35756 7634 35812 7644
rect 35532 7534 35534 7586
rect 35586 7534 35588 7586
rect 35532 7476 35588 7534
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35532 6692 35588 7420
rect 35420 5908 35476 5918
rect 35532 5908 35588 6636
rect 35420 5906 35588 5908
rect 35420 5854 35422 5906
rect 35474 5854 35588 5906
rect 35420 5852 35588 5854
rect 35420 5842 35476 5852
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35420 5348 35476 5358
rect 35308 5236 35364 5246
rect 35084 5070 35086 5122
rect 35138 5070 35140 5122
rect 35084 5058 35140 5070
rect 35196 5180 35308 5236
rect 33964 4722 34020 4732
rect 34076 5012 34132 5022
rect 33516 4398 33518 4450
rect 33570 4398 33572 4450
rect 33516 4386 33572 4398
rect 34076 4340 34132 4956
rect 34860 4898 34916 4910
rect 34860 4846 34862 4898
rect 34914 4846 34916 4898
rect 34860 4564 34916 4846
rect 34860 4498 34916 4508
rect 34972 4900 35028 4910
rect 35196 4900 35252 5180
rect 35308 5170 35364 5180
rect 35308 5012 35364 5022
rect 35420 5012 35476 5292
rect 35308 5010 35476 5012
rect 35308 4958 35310 5010
rect 35362 4958 35476 5010
rect 35308 4956 35476 4958
rect 35532 5012 35588 5852
rect 35756 6690 35812 6702
rect 35756 6638 35758 6690
rect 35810 6638 35812 6690
rect 35756 5236 35812 6638
rect 35756 5170 35812 5180
rect 35868 6468 35924 6478
rect 35868 5234 35924 6412
rect 35868 5182 35870 5234
rect 35922 5182 35924 5234
rect 35868 5170 35924 5182
rect 35644 5124 35700 5134
rect 35644 5030 35700 5068
rect 35308 4946 35364 4956
rect 35532 4946 35588 4956
rect 35868 5012 35924 5022
rect 35980 5012 36036 9548
rect 36092 9602 36148 9614
rect 36092 9550 36094 9602
rect 36146 9550 36148 9602
rect 36092 9268 36148 9550
rect 36316 9604 36372 13020
rect 36876 12852 36932 16044
rect 36988 15426 37044 16828
rect 37100 16098 37156 18396
rect 37324 19234 37380 22652
rect 37548 22036 37604 22046
rect 37436 21812 37492 21822
rect 37436 21586 37492 21756
rect 37436 21534 37438 21586
rect 37490 21534 37492 21586
rect 37436 21522 37492 21534
rect 37324 19182 37326 19234
rect 37378 19182 37380 19234
rect 37212 17780 37268 17790
rect 37324 17780 37380 19182
rect 37212 17778 37380 17780
rect 37212 17726 37214 17778
rect 37266 17726 37380 17778
rect 37212 17724 37380 17726
rect 37212 17714 37268 17724
rect 37100 16046 37102 16098
rect 37154 16046 37156 16098
rect 37100 16034 37156 16046
rect 37436 17108 37492 17118
rect 36988 15374 36990 15426
rect 37042 15374 37044 15426
rect 36988 15362 37044 15374
rect 37100 15652 37156 15662
rect 37100 15204 37156 15596
rect 36876 12786 36932 12796
rect 36988 15148 37156 15204
rect 37212 15428 37268 15438
rect 36988 12404 37044 15148
rect 37212 14756 37268 15372
rect 37100 14700 37268 14756
rect 37436 15314 37492 17052
rect 37436 15262 37438 15314
rect 37490 15262 37492 15314
rect 37100 14418 37156 14700
rect 37212 14532 37268 14542
rect 37212 14438 37268 14476
rect 37100 14366 37102 14418
rect 37154 14366 37156 14418
rect 37100 13524 37156 14366
rect 37324 14420 37380 14430
rect 37324 14326 37380 14364
rect 37436 14308 37492 15262
rect 37436 13636 37492 14252
rect 37436 13570 37492 13580
rect 37100 13458 37156 13468
rect 37324 13188 37380 13198
rect 36988 12348 37268 12404
rect 37100 12180 37156 12190
rect 36652 12066 36708 12078
rect 36652 12014 36654 12066
rect 36706 12014 36708 12066
rect 36540 11954 36596 11966
rect 36540 11902 36542 11954
rect 36594 11902 36596 11954
rect 36428 11394 36484 11406
rect 36428 11342 36430 11394
rect 36482 11342 36484 11394
rect 36428 10836 36484 11342
rect 36428 10770 36484 10780
rect 36428 10612 36484 10622
rect 36540 10612 36596 11902
rect 36652 11172 36708 12014
rect 36988 12068 37044 12078
rect 36988 11394 37044 12012
rect 36988 11342 36990 11394
rect 37042 11342 37044 11394
rect 36988 11330 37044 11342
rect 37100 11508 37156 12124
rect 37100 11282 37156 11452
rect 37100 11230 37102 11282
rect 37154 11230 37156 11282
rect 37100 11218 37156 11230
rect 36652 11106 36708 11116
rect 36428 10610 36596 10612
rect 36428 10558 36430 10610
rect 36482 10558 36596 10610
rect 36428 10556 36596 10558
rect 36652 10724 36708 10734
rect 36428 10546 36484 10556
rect 36428 9828 36484 9838
rect 36428 9734 36484 9772
rect 36316 9548 36596 9604
rect 36092 9202 36148 9212
rect 36204 9156 36260 9166
rect 36428 9156 36484 9166
rect 36260 9154 36484 9156
rect 36260 9102 36430 9154
rect 36482 9102 36484 9154
rect 36260 9100 36484 9102
rect 36204 9090 36260 9100
rect 36428 9090 36484 9100
rect 36540 8484 36596 9548
rect 36428 8260 36484 8270
rect 36540 8260 36596 8428
rect 36428 8258 36596 8260
rect 36428 8206 36430 8258
rect 36482 8206 36596 8258
rect 36428 8204 36596 8206
rect 36652 8372 36708 10668
rect 37100 10612 37156 10622
rect 37100 10518 37156 10556
rect 37212 10052 37268 12348
rect 37324 12180 37380 13132
rect 37548 12292 37604 21980
rect 37660 15876 37716 25452
rect 37772 25282 37828 26852
rect 38444 26514 38500 26852
rect 38444 26462 38446 26514
rect 38498 26462 38500 26514
rect 38444 26450 38500 26462
rect 38332 26292 38388 26302
rect 38780 26292 38836 27020
rect 39228 27074 39284 27086
rect 39228 27022 39230 27074
rect 39282 27022 39284 27074
rect 39228 26964 39284 27022
rect 39340 27076 39396 27086
rect 39340 26982 39396 27020
rect 39564 27076 39620 27086
rect 39900 27076 39956 28028
rect 40124 27972 40180 29372
rect 40236 29316 40292 29326
rect 40236 29222 40292 29260
rect 40348 28420 40404 28430
rect 40348 28082 40404 28364
rect 41132 28196 41188 30716
rect 41244 29540 41300 29550
rect 41300 29484 41412 29540
rect 41244 29446 41300 29484
rect 40348 28030 40350 28082
rect 40402 28030 40404 28082
rect 40348 28018 40404 28030
rect 40908 28140 41188 28196
rect 41244 28420 41300 28430
rect 40236 27972 40292 27982
rect 39564 27074 39956 27076
rect 39564 27022 39566 27074
rect 39618 27022 39956 27074
rect 39564 27020 39956 27022
rect 40012 27970 40292 27972
rect 40012 27918 40238 27970
rect 40290 27918 40292 27970
rect 40012 27916 40292 27918
rect 39564 27010 39620 27020
rect 40012 26908 40068 27916
rect 40236 27906 40292 27916
rect 40684 27188 40740 27198
rect 40460 27186 40740 27188
rect 40460 27134 40686 27186
rect 40738 27134 40740 27186
rect 40460 27132 40740 27134
rect 40348 27076 40404 27114
rect 40348 27010 40404 27020
rect 39228 26898 39284 26908
rect 39452 26850 39508 26862
rect 39452 26798 39454 26850
rect 39506 26798 39508 26850
rect 39452 26516 39508 26798
rect 39676 26852 40068 26908
rect 40124 26964 40180 27002
rect 40460 26908 40516 27132
rect 40684 27122 40740 27132
rect 40908 26964 40964 28140
rect 41244 28082 41300 28364
rect 41244 28030 41246 28082
rect 41298 28030 41300 28082
rect 41244 28018 41300 28030
rect 40124 26898 40180 26908
rect 40236 26852 40516 26908
rect 40572 26908 40964 26964
rect 41020 27860 41076 27870
rect 41020 26962 41076 27804
rect 41132 27860 41188 27870
rect 41356 27860 41412 29484
rect 41692 29314 41748 30940
rect 42364 30996 42420 31838
rect 42476 31780 42532 33966
rect 42476 31714 42532 31724
rect 42924 33684 42980 33694
rect 43708 33684 43764 34636
rect 44044 34468 44100 34478
rect 43932 34132 43988 34142
rect 43708 33628 43876 33684
rect 42924 31668 42980 33628
rect 43708 33460 43764 33470
rect 43708 32564 43764 33404
rect 43708 32498 43764 32508
rect 43372 32002 43428 32014
rect 43372 31950 43374 32002
rect 43426 31950 43428 32002
rect 43036 31892 43092 31902
rect 43036 31798 43092 31836
rect 42924 31220 42980 31612
rect 43148 31666 43204 31678
rect 43148 31614 43150 31666
rect 43202 31614 43204 31666
rect 43036 31220 43092 31230
rect 42924 31218 43092 31220
rect 42924 31166 43038 31218
rect 43090 31166 43092 31218
rect 42924 31164 43092 31166
rect 43036 31154 43092 31164
rect 43148 31218 43204 31614
rect 43148 31166 43150 31218
rect 43202 31166 43204 31218
rect 43148 31154 43204 31166
rect 43260 31556 43316 31566
rect 43260 31218 43316 31500
rect 43260 31166 43262 31218
rect 43314 31166 43316 31218
rect 43260 31108 43316 31166
rect 43260 31042 43316 31052
rect 42364 30930 42420 30940
rect 42812 30996 42868 31006
rect 42028 30884 42084 30894
rect 42028 30790 42084 30828
rect 42476 30882 42532 30894
rect 42476 30830 42478 30882
rect 42530 30830 42532 30882
rect 42476 30772 42532 30830
rect 42476 30706 42532 30716
rect 42812 30436 42868 30940
rect 42812 30370 42868 30380
rect 43372 30994 43428 31950
rect 43708 31892 43764 31902
rect 43372 30942 43374 30994
rect 43426 30942 43428 30994
rect 42364 30324 42420 30334
rect 41692 29262 41694 29314
rect 41746 29262 41748 29314
rect 41580 29202 41636 29214
rect 41580 29150 41582 29202
rect 41634 29150 41636 29202
rect 41468 28084 41524 28094
rect 41468 27990 41524 28028
rect 41580 28082 41636 29150
rect 41692 28420 41748 29262
rect 41804 30212 41860 30222
rect 41804 30098 41860 30156
rect 41804 30046 41806 30098
rect 41858 30046 41860 30098
rect 41804 28642 41860 30046
rect 41804 28590 41806 28642
rect 41858 28590 41860 28642
rect 41804 28578 41860 28590
rect 41692 28364 42308 28420
rect 41580 28030 41582 28082
rect 41634 28030 41636 28082
rect 41580 28018 41636 28030
rect 42140 28084 42196 28094
rect 42140 27990 42196 28028
rect 41132 27858 41412 27860
rect 41132 27806 41134 27858
rect 41186 27806 41412 27858
rect 41132 27804 41412 27806
rect 41132 27794 41188 27804
rect 41580 27746 41636 27758
rect 41580 27694 41582 27746
rect 41634 27694 41636 27746
rect 41356 27076 41412 27086
rect 41356 26982 41412 27020
rect 41020 26910 41022 26962
rect 41074 26910 41076 26962
rect 39676 26850 39732 26852
rect 39676 26798 39678 26850
rect 39730 26798 39732 26850
rect 39676 26786 39732 26798
rect 40124 26740 40180 26750
rect 39452 26450 39508 26460
rect 39788 26684 40124 26740
rect 39788 26514 39844 26684
rect 40124 26674 40180 26684
rect 39788 26462 39790 26514
rect 39842 26462 39844 26514
rect 39788 26450 39844 26462
rect 39228 26402 39284 26414
rect 39228 26350 39230 26402
rect 39282 26350 39284 26402
rect 38332 26290 38836 26292
rect 38332 26238 38334 26290
rect 38386 26238 38782 26290
rect 38834 26238 38836 26290
rect 38332 26236 38836 26238
rect 38332 26226 38388 26236
rect 38780 26198 38836 26236
rect 38892 26292 38948 26302
rect 37772 25230 37774 25282
rect 37826 25230 37828 25282
rect 37772 23044 37828 25230
rect 37884 26178 37940 26190
rect 37884 26126 37886 26178
rect 37938 26126 37940 26178
rect 37884 24612 37940 26126
rect 37996 26066 38052 26078
rect 37996 26014 37998 26066
rect 38050 26014 38052 26066
rect 37996 25732 38052 26014
rect 37996 25666 38052 25676
rect 38780 25732 38836 25742
rect 38780 25638 38836 25676
rect 38108 25396 38164 25406
rect 38108 25302 38164 25340
rect 38444 25394 38500 25406
rect 38444 25342 38446 25394
rect 38498 25342 38500 25394
rect 38332 24724 38388 24734
rect 37940 24556 38052 24612
rect 37884 24546 37940 24556
rect 37996 24050 38052 24556
rect 37996 23998 37998 24050
rect 38050 23998 38052 24050
rect 37996 23986 38052 23998
rect 38332 24050 38388 24668
rect 38332 23998 38334 24050
rect 38386 23998 38388 24050
rect 38332 23986 38388 23998
rect 37884 23940 37940 23950
rect 37884 23846 37940 23884
rect 38444 23940 38500 25342
rect 38444 23874 38500 23884
rect 38668 23716 38724 23726
rect 38780 23716 38836 23726
rect 38724 23714 38836 23716
rect 38724 23662 38782 23714
rect 38834 23662 38836 23714
rect 38724 23660 38836 23662
rect 38892 23716 38948 26236
rect 39004 26290 39060 26302
rect 39004 26238 39006 26290
rect 39058 26238 39060 26290
rect 39004 25396 39060 26238
rect 39228 25844 39284 26350
rect 39340 26292 39396 26302
rect 39340 26198 39396 26236
rect 39228 25788 39956 25844
rect 39116 25620 39172 25630
rect 39116 25618 39284 25620
rect 39116 25566 39118 25618
rect 39170 25566 39284 25618
rect 39116 25564 39284 25566
rect 39116 25554 39172 25564
rect 39228 25508 39284 25564
rect 39564 25564 39844 25620
rect 39564 25508 39620 25564
rect 39228 25452 39620 25508
rect 39788 25506 39844 25564
rect 39788 25454 39790 25506
rect 39842 25454 39844 25506
rect 39788 25442 39844 25454
rect 39004 25302 39060 25340
rect 39676 25396 39732 25406
rect 39676 25302 39732 25340
rect 39452 25284 39508 25294
rect 39452 24722 39508 25228
rect 39564 25282 39620 25294
rect 39564 25230 39566 25282
rect 39618 25230 39620 25282
rect 39564 24948 39620 25230
rect 39788 24948 39844 24958
rect 39564 24946 39844 24948
rect 39564 24894 39790 24946
rect 39842 24894 39844 24946
rect 39564 24892 39844 24894
rect 39452 24670 39454 24722
rect 39506 24670 39508 24722
rect 39228 24610 39284 24622
rect 39228 24558 39230 24610
rect 39282 24558 39284 24610
rect 39228 23940 39284 24558
rect 39228 23874 39284 23884
rect 39340 23940 39396 23950
rect 39452 23940 39508 24670
rect 39340 23938 39508 23940
rect 39340 23886 39342 23938
rect 39394 23886 39508 23938
rect 39340 23884 39508 23886
rect 39788 23940 39844 24892
rect 39340 23874 39396 23884
rect 39788 23874 39844 23884
rect 39900 24834 39956 25788
rect 40236 25508 40292 26852
rect 39900 24782 39902 24834
rect 39954 24782 39956 24834
rect 38892 23660 39396 23716
rect 38444 23380 38500 23390
rect 37772 22978 37828 22988
rect 37884 23042 37940 23054
rect 37884 22990 37886 23042
rect 37938 22990 37940 23042
rect 37884 22932 37940 22990
rect 37884 22866 37940 22876
rect 38444 22708 38500 23324
rect 38444 22642 38500 22652
rect 37772 22260 37828 22270
rect 37772 22258 38164 22260
rect 37772 22206 37774 22258
rect 37826 22206 38164 22258
rect 37772 22204 38164 22206
rect 37772 22194 37828 22204
rect 38108 21810 38164 22204
rect 38108 21758 38110 21810
rect 38162 21758 38164 21810
rect 38108 21746 38164 21758
rect 38332 21586 38388 21598
rect 38332 21534 38334 21586
rect 38386 21534 38388 21586
rect 37772 21476 37828 21486
rect 38332 21476 38388 21534
rect 37772 21474 38388 21476
rect 37772 21422 37774 21474
rect 37826 21422 38388 21474
rect 37772 21420 38388 21422
rect 37772 21410 37828 21420
rect 38668 18564 38724 23660
rect 38780 23650 38836 23660
rect 38780 23156 38836 23166
rect 39116 23156 39172 23166
rect 38836 23154 39172 23156
rect 38836 23102 39118 23154
rect 39170 23102 39172 23154
rect 38836 23100 39172 23102
rect 38780 23062 38836 23100
rect 38780 21812 38836 21822
rect 38780 21718 38836 21756
rect 39116 21698 39172 23100
rect 39340 22596 39396 23660
rect 39452 23714 39508 23726
rect 39452 23662 39454 23714
rect 39506 23662 39508 23714
rect 39452 23492 39508 23662
rect 39452 23426 39508 23436
rect 39564 23716 39620 23726
rect 39452 23266 39508 23278
rect 39452 23214 39454 23266
rect 39506 23214 39508 23266
rect 39452 23156 39508 23214
rect 39564 23268 39620 23660
rect 39564 23202 39620 23212
rect 39452 23090 39508 23100
rect 39340 22540 39732 22596
rect 39116 21646 39118 21698
rect 39170 21646 39172 21698
rect 39116 21634 39172 21646
rect 38556 18508 38724 18564
rect 39340 19906 39396 19918
rect 39340 19854 39342 19906
rect 39394 19854 39396 19906
rect 39340 19796 39396 19854
rect 39340 18564 39396 19740
rect 37772 18340 37828 18350
rect 37772 18246 37828 18284
rect 37884 17666 37940 17678
rect 37884 17614 37886 17666
rect 37938 17614 37940 17666
rect 37884 16884 37940 17614
rect 37884 16790 37940 16828
rect 38556 16884 38612 18508
rect 39340 18498 39396 18508
rect 38668 17108 38724 17118
rect 38668 16994 38724 17052
rect 38668 16942 38670 16994
rect 38722 16942 38724 16994
rect 38668 16930 38724 16942
rect 38556 16818 38612 16828
rect 38892 16882 38948 16894
rect 38892 16830 38894 16882
rect 38946 16830 38948 16882
rect 37772 16212 37828 16222
rect 37772 16118 37828 16156
rect 38892 16212 38948 16830
rect 37772 15876 37828 15886
rect 37660 15820 37772 15876
rect 37660 15204 37716 15214
rect 37660 14756 37716 15148
rect 37772 15202 37828 15820
rect 38332 15426 38388 15438
rect 38332 15374 38334 15426
rect 38386 15374 38388 15426
rect 38332 15316 38388 15374
rect 38556 15316 38612 15326
rect 38332 15250 38388 15260
rect 38444 15314 38612 15316
rect 38444 15262 38558 15314
rect 38610 15262 38612 15314
rect 38444 15260 38612 15262
rect 37772 15150 37774 15202
rect 37826 15150 37828 15202
rect 37772 15138 37828 15150
rect 38444 15148 38500 15260
rect 38556 15250 38612 15260
rect 38892 15148 38948 16156
rect 39564 16882 39620 16894
rect 39564 16830 39566 16882
rect 39618 16830 39620 16882
rect 39116 15876 39172 15886
rect 39116 15538 39172 15820
rect 39564 15764 39620 16830
rect 39564 15698 39620 15708
rect 39116 15486 39118 15538
rect 39170 15486 39172 15538
rect 39116 15474 39172 15486
rect 39340 15260 39620 15316
rect 39340 15148 39396 15260
rect 38108 15092 38500 15148
rect 38780 15092 38948 15148
rect 39116 15092 39396 15148
rect 39564 15204 39620 15260
rect 39564 15138 39620 15148
rect 37660 14700 38052 14756
rect 37996 14530 38052 14700
rect 37996 14478 37998 14530
rect 38050 14478 38052 14530
rect 37996 14466 38052 14478
rect 37772 14308 37828 14318
rect 38108 14308 38164 15092
rect 38780 14756 38836 15092
rect 38332 14700 38836 14756
rect 38220 14642 38276 14654
rect 38220 14590 38222 14642
rect 38274 14590 38276 14642
rect 38220 14532 38276 14590
rect 38220 14466 38276 14476
rect 38332 14530 38388 14700
rect 38332 14478 38334 14530
rect 38386 14478 38388 14530
rect 38332 14466 38388 14478
rect 37772 14306 38164 14308
rect 37772 14254 37774 14306
rect 37826 14254 38164 14306
rect 37772 14252 38164 14254
rect 38556 14306 38612 14318
rect 38556 14254 38558 14306
rect 38610 14254 38612 14306
rect 37772 14242 37828 14252
rect 38556 13860 38612 14254
rect 38780 14308 38836 14700
rect 39004 14532 39060 14542
rect 39004 14438 39060 14476
rect 38780 14242 38836 14252
rect 37324 12086 37380 12124
rect 37436 12236 37604 12292
rect 37772 13636 37828 13646
rect 37324 11170 37380 11182
rect 37324 11118 37326 11170
rect 37378 11118 37380 11170
rect 37324 10500 37380 11118
rect 37436 10724 37492 12236
rect 37772 12178 37828 13580
rect 38444 13636 38500 13646
rect 38556 13636 38612 13804
rect 39004 13748 39060 13758
rect 38444 13634 38612 13636
rect 38444 13582 38446 13634
rect 38498 13582 38612 13634
rect 38444 13580 38612 13582
rect 38892 13692 39004 13748
rect 38108 13188 38164 13198
rect 38108 13094 38164 13132
rect 38220 12964 38276 12974
rect 38444 12964 38500 13580
rect 38892 13074 38948 13692
rect 39004 13682 39060 13692
rect 39116 13746 39172 15092
rect 39452 15090 39508 15102
rect 39452 15038 39454 15090
rect 39506 15038 39508 15090
rect 39340 14532 39396 14542
rect 39452 14532 39508 15038
rect 39340 14530 39508 14532
rect 39340 14478 39342 14530
rect 39394 14478 39508 14530
rect 39340 14476 39508 14478
rect 39228 13860 39284 13870
rect 39228 13766 39284 13804
rect 39116 13694 39118 13746
rect 39170 13694 39172 13746
rect 39116 13682 39172 13694
rect 39340 13412 39396 14476
rect 39452 14308 39508 14318
rect 39452 13858 39508 14252
rect 39452 13806 39454 13858
rect 39506 13806 39508 13858
rect 39452 13794 39508 13806
rect 39676 13748 39732 22540
rect 39900 22484 39956 24782
rect 40124 25506 40292 25508
rect 40124 25454 40238 25506
rect 40290 25454 40292 25506
rect 40124 25452 40292 25454
rect 40012 24724 40068 24734
rect 40012 24630 40068 24668
rect 40012 23940 40068 23950
rect 40124 23940 40180 25452
rect 40236 25442 40292 25452
rect 40012 23938 40180 23940
rect 40012 23886 40014 23938
rect 40066 23886 40180 23938
rect 40012 23884 40180 23886
rect 40012 23874 40068 23884
rect 39900 22390 39956 22428
rect 40236 23716 40292 23726
rect 40236 22258 40292 23660
rect 40460 22484 40516 22494
rect 40460 22370 40516 22428
rect 40460 22318 40462 22370
rect 40514 22318 40516 22370
rect 40460 22306 40516 22318
rect 40236 22206 40238 22258
rect 40290 22206 40292 22258
rect 40236 22194 40292 22206
rect 40012 20020 40068 20030
rect 40012 19124 40068 19964
rect 40348 20018 40404 20030
rect 40348 19966 40350 20018
rect 40402 19966 40404 20018
rect 40236 19908 40292 19918
rect 40236 19814 40292 19852
rect 40348 19684 40404 19966
rect 40348 19618 40404 19628
rect 39900 18340 39956 18350
rect 40012 18340 40068 19068
rect 40572 19012 40628 26908
rect 41020 26898 41076 26910
rect 40796 26516 40852 26526
rect 40684 25506 40740 25518
rect 40684 25454 40686 25506
rect 40738 25454 40740 25506
rect 40684 25396 40740 25454
rect 40796 25508 40852 26460
rect 40908 26404 40964 26414
rect 40908 26310 40964 26348
rect 41580 26404 41636 27694
rect 42140 27300 42196 27310
rect 42028 26962 42084 26974
rect 42028 26910 42030 26962
rect 42082 26910 42084 26962
rect 42028 26628 42084 26910
rect 42028 26562 42084 26572
rect 41580 26338 41636 26348
rect 41804 26516 41860 26526
rect 41804 26402 41860 26460
rect 41804 26350 41806 26402
rect 41858 26350 41860 26402
rect 41804 26338 41860 26350
rect 42028 26404 42084 26414
rect 42028 26310 42084 26348
rect 41020 26292 41076 26302
rect 41020 26290 41412 26292
rect 41020 26238 41022 26290
rect 41074 26238 41412 26290
rect 41020 26236 41412 26238
rect 41020 26226 41076 26236
rect 41132 26068 41188 26078
rect 41020 25508 41076 25518
rect 40796 25506 41076 25508
rect 40796 25454 41022 25506
rect 41074 25454 41076 25506
rect 40796 25452 41076 25454
rect 41020 25442 41076 25452
rect 40684 25330 40740 25340
rect 41020 25284 41076 25294
rect 41132 25284 41188 26012
rect 41020 25282 41188 25284
rect 41020 25230 41022 25282
rect 41074 25230 41188 25282
rect 41020 25228 41188 25230
rect 41244 26066 41300 26078
rect 41244 26014 41246 26066
rect 41298 26014 41300 26066
rect 41020 25218 41076 25228
rect 41244 23938 41300 26014
rect 41356 25506 41412 26236
rect 41356 25454 41358 25506
rect 41410 25454 41412 25506
rect 41356 25442 41412 25454
rect 41692 26290 41748 26302
rect 41692 26238 41694 26290
rect 41746 26238 41748 26290
rect 41692 24836 41748 26238
rect 42140 26292 42196 27244
rect 42252 27074 42308 28364
rect 42252 27022 42254 27074
rect 42306 27022 42308 27074
rect 42252 27010 42308 27022
rect 42140 26198 42196 26236
rect 42252 25956 42308 25966
rect 42028 25900 42252 25956
rect 42028 25506 42084 25900
rect 42252 25890 42308 25900
rect 42364 25620 42420 30268
rect 42700 29540 42756 29550
rect 42588 29426 42644 29438
rect 42588 29374 42590 29426
rect 42642 29374 42644 29426
rect 42476 28420 42532 28430
rect 42476 28082 42532 28364
rect 42588 28308 42644 29374
rect 42700 28756 42756 29484
rect 42924 29428 42980 29438
rect 43260 29428 43316 29438
rect 42924 29426 43316 29428
rect 42924 29374 42926 29426
rect 42978 29374 43262 29426
rect 43314 29374 43316 29426
rect 42924 29372 43316 29374
rect 42924 29362 42980 29372
rect 43260 29362 43316 29372
rect 43372 29428 43428 30942
rect 43484 31780 43540 31790
rect 43484 30324 43540 31724
rect 43708 31668 43764 31836
rect 43708 31574 43764 31612
rect 43484 30210 43540 30268
rect 43484 30158 43486 30210
rect 43538 30158 43540 30210
rect 43484 30146 43540 30158
rect 43820 30212 43876 33628
rect 43932 33124 43988 34076
rect 44044 33346 44100 34412
rect 44156 33570 44212 34748
rect 44268 34692 44324 34702
rect 44268 34598 44324 34636
rect 44156 33518 44158 33570
rect 44210 33518 44212 33570
rect 44156 33506 44212 33518
rect 44268 33572 44324 33582
rect 44044 33294 44046 33346
rect 44098 33294 44100 33346
rect 44044 33282 44100 33294
rect 44156 33124 44212 33134
rect 43932 33122 44212 33124
rect 43932 33070 44158 33122
rect 44210 33070 44212 33122
rect 43932 33068 44212 33070
rect 44156 32676 44212 33068
rect 44156 32610 44212 32620
rect 44044 32450 44100 32462
rect 44044 32398 44046 32450
rect 44098 32398 44100 32450
rect 44044 32002 44100 32398
rect 44044 31950 44046 32002
rect 44098 31950 44100 32002
rect 44044 31938 44100 31950
rect 44268 31890 44324 33516
rect 44380 33460 44436 35084
rect 44940 35026 44996 35532
rect 45276 35586 45332 36540
rect 45276 35534 45278 35586
rect 45330 35534 45332 35586
rect 45276 35522 45332 35534
rect 45388 36482 45444 36494
rect 45388 36430 45390 36482
rect 45442 36430 45444 36482
rect 45388 35700 45444 36430
rect 45948 35700 46004 38780
rect 46172 38724 46228 38734
rect 46060 38668 46172 38724
rect 46060 37044 46116 38668
rect 46172 38658 46228 38668
rect 46284 37940 46340 40238
rect 46396 42084 46452 42094
rect 46396 40292 46452 42028
rect 46508 40516 46564 43596
rect 46620 40628 46676 45724
rect 47404 45780 47460 45790
rect 47404 45686 47460 45724
rect 46844 45666 46900 45678
rect 46844 45614 46846 45666
rect 46898 45614 46900 45666
rect 46844 42980 46900 45614
rect 47516 45666 47572 45678
rect 47516 45614 47518 45666
rect 47570 45614 47572 45666
rect 47068 44100 47124 44110
rect 47068 43708 47124 44044
rect 47516 43708 47572 45614
rect 47628 45666 47684 45678
rect 47628 45614 47630 45666
rect 47682 45614 47684 45666
rect 47628 45444 47684 45614
rect 47628 45378 47684 45388
rect 48188 45666 48244 45678
rect 48188 45614 48190 45666
rect 48242 45614 48244 45666
rect 48188 45444 48244 45614
rect 48188 45378 48244 45388
rect 48188 45106 48244 45118
rect 48188 45054 48190 45106
rect 48242 45054 48244 45106
rect 47628 44996 47684 45006
rect 47628 44902 47684 44940
rect 47740 44434 47796 44446
rect 47740 44382 47742 44434
rect 47794 44382 47796 44434
rect 47068 43652 47348 43708
rect 47516 43652 47684 43708
rect 46844 42914 46900 42924
rect 46956 43092 47012 43102
rect 46732 42756 46788 42766
rect 46732 42530 46788 42700
rect 46844 42756 46900 42766
rect 46956 42756 47012 43036
rect 46844 42754 47012 42756
rect 46844 42702 46846 42754
rect 46898 42702 47012 42754
rect 46844 42700 47012 42702
rect 46844 42690 46900 42700
rect 47068 42644 47124 42654
rect 46732 42478 46734 42530
rect 46786 42478 46788 42530
rect 46732 42466 46788 42478
rect 46956 42642 47124 42644
rect 46956 42590 47070 42642
rect 47122 42590 47124 42642
rect 46956 42588 47124 42590
rect 46956 42084 47012 42588
rect 47068 42578 47124 42588
rect 47292 42196 47348 43652
rect 47404 43426 47460 43438
rect 47404 43374 47406 43426
rect 47458 43374 47460 43426
rect 47404 42978 47460 43374
rect 47404 42926 47406 42978
rect 47458 42926 47460 42978
rect 47404 42914 47460 42926
rect 47516 42980 47572 42990
rect 47516 42886 47572 42924
rect 47292 42130 47348 42140
rect 46956 42018 47012 42028
rect 47404 41300 47460 41310
rect 47628 41300 47684 43652
rect 47740 43092 47796 44382
rect 48188 44100 48244 45054
rect 48188 44006 48244 44044
rect 48076 43540 48132 43550
rect 47740 43026 47796 43036
rect 47964 43538 48132 43540
rect 47964 43486 48078 43538
rect 48130 43486 48132 43538
rect 47964 43484 48132 43486
rect 47740 42756 47796 42766
rect 47740 42662 47796 42700
rect 47852 42754 47908 42766
rect 47852 42702 47854 42754
rect 47906 42702 47908 42754
rect 47852 42532 47908 42702
rect 47852 42466 47908 42476
rect 47404 41298 47684 41300
rect 47404 41246 47406 41298
rect 47458 41246 47684 41298
rect 47404 41244 47684 41246
rect 47964 42082 48020 43484
rect 48076 43474 48132 43484
rect 47964 42030 47966 42082
rect 48018 42030 48020 42082
rect 47404 41234 47460 41244
rect 47964 41188 48020 42030
rect 48076 41188 48132 41198
rect 48020 41186 48132 41188
rect 48020 41134 48078 41186
rect 48130 41134 48132 41186
rect 48020 41132 48132 41134
rect 47964 41094 48020 41132
rect 46620 40572 47012 40628
rect 46956 40516 47012 40572
rect 47068 40516 47124 40526
rect 46956 40514 47124 40516
rect 46956 40462 47070 40514
rect 47122 40462 47124 40514
rect 46956 40460 47124 40462
rect 46508 40450 46564 40460
rect 47068 40450 47124 40460
rect 47964 40516 48020 40526
rect 47964 40422 48020 40460
rect 46620 40402 46676 40414
rect 46620 40350 46622 40402
rect 46674 40350 46676 40402
rect 46396 40236 46564 40292
rect 46396 39396 46452 39406
rect 46396 38946 46452 39340
rect 46396 38894 46398 38946
rect 46450 38894 46452 38946
rect 46396 38882 46452 38894
rect 46508 38668 46564 40236
rect 46620 40180 46676 40350
rect 46620 39508 46676 40124
rect 47292 40402 47348 40414
rect 47292 40350 47294 40402
rect 47346 40350 47348 40402
rect 47068 39508 47124 39518
rect 46620 39452 47068 39508
rect 47068 39442 47124 39452
rect 46732 39284 46788 39294
rect 46732 39058 46788 39228
rect 46732 39006 46734 39058
rect 46786 39006 46788 39058
rect 46732 38994 46788 39006
rect 46844 39060 46900 39070
rect 46844 38966 46900 39004
rect 46620 38948 46676 38958
rect 46620 38854 46676 38892
rect 47068 38948 47124 38958
rect 46956 38836 47012 38846
rect 46956 38742 47012 38780
rect 46508 38612 46788 38668
rect 46732 38050 46788 38612
rect 47068 38276 47124 38892
rect 47292 38724 47348 40350
rect 47740 40402 47796 40414
rect 47740 40350 47742 40402
rect 47794 40350 47796 40402
rect 47516 40290 47572 40302
rect 47516 40238 47518 40290
rect 47570 40238 47572 40290
rect 47404 39732 47460 39742
rect 47516 39732 47572 40238
rect 47404 39730 47572 39732
rect 47404 39678 47406 39730
rect 47458 39678 47572 39730
rect 47404 39676 47572 39678
rect 47740 39844 47796 40350
rect 47404 39666 47460 39676
rect 47740 38948 47796 39788
rect 48076 39618 48132 41132
rect 48076 39566 48078 39618
rect 48130 39566 48132 39618
rect 48076 39554 48132 39566
rect 48188 39172 48244 39182
rect 47740 38882 47796 38892
rect 47852 38948 47908 38958
rect 47852 38946 48020 38948
rect 47852 38894 47854 38946
rect 47906 38894 48020 38946
rect 47852 38892 48020 38894
rect 47852 38882 47908 38892
rect 47404 38836 47460 38846
rect 47404 38742 47460 38780
rect 47292 38658 47348 38668
rect 47516 38724 47572 38734
rect 47516 38722 47908 38724
rect 47516 38670 47518 38722
rect 47570 38670 47908 38722
rect 47516 38668 47908 38670
rect 47516 38658 47572 38668
rect 47740 38500 47796 38510
rect 47012 38220 47124 38276
rect 47404 38276 47460 38286
rect 47012 38052 47068 38220
rect 47404 38162 47460 38220
rect 47404 38110 47406 38162
rect 47458 38110 47460 38162
rect 47404 38098 47460 38110
rect 46732 37998 46734 38050
rect 46786 37998 46788 38050
rect 46172 37884 46340 37940
rect 46396 37940 46452 37950
rect 46452 37884 46676 37940
rect 46172 37378 46228 37884
rect 46396 37874 46452 37884
rect 46284 37492 46340 37502
rect 46284 37398 46340 37436
rect 46172 37326 46174 37378
rect 46226 37326 46228 37378
rect 46172 37314 46228 37326
rect 46284 37044 46340 37054
rect 46060 37042 46340 37044
rect 46060 36990 46286 37042
rect 46338 36990 46340 37042
rect 46060 36988 46340 36990
rect 46284 36978 46340 36988
rect 46060 36372 46116 36382
rect 46060 36370 46340 36372
rect 46060 36318 46062 36370
rect 46114 36318 46340 36370
rect 46060 36316 46340 36318
rect 46060 36306 46116 36316
rect 46284 35810 46340 36316
rect 46284 35758 46286 35810
rect 46338 35758 46340 35810
rect 46284 35746 46340 35758
rect 46060 35700 46116 35710
rect 45948 35698 46116 35700
rect 45948 35646 46062 35698
rect 46114 35646 46116 35698
rect 45948 35644 46116 35646
rect 44940 34974 44942 35026
rect 44994 34974 44996 35026
rect 44940 34962 44996 34974
rect 45388 34914 45444 35644
rect 46060 35634 46116 35644
rect 46396 35698 46452 35710
rect 46396 35646 46398 35698
rect 46450 35646 46452 35698
rect 46172 35588 46228 35598
rect 46396 35588 46452 35646
rect 46620 35700 46676 37884
rect 46732 35812 46788 37998
rect 46956 37996 47068 38052
rect 47516 38050 47572 38062
rect 47516 37998 47518 38050
rect 47570 37998 47572 38050
rect 46844 37826 46900 37838
rect 46844 37774 46846 37826
rect 46898 37774 46900 37826
rect 46844 36260 46900 37774
rect 46956 37716 47012 37996
rect 46956 37660 47124 37716
rect 47068 37490 47124 37660
rect 47068 37438 47070 37490
rect 47122 37438 47124 37490
rect 47068 37426 47124 37438
rect 46844 36194 46900 36204
rect 46956 37378 47012 37390
rect 46956 37326 46958 37378
rect 47010 37326 47012 37378
rect 46956 36036 47012 37326
rect 47068 37268 47124 37278
rect 47068 37174 47124 37212
rect 46956 35980 47460 36036
rect 47068 35812 47124 35822
rect 46732 35810 47124 35812
rect 46732 35758 47070 35810
rect 47122 35758 47124 35810
rect 46732 35756 47124 35758
rect 47068 35746 47124 35756
rect 47404 35812 47460 35980
rect 47404 35718 47460 35756
rect 47516 35922 47572 37998
rect 47628 37938 47684 37950
rect 47628 37886 47630 37938
rect 47682 37886 47684 37938
rect 47628 37492 47684 37886
rect 47628 37426 47684 37436
rect 47740 37378 47796 38444
rect 47740 37326 47742 37378
rect 47794 37326 47796 37378
rect 47740 37314 47796 37326
rect 47852 37268 47908 38668
rect 47852 37174 47908 37212
rect 47516 35870 47518 35922
rect 47570 35870 47572 35922
rect 46620 35644 47012 35700
rect 46228 35532 46452 35588
rect 46956 35586 47012 35644
rect 46956 35534 46958 35586
rect 47010 35534 47012 35586
rect 45836 35476 45892 35486
rect 45836 35382 45892 35420
rect 45388 34862 45390 34914
rect 45442 34862 45444 34914
rect 44380 33394 44436 33404
rect 44940 33572 44996 33582
rect 44940 33458 44996 33516
rect 44940 33406 44942 33458
rect 44994 33406 44996 33458
rect 44940 33394 44996 33406
rect 45388 33124 45444 34862
rect 46060 34802 46116 34814
rect 46060 34750 46062 34802
rect 46114 34750 46116 34802
rect 46060 33458 46116 34750
rect 46060 33406 46062 33458
rect 46114 33406 46116 33458
rect 46060 33394 46116 33406
rect 45500 33348 45556 33358
rect 45500 33254 45556 33292
rect 45948 33348 46004 33358
rect 45836 33236 45892 33246
rect 45388 33058 45444 33068
rect 45724 33234 45892 33236
rect 45724 33182 45838 33234
rect 45890 33182 45892 33234
rect 45724 33180 45892 33182
rect 44492 32788 44548 32798
rect 44492 32694 44548 32732
rect 44940 32676 44996 32686
rect 44940 32004 44996 32620
rect 45052 32004 45108 32014
rect 44940 31948 45052 32004
rect 45052 31938 45108 31948
rect 44268 31838 44270 31890
rect 44322 31838 44324 31890
rect 44044 31780 44100 31790
rect 44044 31218 44100 31724
rect 44268 31780 44324 31838
rect 44268 31714 44324 31724
rect 44828 31778 44884 31790
rect 44828 31726 44830 31778
rect 44882 31726 44884 31778
rect 44044 31166 44046 31218
rect 44098 31166 44100 31218
rect 44044 31154 44100 31166
rect 44156 31220 44212 31230
rect 44156 31126 44212 31164
rect 44268 31108 44324 31118
rect 44268 31014 44324 31052
rect 43932 30996 43988 31006
rect 43932 30902 43988 30940
rect 44492 30994 44548 31006
rect 44492 30942 44494 30994
rect 44546 30942 44548 30994
rect 44492 30772 44548 30942
rect 44828 30996 44884 31726
rect 45052 31780 45108 31790
rect 45052 31686 45108 31724
rect 45388 31778 45444 31790
rect 45388 31726 45390 31778
rect 45442 31726 45444 31778
rect 45164 31668 45220 31678
rect 45164 31574 45220 31612
rect 45276 31554 45332 31566
rect 45276 31502 45278 31554
rect 45330 31502 45332 31554
rect 45276 31108 45332 31502
rect 45276 31042 45332 31052
rect 44828 30930 44884 30940
rect 45052 30884 45108 30894
rect 44940 30882 45108 30884
rect 44940 30830 45054 30882
rect 45106 30830 45108 30882
rect 44940 30828 45108 30830
rect 44940 30772 44996 30828
rect 45052 30818 45108 30828
rect 44492 30716 44996 30772
rect 43876 30156 44100 30212
rect 43820 30146 43876 30156
rect 43820 29484 43988 29540
rect 43372 29362 43428 29372
rect 43708 29428 43764 29438
rect 43820 29428 43876 29484
rect 43708 29426 43876 29428
rect 43708 29374 43710 29426
rect 43762 29374 43876 29426
rect 43708 29372 43876 29374
rect 43708 29362 43764 29372
rect 43708 28866 43764 28878
rect 43708 28814 43710 28866
rect 43762 28814 43764 28866
rect 43708 28756 43764 28814
rect 42700 28700 42980 28756
rect 42812 28530 42868 28542
rect 42812 28478 42814 28530
rect 42866 28478 42868 28530
rect 42700 28308 42756 28318
rect 42812 28308 42868 28478
rect 42924 28420 42980 28700
rect 43596 28754 43764 28756
rect 43596 28702 43710 28754
rect 43762 28702 43764 28754
rect 43596 28700 43764 28702
rect 43372 28644 43428 28654
rect 43372 28550 43428 28588
rect 43036 28420 43092 28430
rect 42924 28418 43092 28420
rect 42924 28366 43038 28418
rect 43090 28366 43092 28418
rect 42924 28364 43092 28366
rect 42588 28252 42700 28308
rect 42756 28252 42868 28308
rect 42700 28242 42756 28252
rect 42476 28030 42478 28082
rect 42530 28030 42532 28082
rect 42476 28018 42532 28030
rect 43036 27636 43092 28364
rect 43260 28420 43316 28430
rect 43260 28326 43316 28364
rect 43596 27858 43652 28700
rect 43708 28690 43764 28700
rect 43596 27806 43598 27858
rect 43650 27806 43652 27858
rect 43596 27794 43652 27806
rect 43820 28420 43876 28430
rect 43932 28420 43988 29484
rect 44044 28868 44100 30156
rect 44156 29316 44212 29326
rect 44156 29222 44212 29260
rect 44044 28866 44212 28868
rect 44044 28814 44046 28866
rect 44098 28814 44212 28866
rect 44044 28812 44212 28814
rect 44044 28802 44100 28812
rect 44156 28754 44212 28812
rect 44156 28702 44158 28754
rect 44210 28702 44212 28754
rect 44156 28690 44212 28702
rect 44828 28644 44884 28654
rect 43876 28364 43988 28420
rect 44380 28642 44884 28644
rect 44380 28590 44830 28642
rect 44882 28590 44884 28642
rect 44380 28588 44884 28590
rect 43036 27570 43092 27580
rect 43596 27636 43652 27646
rect 42476 27300 42532 27310
rect 42476 27186 42532 27244
rect 42476 27134 42478 27186
rect 42530 27134 42532 27186
rect 42476 27122 42532 27134
rect 42700 27300 42756 27310
rect 42700 27074 42756 27244
rect 42700 27022 42702 27074
rect 42754 27022 42756 27074
rect 42700 27010 42756 27022
rect 43148 27076 43204 27114
rect 43148 27010 43204 27020
rect 43596 27074 43652 27580
rect 43596 27022 43598 27074
rect 43650 27022 43652 27074
rect 43596 27010 43652 27022
rect 43820 27300 43876 28364
rect 43820 27244 44100 27300
rect 42924 26964 42980 27002
rect 42924 26898 42980 26908
rect 43820 26962 43876 27244
rect 43820 26910 43822 26962
rect 43874 26910 43876 26962
rect 43820 26898 43876 26910
rect 43932 27074 43988 27086
rect 43932 27022 43934 27074
rect 43986 27022 43988 27074
rect 43932 26964 43988 27022
rect 43932 26898 43988 26908
rect 42476 26850 42532 26862
rect 42476 26798 42478 26850
rect 42530 26798 42532 26850
rect 42476 26740 42532 26798
rect 42476 26674 42532 26684
rect 43932 26628 43988 26638
rect 43932 26514 43988 26572
rect 43932 26462 43934 26514
rect 43986 26462 43988 26514
rect 43932 26450 43988 26462
rect 42812 26404 42868 26414
rect 42812 26310 42868 26348
rect 43036 26402 43092 26414
rect 43036 26350 43038 26402
rect 43090 26350 43092 26402
rect 42588 26290 42644 26302
rect 42588 26238 42590 26290
rect 42642 26238 42644 26290
rect 42588 26068 42644 26238
rect 42588 26002 42644 26012
rect 42700 26178 42756 26190
rect 42700 26126 42702 26178
rect 42754 26126 42756 26178
rect 42700 25956 42756 26126
rect 42700 25890 42756 25900
rect 43036 25844 43092 26350
rect 43484 26404 43540 26414
rect 43484 26310 43540 26348
rect 44044 26402 44100 27244
rect 44380 26740 44436 28588
rect 44828 28578 44884 28588
rect 44940 27300 44996 30716
rect 45276 30324 45332 30334
rect 45388 30324 45444 31726
rect 45724 31778 45780 33180
rect 45836 33170 45892 33180
rect 45724 31726 45726 31778
rect 45778 31726 45780 31778
rect 45724 31714 45780 31726
rect 45948 32562 46004 33292
rect 46060 33236 46116 33246
rect 46172 33236 46228 35532
rect 46956 35522 47012 35534
rect 46508 35476 46564 35486
rect 46396 35252 46452 35262
rect 46396 33570 46452 35196
rect 46396 33518 46398 33570
rect 46450 33518 46452 33570
rect 46396 33506 46452 33518
rect 46508 33572 46564 35420
rect 46620 35474 46676 35486
rect 46620 35422 46622 35474
rect 46674 35422 46676 35474
rect 46620 34244 46676 35422
rect 47516 35252 47572 35870
rect 47516 35186 47572 35196
rect 47852 35810 47908 35822
rect 47852 35758 47854 35810
rect 47906 35758 47908 35810
rect 47852 34356 47908 35758
rect 46620 34178 46676 34188
rect 47516 34300 47908 34356
rect 46956 34018 47012 34030
rect 46956 33966 46958 34018
rect 47010 33966 47012 34018
rect 46620 33572 46676 33582
rect 46508 33570 46676 33572
rect 46508 33518 46622 33570
rect 46674 33518 46676 33570
rect 46508 33516 46676 33518
rect 46620 33506 46676 33516
rect 46060 33234 46228 33236
rect 46060 33182 46062 33234
rect 46114 33182 46228 33234
rect 46060 33180 46228 33182
rect 46060 33170 46116 33180
rect 46956 33124 47012 33966
rect 46956 33058 47012 33068
rect 47068 33346 47124 33358
rect 47068 33294 47070 33346
rect 47122 33294 47124 33346
rect 45948 32510 45950 32562
rect 46002 32510 46004 32562
rect 45948 31666 46004 32510
rect 46060 33012 46116 33022
rect 46060 31778 46116 32956
rect 47068 31892 47124 33294
rect 47516 33348 47572 34300
rect 47964 33460 48020 38892
rect 48188 38836 48244 39116
rect 48188 38834 48468 38836
rect 48188 38782 48190 38834
rect 48242 38782 48468 38834
rect 48188 38780 48468 38782
rect 48188 38770 48244 38780
rect 48188 37268 48244 37278
rect 48188 36594 48244 37212
rect 48412 37268 48468 38780
rect 48412 37202 48468 37212
rect 48188 36542 48190 36594
rect 48242 36542 48244 36594
rect 48188 36530 48244 36542
rect 48188 35924 48244 35934
rect 48244 35868 48356 35924
rect 48188 35830 48244 35868
rect 48076 35812 48132 35822
rect 48076 35028 48132 35756
rect 48188 35028 48244 35038
rect 48076 35026 48244 35028
rect 48076 34974 48190 35026
rect 48242 34974 48244 35026
rect 48076 34972 48244 34974
rect 48188 34962 48244 34972
rect 48076 34244 48132 34254
rect 48076 33570 48132 34188
rect 48076 33518 48078 33570
rect 48130 33518 48132 33570
rect 48076 33506 48132 33518
rect 47516 33282 47572 33292
rect 47628 33404 48020 33460
rect 47628 33346 47684 33404
rect 47628 33294 47630 33346
rect 47682 33294 47684 33346
rect 47628 33282 47684 33294
rect 47964 33348 48020 33404
rect 47964 33292 48132 33348
rect 48076 33236 48132 33292
rect 48076 33234 48244 33236
rect 47964 33178 48020 33190
rect 47852 33124 47908 33134
rect 47068 31826 47124 31836
rect 47628 32004 47684 32014
rect 46060 31726 46062 31778
rect 46114 31726 46116 31778
rect 46060 31714 46116 31726
rect 46172 31780 46228 31790
rect 46228 31724 46340 31780
rect 46172 31714 46228 31724
rect 45948 31614 45950 31666
rect 46002 31614 46004 31666
rect 45948 31602 46004 31614
rect 45164 30322 45444 30324
rect 45164 30270 45278 30322
rect 45330 30270 45444 30322
rect 45164 30268 45444 30270
rect 45052 28644 45108 28654
rect 45052 28550 45108 28588
rect 44940 27234 44996 27244
rect 45052 28420 45108 28430
rect 44380 26514 44436 26684
rect 44380 26462 44382 26514
rect 44434 26462 44436 26514
rect 44380 26450 44436 26462
rect 44492 26964 44548 26974
rect 44044 26350 44046 26402
rect 44098 26350 44100 26402
rect 44044 26338 44100 26350
rect 44492 26402 44548 26908
rect 44492 26350 44494 26402
rect 44546 26350 44548 26402
rect 44492 26338 44548 26350
rect 44828 26852 44884 26862
rect 43596 26292 43652 26302
rect 43596 26198 43652 26236
rect 44828 26292 44884 26796
rect 44940 26516 44996 26526
rect 44940 26422 44996 26460
rect 44828 26290 44996 26292
rect 44828 26238 44830 26290
rect 44882 26238 44996 26290
rect 44828 26236 44996 26238
rect 44828 26226 44884 26236
rect 43148 25844 43204 25854
rect 43036 25788 43148 25844
rect 42364 25564 42532 25620
rect 42028 25454 42030 25506
rect 42082 25454 42084 25506
rect 42028 25442 42084 25454
rect 42364 25394 42420 25406
rect 42364 25342 42366 25394
rect 42418 25342 42420 25394
rect 41692 24770 41748 24780
rect 42252 25282 42308 25294
rect 42252 25230 42254 25282
rect 42306 25230 42308 25282
rect 41916 24164 41972 24174
rect 41244 23886 41246 23938
rect 41298 23886 41300 23938
rect 41244 23874 41300 23886
rect 41804 23940 41860 23950
rect 41804 23846 41860 23884
rect 41692 23826 41748 23838
rect 41692 23774 41694 23826
rect 41746 23774 41748 23826
rect 41020 23716 41076 23726
rect 41020 23714 41300 23716
rect 41020 23662 41022 23714
rect 41074 23662 41300 23714
rect 41020 23660 41300 23662
rect 41020 23650 41076 23660
rect 41244 22372 41300 23660
rect 41580 23492 41636 23502
rect 41468 23156 41524 23166
rect 41580 23156 41636 23436
rect 41692 23380 41748 23774
rect 41804 23380 41860 23390
rect 41692 23378 41860 23380
rect 41692 23326 41806 23378
rect 41858 23326 41860 23378
rect 41692 23324 41860 23326
rect 41804 23314 41860 23324
rect 41692 23156 41748 23166
rect 41580 23154 41748 23156
rect 41580 23102 41694 23154
rect 41746 23102 41748 23154
rect 41580 23100 41748 23102
rect 41468 23062 41524 23100
rect 41692 23090 41748 23100
rect 41916 23154 41972 24108
rect 42028 23938 42084 23950
rect 42028 23886 42030 23938
rect 42082 23886 42084 23938
rect 42028 23380 42084 23886
rect 42084 23324 42196 23380
rect 42028 23314 42084 23324
rect 41916 23102 41918 23154
rect 41970 23102 41972 23154
rect 41916 23090 41972 23102
rect 41356 22372 41412 22382
rect 41244 22370 41412 22372
rect 41244 22318 41358 22370
rect 41410 22318 41412 22370
rect 41244 22316 41412 22318
rect 41356 22306 41412 22316
rect 42028 22370 42084 22382
rect 42028 22318 42030 22370
rect 42082 22318 42084 22370
rect 41804 22260 41860 22270
rect 41468 22148 41524 22158
rect 41468 22054 41524 22092
rect 41804 21810 41860 22204
rect 41804 21758 41806 21810
rect 41858 21758 41860 21810
rect 41804 21746 41860 21758
rect 41916 21924 41972 21934
rect 41916 21810 41972 21868
rect 41916 21758 41918 21810
rect 41970 21758 41972 21810
rect 41916 21746 41972 21758
rect 41468 21586 41524 21598
rect 41692 21588 41748 21598
rect 41468 21534 41470 21586
rect 41522 21534 41524 21586
rect 41468 20916 41524 21534
rect 41132 20860 41524 20916
rect 41580 21586 41748 21588
rect 41580 21534 41694 21586
rect 41746 21534 41748 21586
rect 41580 21532 41748 21534
rect 41020 20580 41076 20590
rect 41132 20580 41188 20860
rect 41244 20692 41300 20702
rect 41244 20598 41300 20636
rect 41356 20690 41412 20702
rect 41356 20638 41358 20690
rect 41410 20638 41412 20690
rect 41020 20578 41188 20580
rect 41020 20526 41022 20578
rect 41074 20526 41188 20578
rect 41020 20524 41188 20526
rect 41020 20132 41076 20524
rect 41356 20356 41412 20638
rect 41580 20692 41636 21532
rect 41692 21522 41748 21532
rect 41804 21476 41860 21486
rect 41804 20914 41860 21420
rect 42028 21028 42084 22318
rect 42140 21924 42196 23324
rect 42252 23378 42308 25230
rect 42364 25284 42420 25342
rect 42364 25218 42420 25228
rect 42476 25060 42532 25564
rect 43148 25506 43204 25788
rect 44940 25620 44996 26236
rect 45052 26290 45108 28364
rect 45052 26238 45054 26290
rect 45106 26238 45108 26290
rect 45052 26226 45108 26238
rect 45164 26292 45220 30268
rect 45276 30258 45332 30268
rect 45388 29428 45444 29438
rect 45388 29426 45556 29428
rect 45388 29374 45390 29426
rect 45442 29374 45556 29426
rect 45388 29372 45556 29374
rect 45388 29362 45444 29372
rect 45388 28420 45444 28430
rect 45388 28326 45444 28364
rect 45388 27748 45444 27758
rect 45500 27748 45556 29372
rect 45724 29316 45780 29326
rect 45724 28866 45780 29260
rect 45724 28814 45726 28866
rect 45778 28814 45780 28866
rect 45724 28802 45780 28814
rect 46060 29314 46116 29326
rect 46060 29262 46062 29314
rect 46114 29262 46116 29314
rect 46060 28866 46116 29262
rect 46060 28814 46062 28866
rect 46114 28814 46116 28866
rect 46060 28802 46116 28814
rect 45836 28756 45892 28766
rect 45892 28700 46004 28756
rect 45836 28690 45892 28700
rect 45948 28644 46004 28700
rect 46060 28644 46116 28654
rect 45948 28642 46116 28644
rect 45948 28590 46062 28642
rect 46114 28590 46116 28642
rect 45948 28588 46116 28590
rect 45388 27746 45556 27748
rect 45388 27694 45390 27746
rect 45442 27694 45556 27746
rect 45388 27692 45556 27694
rect 45276 27076 45332 27086
rect 45388 27076 45444 27692
rect 45276 27074 45444 27076
rect 45276 27022 45278 27074
rect 45330 27022 45444 27074
rect 45276 27020 45444 27022
rect 45276 27010 45332 27020
rect 44940 25564 45108 25620
rect 43148 25454 43150 25506
rect 43202 25454 43204 25506
rect 43148 25442 43204 25454
rect 43596 25508 43652 25518
rect 42364 25004 42532 25060
rect 42588 25394 42644 25406
rect 42588 25342 42590 25394
rect 42642 25342 42644 25394
rect 42364 23604 42420 25004
rect 42588 24946 42644 25342
rect 43372 25396 43428 25406
rect 42588 24894 42590 24946
rect 42642 24894 42644 24946
rect 42588 24882 42644 24894
rect 42812 25282 42868 25294
rect 42812 25230 42814 25282
rect 42866 25230 42868 25282
rect 42476 24836 42532 24846
rect 42476 24052 42532 24780
rect 42812 24164 42868 25230
rect 43036 25284 43092 25294
rect 43036 25190 43092 25228
rect 43148 24836 43204 24846
rect 43148 24742 43204 24780
rect 43036 24500 43092 24510
rect 42812 24098 42868 24108
rect 42924 24498 43092 24500
rect 42924 24446 43038 24498
rect 43090 24446 43092 24498
rect 42924 24444 43092 24446
rect 42588 24052 42644 24062
rect 42476 24050 42644 24052
rect 42476 23998 42590 24050
rect 42642 23998 42644 24050
rect 42476 23996 42644 23998
rect 42588 23986 42644 23996
rect 42924 23826 42980 24444
rect 43036 24434 43092 24444
rect 43148 23940 43204 23950
rect 43148 23846 43204 23884
rect 42924 23774 42926 23826
rect 42978 23774 42980 23826
rect 42924 23762 42980 23774
rect 42364 23538 42420 23548
rect 42588 23714 42644 23726
rect 42588 23662 42590 23714
rect 42642 23662 42644 23714
rect 42252 23326 42254 23378
rect 42306 23326 42308 23378
rect 42252 23314 42308 23326
rect 42476 23156 42532 23166
rect 42364 23042 42420 23054
rect 42364 22990 42366 23042
rect 42418 22990 42420 23042
rect 42364 22258 42420 22990
rect 42476 22596 42532 23100
rect 42588 22820 42644 23662
rect 42700 23716 42756 23726
rect 42700 23714 42868 23716
rect 42700 23662 42702 23714
rect 42754 23662 42868 23714
rect 42700 23660 42868 23662
rect 42700 23650 42756 23660
rect 42812 23492 42868 23660
rect 42812 23426 42868 23436
rect 42700 23380 42756 23390
rect 42700 23286 42756 23324
rect 42588 22764 43204 22820
rect 42476 22540 42756 22596
rect 42700 22372 42756 22540
rect 43036 22484 43092 22494
rect 42812 22372 42868 22382
rect 42700 22370 42868 22372
rect 42700 22318 42814 22370
rect 42866 22318 42868 22370
rect 42700 22316 42868 22318
rect 42812 22306 42868 22316
rect 42364 22206 42366 22258
rect 42418 22206 42420 22258
rect 42364 22194 42420 22206
rect 42924 22260 42980 22270
rect 42924 22166 42980 22204
rect 42140 21868 42532 21924
rect 42476 21812 42532 21868
rect 42476 21756 42644 21812
rect 42140 21586 42196 21598
rect 42140 21534 42142 21586
rect 42194 21534 42196 21586
rect 42140 21252 42196 21534
rect 42476 21476 42532 21486
rect 42476 21382 42532 21420
rect 42588 21474 42644 21756
rect 43036 21586 43092 22428
rect 43148 22372 43204 22764
rect 43372 22596 43428 25340
rect 43596 24836 43652 25452
rect 44044 25508 44100 25518
rect 44044 25414 44100 25452
rect 44268 25396 44324 25406
rect 44828 25396 44884 25406
rect 44268 25394 44884 25396
rect 44268 25342 44270 25394
rect 44322 25342 44830 25394
rect 44882 25342 44884 25394
rect 44268 25340 44884 25342
rect 44268 25330 44324 25340
rect 43820 25282 43876 25294
rect 43820 25230 43822 25282
rect 43874 25230 43876 25282
rect 43820 25060 43876 25230
rect 43932 25284 43988 25294
rect 43932 25190 43988 25228
rect 43820 25004 44100 25060
rect 44044 24946 44100 25004
rect 44044 24894 44046 24946
rect 44098 24894 44100 24946
rect 44044 24882 44100 24894
rect 43596 24770 43652 24780
rect 44828 24722 44884 25340
rect 44828 24670 44830 24722
rect 44882 24670 44884 24722
rect 44828 24658 44884 24670
rect 44940 25396 44996 25406
rect 44156 24610 44212 24622
rect 44156 24558 44158 24610
rect 44210 24558 44212 24610
rect 43596 23940 43652 23950
rect 43596 23846 43652 23884
rect 44156 23940 44212 24558
rect 44156 23874 44212 23884
rect 43708 23826 43764 23838
rect 43708 23774 43710 23826
rect 43762 23774 43764 23826
rect 43708 23716 43764 23774
rect 43820 23828 43876 23838
rect 44044 23828 44100 23838
rect 43820 23826 44044 23828
rect 43820 23774 43822 23826
rect 43874 23774 44044 23826
rect 43820 23772 44044 23774
rect 43820 23762 43876 23772
rect 44044 23762 44100 23772
rect 43708 23650 43764 23660
rect 44268 23714 44324 23726
rect 44268 23662 44270 23714
rect 44322 23662 44324 23714
rect 43596 23604 43652 23614
rect 43372 22530 43428 22540
rect 43484 22708 43540 22718
rect 43260 22372 43316 22382
rect 43148 22370 43316 22372
rect 43148 22318 43262 22370
rect 43314 22318 43316 22370
rect 43148 22316 43316 22318
rect 43260 22306 43316 22316
rect 43372 22258 43428 22270
rect 43372 22206 43374 22258
rect 43426 22206 43428 22258
rect 43372 21924 43428 22206
rect 43372 21858 43428 21868
rect 43036 21534 43038 21586
rect 43090 21534 43092 21586
rect 43036 21522 43092 21534
rect 42588 21422 42590 21474
rect 42642 21422 42644 21474
rect 42588 21410 42644 21422
rect 42924 21364 42980 21374
rect 42700 21362 42980 21364
rect 42700 21310 42926 21362
rect 42978 21310 42980 21362
rect 42700 21308 42980 21310
rect 42700 21252 42756 21308
rect 42924 21298 42980 21308
rect 42140 21196 42756 21252
rect 42028 20972 42532 21028
rect 41804 20862 41806 20914
rect 41858 20862 41860 20914
rect 41804 20850 41860 20862
rect 41580 20626 41636 20636
rect 41692 20802 41748 20814
rect 41692 20750 41694 20802
rect 41746 20750 41748 20802
rect 41244 20244 41300 20254
rect 41356 20244 41412 20300
rect 41244 20242 41412 20244
rect 41244 20190 41246 20242
rect 41298 20190 41412 20242
rect 41244 20188 41412 20190
rect 41468 20580 41524 20590
rect 41244 20178 41300 20188
rect 41468 20132 41524 20524
rect 41020 20066 41076 20076
rect 41356 20076 41524 20132
rect 41580 20132 41636 20142
rect 40908 20018 40964 20030
rect 40908 19966 40910 20018
rect 40962 19966 40964 20018
rect 40908 19684 40964 19966
rect 41132 20020 41188 20030
rect 41132 19926 41188 19964
rect 41356 20018 41412 20076
rect 41580 20020 41636 20076
rect 41356 19966 41358 20018
rect 41410 19966 41412 20018
rect 41356 19954 41412 19966
rect 41468 20018 41636 20020
rect 41468 19966 41582 20018
rect 41634 19966 41636 20018
rect 41468 19964 41636 19966
rect 41468 19796 41524 19964
rect 41580 19954 41636 19964
rect 41468 19730 41524 19740
rect 40908 19236 40964 19628
rect 41020 19236 41076 19246
rect 40908 19180 41020 19236
rect 41020 19170 41076 19180
rect 40572 18946 40628 18956
rect 41132 19012 41188 19022
rect 40908 18452 40964 18462
rect 39900 18338 40068 18340
rect 39900 18286 39902 18338
rect 39954 18286 40068 18338
rect 39900 18284 40068 18286
rect 40236 18338 40292 18350
rect 40236 18286 40238 18338
rect 40290 18286 40292 18338
rect 39900 18274 39956 18284
rect 39900 16994 39956 17006
rect 39900 16942 39902 16994
rect 39954 16942 39956 16994
rect 39900 16660 39956 16942
rect 40236 16772 40292 18286
rect 40348 18228 40404 18238
rect 40348 18134 40404 18172
rect 40908 17778 40964 18396
rect 40908 17726 40910 17778
rect 40962 17726 40964 17778
rect 40908 17714 40964 17726
rect 40236 16706 40292 16716
rect 40348 17108 40404 17118
rect 39900 16594 39956 16604
rect 39900 16236 39956 16248
rect 39788 16212 39844 16222
rect 39900 16212 39902 16236
rect 39844 16184 39902 16212
rect 39954 16184 39956 16236
rect 39844 16156 39956 16184
rect 39788 16146 39844 16156
rect 40236 15874 40292 15886
rect 40236 15822 40238 15874
rect 40290 15822 40292 15874
rect 40012 15540 40068 15550
rect 40236 15540 40292 15822
rect 40068 15484 40292 15540
rect 40012 15446 40068 15484
rect 39900 14532 39956 14542
rect 39900 14438 39956 14476
rect 40236 14530 40292 14542
rect 40236 14478 40238 14530
rect 40290 14478 40292 14530
rect 40236 14084 40292 14478
rect 40236 14018 40292 14028
rect 39676 13654 39732 13692
rect 40124 13636 40180 13646
rect 40124 13542 40180 13580
rect 38892 13022 38894 13074
rect 38946 13022 38948 13074
rect 38892 13010 38948 13022
rect 39228 13356 39396 13412
rect 38220 12962 38500 12964
rect 38220 12910 38222 12962
rect 38274 12910 38500 12962
rect 38220 12908 38500 12910
rect 38220 12898 38276 12908
rect 37772 12126 37774 12178
rect 37826 12126 37828 12178
rect 37548 12068 37604 12078
rect 37548 11974 37604 12012
rect 37660 11396 37716 11406
rect 37660 11282 37716 11340
rect 37772 11394 37828 12126
rect 37996 12178 38052 12190
rect 37996 12126 37998 12178
rect 38050 12126 38052 12178
rect 37772 11342 37774 11394
rect 37826 11342 37828 11394
rect 37772 11330 37828 11342
rect 37884 12066 37940 12078
rect 37884 12014 37886 12066
rect 37938 12014 37940 12066
rect 37660 11230 37662 11282
rect 37714 11230 37716 11282
rect 37660 11218 37716 11230
rect 37660 10836 37716 10846
rect 37660 10742 37716 10780
rect 37884 10724 37940 12014
rect 37996 11396 38052 12126
rect 38668 12180 38724 12190
rect 37996 11330 38052 11340
rect 38444 12068 38500 12078
rect 38444 11394 38500 12012
rect 38668 11508 38724 12124
rect 38444 11342 38446 11394
rect 38498 11342 38500 11394
rect 38444 11330 38500 11342
rect 38556 11452 38724 11508
rect 39004 12178 39060 12190
rect 39004 12126 39006 12178
rect 39058 12126 39060 12178
rect 38220 11170 38276 11182
rect 38220 11118 38222 11170
rect 38274 11118 38276 11170
rect 38220 11060 38276 11118
rect 38220 10994 38276 11004
rect 38332 11172 38388 11182
rect 38556 11172 38612 11452
rect 38332 10834 38388 11116
rect 38332 10782 38334 10834
rect 38386 10782 38388 10834
rect 38332 10770 38388 10782
rect 38444 11116 38612 11172
rect 38668 11282 38724 11294
rect 38668 11230 38670 11282
rect 38722 11230 38724 11282
rect 37436 10668 37604 10724
rect 37436 10500 37492 10510
rect 37324 10498 37492 10500
rect 37324 10446 37438 10498
rect 37490 10446 37492 10498
rect 37324 10444 37492 10446
rect 37436 10434 37492 10444
rect 37548 10276 37604 10668
rect 37884 10658 37940 10668
rect 38220 10724 38276 10734
rect 37996 10610 38052 10622
rect 37996 10558 37998 10610
rect 38050 10558 38052 10610
rect 37884 10388 37940 10398
rect 37996 10388 38052 10558
rect 38220 10612 38276 10668
rect 38332 10612 38388 10622
rect 38220 10610 38388 10612
rect 38220 10558 38334 10610
rect 38386 10558 38388 10610
rect 38220 10556 38388 10558
rect 37884 10386 38052 10388
rect 37884 10334 37886 10386
rect 37938 10334 38052 10386
rect 37884 10332 38052 10334
rect 37884 10322 37940 10332
rect 36428 8194 36484 8204
rect 36092 8036 36148 8046
rect 36652 8036 36708 8316
rect 36988 10050 37268 10052
rect 36988 9998 37214 10050
rect 37266 9998 37268 10050
rect 36988 9996 37268 9998
rect 36988 8258 37044 9996
rect 37212 9986 37268 9996
rect 37436 10220 37604 10276
rect 37100 9604 37156 9614
rect 37100 8596 37156 9548
rect 37100 8530 37156 8540
rect 37212 8372 37268 8382
rect 37212 8278 37268 8316
rect 37436 8372 37492 10220
rect 37548 10050 37604 10062
rect 37548 9998 37550 10050
rect 37602 9998 37604 10050
rect 37548 9938 37604 9998
rect 37548 9886 37550 9938
rect 37602 9886 37604 9938
rect 37548 9874 37604 9886
rect 38332 9940 38388 10556
rect 38332 9874 38388 9884
rect 38444 9828 38500 11116
rect 38668 10610 38724 11230
rect 38668 10558 38670 10610
rect 38722 10558 38724 10610
rect 38668 10276 38724 10558
rect 39004 10500 39060 12126
rect 39228 12178 39284 13356
rect 40012 12850 40068 12862
rect 40012 12798 40014 12850
rect 40066 12798 40068 12850
rect 40012 12404 40068 12798
rect 40124 12740 40180 12750
rect 40124 12646 40180 12684
rect 39564 12348 40068 12404
rect 40236 12628 40292 12638
rect 39228 12126 39230 12178
rect 39282 12126 39284 12178
rect 39228 10834 39284 12126
rect 39452 12180 39508 12190
rect 39564 12180 39620 12348
rect 40124 12292 40180 12302
rect 40236 12292 40292 12572
rect 40124 12290 40292 12292
rect 40124 12238 40126 12290
rect 40178 12238 40292 12290
rect 40124 12236 40292 12238
rect 40124 12226 40180 12236
rect 39508 12124 39620 12180
rect 39676 12180 39732 12190
rect 40012 12180 40068 12190
rect 39676 12178 40068 12180
rect 39676 12126 39678 12178
rect 39730 12126 40014 12178
rect 40066 12126 40068 12178
rect 39676 12124 40068 12126
rect 39452 12086 39508 12124
rect 39676 12114 39732 12124
rect 40012 12114 40068 12124
rect 39340 12066 39396 12078
rect 39340 12014 39342 12066
rect 39394 12014 39396 12066
rect 39340 11620 39396 12014
rect 40348 12068 40404 17052
rect 41132 17106 41188 18956
rect 41692 19012 41748 20750
rect 42140 20690 42196 20702
rect 42140 20638 42142 20690
rect 42194 20638 42196 20690
rect 41804 20356 41860 20366
rect 41860 20300 41972 20356
rect 41804 20290 41860 20300
rect 41916 20130 41972 20300
rect 42140 20244 42196 20638
rect 42140 20178 42196 20188
rect 42252 20578 42308 20590
rect 42252 20526 42254 20578
rect 42306 20526 42308 20578
rect 41916 20078 41918 20130
rect 41970 20078 41972 20130
rect 41916 20066 41972 20078
rect 42028 20020 42084 20030
rect 42028 19348 42084 19964
rect 42140 20020 42196 20030
rect 42252 20020 42308 20526
rect 42364 20580 42420 20590
rect 42364 20486 42420 20524
rect 42140 20018 42420 20020
rect 42140 19966 42142 20018
rect 42194 19966 42420 20018
rect 42140 19964 42420 19966
rect 42140 19954 42196 19964
rect 42028 19346 42196 19348
rect 42028 19294 42030 19346
rect 42082 19294 42196 19346
rect 42028 19292 42196 19294
rect 42028 19282 42084 19292
rect 41692 18946 41748 18956
rect 41692 18338 41748 18350
rect 41692 18286 41694 18338
rect 41746 18286 41748 18338
rect 41468 18228 41524 18238
rect 41692 18228 41748 18286
rect 41524 18172 41748 18228
rect 41468 18162 41524 18172
rect 41132 17054 41134 17106
rect 41186 17054 41188 17106
rect 40908 16884 40964 16894
rect 40572 16882 40964 16884
rect 40572 16830 40910 16882
rect 40962 16830 40964 16882
rect 40572 16828 40964 16830
rect 40572 15986 40628 16828
rect 40908 16818 40964 16828
rect 41020 16772 41076 16782
rect 41020 16678 41076 16716
rect 41132 16210 41188 17054
rect 41580 17668 41636 17678
rect 41580 16996 41636 17612
rect 41916 17108 41972 17118
rect 42140 17108 42196 19292
rect 42364 19236 42420 19964
rect 42476 19906 42532 20972
rect 42924 20916 42980 20926
rect 42924 20822 42980 20860
rect 42812 20692 42868 20702
rect 42812 20598 42868 20636
rect 43372 20578 43428 20590
rect 43372 20526 43374 20578
rect 43426 20526 43428 20578
rect 43372 20020 43428 20526
rect 43372 19926 43428 19964
rect 42476 19854 42478 19906
rect 42530 19854 42532 19906
rect 42476 19842 42532 19854
rect 42588 19908 42644 19918
rect 42588 19458 42644 19852
rect 42588 19406 42590 19458
rect 42642 19406 42644 19458
rect 42588 19394 42644 19406
rect 42364 19180 42868 19236
rect 42812 19122 42868 19180
rect 42812 19070 42814 19122
rect 42866 19070 42868 19122
rect 42812 19058 42868 19070
rect 43260 19122 43316 19134
rect 43260 19070 43262 19122
rect 43314 19070 43316 19122
rect 42700 19012 42756 19022
rect 42700 18918 42756 18956
rect 43260 18676 43316 19070
rect 43260 18610 43316 18620
rect 43484 18564 43540 22652
rect 43372 18508 43540 18564
rect 43372 17666 43428 18508
rect 43596 18340 43652 23548
rect 43708 23492 43764 23502
rect 43708 22484 43764 23436
rect 44268 22932 44324 23662
rect 44940 23604 44996 25340
rect 44940 23538 44996 23548
rect 45052 24610 45108 25564
rect 45164 25508 45220 26236
rect 45164 25442 45220 25452
rect 45276 26066 45332 26078
rect 45276 26014 45278 26066
rect 45330 26014 45332 26066
rect 45052 24558 45054 24610
rect 45106 24558 45108 24610
rect 45052 23828 45108 24558
rect 45276 24276 45332 26014
rect 45388 25506 45444 27020
rect 45948 26962 46004 26974
rect 45948 26910 45950 26962
rect 46002 26910 46004 26962
rect 45948 26908 46004 26910
rect 45836 26852 46004 26908
rect 46060 26908 46116 28588
rect 46284 26908 46340 31724
rect 47404 31778 47460 31790
rect 47404 31726 47406 31778
rect 47458 31726 47460 31778
rect 46396 31666 46452 31678
rect 46396 31614 46398 31666
rect 46450 31614 46452 31666
rect 46396 31220 46452 31614
rect 46844 31668 46900 31678
rect 46844 31574 46900 31612
rect 46508 31556 46564 31566
rect 46508 31462 46564 31500
rect 46956 31554 47012 31566
rect 46956 31502 46958 31554
rect 47010 31502 47012 31554
rect 46396 31154 46452 31164
rect 46956 30212 47012 31502
rect 47180 31556 47236 31566
rect 47180 31106 47236 31500
rect 47404 31444 47460 31726
rect 47404 31378 47460 31388
rect 47180 31054 47182 31106
rect 47234 31054 47236 31106
rect 47180 31042 47236 31054
rect 47404 30212 47460 30222
rect 46956 30210 47460 30212
rect 46956 30158 47406 30210
rect 47458 30158 47460 30210
rect 46956 30156 47460 30158
rect 47404 30146 47460 30156
rect 47628 28754 47684 31948
rect 47852 30996 47908 33068
rect 47964 33126 47966 33178
rect 48018 33126 48020 33178
rect 48076 33182 48078 33234
rect 48130 33182 48244 33234
rect 48076 33180 48244 33182
rect 48076 33170 48132 33180
rect 47964 33012 48020 33126
rect 47964 32946 48020 32956
rect 48076 32674 48132 32686
rect 48076 32622 48078 32674
rect 48130 32622 48132 32674
rect 47964 31554 48020 31566
rect 47964 31502 47966 31554
rect 48018 31502 48020 31554
rect 47964 31220 48020 31502
rect 48076 31220 48132 32622
rect 48188 32562 48244 33180
rect 48300 32676 48356 35868
rect 48300 32610 48356 32620
rect 48188 32510 48190 32562
rect 48242 32510 48244 32562
rect 48188 32498 48244 32510
rect 48524 31892 48580 31902
rect 47964 31164 48356 31220
rect 47964 30996 48020 31006
rect 47852 30994 48020 30996
rect 47852 30942 47966 30994
rect 48018 30942 48020 30994
rect 47852 30940 48020 30942
rect 47964 30212 48020 30940
rect 48076 30212 48132 30222
rect 47964 30210 48132 30212
rect 47964 30158 48078 30210
rect 48130 30158 48132 30210
rect 47964 30156 48132 30158
rect 48076 30146 48132 30156
rect 48188 29316 48244 29326
rect 47628 28702 47630 28754
rect 47682 28702 47684 28754
rect 47628 28690 47684 28702
rect 48076 29314 48244 29316
rect 48076 29262 48190 29314
rect 48242 29262 48244 29314
rect 48076 29260 48244 29262
rect 47404 28644 47460 28654
rect 47404 28550 47460 28588
rect 48076 28084 48132 29260
rect 48188 29250 48244 29260
rect 48076 28018 48132 28028
rect 48188 28644 48244 28654
rect 48188 27412 48244 28588
rect 48188 27346 48244 27356
rect 48076 27186 48132 27198
rect 48076 27134 48078 27186
rect 48130 27134 48132 27186
rect 47628 26964 47684 26974
rect 48076 26908 48132 27134
rect 46060 26852 46228 26908
rect 46284 26852 46452 26908
rect 45836 26516 45892 26852
rect 45836 26450 45892 26460
rect 45388 25454 45390 25506
rect 45442 25454 45444 25506
rect 45388 25442 45444 25454
rect 46060 25396 46116 25406
rect 45948 25394 46116 25396
rect 45948 25342 46062 25394
rect 46114 25342 46116 25394
rect 45948 25340 46116 25342
rect 45948 24946 46004 25340
rect 46060 25330 46116 25340
rect 45948 24894 45950 24946
rect 46002 24894 46004 24946
rect 45948 24882 46004 24894
rect 46060 24836 46116 24846
rect 46172 24836 46228 26852
rect 46060 24834 46228 24836
rect 46060 24782 46062 24834
rect 46114 24782 46228 24834
rect 46060 24780 46228 24782
rect 45500 24612 45556 24622
rect 45836 24612 45892 24622
rect 45500 24610 45892 24612
rect 45500 24558 45502 24610
rect 45554 24558 45838 24610
rect 45890 24558 45892 24610
rect 45500 24556 45892 24558
rect 45500 24546 45556 24556
rect 45836 24546 45892 24556
rect 45164 24220 45332 24276
rect 45164 23828 45220 24220
rect 45276 24052 45332 24062
rect 45276 24050 45444 24052
rect 45276 23998 45278 24050
rect 45330 23998 45444 24050
rect 45276 23996 45444 23998
rect 45276 23986 45332 23996
rect 45388 23940 45444 23996
rect 45164 23772 45332 23828
rect 44492 23492 44548 23502
rect 44492 23378 44548 23436
rect 44492 23326 44494 23378
rect 44546 23326 44548 23378
rect 44492 23314 44548 23326
rect 44940 23268 44996 23278
rect 45052 23268 45108 23772
rect 44940 23266 45108 23268
rect 44940 23214 44942 23266
rect 44994 23214 45108 23266
rect 44940 23212 45108 23214
rect 45164 23604 45220 23614
rect 44940 23202 44996 23212
rect 45164 23154 45220 23548
rect 45164 23102 45166 23154
rect 45218 23102 45220 23154
rect 45164 23090 45220 23102
rect 45052 23044 45108 23054
rect 45052 22950 45108 22988
rect 43932 22876 44268 22932
rect 43932 22594 43988 22876
rect 44268 22838 44324 22876
rect 44604 22932 44660 22942
rect 44604 22930 44996 22932
rect 44604 22878 44606 22930
rect 44658 22878 44996 22930
rect 44604 22876 44996 22878
rect 44604 22866 44660 22876
rect 43932 22542 43934 22594
rect 43986 22542 43988 22594
rect 43932 22530 43988 22542
rect 43708 22390 43764 22428
rect 44268 22146 44324 22158
rect 44268 22094 44270 22146
rect 44322 22094 44324 22146
rect 44268 21476 44324 22094
rect 44492 21700 44548 21710
rect 43932 21420 44268 21476
rect 43932 21026 43988 21420
rect 44268 21410 44324 21420
rect 44380 21644 44492 21700
rect 44268 21028 44324 21038
rect 44380 21028 44436 21644
rect 44492 21606 44548 21644
rect 44604 21700 44660 21710
rect 44604 21698 44772 21700
rect 44604 21646 44606 21698
rect 44658 21646 44772 21698
rect 44604 21644 44772 21646
rect 44604 21634 44660 21644
rect 43932 20974 43934 21026
rect 43986 20974 43988 21026
rect 43932 20962 43988 20974
rect 44156 21026 44436 21028
rect 44156 20974 44270 21026
rect 44322 20974 44436 21026
rect 44156 20972 44436 20974
rect 43708 20916 43764 20926
rect 43708 20822 43764 20860
rect 44156 19346 44212 20972
rect 44268 20962 44324 20972
rect 44716 19684 44772 21644
rect 44828 21588 44884 21598
rect 44940 21588 44996 22876
rect 45276 22708 45332 23772
rect 45388 23154 45444 23884
rect 46060 23268 46116 24780
rect 46396 24052 46452 26852
rect 47628 26852 48132 26908
rect 48188 27188 48244 27198
rect 47628 26402 47684 26852
rect 47628 26350 47630 26402
rect 47682 26350 47684 26402
rect 47628 26338 47684 26350
rect 48076 26404 48132 26414
rect 48188 26404 48244 27132
rect 48076 26402 48244 26404
rect 48076 26350 48078 26402
rect 48130 26350 48244 26402
rect 48076 26348 48244 26350
rect 48076 26338 48132 26348
rect 46508 26292 46564 26302
rect 46508 26198 46564 26236
rect 46620 26292 46676 26302
rect 46956 26292 47012 26302
rect 46620 26290 47012 26292
rect 46620 26238 46622 26290
rect 46674 26238 46958 26290
rect 47010 26238 47012 26290
rect 46620 26236 47012 26238
rect 46620 26226 46676 26236
rect 46956 26226 47012 26236
rect 47180 26290 47236 26302
rect 47180 26238 47182 26290
rect 47234 26238 47236 26290
rect 47068 26178 47124 26190
rect 47068 26126 47070 26178
rect 47122 26126 47124 26178
rect 47068 25844 47124 26126
rect 47068 25778 47124 25788
rect 47180 25396 47236 26238
rect 47404 26292 47460 26302
rect 47404 26290 47572 26292
rect 47404 26238 47406 26290
rect 47458 26238 47572 26290
rect 47404 26236 47572 26238
rect 47404 26226 47460 26236
rect 47516 26180 47572 26236
rect 47964 26180 48020 26190
rect 47516 26178 48020 26180
rect 47516 26126 47966 26178
rect 48018 26126 48020 26178
rect 47516 26124 48020 26126
rect 47964 26114 48020 26124
rect 47180 25330 47236 25340
rect 48188 25618 48244 25630
rect 48188 25566 48190 25618
rect 48242 25566 48244 25618
rect 48188 25396 48244 25566
rect 48188 25330 48244 25340
rect 48300 25172 48356 31164
rect 47852 25116 48356 25172
rect 46396 23996 46564 24052
rect 46060 23202 46116 23212
rect 46396 23828 46452 23838
rect 46396 23266 46452 23772
rect 46396 23214 46398 23266
rect 46450 23214 46452 23266
rect 46396 23202 46452 23214
rect 45388 23102 45390 23154
rect 45442 23102 45444 23154
rect 45388 23090 45444 23102
rect 45836 23154 45892 23166
rect 45836 23102 45838 23154
rect 45890 23102 45892 23154
rect 45836 23044 45892 23102
rect 45836 22978 45892 22988
rect 46060 22932 46116 22942
rect 46060 22838 46116 22876
rect 46284 22930 46340 22942
rect 46284 22878 46286 22930
rect 46338 22878 46340 22930
rect 45276 22642 45332 22652
rect 45276 22484 45332 22494
rect 45276 22390 45332 22428
rect 45612 22260 45668 22270
rect 45388 21924 45444 21934
rect 45052 21588 45108 21598
rect 44940 21586 45108 21588
rect 44940 21534 45054 21586
rect 45106 21534 45108 21586
rect 44940 21532 45108 21534
rect 44828 21494 44884 21532
rect 45052 21522 45108 21532
rect 45276 21476 45332 21486
rect 45276 21382 45332 21420
rect 45388 20802 45444 21868
rect 45500 21812 45556 21822
rect 45500 21586 45556 21756
rect 45612 21698 45668 22204
rect 45612 21646 45614 21698
rect 45666 21646 45668 21698
rect 45612 21634 45668 21646
rect 46060 21812 46116 21822
rect 46284 21812 46340 22878
rect 46116 21756 46340 21812
rect 45500 21534 45502 21586
rect 45554 21534 45556 21586
rect 45500 21522 45556 21534
rect 46060 21586 46116 21756
rect 46060 21534 46062 21586
rect 46114 21534 46116 21586
rect 46060 21522 46116 21534
rect 46396 21700 46452 21710
rect 46396 21586 46452 21644
rect 46396 21534 46398 21586
rect 46450 21534 46452 21586
rect 46396 21522 46452 21534
rect 45948 21362 46004 21374
rect 45948 21310 45950 21362
rect 46002 21310 46004 21362
rect 45948 20916 46004 21310
rect 46284 21364 46340 21374
rect 46284 21270 46340 21308
rect 46060 20916 46116 20926
rect 45948 20914 46116 20916
rect 45948 20862 46062 20914
rect 46114 20862 46116 20914
rect 45948 20860 46116 20862
rect 46060 20850 46116 20860
rect 45388 20750 45390 20802
rect 45442 20750 45444 20802
rect 44716 19628 44996 19684
rect 44156 19294 44158 19346
rect 44210 19294 44212 19346
rect 44156 19282 44212 19294
rect 44940 19348 44996 19628
rect 44940 19346 45108 19348
rect 44940 19294 44942 19346
rect 44994 19294 45108 19346
rect 44940 19292 45108 19294
rect 44940 19282 44996 19292
rect 43932 19236 43988 19246
rect 43932 19142 43988 19180
rect 44828 19236 44884 19246
rect 44828 19142 44884 19180
rect 43372 17614 43374 17666
rect 43426 17614 43428 17666
rect 43372 17602 43428 17614
rect 43484 18284 43652 18340
rect 43708 18452 43764 18462
rect 43484 17444 43540 18284
rect 43596 17892 43652 17902
rect 43596 17778 43652 17836
rect 43708 17890 43764 18396
rect 44268 18450 44324 18462
rect 44268 18398 44270 18450
rect 44322 18398 44324 18450
rect 43708 17838 43710 17890
rect 43762 17838 43764 17890
rect 43708 17826 43764 17838
rect 43820 18338 43876 18350
rect 43820 18286 43822 18338
rect 43874 18286 43876 18338
rect 43596 17726 43598 17778
rect 43650 17726 43652 17778
rect 43596 17714 43652 17726
rect 43820 17668 43876 18286
rect 43820 17602 43876 17612
rect 44156 17554 44212 17566
rect 44156 17502 44158 17554
rect 44210 17502 44212 17554
rect 44044 17444 44100 17454
rect 43260 17388 43540 17444
rect 43708 17442 44100 17444
rect 43708 17390 44046 17442
rect 44098 17390 44100 17442
rect 43708 17388 44100 17390
rect 42588 17108 42644 17118
rect 41972 17106 42980 17108
rect 41972 17054 42142 17106
rect 42194 17054 42590 17106
rect 42642 17054 42980 17106
rect 41972 17052 42980 17054
rect 41916 17042 41972 17052
rect 42140 17042 42196 17052
rect 42588 17042 42644 17052
rect 41580 16994 41860 16996
rect 41580 16942 41582 16994
rect 41634 16942 41860 16994
rect 41580 16940 41860 16942
rect 41580 16930 41636 16940
rect 41356 16882 41412 16894
rect 41356 16830 41358 16882
rect 41410 16830 41412 16882
rect 41356 16660 41412 16830
rect 41356 16436 41412 16604
rect 41356 16380 41636 16436
rect 41132 16158 41134 16210
rect 41186 16158 41188 16210
rect 41132 16146 41188 16158
rect 41356 16210 41412 16222
rect 41356 16158 41358 16210
rect 41410 16158 41412 16210
rect 40572 15934 40574 15986
rect 40626 15934 40628 15986
rect 40572 14756 40628 15934
rect 40908 15204 40964 15242
rect 40908 15138 40964 15148
rect 40572 14690 40628 14700
rect 41356 14644 41412 16158
rect 41356 14578 41412 14588
rect 41468 15204 41524 15214
rect 40460 14532 40516 14542
rect 40460 14438 40516 14476
rect 40796 14420 40852 14430
rect 41132 14420 41188 14430
rect 40796 14418 41188 14420
rect 40796 14366 40798 14418
rect 40850 14366 41134 14418
rect 41186 14366 41188 14418
rect 40796 14364 41188 14366
rect 40796 14354 40852 14364
rect 41132 14354 41188 14364
rect 41468 14418 41524 15148
rect 41580 14532 41636 16380
rect 41580 14466 41636 14476
rect 41468 14366 41470 14418
rect 41522 14366 41524 14418
rect 41468 14354 41524 14366
rect 41692 14308 41748 14318
rect 41020 14084 41076 14094
rect 41020 13970 41076 14028
rect 41020 13918 41022 13970
rect 41074 13918 41076 13970
rect 41020 13906 41076 13918
rect 41692 13634 41748 14252
rect 41692 13582 41694 13634
rect 41746 13582 41748 13634
rect 40460 13076 40516 13086
rect 40460 12982 40516 13020
rect 40572 12964 40628 12974
rect 40572 12962 41412 12964
rect 40572 12910 40574 12962
rect 40626 12910 41412 12962
rect 40572 12908 41412 12910
rect 40572 12898 40628 12908
rect 40908 12740 40964 12750
rect 40908 12178 40964 12684
rect 41132 12628 41188 12638
rect 41132 12402 41188 12572
rect 41132 12350 41134 12402
rect 41186 12350 41188 12402
rect 41132 12338 41188 12350
rect 41356 12402 41412 12908
rect 41356 12350 41358 12402
rect 41410 12350 41412 12402
rect 41356 12338 41412 12350
rect 40908 12126 40910 12178
rect 40962 12126 40964 12178
rect 40908 12114 40964 12126
rect 41580 12178 41636 12190
rect 41580 12126 41582 12178
rect 41634 12126 41636 12178
rect 40348 12012 40740 12068
rect 39340 11564 39956 11620
rect 39340 11396 39396 11406
rect 39340 11302 39396 11340
rect 39788 11396 39844 11406
rect 39228 10782 39230 10834
rect 39282 10782 39284 10834
rect 39228 10770 39284 10782
rect 39788 10834 39844 11340
rect 39788 10782 39790 10834
rect 39842 10782 39844 10834
rect 39788 10770 39844 10782
rect 39900 10724 39956 11564
rect 40236 11284 40292 11294
rect 40236 11190 40292 11228
rect 40124 11172 40180 11182
rect 40124 11078 40180 11116
rect 40348 11170 40404 11182
rect 40348 11118 40350 11170
rect 40402 11118 40404 11170
rect 40348 10948 40404 11118
rect 40348 10892 40628 10948
rect 40236 10724 40292 10734
rect 39900 10722 40292 10724
rect 39900 10670 39902 10722
rect 39954 10670 40238 10722
rect 40290 10670 40292 10722
rect 39900 10668 40292 10670
rect 39900 10658 39956 10668
rect 40236 10658 40292 10668
rect 39564 10612 39620 10622
rect 40572 10612 40628 10892
rect 40684 10724 40740 12012
rect 41020 12066 41076 12078
rect 41020 12014 41022 12066
rect 41074 12014 41076 12066
rect 41020 11508 41076 12014
rect 41580 12068 41636 12126
rect 41580 12002 41636 12012
rect 40796 11452 41076 11508
rect 40796 11396 40852 11452
rect 40796 11302 40852 11340
rect 40684 10658 40740 10668
rect 40908 11284 40964 11294
rect 40908 10722 40964 11228
rect 41020 11060 41076 11070
rect 41076 11004 41188 11060
rect 41020 10994 41076 11004
rect 40908 10670 40910 10722
rect 40962 10670 40964 10722
rect 40908 10658 40964 10670
rect 39452 10610 39620 10612
rect 39452 10558 39566 10610
rect 39618 10558 39620 10610
rect 39452 10556 39620 10558
rect 39004 10406 39060 10444
rect 39116 10498 39172 10510
rect 39116 10446 39118 10498
rect 39170 10446 39172 10498
rect 39116 10276 39172 10446
rect 38668 10220 39172 10276
rect 39340 10052 39396 10062
rect 39452 10052 39508 10556
rect 39564 10546 39620 10556
rect 40460 10556 40628 10612
rect 40348 10500 40404 10510
rect 40460 10500 40516 10556
rect 40348 10498 40516 10500
rect 40348 10446 40350 10498
rect 40402 10446 40516 10498
rect 40348 10444 40516 10446
rect 41020 10498 41076 10510
rect 41020 10446 41022 10498
rect 41074 10446 41076 10498
rect 40348 10434 40404 10444
rect 39340 10050 39508 10052
rect 39340 9998 39342 10050
rect 39394 9998 39508 10050
rect 39340 9996 39508 9998
rect 39340 9986 39396 9996
rect 38892 9940 38948 9950
rect 41020 9940 41076 10446
rect 38892 9846 38948 9884
rect 40908 9884 41076 9940
rect 38444 8932 38500 9772
rect 39116 9828 39172 9838
rect 40796 9828 40852 9838
rect 39116 9826 39620 9828
rect 39116 9774 39118 9826
rect 39170 9774 39620 9826
rect 39116 9772 39620 9774
rect 39116 9762 39172 9772
rect 39564 9266 39620 9772
rect 40236 9826 40852 9828
rect 40236 9774 40798 9826
rect 40850 9774 40852 9826
rect 40236 9772 40852 9774
rect 39564 9214 39566 9266
rect 39618 9214 39620 9266
rect 39564 9202 39620 9214
rect 39788 9602 39844 9614
rect 39788 9550 39790 9602
rect 39842 9550 39844 9602
rect 39676 9044 39732 9054
rect 39676 8950 39732 8988
rect 38556 8932 38612 8942
rect 38444 8930 38612 8932
rect 38444 8878 38558 8930
rect 38610 8878 38612 8930
rect 38444 8876 38612 8878
rect 38556 8866 38612 8876
rect 38668 8596 38724 8606
rect 37436 8278 37492 8316
rect 38332 8372 38388 8382
rect 36988 8206 36990 8258
rect 37042 8206 37044 8258
rect 36988 8194 37044 8206
rect 37660 8148 37716 8158
rect 37660 8054 37716 8092
rect 37884 8148 37940 8158
rect 37884 8054 37940 8092
rect 36092 8034 36708 8036
rect 36092 7982 36094 8034
rect 36146 7982 36708 8034
rect 36092 7980 36708 7982
rect 37548 8034 37604 8046
rect 37548 7982 37550 8034
rect 37602 7982 37604 8034
rect 36092 7970 36148 7980
rect 37548 7700 37604 7982
rect 37548 7644 37828 7700
rect 37660 7474 37716 7486
rect 37660 7422 37662 7474
rect 37714 7422 37716 7474
rect 37660 7364 37716 7422
rect 37660 6804 37716 7308
rect 37660 6738 37716 6748
rect 37772 6802 37828 7644
rect 38332 7140 38388 8316
rect 38332 7074 38388 7084
rect 37772 6750 37774 6802
rect 37826 6750 37828 6802
rect 37772 6738 37828 6750
rect 36988 6692 37044 6702
rect 36988 6598 37044 6636
rect 36092 6580 36148 6590
rect 36092 6018 36148 6524
rect 38668 6130 38724 8540
rect 39788 8372 39844 9550
rect 40236 9266 40292 9772
rect 40796 9762 40852 9772
rect 40236 9214 40238 9266
rect 40290 9214 40292 9266
rect 40236 9202 40292 9214
rect 40908 9266 40964 9884
rect 41020 9716 41076 9726
rect 41132 9716 41188 11004
rect 41468 10836 41524 10846
rect 41468 10722 41524 10780
rect 41468 10670 41470 10722
rect 41522 10670 41524 10722
rect 41468 10658 41524 10670
rect 41244 10610 41300 10622
rect 41244 10558 41246 10610
rect 41298 10558 41300 10610
rect 41244 10388 41300 10558
rect 41580 10388 41636 10398
rect 41244 10386 41636 10388
rect 41244 10334 41582 10386
rect 41634 10334 41636 10386
rect 41244 10332 41636 10334
rect 41580 10322 41636 10332
rect 41692 10164 41748 13582
rect 41804 13076 41860 16940
rect 42924 16882 42980 17052
rect 42924 16830 42926 16882
rect 42978 16830 42980 16882
rect 42924 16818 42980 16830
rect 42588 16660 42644 16670
rect 42588 14644 42644 16604
rect 43036 15204 43092 15242
rect 43036 15138 43092 15148
rect 42140 14642 42644 14644
rect 42140 14590 42590 14642
rect 42642 14590 42644 14642
rect 42140 14588 42644 14590
rect 42028 14308 42084 14318
rect 42028 14214 42084 14252
rect 42140 14084 42196 14588
rect 42588 14578 42644 14588
rect 42924 14644 42980 14654
rect 42924 14530 42980 14588
rect 42924 14478 42926 14530
rect 42978 14478 42980 14530
rect 42924 14466 42980 14478
rect 43148 14532 43204 14542
rect 43148 14438 43204 14476
rect 42028 14028 42196 14084
rect 41804 12740 41860 13020
rect 41804 12674 41860 12684
rect 41916 13188 41972 13198
rect 41916 12962 41972 13132
rect 41916 12910 41918 12962
rect 41970 12910 41972 12962
rect 41916 12628 41972 12910
rect 41916 12562 41972 12572
rect 41916 12404 41972 12414
rect 41804 11170 41860 11182
rect 41804 11118 41806 11170
rect 41858 11118 41860 11170
rect 41804 10612 41860 11118
rect 41804 10546 41860 10556
rect 41804 10388 41860 10398
rect 41916 10388 41972 12348
rect 42028 11060 42084 14028
rect 42588 13972 42644 13982
rect 43260 13972 43316 17388
rect 43708 16884 43764 17388
rect 44044 17378 44100 17388
rect 43484 16828 43764 16884
rect 43372 16324 43428 16334
rect 43372 14642 43428 16268
rect 43484 16210 43540 16828
rect 44156 16324 44212 17502
rect 44156 16258 44212 16268
rect 44268 16772 44324 18398
rect 44940 18338 44996 18350
rect 44940 18286 44942 18338
rect 44994 18286 44996 18338
rect 44940 17892 44996 18286
rect 45052 18340 45108 19292
rect 45388 19234 45444 20750
rect 46172 20468 46228 20478
rect 46060 20412 46172 20468
rect 46060 19346 46116 20412
rect 46172 20402 46228 20412
rect 46508 20244 46564 23996
rect 47404 23828 47460 23838
rect 47404 23734 47460 23772
rect 47852 23378 47908 25116
rect 47852 23326 47854 23378
rect 47906 23326 47908 23378
rect 47852 23314 47908 23326
rect 48076 23938 48132 23950
rect 48076 23886 48078 23938
rect 48130 23886 48132 23938
rect 47292 23268 47348 23278
rect 46732 21588 46788 21598
rect 46732 21494 46788 21532
rect 47180 21586 47236 21598
rect 47180 21534 47182 21586
rect 47234 21534 47236 21586
rect 46956 21474 47012 21486
rect 46956 21422 46958 21474
rect 47010 21422 47012 21474
rect 46956 20468 47012 21422
rect 46956 20402 47012 20412
rect 47180 20580 47236 21534
rect 47292 21586 47348 23212
rect 47628 23044 47684 23054
rect 47628 22950 47684 22988
rect 48076 22370 48132 23886
rect 48188 23154 48244 23166
rect 48188 23102 48190 23154
rect 48242 23102 48244 23154
rect 48188 23044 48244 23102
rect 48188 22484 48244 22988
rect 48188 22418 48244 22428
rect 48076 22318 48078 22370
rect 48130 22318 48132 22370
rect 47404 22260 47460 22270
rect 47404 22166 47460 22204
rect 48076 21924 48132 22318
rect 48076 21858 48132 21868
rect 47964 21812 48020 21822
rect 47964 21718 48020 21756
rect 48188 21812 48244 21822
rect 47292 21534 47294 21586
rect 47346 21534 47348 21586
rect 47292 21522 47348 21534
rect 47740 21476 47796 21486
rect 47740 21382 47796 21420
rect 47852 21474 47908 21486
rect 47852 21422 47854 21474
rect 47906 21422 47908 21474
rect 47852 21364 47908 21422
rect 47852 21298 47908 21308
rect 48188 20916 48244 21756
rect 48188 20822 48244 20860
rect 46508 20188 47012 20244
rect 46060 19294 46062 19346
rect 46114 19294 46116 19346
rect 46060 19282 46116 19294
rect 46844 19906 46900 19918
rect 46844 19854 46846 19906
rect 46898 19854 46900 19906
rect 45388 19182 45390 19234
rect 45442 19182 45444 19234
rect 45388 18452 45444 19182
rect 45388 18386 45444 18396
rect 46844 18452 46900 19854
rect 46844 18386 46900 18396
rect 45052 18274 45108 18284
rect 44940 17826 44996 17836
rect 45612 17780 45668 17790
rect 45276 17666 45332 17678
rect 45276 17614 45278 17666
rect 45330 17614 45332 17666
rect 44940 16772 44996 16782
rect 44268 16770 44996 16772
rect 44268 16718 44942 16770
rect 44994 16718 44996 16770
rect 44268 16716 44996 16718
rect 43484 16158 43486 16210
rect 43538 16158 43540 16210
rect 43484 16146 43540 16158
rect 44268 16100 44324 16716
rect 44940 16706 44996 16716
rect 44940 16212 44996 16222
rect 45276 16212 45332 17614
rect 45612 17666 45668 17724
rect 45724 17780 45780 17790
rect 46172 17780 46228 17790
rect 45724 17778 46228 17780
rect 45724 17726 45726 17778
rect 45778 17726 46174 17778
rect 46226 17726 46228 17778
rect 45724 17724 46228 17726
rect 45724 17714 45780 17724
rect 46172 17714 46228 17724
rect 45612 17614 45614 17666
rect 45666 17614 45668 17666
rect 45612 17602 45668 17614
rect 46620 17554 46676 17566
rect 46620 17502 46622 17554
rect 46674 17502 46676 17554
rect 44940 16210 45332 16212
rect 44940 16158 44942 16210
rect 44994 16158 45278 16210
rect 45330 16158 45332 16210
rect 44940 16156 45332 16158
rect 44940 16146 44996 16156
rect 45276 16146 45332 16156
rect 45388 17442 45444 17454
rect 45388 17390 45390 17442
rect 45442 17390 45444 17442
rect 43820 16098 44324 16100
rect 43820 16046 44270 16098
rect 44322 16046 44324 16098
rect 43820 16044 44324 16046
rect 43820 15314 43876 16044
rect 44268 16034 44324 16044
rect 44828 15876 44884 15886
rect 44828 15782 44884 15820
rect 43820 15262 43822 15314
rect 43874 15262 43876 15314
rect 43820 15250 43876 15262
rect 44716 15202 44772 15214
rect 44716 15150 44718 15202
rect 44770 15150 44772 15202
rect 44716 15148 44772 15150
rect 45276 15202 45332 15214
rect 45276 15150 45278 15202
rect 45330 15150 45332 15202
rect 45276 15148 45332 15150
rect 44604 15092 44660 15102
rect 44716 15092 45332 15148
rect 44380 15090 44660 15092
rect 44380 15038 44606 15090
rect 44658 15038 44660 15090
rect 44380 15036 44660 15038
rect 43372 14590 43374 14642
rect 43426 14590 43428 14642
rect 43372 14578 43428 14590
rect 43484 14756 43540 14766
rect 43484 14530 43540 14700
rect 43484 14478 43486 14530
rect 43538 14478 43540 14530
rect 43484 14466 43540 14478
rect 43596 14644 43652 14654
rect 43372 14306 43428 14318
rect 43372 14254 43374 14306
rect 43426 14254 43428 14306
rect 43372 13972 43428 14254
rect 42588 13970 43428 13972
rect 42588 13918 42590 13970
rect 42642 13918 43428 13970
rect 42588 13916 43428 13918
rect 42588 13906 42644 13916
rect 42812 13748 42868 13758
rect 42700 13692 42812 13748
rect 42476 13636 42532 13646
rect 42476 12962 42532 13580
rect 42476 12910 42478 12962
rect 42530 12910 42532 12962
rect 42476 12898 42532 12910
rect 42588 13524 42644 13534
rect 42140 12738 42196 12750
rect 42140 12686 42142 12738
rect 42194 12686 42196 12738
rect 42140 12628 42196 12686
rect 42140 12562 42196 12572
rect 42252 12740 42308 12750
rect 42252 12402 42308 12684
rect 42252 12350 42254 12402
rect 42306 12350 42308 12402
rect 42252 12338 42308 12350
rect 42476 12404 42532 12414
rect 42476 12310 42532 12348
rect 42252 12180 42308 12190
rect 42140 12068 42196 12078
rect 42140 11506 42196 12012
rect 42252 11618 42308 12124
rect 42252 11566 42254 11618
rect 42306 11566 42308 11618
rect 42252 11554 42308 11566
rect 42140 11454 42142 11506
rect 42194 11454 42196 11506
rect 42140 11442 42196 11454
rect 42140 11060 42196 11070
rect 42588 11060 42644 13468
rect 42700 12962 42756 13692
rect 42812 13654 42868 13692
rect 43372 13748 43428 13758
rect 43036 13636 43092 13646
rect 43092 13580 43204 13636
rect 43036 13542 43092 13580
rect 42700 12910 42702 12962
rect 42754 12910 42756 12962
rect 42700 12628 42756 12910
rect 42700 12562 42756 12572
rect 42812 12964 42868 12974
rect 42700 12180 42756 12190
rect 42812 12180 42868 12908
rect 42756 12124 42868 12180
rect 42924 12738 42980 12750
rect 42924 12686 42926 12738
rect 42978 12686 42980 12738
rect 42700 12086 42756 12124
rect 42924 12068 42980 12686
rect 43036 12740 43092 12778
rect 43036 12674 43092 12684
rect 42812 12012 42924 12068
rect 42700 11394 42756 11406
rect 42700 11342 42702 11394
rect 42754 11342 42756 11394
rect 42700 11284 42756 11342
rect 42812 11394 42868 12012
rect 42924 12002 42980 12012
rect 43036 12516 43092 12526
rect 42812 11342 42814 11394
rect 42866 11342 42868 11394
rect 42812 11330 42868 11342
rect 42700 11218 42756 11228
rect 43036 11282 43092 12460
rect 43148 11394 43204 13580
rect 43372 13634 43428 13692
rect 43372 13582 43374 13634
rect 43426 13582 43428 13634
rect 43372 13570 43428 13582
rect 43596 13188 43652 14588
rect 43932 14420 43988 14430
rect 43708 14418 43988 14420
rect 43708 14366 43934 14418
rect 43986 14366 43988 14418
rect 43708 14364 43988 14366
rect 43708 13636 43764 14364
rect 43932 14354 43988 14364
rect 44044 14306 44100 14318
rect 44044 14254 44046 14306
rect 44098 14254 44100 14306
rect 44044 13972 44100 14254
rect 44044 13906 44100 13916
rect 44268 14306 44324 14318
rect 44268 14254 44270 14306
rect 44322 14254 44324 14306
rect 43708 13570 43764 13580
rect 43820 13746 43876 13758
rect 43820 13694 43822 13746
rect 43874 13694 43876 13746
rect 43820 13524 43876 13694
rect 43932 13748 43988 13758
rect 43932 13654 43988 13692
rect 44044 13748 44100 13758
rect 44268 13748 44324 14254
rect 44044 13746 44324 13748
rect 44044 13694 44046 13746
rect 44098 13694 44324 13746
rect 44044 13692 44324 13694
rect 43820 13458 43876 13468
rect 43148 11342 43150 11394
rect 43202 11342 43204 11394
rect 43148 11330 43204 11342
rect 43484 13132 43652 13188
rect 43484 12178 43540 13132
rect 43596 12964 43652 12974
rect 43596 12870 43652 12908
rect 44044 12962 44100 13692
rect 44044 12910 44046 12962
rect 44098 12910 44100 12962
rect 44044 12898 44100 12910
rect 44268 12964 44324 12974
rect 44268 12870 44324 12908
rect 44268 12740 44324 12750
rect 43596 12292 43652 12302
rect 43596 12290 43988 12292
rect 43596 12238 43598 12290
rect 43650 12238 43988 12290
rect 43596 12236 43988 12238
rect 43596 12226 43652 12236
rect 43484 12126 43486 12178
rect 43538 12126 43540 12178
rect 43036 11230 43038 11282
rect 43090 11230 43092 11282
rect 43036 11218 43092 11230
rect 42028 11004 42140 11060
rect 42140 10994 42196 11004
rect 42364 11004 42644 11060
rect 42028 10836 42084 10846
rect 42028 10742 42084 10780
rect 41804 10386 41972 10388
rect 41804 10334 41806 10386
rect 41858 10334 41972 10386
rect 41804 10332 41972 10334
rect 41804 10322 41860 10332
rect 41692 10098 41748 10108
rect 41580 10050 41636 10062
rect 41580 9998 41582 10050
rect 41634 9998 41636 10050
rect 41020 9714 41188 9716
rect 41020 9662 41022 9714
rect 41074 9662 41188 9714
rect 41020 9660 41188 9662
rect 41468 9826 41524 9838
rect 41468 9774 41470 9826
rect 41522 9774 41524 9826
rect 41020 9650 41076 9660
rect 41468 9604 41524 9774
rect 41468 9538 41524 9548
rect 40908 9214 40910 9266
rect 40962 9214 40964 9266
rect 40908 9202 40964 9214
rect 40348 9156 40404 9166
rect 40348 9062 40404 9100
rect 41132 9156 41188 9166
rect 41132 9062 41188 9100
rect 41356 9154 41412 9166
rect 41356 9102 41358 9154
rect 41410 9102 41412 9154
rect 39788 8306 39844 8316
rect 40012 9042 40068 9054
rect 40012 8990 40014 9042
rect 40066 8990 40068 9042
rect 38780 8260 38836 8270
rect 38780 8166 38836 8204
rect 39452 8148 39508 8158
rect 39452 7700 39508 8092
rect 38668 6078 38670 6130
rect 38722 6078 38724 6130
rect 38668 6066 38724 6078
rect 39340 7698 39508 7700
rect 39340 7646 39454 7698
rect 39506 7646 39508 7698
rect 39340 7644 39508 7646
rect 39340 6130 39396 7644
rect 39452 7634 39508 7644
rect 40012 7700 40068 8990
rect 41356 9044 41412 9102
rect 41356 8978 41412 8988
rect 41020 8930 41076 8942
rect 41020 8878 41022 8930
rect 41074 8878 41076 8930
rect 40348 8484 40404 8494
rect 40348 8390 40404 8428
rect 40236 8370 40292 8382
rect 40236 8318 40238 8370
rect 40290 8318 40292 8370
rect 40124 8258 40180 8270
rect 40124 8206 40126 8258
rect 40178 8206 40180 8258
rect 40124 8148 40180 8206
rect 40124 8082 40180 8092
rect 40012 7634 40068 7644
rect 39564 7364 39620 7374
rect 40012 7364 40068 7374
rect 39564 7362 39956 7364
rect 39564 7310 39566 7362
rect 39618 7310 39956 7362
rect 39564 7308 39956 7310
rect 39564 7298 39620 7308
rect 39900 6802 39956 7308
rect 40012 7270 40068 7308
rect 40236 6914 40292 8318
rect 40908 8372 40964 8382
rect 40908 8258 40964 8316
rect 40908 8206 40910 8258
rect 40962 8206 40964 8258
rect 40908 8194 40964 8206
rect 41020 8260 41076 8878
rect 41580 8370 41636 9998
rect 41916 9828 41972 10332
rect 42140 10498 42196 10510
rect 42140 10446 42142 10498
rect 42194 10446 42196 10498
rect 42028 9828 42084 9838
rect 41916 9826 42084 9828
rect 41916 9774 42030 9826
rect 42082 9774 42084 9826
rect 41916 9772 42084 9774
rect 42028 9762 42084 9772
rect 42140 9604 42196 10446
rect 42140 9538 42196 9548
rect 41580 8318 41582 8370
rect 41634 8318 41636 8370
rect 41580 8306 41636 8318
rect 41916 9042 41972 9054
rect 41916 8990 41918 9042
rect 41970 8990 41972 9042
rect 41020 8194 41076 8204
rect 41244 8258 41300 8270
rect 41244 8206 41246 8258
rect 41298 8206 41300 8258
rect 41244 8036 41300 8206
rect 40236 6862 40238 6914
rect 40290 6862 40292 6914
rect 40236 6850 40292 6862
rect 41020 6916 41076 6926
rect 41244 6916 41300 7980
rect 41468 7700 41524 7710
rect 41468 7606 41524 7644
rect 41020 6914 41300 6916
rect 41020 6862 41022 6914
rect 41074 6862 41300 6914
rect 41020 6860 41300 6862
rect 41356 7474 41412 7486
rect 41356 7422 41358 7474
rect 41410 7422 41412 7474
rect 41020 6850 41076 6860
rect 39900 6750 39902 6802
rect 39954 6750 39956 6802
rect 39900 6738 39956 6750
rect 40236 6690 40292 6702
rect 40236 6638 40238 6690
rect 40290 6638 40292 6690
rect 39340 6078 39342 6130
rect 39394 6078 39396 6130
rect 36092 5966 36094 6018
rect 36146 5966 36148 6018
rect 36092 5954 36148 5966
rect 39228 5908 39284 5918
rect 38220 5794 38276 5806
rect 38220 5742 38222 5794
rect 38274 5742 38276 5794
rect 36988 5684 37044 5694
rect 36316 5460 36372 5470
rect 36316 5122 36372 5404
rect 36316 5070 36318 5122
rect 36370 5070 36372 5122
rect 36316 5058 36372 5070
rect 36876 5348 36932 5358
rect 35868 5010 36036 5012
rect 35868 4958 35870 5010
rect 35922 4958 36036 5010
rect 35868 4956 36036 4958
rect 35868 4946 35924 4956
rect 34076 4246 34132 4284
rect 34748 4226 34804 4238
rect 34748 4174 34750 4226
rect 34802 4174 34804 4226
rect 33628 4116 33684 4126
rect 34748 4116 34804 4174
rect 33628 4114 34804 4116
rect 33628 4062 33630 4114
rect 33682 4062 34804 4114
rect 33628 4060 34804 4062
rect 33628 4050 33684 4060
rect 34972 800 35028 4844
rect 35084 4844 35252 4900
rect 36092 4898 36148 4910
rect 36092 4846 36094 4898
rect 36146 4846 36148 4898
rect 35084 3666 35140 4844
rect 36092 4788 36148 4846
rect 36092 4722 36148 4732
rect 36876 4226 36932 5292
rect 36988 5122 37044 5628
rect 38220 5460 38276 5742
rect 38220 5394 38276 5404
rect 39228 5348 39284 5852
rect 39228 5282 39284 5292
rect 39340 5236 39396 6078
rect 39452 6132 39508 6142
rect 39452 6038 39508 6076
rect 40236 6132 40292 6638
rect 40236 6066 40292 6076
rect 40572 6578 40628 6590
rect 40572 6526 40574 6578
rect 40626 6526 40628 6578
rect 39564 5906 39620 5918
rect 39564 5854 39566 5906
rect 39618 5854 39620 5906
rect 39564 5684 39620 5854
rect 39564 5618 39620 5628
rect 39788 5906 39844 5918
rect 39788 5854 39790 5906
rect 39842 5854 39844 5906
rect 39788 5460 39844 5854
rect 39788 5394 39844 5404
rect 39900 5908 39956 5918
rect 39900 5346 39956 5852
rect 40124 5794 40180 5806
rect 40124 5742 40126 5794
rect 40178 5742 40180 5794
rect 40124 5684 40180 5742
rect 40236 5796 40292 5806
rect 40236 5702 40292 5740
rect 40124 5618 40180 5628
rect 39900 5294 39902 5346
rect 39954 5294 39956 5346
rect 39900 5282 39956 5294
rect 40236 5348 40292 5358
rect 40236 5254 40292 5292
rect 40572 5348 40628 6526
rect 41132 6580 41188 6590
rect 41132 6578 41300 6580
rect 41132 6526 41134 6578
rect 41186 6526 41300 6578
rect 41132 6524 41300 6526
rect 41132 6514 41188 6524
rect 41020 6466 41076 6478
rect 41020 6414 41022 6466
rect 41074 6414 41076 6466
rect 41020 6132 41076 6414
rect 41020 6066 41076 6076
rect 41244 6130 41300 6524
rect 41244 6078 41246 6130
rect 41298 6078 41300 6130
rect 41244 6066 41300 6078
rect 41132 6020 41188 6030
rect 40796 5908 40852 5918
rect 40572 5282 40628 5292
rect 40684 5906 40852 5908
rect 40684 5854 40798 5906
rect 40850 5854 40852 5906
rect 40684 5852 40852 5854
rect 41132 5908 41188 5964
rect 41356 5908 41412 7422
rect 41580 7474 41636 7486
rect 41580 7422 41582 7474
rect 41634 7422 41636 7474
rect 41580 6692 41636 7422
rect 41692 7476 41748 7486
rect 41692 7382 41748 7420
rect 41916 7252 41972 8990
rect 42028 9042 42084 9054
rect 42028 8990 42030 9042
rect 42082 8990 42084 9042
rect 42028 7588 42084 8990
rect 42140 9044 42196 9054
rect 42140 8950 42196 8988
rect 42252 9042 42308 9054
rect 42252 8990 42254 9042
rect 42306 8990 42308 9042
rect 42252 8932 42308 8990
rect 42252 8484 42308 8876
rect 42364 8820 42420 11004
rect 43484 10836 43540 12126
rect 43820 11618 43876 12236
rect 43932 12178 43988 12236
rect 43932 12126 43934 12178
rect 43986 12126 43988 12178
rect 43932 12114 43988 12126
rect 44156 12180 44212 12190
rect 44268 12180 44324 12684
rect 44156 12178 44324 12180
rect 44156 12126 44158 12178
rect 44210 12126 44324 12178
rect 44156 12124 44324 12126
rect 44156 12114 44212 12124
rect 43820 11566 43822 11618
rect 43874 11566 43876 11618
rect 43820 11554 43876 11566
rect 43932 11284 43988 11294
rect 43596 11172 43652 11182
rect 43596 11078 43652 11116
rect 42476 10780 43540 10836
rect 42476 10722 42532 10780
rect 42476 10670 42478 10722
rect 42530 10670 42532 10722
rect 42476 10658 42532 10670
rect 43484 10612 43540 10622
rect 42588 10388 42644 10398
rect 42588 10386 42980 10388
rect 42588 10334 42590 10386
rect 42642 10334 42980 10386
rect 42588 10332 42980 10334
rect 42588 10322 42644 10332
rect 42924 9602 42980 10332
rect 43372 9940 43428 9950
rect 43372 9826 43428 9884
rect 43372 9774 43374 9826
rect 43426 9774 43428 9826
rect 43372 9762 43428 9774
rect 42924 9550 42926 9602
rect 42978 9550 42980 9602
rect 42924 9538 42980 9550
rect 43148 9604 43204 9614
rect 43148 9510 43204 9548
rect 43372 9604 43428 9614
rect 42476 9268 42532 9278
rect 42476 9042 42532 9212
rect 42924 9268 42980 9278
rect 42924 9174 42980 9212
rect 43036 9156 43092 9166
rect 43036 9062 43092 9100
rect 42476 8990 42478 9042
rect 42530 8990 42532 9042
rect 42476 8978 42532 8990
rect 43148 9044 43204 9054
rect 43204 8988 43316 9044
rect 43148 8950 43204 8988
rect 42364 8764 43092 8820
rect 42252 8428 42532 8484
rect 42140 8260 42196 8270
rect 42140 8166 42196 8204
rect 42364 8148 42420 8158
rect 42364 8054 42420 8092
rect 42028 7522 42084 7532
rect 42252 7924 42308 7934
rect 42028 7252 42084 7262
rect 41916 7196 42028 7252
rect 42028 7158 42084 7196
rect 42252 6914 42308 7868
rect 42476 7698 42532 8428
rect 42588 8148 42644 8158
rect 42588 8054 42644 8092
rect 42812 8146 42868 8158
rect 42812 8094 42814 8146
rect 42866 8094 42868 8146
rect 42700 8036 42756 8046
rect 42812 8036 42868 8094
rect 42756 7980 42868 8036
rect 42700 7970 42756 7980
rect 42476 7646 42478 7698
rect 42530 7646 42532 7698
rect 42476 7634 42532 7646
rect 42812 7698 42868 7710
rect 42812 7646 42814 7698
rect 42866 7646 42868 7698
rect 42812 7588 42868 7646
rect 42924 7588 42980 7598
rect 42812 7532 42924 7588
rect 42924 7522 42980 7532
rect 42252 6862 42254 6914
rect 42306 6862 42308 6914
rect 42252 6850 42308 6862
rect 41580 6636 42084 6692
rect 41580 6468 41636 6478
rect 41916 6468 41972 6478
rect 41580 6466 41748 6468
rect 41580 6414 41582 6466
rect 41634 6414 41748 6466
rect 41580 6412 41748 6414
rect 41580 6402 41636 6412
rect 41132 5852 41412 5908
rect 41692 6356 41748 6412
rect 39340 5180 39844 5236
rect 36988 5070 36990 5122
rect 37042 5070 37044 5122
rect 36988 5058 37044 5070
rect 37436 5124 37492 5134
rect 39788 5124 39844 5180
rect 40236 5124 40292 5134
rect 39788 5122 40292 5124
rect 39788 5070 40238 5122
rect 40290 5070 40292 5122
rect 39788 5068 40292 5070
rect 36876 4174 36878 4226
rect 36930 4174 36932 4226
rect 36876 4162 36932 4174
rect 37436 4226 37492 5068
rect 40236 5058 40292 5068
rect 40684 5124 40740 5852
rect 40796 5842 40852 5852
rect 41580 5796 41636 5806
rect 41580 5702 41636 5740
rect 41244 5684 41300 5694
rect 40684 5030 40740 5068
rect 41020 5124 41076 5134
rect 41020 5010 41076 5068
rect 41020 4958 41022 5010
rect 41074 4958 41076 5010
rect 41020 4946 41076 4958
rect 37996 4900 38052 4910
rect 37996 4806 38052 4844
rect 39564 4452 39620 4462
rect 39564 4358 39620 4396
rect 40908 4452 40964 4462
rect 40908 4358 40964 4396
rect 41244 4450 41300 5628
rect 41356 5682 41412 5694
rect 41356 5630 41358 5682
rect 41410 5630 41412 5682
rect 41356 5348 41412 5630
rect 41356 5282 41412 5292
rect 41580 5572 41636 5582
rect 41580 5346 41636 5516
rect 41580 5294 41582 5346
rect 41634 5294 41636 5346
rect 41580 5282 41636 5294
rect 41692 5236 41748 6300
rect 41804 6466 41972 6468
rect 41804 6414 41918 6466
rect 41970 6414 41972 6466
rect 41804 6412 41972 6414
rect 41804 5906 41860 6412
rect 41916 6402 41972 6412
rect 42028 6468 42084 6636
rect 42364 6580 42420 6590
rect 42140 6468 42196 6478
rect 42028 6412 42140 6468
rect 41804 5854 41806 5906
rect 41858 5854 41860 5906
rect 41804 5348 41860 5854
rect 41804 5282 41860 5292
rect 41916 5908 41972 5918
rect 41916 5346 41972 5852
rect 41916 5294 41918 5346
rect 41970 5294 41972 5346
rect 41916 5282 41972 5294
rect 41692 5170 41748 5180
rect 41356 5124 41412 5134
rect 41356 5030 41412 5068
rect 42028 5124 42084 6412
rect 42140 6374 42196 6412
rect 42252 5684 42308 5694
rect 42252 5590 42308 5628
rect 42364 5572 42420 6524
rect 42924 6580 42980 6590
rect 42924 6486 42980 6524
rect 42588 6466 42644 6478
rect 42588 6414 42590 6466
rect 42642 6414 42644 6466
rect 42588 5908 42644 6414
rect 42812 6468 42868 6478
rect 42812 6374 42868 6412
rect 42700 5908 42756 5918
rect 42588 5906 42756 5908
rect 42588 5854 42702 5906
rect 42754 5854 42756 5906
rect 42588 5852 42756 5854
rect 42364 5506 42420 5516
rect 42252 5460 42308 5470
rect 42028 5058 42084 5068
rect 42140 5348 42196 5358
rect 41244 4398 41246 4450
rect 41298 4398 41300 4450
rect 41244 4386 41300 4398
rect 41580 4450 41636 4462
rect 41580 4398 41582 4450
rect 41634 4398 41636 4450
rect 40348 4340 40404 4350
rect 40348 4246 40404 4284
rect 37436 4174 37438 4226
rect 37490 4174 37492 4226
rect 37436 4162 37492 4174
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 39676 3892 39732 3902
rect 35084 3614 35086 3666
rect 35138 3614 35140 3666
rect 35084 3602 35140 3614
rect 36540 3780 36596 3790
rect 35980 3556 36036 3566
rect 35980 3462 36036 3500
rect 36540 800 36596 3724
rect 36988 3668 37044 3678
rect 36988 3574 37044 3612
rect 38108 3332 38164 3342
rect 38108 800 38164 3276
rect 38892 3332 38948 3342
rect 38892 3238 38948 3276
rect 39676 800 39732 3836
rect 41580 3892 41636 4398
rect 42140 4450 42196 5292
rect 42140 4398 42142 4450
rect 42194 4398 42196 4450
rect 42140 4386 42196 4398
rect 42028 4228 42084 4238
rect 42252 4228 42308 5404
rect 42028 4226 42308 4228
rect 42028 4174 42030 4226
rect 42082 4174 42308 4226
rect 42028 4172 42308 4174
rect 42364 5236 42420 5246
rect 42028 4162 42084 4172
rect 41580 3826 41636 3836
rect 40012 3780 40068 3790
rect 40012 3686 40068 3724
rect 42364 3554 42420 5180
rect 42700 5234 42756 5852
rect 42812 5908 42868 5918
rect 42812 5814 42868 5852
rect 43036 5908 43092 8764
rect 43260 8372 43316 8988
rect 43372 9042 43428 9548
rect 43372 8990 43374 9042
rect 43426 8990 43428 9042
rect 43372 8978 43428 8990
rect 43260 8316 43428 8372
rect 43148 8148 43204 8158
rect 43148 8054 43204 8092
rect 43260 8146 43316 8158
rect 43260 8094 43262 8146
rect 43314 8094 43316 8146
rect 43260 7924 43316 8094
rect 43260 7858 43316 7868
rect 43372 7588 43428 8316
rect 43260 7474 43316 7486
rect 43260 7422 43262 7474
rect 43314 7422 43316 7474
rect 43260 7252 43316 7422
rect 43260 7186 43316 7196
rect 43372 6692 43428 7532
rect 43484 7364 43540 10556
rect 43932 9940 43988 11228
rect 43932 9874 43988 9884
rect 44268 9828 44324 9838
rect 44380 9828 44436 15036
rect 44604 15026 44660 15036
rect 45276 14530 45332 15092
rect 45276 14478 45278 14530
rect 45330 14478 45332 14530
rect 45276 14466 45332 14478
rect 45388 14532 45444 17390
rect 45724 17442 45780 17454
rect 45724 17390 45726 17442
rect 45778 17390 45780 17442
rect 45724 15148 45780 17390
rect 46284 17442 46340 17454
rect 46284 17390 46286 17442
rect 46338 17390 46340 17442
rect 46284 16212 46340 17390
rect 46284 16146 46340 16156
rect 46620 15148 46676 17502
rect 46732 17442 46788 17454
rect 46732 17390 46734 17442
rect 46786 17390 46788 17442
rect 46732 15428 46788 17390
rect 46732 15362 46788 15372
rect 45388 14438 45444 14476
rect 45500 15092 45780 15148
rect 45836 15092 46676 15148
rect 45500 14756 45556 15092
rect 44492 14420 44548 14430
rect 44492 13970 44548 14364
rect 45500 14308 45556 14700
rect 45724 14644 45780 14654
rect 45836 14644 45892 15092
rect 45724 14642 45892 14644
rect 45724 14590 45726 14642
rect 45778 14590 45892 14642
rect 45724 14588 45892 14590
rect 45724 14578 45780 14588
rect 45612 14532 45668 14542
rect 45612 14438 45668 14476
rect 46732 14532 46788 14542
rect 46956 14532 47012 20188
rect 47180 18676 47236 20524
rect 48188 19348 48244 19358
rect 47628 19346 48244 19348
rect 47628 19294 48190 19346
rect 48242 19294 48244 19346
rect 47628 19292 48244 19294
rect 47516 18676 47572 18686
rect 47180 18674 47572 18676
rect 47180 18622 47518 18674
rect 47570 18622 47572 18674
rect 47180 18620 47572 18622
rect 47516 18610 47572 18620
rect 47628 18562 47684 19292
rect 48188 19282 48244 19292
rect 47628 18510 47630 18562
rect 47682 18510 47684 18562
rect 47628 18498 47684 18510
rect 48076 18452 48132 18462
rect 47068 18340 47124 18350
rect 47068 18246 47124 18284
rect 47852 18116 47908 18126
rect 47180 17780 47236 17790
rect 47180 17686 47236 17724
rect 47852 17554 47908 18060
rect 47852 17502 47854 17554
rect 47906 17502 47908 17554
rect 47852 17490 47908 17502
rect 47404 16212 47460 16222
rect 47404 16118 47460 16156
rect 48076 16098 48132 18396
rect 48188 18338 48244 18350
rect 48188 18286 48190 18338
rect 48242 18286 48244 18338
rect 48188 17556 48244 18286
rect 48524 17780 48580 31836
rect 48524 17714 48580 17724
rect 48188 17462 48244 17500
rect 48076 16046 48078 16098
rect 48130 16046 48132 16098
rect 47404 15428 47460 15438
rect 47404 15334 47460 15372
rect 48076 15314 48132 16046
rect 48076 15262 48078 15314
rect 48130 15262 48132 15314
rect 48076 15250 48132 15262
rect 46788 14530 47012 14532
rect 46788 14478 46958 14530
rect 47010 14478 47012 14530
rect 46788 14476 47012 14478
rect 46732 14466 46788 14476
rect 46956 14466 47012 14476
rect 46172 14420 46228 14430
rect 46172 14326 46228 14364
rect 45724 14308 45780 14318
rect 45500 14306 45780 14308
rect 45500 14254 45726 14306
rect 45778 14254 45780 14306
rect 45500 14252 45780 14254
rect 45724 14242 45780 14252
rect 46508 14308 46564 14318
rect 46508 14214 46564 14252
rect 47404 14308 47460 14318
rect 44492 13918 44494 13970
rect 44546 13918 44548 13970
rect 44492 13906 44548 13918
rect 45164 14084 45220 14094
rect 45164 12962 45220 14028
rect 47404 13858 47460 14252
rect 47404 13806 47406 13858
rect 47458 13806 47460 13858
rect 47404 13794 47460 13806
rect 48076 13746 48132 13758
rect 48076 13694 48078 13746
rect 48130 13694 48132 13746
rect 45276 13634 45332 13646
rect 45276 13582 45278 13634
rect 45330 13582 45332 13634
rect 45276 13188 45332 13582
rect 45276 13122 45332 13132
rect 45164 12910 45166 12962
rect 45218 12910 45220 12962
rect 44940 12068 44996 12078
rect 45164 12068 45220 12910
rect 45388 12964 45444 12974
rect 45388 12870 45444 12908
rect 45724 12852 45780 12862
rect 46060 12852 46116 12862
rect 45724 12850 46116 12852
rect 45724 12798 45726 12850
rect 45778 12798 46062 12850
rect 46114 12798 46116 12850
rect 45724 12796 46116 12798
rect 45724 12786 45780 12796
rect 46060 12786 46116 12796
rect 47852 12852 47908 12862
rect 47852 12758 47908 12796
rect 46396 12740 46452 12750
rect 46396 12646 46452 12684
rect 47404 12740 47460 12750
rect 47404 12290 47460 12684
rect 47628 12738 47684 12750
rect 47628 12686 47630 12738
rect 47682 12686 47684 12738
rect 47628 12628 47684 12686
rect 47628 12562 47684 12572
rect 47404 12238 47406 12290
rect 47458 12238 47460 12290
rect 47404 12226 47460 12238
rect 48076 12178 48132 13694
rect 48188 12738 48244 12750
rect 48188 12686 48190 12738
rect 48242 12686 48244 12738
rect 48188 12628 48244 12686
rect 48188 12562 48244 12572
rect 48076 12126 48078 12178
rect 48130 12126 48132 12178
rect 44492 12012 44884 12068
rect 44492 11954 44548 12012
rect 44492 11902 44494 11954
rect 44546 11902 44548 11954
rect 44492 11890 44548 11902
rect 44604 11788 44660 11798
rect 44828 11788 44884 12012
rect 44940 12066 45220 12068
rect 44940 12014 44942 12066
rect 44994 12014 45220 12066
rect 44940 12012 45220 12014
rect 44940 12002 44996 12012
rect 44828 11732 45108 11788
rect 44268 9826 44436 9828
rect 44268 9774 44270 9826
rect 44322 9774 44436 9826
rect 44268 9772 44436 9774
rect 44492 11396 44548 11406
rect 43820 9714 43876 9726
rect 43820 9662 43822 9714
rect 43874 9662 43876 9714
rect 43596 8820 43652 8830
rect 43820 8820 43876 9662
rect 44268 9604 44324 9772
rect 44268 9538 44324 9548
rect 44268 9044 44324 9054
rect 44268 8950 44324 8988
rect 43596 8818 43876 8820
rect 43596 8766 43598 8818
rect 43650 8766 43876 8818
rect 43596 8764 43876 8766
rect 44156 8930 44212 8942
rect 44156 8878 44158 8930
rect 44210 8878 44212 8930
rect 43596 8258 43652 8764
rect 44156 8484 44212 8878
rect 43932 8482 44212 8484
rect 43932 8430 44158 8482
rect 44210 8430 44212 8482
rect 43932 8428 44212 8430
rect 43820 8372 43876 8382
rect 43820 8278 43876 8316
rect 43596 8206 43598 8258
rect 43650 8206 43652 8258
rect 43596 8036 43652 8206
rect 43596 7970 43652 7980
rect 43596 7476 43652 7486
rect 43820 7476 43876 7486
rect 43932 7476 43988 8428
rect 44156 8418 44212 8428
rect 43596 7382 43652 7420
rect 43708 7474 43988 7476
rect 43708 7422 43822 7474
rect 43874 7422 43988 7474
rect 43708 7420 43988 7422
rect 43484 7252 43540 7308
rect 43484 7196 43652 7252
rect 43372 6626 43428 6636
rect 43260 6580 43316 6590
rect 43260 6486 43316 6524
rect 43484 5908 43540 5918
rect 43036 5906 43540 5908
rect 43036 5854 43038 5906
rect 43090 5854 43486 5906
rect 43538 5854 43540 5906
rect 43036 5852 43540 5854
rect 43036 5842 43092 5852
rect 43484 5842 43540 5852
rect 42700 5182 42702 5234
rect 42754 5182 42756 5234
rect 42700 5170 42756 5182
rect 42812 5460 42868 5470
rect 42812 5122 42868 5404
rect 43484 5236 43540 5246
rect 43484 5142 43540 5180
rect 42812 5070 42814 5122
rect 42866 5070 42868 5122
rect 42812 5058 42868 5070
rect 43596 4338 43652 7196
rect 43708 6690 43764 7420
rect 43820 7410 43876 7420
rect 43932 7364 43988 7420
rect 44380 7476 44436 7486
rect 44492 7476 44548 11340
rect 44604 9268 44660 11732
rect 45052 11618 45108 11732
rect 45052 11566 45054 11618
rect 45106 11566 45108 11618
rect 45052 11554 45108 11566
rect 45164 11620 45220 12012
rect 45276 12068 45332 12078
rect 45276 11974 45332 12012
rect 45164 11554 45220 11564
rect 44828 11396 44884 11406
rect 44604 9202 44660 9212
rect 44716 11394 44884 11396
rect 44716 11342 44830 11394
rect 44882 11342 44884 11394
rect 44716 11340 44884 11342
rect 44716 11172 44772 11340
rect 44828 11330 44884 11340
rect 45276 11396 45332 11406
rect 45276 11302 45332 11340
rect 45500 11394 45556 11406
rect 45500 11342 45502 11394
rect 45554 11342 45556 11394
rect 45500 11172 45556 11342
rect 46732 11396 46788 11406
rect 46732 11302 46788 11340
rect 45612 11284 45668 11294
rect 45948 11284 46004 11294
rect 45612 11282 46004 11284
rect 45612 11230 45614 11282
rect 45666 11230 45950 11282
rect 46002 11230 46004 11282
rect 45612 11228 46004 11230
rect 45612 11218 45668 11228
rect 45948 11218 46004 11228
rect 44716 8372 44772 11116
rect 45164 11116 45556 11172
rect 46284 11170 46340 11182
rect 46284 11118 46286 11170
rect 46338 11118 46340 11170
rect 45164 11060 45220 11116
rect 45052 9940 45108 9950
rect 45164 9940 45220 11004
rect 45052 9938 45220 9940
rect 45052 9886 45054 9938
rect 45106 9886 45220 9938
rect 45052 9884 45220 9886
rect 45276 9940 45332 9950
rect 45052 9874 45108 9884
rect 45276 9846 45332 9884
rect 46284 9940 46340 11118
rect 47964 10724 48020 10734
rect 48076 10724 48132 12126
rect 47964 10722 48132 10724
rect 47964 10670 47966 10722
rect 48018 10670 48132 10722
rect 47964 10668 48132 10670
rect 47964 10658 48020 10668
rect 46284 9874 46340 9884
rect 47404 9940 47460 9950
rect 47404 9846 47460 9884
rect 48076 9826 48132 10668
rect 48076 9774 48078 9826
rect 48130 9774 48132 9826
rect 48076 9042 48132 9774
rect 48076 8990 48078 9042
rect 48130 8990 48132 9042
rect 44940 8932 44996 8942
rect 45276 8932 45332 8942
rect 44940 8930 45220 8932
rect 44940 8878 44942 8930
rect 44994 8878 45220 8930
rect 44940 8876 45220 8878
rect 44940 8866 44996 8876
rect 45164 8596 45220 8876
rect 45276 8838 45332 8876
rect 46508 8932 46564 8942
rect 45164 8540 45332 8596
rect 44716 8306 44772 8316
rect 44828 8484 44884 8494
rect 45276 8484 45332 8540
rect 45276 8428 45444 8484
rect 44716 8148 44772 8158
rect 44716 7698 44772 8092
rect 44716 7646 44718 7698
rect 44770 7646 44772 7698
rect 44716 7634 44772 7646
rect 44380 7474 44548 7476
rect 44380 7422 44382 7474
rect 44434 7422 44548 7474
rect 44380 7420 44548 7422
rect 44380 7410 44436 7420
rect 43932 7298 43988 7308
rect 44044 7252 44100 7262
rect 43708 6638 43710 6690
rect 43762 6638 43764 6690
rect 43708 6626 43764 6638
rect 43820 6692 43876 6702
rect 43820 6598 43876 6636
rect 44044 6690 44100 7196
rect 44156 7250 44212 7262
rect 44156 7198 44158 7250
rect 44210 7198 44212 7250
rect 44156 7140 44212 7198
rect 44212 7084 44324 7140
rect 44156 7074 44212 7084
rect 44044 6638 44046 6690
rect 44098 6638 44100 6690
rect 44044 6580 44100 6638
rect 44156 6580 44212 6590
rect 44044 6578 44212 6580
rect 44044 6526 44158 6578
rect 44210 6526 44212 6578
rect 44044 6524 44212 6526
rect 44156 6514 44212 6524
rect 43708 5682 43764 5694
rect 44044 5684 44100 5694
rect 43708 5630 43710 5682
rect 43762 5630 43764 5682
rect 43708 5236 43764 5630
rect 43708 5170 43764 5180
rect 43932 5682 44100 5684
rect 43932 5630 44046 5682
rect 44098 5630 44100 5682
rect 43932 5628 44100 5630
rect 43596 4286 43598 4338
rect 43650 4286 43652 4338
rect 43596 3668 43652 4286
rect 43596 3602 43652 3612
rect 42364 3502 42366 3554
rect 42418 3502 42420 3554
rect 42364 3490 42420 3502
rect 43932 3554 43988 5628
rect 44044 5618 44100 5628
rect 44268 5236 44324 7084
rect 44492 6916 44548 7420
rect 44828 7474 44884 8428
rect 45388 8372 45444 8428
rect 45500 8372 45556 8382
rect 45388 8370 45556 8372
rect 45276 8314 45332 8326
rect 45388 8318 45502 8370
rect 45554 8318 45556 8370
rect 45388 8316 45556 8318
rect 45164 8260 45220 8270
rect 45276 8262 45278 8314
rect 45330 8262 45332 8314
rect 45500 8306 45556 8316
rect 45276 8260 45332 8262
rect 45220 8204 45332 8260
rect 44828 7422 44830 7474
rect 44882 7422 44884 7474
rect 44828 7410 44884 7422
rect 44940 8034 44996 8046
rect 44940 7982 44942 8034
rect 44994 7982 44996 8034
rect 44604 7364 44660 7374
rect 44604 7270 44660 7308
rect 44940 7140 44996 7982
rect 44940 7074 44996 7084
rect 45052 7476 45108 7486
rect 44548 6860 44660 6916
rect 44492 6850 44548 6860
rect 44380 6578 44436 6590
rect 44380 6526 44382 6578
rect 44434 6526 44436 6578
rect 44380 5682 44436 6526
rect 44604 6130 44660 6860
rect 45052 6914 45108 7420
rect 45052 6862 45054 6914
rect 45106 6862 45108 6914
rect 45052 6850 45108 6862
rect 44828 6690 44884 6702
rect 44828 6638 44830 6690
rect 44882 6638 44884 6690
rect 44828 6580 44884 6638
rect 44828 6514 44884 6524
rect 44604 6078 44606 6130
rect 44658 6078 44660 6130
rect 44604 6066 44660 6078
rect 45052 6132 45108 6142
rect 45164 6132 45220 8204
rect 45836 8148 45892 8158
rect 46172 8148 46228 8158
rect 45836 8146 46228 8148
rect 45836 8094 45838 8146
rect 45890 8094 46174 8146
rect 46226 8094 46228 8146
rect 45836 8092 46228 8094
rect 45836 8082 45892 8092
rect 46172 8082 46228 8092
rect 46508 8146 46564 8876
rect 47404 8932 47460 8942
rect 47404 8838 47460 8876
rect 47180 8484 47236 8494
rect 47180 8390 47236 8428
rect 46844 8372 46900 8382
rect 46844 8278 46900 8316
rect 46508 8094 46510 8146
rect 46562 8094 46564 8146
rect 46508 8082 46564 8094
rect 47852 8148 47908 8158
rect 47852 8054 47908 8092
rect 45276 8036 45332 8046
rect 45276 7362 45332 7980
rect 47068 8036 47124 8046
rect 47516 8036 47572 8046
rect 47068 7942 47124 7980
rect 47404 8034 47572 8036
rect 47404 7982 47518 8034
rect 47570 7982 47572 8034
rect 47404 7980 47572 7982
rect 47404 7586 47460 7980
rect 47516 7970 47572 7980
rect 47404 7534 47406 7586
rect 47458 7534 47460 7586
rect 47404 7522 47460 7534
rect 45276 7310 45278 7362
rect 45330 7310 45332 7362
rect 45276 7298 45332 7310
rect 48076 7474 48132 8990
rect 48076 7422 48078 7474
rect 48130 7422 48132 7474
rect 45500 7140 45556 7150
rect 45276 6916 45332 6926
rect 45276 6822 45332 6860
rect 45500 6914 45556 7084
rect 45500 6862 45502 6914
rect 45554 6862 45556 6914
rect 45500 6850 45556 6862
rect 46732 6916 46788 6926
rect 46732 6802 46788 6860
rect 46732 6750 46734 6802
rect 46786 6750 46788 6802
rect 46732 6738 46788 6750
rect 47852 6804 47908 6814
rect 47628 6692 47684 6702
rect 47628 6598 47684 6636
rect 45612 6580 45668 6590
rect 45948 6580 46004 6590
rect 45612 6578 46004 6580
rect 45612 6526 45614 6578
rect 45666 6526 45950 6578
rect 46002 6526 46004 6578
rect 45612 6524 46004 6526
rect 45612 6514 45668 6524
rect 45948 6514 46004 6524
rect 47852 6578 47908 6748
rect 47852 6526 47854 6578
rect 47906 6526 47908 6578
rect 47852 6514 47908 6526
rect 46284 6468 46340 6478
rect 46284 6374 46340 6412
rect 47404 6468 47460 6478
rect 45052 6130 45220 6132
rect 45052 6078 45054 6130
rect 45106 6078 45220 6130
rect 45052 6076 45220 6078
rect 45052 6066 45108 6076
rect 47404 6018 47460 6412
rect 47404 5966 47406 6018
rect 47458 5966 47460 6018
rect 47404 5954 47460 5966
rect 48076 5906 48132 7422
rect 48188 7700 48244 7710
rect 48188 6692 48244 7644
rect 48188 6598 48244 6636
rect 48076 5854 48078 5906
rect 48130 5854 48132 5906
rect 48076 5842 48132 5854
rect 45276 5794 45332 5806
rect 45276 5742 45278 5794
rect 45330 5742 45332 5794
rect 44380 5630 44382 5682
rect 44434 5630 44436 5682
rect 44380 5618 44436 5630
rect 45052 5684 45108 5694
rect 45276 5684 45332 5742
rect 45052 5682 45332 5684
rect 45052 5630 45054 5682
rect 45106 5630 45332 5682
rect 45052 5628 45332 5630
rect 45052 5618 45108 5628
rect 44828 5348 44884 5358
rect 44380 5236 44436 5246
rect 44268 5234 44436 5236
rect 44268 5182 44382 5234
rect 44434 5182 44436 5234
rect 44268 5180 44436 5182
rect 44380 5170 44436 5180
rect 44828 5234 44884 5292
rect 44828 5182 44830 5234
rect 44882 5182 44884 5234
rect 44828 5170 44884 5182
rect 43932 3502 43934 3554
rect 43986 3502 43988 3554
rect 43932 3490 43988 3502
rect 44156 5124 44212 5134
rect 44156 3442 44212 5068
rect 46956 5124 47012 5134
rect 46956 5030 47012 5068
rect 47628 5122 47684 5134
rect 47628 5070 47630 5122
rect 47682 5070 47684 5122
rect 45388 4450 45444 4462
rect 45388 4398 45390 4450
rect 45442 4398 45444 4450
rect 45388 4340 45444 4398
rect 45388 4274 45444 4284
rect 47628 4340 47684 5070
rect 47628 4274 47684 4284
rect 45500 3668 45556 3678
rect 45500 3574 45556 3612
rect 44156 3390 44158 3442
rect 44210 3390 44212 3442
rect 44156 3378 44212 3390
rect 47628 3554 47684 3566
rect 47628 3502 47630 3554
rect 47682 3502 47684 3554
rect 42700 3330 42756 3342
rect 42700 3278 42702 3330
rect 42754 3278 42756 3330
rect 41244 1764 41300 1774
rect 41244 800 41300 1708
rect 42700 1764 42756 3278
rect 42700 1698 42756 1708
rect 42812 3332 42868 3342
rect 42812 800 42868 3276
rect 44492 3332 44548 3342
rect 44940 3332 44996 3342
rect 46172 3332 46228 3342
rect 44492 3238 44548 3276
rect 44604 3330 44996 3332
rect 44604 3278 44942 3330
rect 44994 3278 44996 3330
rect 44604 3276 44996 3278
rect 44604 980 44660 3276
rect 44940 3266 44996 3276
rect 45948 3330 46228 3332
rect 45948 3278 46174 3330
rect 46226 3278 46228 3330
rect 45948 3276 46228 3278
rect 44380 924 44660 980
rect 44380 800 44436 924
rect 45948 800 46004 3276
rect 46172 3266 46228 3276
rect 47628 3332 47684 3502
rect 47852 3444 47908 3482
rect 47852 3378 47908 3388
rect 48188 3442 48244 3454
rect 48188 3390 48190 3442
rect 48242 3390 48244 3442
rect 47628 3266 47684 3276
rect 48188 3332 48244 3390
rect 48188 2772 48244 3276
rect 48188 2706 48244 2716
rect 15372 700 15876 756
rect 16128 0 16240 800
rect 17696 0 17808 800
rect 19264 0 19376 800
rect 20832 0 20944 800
rect 22400 0 22512 800
rect 23968 0 24080 800
rect 25536 0 25648 800
rect 27104 0 27216 800
rect 28672 0 28784 800
rect 30240 0 30352 800
rect 31808 0 31920 800
rect 33376 0 33488 800
rect 34944 0 35056 800
rect 36512 0 36624 800
rect 38080 0 38192 800
rect 39648 0 39760 800
rect 41216 0 41328 800
rect 42784 0 42896 800
rect 44352 0 44464 800
rect 45920 0 46032 800
<< via2 >>
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 4620 41244 4676 41300
rect 6076 41298 6132 41300
rect 6076 41246 6078 41298
rect 6078 41246 6130 41298
rect 6130 41246 6132 41298
rect 6076 41244 6132 41246
rect 1708 39452 1764 39508
rect 3052 39394 3108 39396
rect 3052 39342 3054 39394
rect 3054 39342 3106 39394
rect 3106 39342 3108 39394
rect 3052 39340 3108 39342
rect 3388 39506 3444 39508
rect 3388 39454 3390 39506
rect 3390 39454 3442 39506
rect 3442 39454 3444 39506
rect 3388 39452 3444 39454
rect 2828 38780 2884 38836
rect 2716 38668 2772 38724
rect 1708 37996 1764 38052
rect 3388 38780 3444 38836
rect 2604 37826 2660 37828
rect 2604 37774 2606 37826
rect 2606 37774 2658 37826
rect 2658 37774 2660 37826
rect 2604 37772 2660 37774
rect 3276 37772 3332 37828
rect 2940 36540 2996 36596
rect 1708 35756 1764 35812
rect 3276 34860 3332 34916
rect 2940 34802 2996 34804
rect 2940 34750 2942 34802
rect 2942 34750 2994 34802
rect 2994 34750 2996 34802
rect 2940 34748 2996 34750
rect 2380 34636 2436 34692
rect 3276 34636 3332 34692
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 4060 39452 4116 39508
rect 3948 39228 4004 39284
rect 3836 38722 3892 38724
rect 3836 38670 3838 38722
rect 3838 38670 3890 38722
rect 3890 38670 3892 38722
rect 3836 38668 3892 38670
rect 3836 38050 3892 38052
rect 3836 37998 3838 38050
rect 3838 37998 3890 38050
rect 3890 37998 3892 38050
rect 3836 37996 3892 37998
rect 3500 35084 3556 35140
rect 3836 36594 3892 36596
rect 3836 36542 3838 36594
rect 3838 36542 3890 36594
rect 3890 36542 3892 36594
rect 3836 36540 3892 36542
rect 3724 35810 3780 35812
rect 3724 35758 3726 35810
rect 3726 35758 3778 35810
rect 3778 35758 3780 35810
rect 3724 35756 3780 35758
rect 4508 39340 4564 39396
rect 4620 39228 4676 39284
rect 6076 38946 6132 38948
rect 6076 38894 6078 38946
rect 6078 38894 6130 38946
rect 6130 38894 6132 38946
rect 6076 38892 6132 38894
rect 10444 44492 10500 44548
rect 7644 44434 7700 44436
rect 7644 44382 7646 44434
rect 7646 44382 7698 44434
rect 7698 44382 7700 44434
rect 7644 44380 7700 44382
rect 9772 43484 9828 43540
rect 9884 43596 9940 43652
rect 6636 43426 6692 43428
rect 6636 43374 6638 43426
rect 6638 43374 6690 43426
rect 6690 43374 6692 43426
rect 6636 43372 6692 43374
rect 8876 43148 8932 43204
rect 9548 43148 9604 43204
rect 10780 44156 10836 44212
rect 17500 45836 17556 45892
rect 11564 44380 11620 44436
rect 12012 44434 12068 44436
rect 12012 44382 12014 44434
rect 12014 44382 12066 44434
rect 12066 44382 12068 44434
rect 12012 44380 12068 44382
rect 11340 44044 11396 44100
rect 11452 44210 11508 44212
rect 11452 44158 11454 44210
rect 11454 44158 11506 44210
rect 11506 44158 11508 44210
rect 11452 44156 11508 44158
rect 11676 43708 11732 43764
rect 10892 43596 10948 43652
rect 10444 43426 10500 43428
rect 10444 43374 10446 43426
rect 10446 43374 10498 43426
rect 10498 43374 10500 43426
rect 10444 43372 10500 43374
rect 11900 43538 11956 43540
rect 11900 43486 11902 43538
rect 11902 43486 11954 43538
rect 11954 43486 11956 43538
rect 11900 43484 11956 43486
rect 11004 43372 11060 43428
rect 11564 43426 11620 43428
rect 11564 43374 11566 43426
rect 11566 43374 11618 43426
rect 11618 43374 11620 43426
rect 11564 43372 11620 43374
rect 6860 42028 6916 42084
rect 8988 41580 9044 41636
rect 10780 43314 10836 43316
rect 10780 43262 10782 43314
rect 10782 43262 10834 43314
rect 10834 43262 10836 43314
rect 10780 43260 10836 43262
rect 10556 43036 10612 43092
rect 10332 41916 10388 41972
rect 10444 41858 10500 41860
rect 10444 41806 10446 41858
rect 10446 41806 10498 41858
rect 10498 41806 10500 41858
rect 10444 41804 10500 41806
rect 10780 42082 10836 42084
rect 10780 42030 10782 42082
rect 10782 42030 10834 42082
rect 10834 42030 10836 42082
rect 10780 42028 10836 42030
rect 11788 43036 11844 43092
rect 12236 43426 12292 43428
rect 12236 43374 12238 43426
rect 12238 43374 12290 43426
rect 12290 43374 12292 43426
rect 12236 43372 12292 43374
rect 12572 43372 12628 43428
rect 12348 43260 12404 43316
rect 12124 43036 12180 43092
rect 16716 44994 16772 44996
rect 16716 44942 16718 44994
rect 16718 44942 16770 44994
rect 16770 44942 16772 44994
rect 16716 44940 16772 44942
rect 14588 44492 14644 44548
rect 16156 44546 16212 44548
rect 16156 44494 16158 44546
rect 16158 44494 16210 44546
rect 16210 44494 16212 44546
rect 16156 44492 16212 44494
rect 13580 43650 13636 43652
rect 13580 43598 13582 43650
rect 13582 43598 13634 43650
rect 13634 43598 13636 43650
rect 13580 43596 13636 43598
rect 12684 42252 12740 42308
rect 10892 41916 10948 41972
rect 11676 41970 11732 41972
rect 11676 41918 11678 41970
rect 11678 41918 11730 41970
rect 11730 41918 11732 41970
rect 11676 41916 11732 41918
rect 11228 41858 11284 41860
rect 11228 41806 11230 41858
rect 11230 41806 11282 41858
rect 11282 41806 11284 41858
rect 11228 41804 11284 41806
rect 9884 41580 9940 41636
rect 10332 41132 10388 41188
rect 11116 41746 11172 41748
rect 11116 41694 11118 41746
rect 11118 41694 11170 41746
rect 11170 41694 11172 41746
rect 11116 41692 11172 41694
rect 11788 41692 11844 41748
rect 11900 41580 11956 41636
rect 12012 41804 12068 41860
rect 12460 41804 12516 41860
rect 11340 40962 11396 40964
rect 11340 40910 11342 40962
rect 11342 40910 11394 40962
rect 11394 40910 11396 40962
rect 11340 40908 11396 40910
rect 12348 40572 12404 40628
rect 15820 44322 15876 44324
rect 15820 44270 15822 44322
rect 15822 44270 15874 44322
rect 15874 44270 15876 44322
rect 15820 44268 15876 44270
rect 15036 44210 15092 44212
rect 15036 44158 15038 44210
rect 15038 44158 15090 44210
rect 15090 44158 15092 44210
rect 15036 44156 15092 44158
rect 14364 44044 14420 44100
rect 15820 44044 15876 44100
rect 16044 44044 16100 44100
rect 15260 43708 15316 43764
rect 17388 44434 17444 44436
rect 17388 44382 17390 44434
rect 17390 44382 17442 44434
rect 17442 44382 17444 44434
rect 17388 44380 17444 44382
rect 16604 44156 16660 44212
rect 16044 43762 16100 43764
rect 16044 43710 16046 43762
rect 16046 43710 16098 43762
rect 16098 43710 16100 43762
rect 16044 43708 16100 43710
rect 17276 44268 17332 44324
rect 17052 44210 17108 44212
rect 17052 44158 17054 44210
rect 17054 44158 17106 44210
rect 17106 44158 17108 44210
rect 17052 44156 17108 44158
rect 16940 44044 16996 44100
rect 16604 43650 16660 43652
rect 16604 43598 16606 43650
rect 16606 43598 16658 43650
rect 16658 43598 16660 43650
rect 16604 43596 16660 43598
rect 14140 43260 14196 43316
rect 13132 41858 13188 41860
rect 13132 41806 13134 41858
rect 13134 41806 13186 41858
rect 13186 41806 13188 41858
rect 13132 41804 13188 41806
rect 12908 41074 12964 41076
rect 12908 41022 12910 41074
rect 12910 41022 12962 41074
rect 12962 41022 12964 41074
rect 12908 41020 12964 41022
rect 13804 42252 13860 42308
rect 16044 42028 16100 42084
rect 13692 41244 13748 41300
rect 13580 41186 13636 41188
rect 13580 41134 13582 41186
rect 13582 41134 13634 41186
rect 13634 41134 13636 41186
rect 13580 41132 13636 41134
rect 13468 41074 13524 41076
rect 13468 41022 13470 41074
rect 13470 41022 13522 41074
rect 13522 41022 13524 41074
rect 13468 41020 13524 41022
rect 14140 41970 14196 41972
rect 14140 41918 14142 41970
rect 14142 41918 14194 41970
rect 14194 41918 14196 41970
rect 14140 41916 14196 41918
rect 15372 41970 15428 41972
rect 15372 41918 15374 41970
rect 15374 41918 15426 41970
rect 15426 41918 15428 41970
rect 15372 41916 15428 41918
rect 16716 43538 16772 43540
rect 16716 43486 16718 43538
rect 16718 43486 16770 43538
rect 16770 43486 16772 43538
rect 16716 43484 16772 43486
rect 16940 43596 16996 43652
rect 18060 45836 18116 45892
rect 17836 44380 17892 44436
rect 17836 43650 17892 43652
rect 17836 43598 17838 43650
rect 17838 43598 17890 43650
rect 17890 43598 17892 43650
rect 17836 43596 17892 43598
rect 18396 45106 18452 45108
rect 18396 45054 18398 45106
rect 18398 45054 18450 45106
rect 18450 45054 18452 45106
rect 18396 45052 18452 45054
rect 18172 44940 18228 44996
rect 17500 43484 17556 43540
rect 16716 42642 16772 42644
rect 16716 42590 16718 42642
rect 16718 42590 16770 42642
rect 16770 42590 16772 42642
rect 16716 42588 16772 42590
rect 16716 42028 16772 42084
rect 17612 42642 17668 42644
rect 17612 42590 17614 42642
rect 17614 42590 17666 42642
rect 17666 42590 17668 42642
rect 17612 42588 17668 42590
rect 19628 45890 19684 45892
rect 19628 45838 19630 45890
rect 19630 45838 19682 45890
rect 19682 45838 19684 45890
rect 19628 45836 19684 45838
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 19068 44940 19124 44996
rect 18172 42700 18228 42756
rect 17164 42140 17220 42196
rect 14476 41298 14532 41300
rect 14476 41246 14478 41298
rect 14478 41246 14530 41298
rect 14530 41246 14532 41298
rect 14476 41244 14532 41246
rect 13132 40908 13188 40964
rect 13580 40908 13636 40964
rect 10892 40236 10948 40292
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 6076 37772 6132 37828
rect 5068 37266 5124 37268
rect 5068 37214 5070 37266
rect 5070 37214 5122 37266
rect 5122 37214 5124 37266
rect 5068 37212 5124 37214
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 5740 36370 5796 36372
rect 5740 36318 5742 36370
rect 5742 36318 5794 36370
rect 5794 36318 5796 36370
rect 5740 36316 5796 36318
rect 4396 35810 4452 35812
rect 4396 35758 4398 35810
rect 4398 35758 4450 35810
rect 4450 35758 4452 35810
rect 4396 35756 4452 35758
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 3500 34636 3556 34692
rect 4396 34914 4452 34916
rect 4396 34862 4398 34914
rect 4398 34862 4450 34914
rect 4450 34862 4452 34914
rect 4396 34860 4452 34862
rect 4732 35084 4788 35140
rect 5404 35084 5460 35140
rect 5068 34860 5124 34916
rect 3612 34748 3668 34804
rect 6412 35868 6468 35924
rect 5628 34972 5684 35028
rect 4620 34412 4676 34468
rect 5964 34412 6020 34468
rect 5964 34242 6020 34244
rect 5964 34190 5966 34242
rect 5966 34190 6018 34242
rect 6018 34190 6020 34242
rect 5964 34188 6020 34190
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 3724 31836 3780 31892
rect 2492 31666 2548 31668
rect 2492 31614 2494 31666
rect 2494 31614 2546 31666
rect 2546 31614 2548 31666
rect 2492 31612 2548 31614
rect 1820 31276 1876 31332
rect 3724 31276 3780 31332
rect 4396 31500 4452 31556
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 2492 30098 2548 30100
rect 2492 30046 2494 30098
rect 2494 30046 2546 30098
rect 2546 30046 2548 30098
rect 2492 30044 2548 30046
rect 4956 31836 5012 31892
rect 5964 33068 6020 33124
rect 7532 39506 7588 39508
rect 7532 39454 7534 39506
rect 7534 39454 7586 39506
rect 7586 39454 7588 39506
rect 7532 39452 7588 39454
rect 8540 39340 8596 39396
rect 8540 39058 8596 39060
rect 8540 39006 8542 39058
rect 8542 39006 8594 39058
rect 8594 39006 8596 39058
rect 8540 39004 8596 39006
rect 7308 38108 7364 38164
rect 10108 39506 10164 39508
rect 10108 39454 10110 39506
rect 10110 39454 10162 39506
rect 10162 39454 10164 39506
rect 10108 39452 10164 39454
rect 9996 39394 10052 39396
rect 9996 39342 9998 39394
rect 9998 39342 10050 39394
rect 10050 39342 10052 39394
rect 9996 39340 10052 39342
rect 10444 39004 10500 39060
rect 9772 38892 9828 38948
rect 10332 38946 10388 38948
rect 10332 38894 10334 38946
rect 10334 38894 10386 38946
rect 10386 38894 10388 38946
rect 10332 38892 10388 38894
rect 8092 38050 8148 38052
rect 8092 37998 8094 38050
rect 8094 37998 8146 38050
rect 8146 37998 8148 38050
rect 8092 37996 8148 37998
rect 7868 37938 7924 37940
rect 7868 37886 7870 37938
rect 7870 37886 7922 37938
rect 7922 37886 7924 37938
rect 7868 37884 7924 37886
rect 8764 38050 8820 38052
rect 8764 37998 8766 38050
rect 8766 37998 8818 38050
rect 8818 37998 8820 38050
rect 8764 37996 8820 37998
rect 8428 37884 8484 37940
rect 6748 37212 6804 37268
rect 6972 37826 7028 37828
rect 6972 37774 6974 37826
rect 6974 37774 7026 37826
rect 7026 37774 7028 37826
rect 6972 37772 7028 37774
rect 6860 36316 6916 36372
rect 6860 35756 6916 35812
rect 6636 34860 6692 34916
rect 7308 36428 7364 36484
rect 7196 35922 7252 35924
rect 7196 35870 7198 35922
rect 7198 35870 7250 35922
rect 7250 35870 7252 35922
rect 7196 35868 7252 35870
rect 8540 37378 8596 37380
rect 8540 37326 8542 37378
rect 8542 37326 8594 37378
rect 8594 37326 8596 37378
rect 8540 37324 8596 37326
rect 8204 36428 8260 36484
rect 8876 36204 8932 36260
rect 7084 35196 7140 35252
rect 8652 35810 8708 35812
rect 8652 35758 8654 35810
rect 8654 35758 8706 35810
rect 8706 35758 8708 35810
rect 8652 35756 8708 35758
rect 7868 35308 7924 35364
rect 7756 35084 7812 35140
rect 7756 34802 7812 34804
rect 7756 34750 7758 34802
rect 7758 34750 7810 34802
rect 7810 34750 7812 34802
rect 7756 34748 7812 34750
rect 8204 35308 8260 35364
rect 6860 34188 6916 34244
rect 7756 34412 7812 34468
rect 8764 34914 8820 34916
rect 8764 34862 8766 34914
rect 8766 34862 8818 34914
rect 8818 34862 8820 34914
rect 8764 34860 8820 34862
rect 8204 34802 8260 34804
rect 8204 34750 8206 34802
rect 8206 34750 8258 34802
rect 8258 34750 8260 34802
rect 8204 34748 8260 34750
rect 8876 34748 8932 34804
rect 9884 38108 9940 38164
rect 11004 39004 11060 39060
rect 10556 38556 10612 38612
rect 10780 38722 10836 38724
rect 10780 38670 10782 38722
rect 10782 38670 10834 38722
rect 10834 38670 10836 38722
rect 10780 38668 10836 38670
rect 9772 37884 9828 37940
rect 10332 37938 10388 37940
rect 10332 37886 10334 37938
rect 10334 37886 10386 37938
rect 10386 37886 10388 37938
rect 10332 37884 10388 37886
rect 9884 37324 9940 37380
rect 9660 35532 9716 35588
rect 9660 35196 9716 35252
rect 9772 37266 9828 37268
rect 9772 37214 9774 37266
rect 9774 37214 9826 37266
rect 9826 37214 9828 37266
rect 9772 37212 9828 37214
rect 9100 34636 9156 34692
rect 10556 35308 10612 35364
rect 11564 39004 11620 39060
rect 11340 38556 11396 38612
rect 11676 38668 11732 38724
rect 13132 40572 13188 40628
rect 12908 39340 12964 39396
rect 13132 38946 13188 38948
rect 13132 38894 13134 38946
rect 13134 38894 13186 38946
rect 13186 38894 13188 38946
rect 13132 38892 13188 38894
rect 14140 40514 14196 40516
rect 14140 40462 14142 40514
rect 14142 40462 14194 40514
rect 14194 40462 14196 40514
rect 14140 40460 14196 40462
rect 14476 40460 14532 40516
rect 13804 38892 13860 38948
rect 14140 40236 14196 40292
rect 15932 40514 15988 40516
rect 15932 40462 15934 40514
rect 15934 40462 15986 40514
rect 15986 40462 15988 40514
rect 15932 40460 15988 40462
rect 15708 40402 15764 40404
rect 15708 40350 15710 40402
rect 15710 40350 15762 40402
rect 15762 40350 15764 40402
rect 15708 40348 15764 40350
rect 16604 40460 16660 40516
rect 13580 38834 13636 38836
rect 13580 38782 13582 38834
rect 13582 38782 13634 38834
rect 13634 38782 13636 38834
rect 13580 38780 13636 38782
rect 12684 38722 12740 38724
rect 12684 38670 12686 38722
rect 12686 38670 12738 38722
rect 12738 38670 12740 38722
rect 12684 38668 12740 38670
rect 11900 38108 11956 38164
rect 11340 37324 11396 37380
rect 10892 35586 10948 35588
rect 10892 35534 10894 35586
rect 10894 35534 10946 35586
rect 10946 35534 10948 35586
rect 10892 35532 10948 35534
rect 10892 35196 10948 35252
rect 10780 35084 10836 35140
rect 11676 35084 11732 35140
rect 9996 34914 10052 34916
rect 9996 34862 9998 34914
rect 9998 34862 10050 34914
rect 10050 34862 10052 34914
rect 9996 34860 10052 34862
rect 11452 34914 11508 34916
rect 11452 34862 11454 34914
rect 11454 34862 11506 34914
rect 11506 34862 11508 34914
rect 11452 34860 11508 34862
rect 11228 34802 11284 34804
rect 11228 34750 11230 34802
rect 11230 34750 11282 34802
rect 11282 34750 11284 34802
rect 11228 34748 11284 34750
rect 9884 34636 9940 34692
rect 9884 33852 9940 33908
rect 11228 33964 11284 34020
rect 10332 33458 10388 33460
rect 10332 33406 10334 33458
rect 10334 33406 10386 33458
rect 10386 33406 10388 33458
rect 10332 33404 10388 33406
rect 6748 33122 6804 33124
rect 6748 33070 6750 33122
rect 6750 33070 6802 33122
rect 6802 33070 6804 33122
rect 6748 33068 6804 33070
rect 6636 31836 6692 31892
rect 5740 31666 5796 31668
rect 5740 31614 5742 31666
rect 5742 31614 5794 31666
rect 5794 31614 5796 31666
rect 5740 31612 5796 31614
rect 6188 31666 6244 31668
rect 6188 31614 6190 31666
rect 6190 31614 6242 31666
rect 6242 31614 6244 31666
rect 6188 31612 6244 31614
rect 5628 30210 5684 30212
rect 5628 30158 5630 30210
rect 5630 30158 5682 30210
rect 5682 30158 5684 30210
rect 5628 30156 5684 30158
rect 5740 30098 5796 30100
rect 5740 30046 5742 30098
rect 5742 30046 5794 30098
rect 5794 30046 5796 30098
rect 5740 30044 5796 30046
rect 4844 29932 4900 29988
rect 5740 29820 5796 29876
rect 4620 29596 4676 29652
rect 5068 29650 5124 29652
rect 5068 29598 5070 29650
rect 5070 29598 5122 29650
rect 5122 29598 5124 29650
rect 5068 29596 5124 29598
rect 3164 29372 3220 29428
rect 2492 29314 2548 29316
rect 2492 29262 2494 29314
rect 2494 29262 2546 29314
rect 2546 29262 2548 29314
rect 2492 29260 2548 29262
rect 3052 28812 3108 28868
rect 1820 27692 1876 27748
rect 2492 28588 2548 28644
rect 1708 25228 1764 25284
rect 4620 29372 4676 29428
rect 3724 29260 3780 29316
rect 3612 29148 3668 29204
rect 3500 28588 3556 28644
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 6636 31554 6692 31556
rect 6636 31502 6638 31554
rect 6638 31502 6690 31554
rect 6690 31502 6692 31554
rect 6636 31500 6692 31502
rect 7084 31666 7140 31668
rect 7084 31614 7086 31666
rect 7086 31614 7138 31666
rect 7138 31614 7140 31666
rect 7084 31612 7140 31614
rect 7084 30940 7140 30996
rect 7196 31276 7252 31332
rect 5964 30098 6020 30100
rect 5964 30046 5966 30098
rect 5966 30046 6018 30098
rect 6018 30046 6020 30098
rect 5964 30044 6020 30046
rect 7196 30716 7252 30772
rect 7756 32620 7812 32676
rect 8764 32674 8820 32676
rect 8764 32622 8766 32674
rect 8766 32622 8818 32674
rect 8818 32622 8820 32674
rect 8764 32620 8820 32622
rect 8316 32396 8372 32452
rect 7756 31276 7812 31332
rect 8652 31612 8708 31668
rect 6188 29932 6244 29988
rect 6636 29932 6692 29988
rect 6188 29708 6244 29764
rect 5628 29372 5684 29428
rect 5628 29202 5684 29204
rect 5628 29150 5630 29202
rect 5630 29150 5682 29202
rect 5682 29150 5684 29202
rect 5628 29148 5684 29150
rect 5180 28812 5236 28868
rect 3836 28700 3892 28756
rect 5068 28700 5124 28756
rect 4172 27692 4228 27748
rect 4172 26908 4228 26964
rect 3724 26236 3780 26292
rect 3836 26178 3892 26180
rect 3836 26126 3838 26178
rect 3838 26126 3890 26178
rect 3890 26126 3892 26178
rect 3836 26124 3892 26126
rect 4172 25676 4228 25732
rect 4732 28642 4788 28644
rect 4732 28590 4734 28642
rect 4734 28590 4786 28642
rect 4786 28590 4788 28642
rect 4732 28588 4788 28590
rect 4620 28476 4676 28532
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4620 27244 4676 27300
rect 4620 26908 4676 26964
rect 5404 28364 5460 28420
rect 5628 27244 5684 27300
rect 6300 29538 6356 29540
rect 6300 29486 6302 29538
rect 6302 29486 6354 29538
rect 6354 29486 6356 29538
rect 6300 29484 6356 29486
rect 6972 30098 7028 30100
rect 6972 30046 6974 30098
rect 6974 30046 7026 30098
rect 7026 30046 7028 30098
rect 6972 30044 7028 30046
rect 7420 30716 7476 30772
rect 7196 29708 7252 29764
rect 6860 29484 6916 29540
rect 6076 29372 6132 29428
rect 4844 26290 4900 26292
rect 4844 26238 4846 26290
rect 4846 26238 4898 26290
rect 4898 26238 4900 26290
rect 4844 26236 4900 26238
rect 5068 26178 5124 26180
rect 5068 26126 5070 26178
rect 5070 26126 5122 26178
rect 5122 26126 5124 26178
rect 5068 26124 5124 26126
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 3052 25506 3108 25508
rect 3052 25454 3054 25506
rect 3054 25454 3106 25506
rect 3106 25454 3108 25506
rect 3052 25452 3108 25454
rect 3948 25506 4004 25508
rect 3948 25454 3950 25506
rect 3950 25454 4002 25506
rect 4002 25454 4004 25506
rect 3948 25452 4004 25454
rect 5180 25676 5236 25732
rect 3612 25394 3668 25396
rect 3612 25342 3614 25394
rect 3614 25342 3666 25394
rect 3666 25342 3668 25394
rect 3612 25340 3668 25342
rect 4732 25506 4788 25508
rect 4732 25454 4734 25506
rect 4734 25454 4786 25506
rect 4786 25454 4788 25506
rect 4732 25452 4788 25454
rect 2940 25282 2996 25284
rect 2940 25230 2942 25282
rect 2942 25230 2994 25282
rect 2994 25230 2996 25282
rect 2940 25228 2996 25230
rect 3500 25282 3556 25284
rect 3500 25230 3502 25282
rect 3502 25230 3554 25282
rect 3554 25230 3556 25282
rect 3500 25228 3556 25230
rect 2716 24780 2772 24836
rect 2492 24610 2548 24612
rect 2492 24558 2494 24610
rect 2494 24558 2546 24610
rect 2546 24558 2548 24610
rect 2492 24556 2548 24558
rect 3276 23660 3332 23716
rect 5964 28364 6020 28420
rect 6636 28418 6692 28420
rect 6636 28366 6638 28418
rect 6638 28366 6690 28418
rect 6690 28366 6692 28418
rect 6636 28364 6692 28366
rect 7308 29932 7364 29988
rect 8316 30994 8372 30996
rect 8316 30942 8318 30994
rect 8318 30942 8370 30994
rect 8370 30942 8372 30994
rect 8316 30940 8372 30942
rect 7532 30098 7588 30100
rect 7532 30046 7534 30098
rect 7534 30046 7586 30098
rect 7586 30046 7588 30098
rect 7532 30044 7588 30046
rect 7868 29932 7924 29988
rect 8428 30098 8484 30100
rect 8428 30046 8430 30098
rect 8430 30046 8482 30098
rect 8482 30046 8484 30098
rect 8428 30044 8484 30046
rect 7644 29596 7700 29652
rect 7868 29484 7924 29540
rect 8092 28476 8148 28532
rect 8540 29484 8596 29540
rect 9212 30210 9268 30212
rect 9212 30158 9214 30210
rect 9214 30158 9266 30210
rect 9266 30158 9268 30210
rect 9212 30156 9268 30158
rect 8540 29314 8596 29316
rect 8540 29262 8542 29314
rect 8542 29262 8594 29314
rect 8594 29262 8596 29314
rect 8540 29260 8596 29262
rect 7084 28252 7140 28308
rect 6076 26908 6132 26964
rect 6860 26460 6916 26516
rect 5628 25452 5684 25508
rect 6748 25394 6804 25396
rect 6748 25342 6750 25394
rect 6750 25342 6802 25394
rect 6802 25342 6804 25394
rect 6748 25340 6804 25342
rect 6412 25282 6468 25284
rect 6412 25230 6414 25282
rect 6414 25230 6466 25282
rect 6466 25230 6468 25282
rect 6412 25228 6468 25230
rect 5180 24780 5236 24836
rect 4172 23660 4228 23716
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 5068 24610 5124 24612
rect 5068 24558 5070 24610
rect 5070 24558 5122 24610
rect 5122 24558 5124 24610
rect 5068 24556 5124 24558
rect 6748 23996 6804 24052
rect 6188 23884 6244 23940
rect 5852 23772 5908 23828
rect 3612 23548 3668 23604
rect 4508 23548 4564 23604
rect 2492 21756 2548 21812
rect 3388 22540 3444 22596
rect 2492 21420 2548 21476
rect 3500 21698 3556 21700
rect 3500 21646 3502 21698
rect 3502 21646 3554 21698
rect 3554 21646 3556 21698
rect 3500 21644 3556 21646
rect 4060 23154 4116 23156
rect 4060 23102 4062 23154
rect 4062 23102 4114 23154
rect 4114 23102 4116 23154
rect 4060 23100 4116 23102
rect 5628 23548 5684 23604
rect 3836 21810 3892 21812
rect 3836 21758 3838 21810
rect 3838 21758 3890 21810
rect 3890 21758 3892 21810
rect 3836 21756 3892 21758
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4620 22540 4676 22596
rect 5404 22540 5460 22596
rect 5628 23100 5684 23156
rect 5628 22370 5684 22372
rect 5628 22318 5630 22370
rect 5630 22318 5682 22370
rect 5682 22318 5684 22370
rect 5628 22316 5684 22318
rect 4956 22092 5012 22148
rect 4396 21644 4452 21700
rect 4284 21586 4340 21588
rect 4284 21534 4286 21586
rect 4286 21534 4338 21586
rect 4338 21534 4340 21586
rect 4284 21532 4340 21534
rect 5180 21586 5236 21588
rect 5180 21534 5182 21586
rect 5182 21534 5234 21586
rect 5234 21534 5236 21586
rect 5180 21532 5236 21534
rect 4732 21474 4788 21476
rect 4732 21422 4734 21474
rect 4734 21422 4786 21474
rect 4786 21422 4788 21474
rect 4732 21420 4788 21422
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 3276 20972 3332 21028
rect 4620 20972 4676 21028
rect 6076 22146 6132 22148
rect 6076 22094 6078 22146
rect 6078 22094 6130 22146
rect 6130 22094 6132 22146
rect 6076 22092 6132 22094
rect 5852 21586 5908 21588
rect 5852 21534 5854 21586
rect 5854 21534 5906 21586
rect 5906 21534 5908 21586
rect 5852 21532 5908 21534
rect 5740 20972 5796 21028
rect 4956 20524 5012 20580
rect 1820 19234 1876 19236
rect 1820 19182 1822 19234
rect 1822 19182 1874 19234
rect 1874 19182 1876 19234
rect 1820 19180 1876 19182
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 3388 19180 3444 19236
rect 2492 19122 2548 19124
rect 2492 19070 2494 19122
rect 2494 19070 2546 19122
rect 2546 19070 2548 19122
rect 2492 19068 2548 19070
rect 3612 18620 3668 18676
rect 3164 18450 3220 18452
rect 3164 18398 3166 18450
rect 3166 18398 3218 18450
rect 3218 18398 3220 18450
rect 3164 18396 3220 18398
rect 4508 19068 4564 19124
rect 4620 18674 4676 18676
rect 4620 18622 4622 18674
rect 4622 18622 4674 18674
rect 4674 18622 4676 18674
rect 4620 18620 4676 18622
rect 5292 19180 5348 19236
rect 4956 18396 5012 18452
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4060 17388 4116 17444
rect 3388 16994 3444 16996
rect 3388 16942 3390 16994
rect 3390 16942 3442 16994
rect 3442 16942 3444 16994
rect 3388 16940 3444 16942
rect 3724 16716 3780 16772
rect 4284 16882 4340 16884
rect 4284 16830 4286 16882
rect 4286 16830 4338 16882
rect 4338 16830 4340 16882
rect 4284 16828 4340 16830
rect 4396 16770 4452 16772
rect 4396 16718 4398 16770
rect 4398 16718 4450 16770
rect 4450 16718 4452 16770
rect 4396 16716 4452 16718
rect 4844 16994 4900 16996
rect 4844 16942 4846 16994
rect 4846 16942 4898 16994
rect 4898 16942 4900 16994
rect 4844 16940 4900 16942
rect 4620 16828 4676 16884
rect 3388 16098 3444 16100
rect 3388 16046 3390 16098
rect 3390 16046 3442 16098
rect 3442 16046 3444 16098
rect 3388 16044 3444 16046
rect 3836 16098 3892 16100
rect 3836 16046 3838 16098
rect 3838 16046 3890 16098
rect 3890 16046 3892 16098
rect 3836 16044 3892 16046
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4844 16380 4900 16436
rect 1820 15148 1876 15204
rect 2492 13132 2548 13188
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4396 14530 4452 14532
rect 4396 14478 4398 14530
rect 4398 14478 4450 14530
rect 4450 14478 4452 14530
rect 4396 14476 4452 14478
rect 5740 19180 5796 19236
rect 5628 19122 5684 19124
rect 5628 19070 5630 19122
rect 5630 19070 5682 19122
rect 5682 19070 5684 19122
rect 5628 19068 5684 19070
rect 5740 19010 5796 19012
rect 5740 18958 5742 19010
rect 5742 18958 5794 19010
rect 5794 18958 5796 19010
rect 5740 18956 5796 18958
rect 5628 18396 5684 18452
rect 5628 17442 5684 17444
rect 5628 17390 5630 17442
rect 5630 17390 5682 17442
rect 5682 17390 5684 17442
rect 5628 17388 5684 17390
rect 5404 16882 5460 16884
rect 5404 16830 5406 16882
rect 5406 16830 5458 16882
rect 5458 16830 5460 16882
rect 5404 16828 5460 16830
rect 5180 16380 5236 16436
rect 5852 16380 5908 16436
rect 5964 16044 6020 16100
rect 5516 15314 5572 15316
rect 5516 15262 5518 15314
rect 5518 15262 5570 15314
rect 5570 15262 5572 15314
rect 5516 15260 5572 15262
rect 6748 23548 6804 23604
rect 6300 22540 6356 22596
rect 6412 22370 6468 22372
rect 6412 22318 6414 22370
rect 6414 22318 6466 22370
rect 6466 22318 6468 22370
rect 6412 22316 6468 22318
rect 6972 25340 7028 25396
rect 6860 21810 6916 21812
rect 6860 21758 6862 21810
rect 6862 21758 6914 21810
rect 6914 21758 6916 21810
rect 6860 21756 6916 21758
rect 6524 19740 6580 19796
rect 7084 25228 7140 25284
rect 7308 25676 7364 25732
rect 9100 28530 9156 28532
rect 9100 28478 9102 28530
rect 9102 28478 9154 28530
rect 9154 28478 9156 28530
rect 9100 28476 9156 28478
rect 8316 28252 8372 28308
rect 8652 28028 8708 28084
rect 8204 27132 8260 27188
rect 8428 26514 8484 26516
rect 8428 26462 8430 26514
rect 8430 26462 8482 26514
rect 8482 26462 8484 26514
rect 8428 26460 8484 26462
rect 7644 25452 7700 25508
rect 7420 25394 7476 25396
rect 7420 25342 7422 25394
rect 7422 25342 7474 25394
rect 7474 25342 7476 25394
rect 7420 25340 7476 25342
rect 7756 25282 7812 25284
rect 7756 25230 7758 25282
rect 7758 25230 7810 25282
rect 7810 25230 7812 25282
rect 7756 25228 7812 25230
rect 7196 23884 7252 23940
rect 8540 25676 8596 25732
rect 8652 25452 8708 25508
rect 8092 25282 8148 25284
rect 8092 25230 8094 25282
rect 8094 25230 8146 25282
rect 8146 25230 8148 25282
rect 8092 25228 8148 25230
rect 7868 24780 7924 24836
rect 8316 24722 8372 24724
rect 8316 24670 8318 24722
rect 8318 24670 8370 24722
rect 8370 24670 8372 24722
rect 8316 24668 8372 24670
rect 8540 25228 8596 25284
rect 8316 23996 8372 24052
rect 7420 22370 7476 22372
rect 7420 22318 7422 22370
rect 7422 22318 7474 22370
rect 7474 22318 7476 22370
rect 7420 22316 7476 22318
rect 7420 21756 7476 21812
rect 7756 21644 7812 21700
rect 7532 21532 7588 21588
rect 7868 21308 7924 21364
rect 7420 19740 7476 19796
rect 6636 19010 6692 19012
rect 6636 18958 6638 19010
rect 6638 18958 6690 19010
rect 6690 18958 6692 19010
rect 6636 18956 6692 18958
rect 8204 21586 8260 21588
rect 8204 21534 8206 21586
rect 8206 21534 8258 21586
rect 8258 21534 8260 21586
rect 8204 21532 8260 21534
rect 8428 23826 8484 23828
rect 8428 23774 8430 23826
rect 8430 23774 8482 23826
rect 8482 23774 8484 23826
rect 8428 23772 8484 23774
rect 8988 28418 9044 28420
rect 8988 28366 8990 28418
rect 8990 28366 9042 28418
rect 9042 28366 9044 28418
rect 8988 28364 9044 28366
rect 8988 27186 9044 27188
rect 8988 27134 8990 27186
rect 8990 27134 9042 27186
rect 9042 27134 9044 27186
rect 8988 27132 9044 27134
rect 8876 25394 8932 25396
rect 8876 25342 8878 25394
rect 8878 25342 8930 25394
rect 8930 25342 8932 25394
rect 8876 25340 8932 25342
rect 8876 25116 8932 25172
rect 8652 23266 8708 23268
rect 8652 23214 8654 23266
rect 8654 23214 8706 23266
rect 8706 23214 8708 23266
rect 8652 23212 8708 23214
rect 8988 23938 9044 23940
rect 8988 23886 8990 23938
rect 8990 23886 9042 23938
rect 9042 23886 9044 23938
rect 8988 23884 9044 23886
rect 8540 21756 8596 21812
rect 8428 21698 8484 21700
rect 8428 21646 8430 21698
rect 8430 21646 8482 21698
rect 8482 21646 8484 21698
rect 8428 21644 8484 21646
rect 8204 21308 8260 21364
rect 9660 32450 9716 32452
rect 9660 32398 9662 32450
rect 9662 32398 9714 32450
rect 9714 32398 9716 32450
rect 9660 32396 9716 32398
rect 9548 30044 9604 30100
rect 10556 31778 10612 31780
rect 10556 31726 10558 31778
rect 10558 31726 10610 31778
rect 10610 31726 10612 31778
rect 10556 31724 10612 31726
rect 9884 31666 9940 31668
rect 9884 31614 9886 31666
rect 9886 31614 9938 31666
rect 9938 31614 9940 31666
rect 9884 31612 9940 31614
rect 11564 32396 11620 32452
rect 11116 31612 11172 31668
rect 10780 30940 10836 30996
rect 11564 30828 11620 30884
rect 9660 28588 9716 28644
rect 10780 28700 10836 28756
rect 9660 28082 9716 28084
rect 9660 28030 9662 28082
rect 9662 28030 9714 28082
rect 9714 28030 9716 28082
rect 9660 28028 9716 28030
rect 10332 28140 10388 28196
rect 9324 27804 9380 27860
rect 11004 28476 11060 28532
rect 10780 28140 10836 28196
rect 12460 38162 12516 38164
rect 12460 38110 12462 38162
rect 12462 38110 12514 38162
rect 12514 38110 12516 38162
rect 12460 38108 12516 38110
rect 12012 36204 12068 36260
rect 12236 38050 12292 38052
rect 12236 37998 12238 38050
rect 12238 37998 12290 38050
rect 12290 37998 12292 38050
rect 12236 37996 12292 37998
rect 13692 38050 13748 38052
rect 13692 37998 13694 38050
rect 13694 37998 13746 38050
rect 13746 37998 13748 38050
rect 13692 37996 13748 37998
rect 15372 39394 15428 39396
rect 15372 39342 15374 39394
rect 15374 39342 15426 39394
rect 15426 39342 15428 39394
rect 15372 39340 15428 39342
rect 15372 39004 15428 39060
rect 14364 38780 14420 38836
rect 14252 38722 14308 38724
rect 14252 38670 14254 38722
rect 14254 38670 14306 38722
rect 14306 38670 14308 38722
rect 14252 38668 14308 38670
rect 15932 38780 15988 38836
rect 16492 38332 16548 38388
rect 17836 41858 17892 41860
rect 17836 41806 17838 41858
rect 17838 41806 17890 41858
rect 17890 41806 17892 41858
rect 17836 41804 17892 41806
rect 17836 41132 17892 41188
rect 17948 40908 18004 40964
rect 18060 41356 18116 41412
rect 19516 44210 19572 44212
rect 19516 44158 19518 44210
rect 19518 44158 19570 44210
rect 19570 44158 19572 44210
rect 19516 44156 19572 44158
rect 20300 44156 20356 44212
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19404 43708 19460 43764
rect 20076 43426 20132 43428
rect 20076 43374 20078 43426
rect 20078 43374 20130 43426
rect 20130 43374 20132 43426
rect 20076 43372 20132 43374
rect 18508 42476 18564 42532
rect 18396 42140 18452 42196
rect 18732 42082 18788 42084
rect 18732 42030 18734 42082
rect 18734 42030 18786 42082
rect 18786 42030 18788 42082
rect 18732 42028 18788 42030
rect 18956 41970 19012 41972
rect 18956 41918 18958 41970
rect 18958 41918 19010 41970
rect 19010 41918 19012 41970
rect 18956 41916 19012 41918
rect 19404 42140 19460 42196
rect 21420 45106 21476 45108
rect 21420 45054 21422 45106
rect 21422 45054 21474 45106
rect 21474 45054 21476 45106
rect 21420 45052 21476 45054
rect 20860 44156 20916 44212
rect 21420 43708 21476 43764
rect 20636 43372 20692 43428
rect 20300 42812 20356 42868
rect 20188 42754 20244 42756
rect 20188 42702 20190 42754
rect 20190 42702 20242 42754
rect 20242 42702 20244 42754
rect 20188 42700 20244 42702
rect 20076 42588 20132 42644
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 20524 41580 20580 41636
rect 19852 41410 19908 41412
rect 19852 41358 19854 41410
rect 19854 41358 19906 41410
rect 19906 41358 19908 41410
rect 19852 41356 19908 41358
rect 19516 41186 19572 41188
rect 19516 41134 19518 41186
rect 19518 41134 19570 41186
rect 19570 41134 19572 41186
rect 19516 41132 19572 41134
rect 18284 39452 18340 39508
rect 18172 39340 18228 39396
rect 16828 38444 16884 38500
rect 17836 38722 17892 38724
rect 17836 38670 17838 38722
rect 17838 38670 17890 38722
rect 17890 38670 17892 38722
rect 17836 38668 17892 38670
rect 18396 39228 18452 39284
rect 16716 38220 16772 38276
rect 12572 36258 12628 36260
rect 12572 36206 12574 36258
rect 12574 36206 12626 36258
rect 12626 36206 12628 36258
rect 12572 36204 12628 36206
rect 13916 37154 13972 37156
rect 13916 37102 13918 37154
rect 13918 37102 13970 37154
rect 13970 37102 13972 37154
rect 13916 37100 13972 37102
rect 15148 37938 15204 37940
rect 15148 37886 15150 37938
rect 15150 37886 15202 37938
rect 15202 37886 15204 37938
rect 15148 37884 15204 37886
rect 16828 37266 16884 37268
rect 16828 37214 16830 37266
rect 16830 37214 16882 37266
rect 16882 37214 16884 37266
rect 16828 37212 16884 37214
rect 16604 36204 16660 36260
rect 13580 35308 13636 35364
rect 13468 35196 13524 35252
rect 12124 34748 12180 34804
rect 12460 34802 12516 34804
rect 12460 34750 12462 34802
rect 12462 34750 12514 34802
rect 12514 34750 12516 34802
rect 12460 34748 12516 34750
rect 12796 34802 12852 34804
rect 12796 34750 12798 34802
rect 12798 34750 12850 34802
rect 12850 34750 12852 34802
rect 12796 34748 12852 34750
rect 13244 34354 13300 34356
rect 13244 34302 13246 34354
rect 13246 34302 13298 34354
rect 13298 34302 13300 34354
rect 13244 34300 13300 34302
rect 14028 35308 14084 35364
rect 13804 34802 13860 34804
rect 13804 34750 13806 34802
rect 13806 34750 13858 34802
rect 13858 34750 13860 34802
rect 13804 34748 13860 34750
rect 13916 34690 13972 34692
rect 13916 34638 13918 34690
rect 13918 34638 13970 34690
rect 13970 34638 13972 34690
rect 13916 34636 13972 34638
rect 13692 34300 13748 34356
rect 13468 34242 13524 34244
rect 13468 34190 13470 34242
rect 13470 34190 13522 34242
rect 13522 34190 13524 34242
rect 13468 34188 13524 34190
rect 13356 34018 13412 34020
rect 13356 33966 13358 34018
rect 13358 33966 13410 34018
rect 13410 33966 13412 34018
rect 13356 33964 13412 33966
rect 12684 33852 12740 33908
rect 12460 33740 12516 33796
rect 13580 33458 13636 33460
rect 13580 33406 13582 33458
rect 13582 33406 13634 33458
rect 13634 33406 13636 33458
rect 13580 33404 13636 33406
rect 14700 34690 14756 34692
rect 14700 34638 14702 34690
rect 14702 34638 14754 34690
rect 14754 34638 14756 34690
rect 14700 34636 14756 34638
rect 14364 34300 14420 34356
rect 14140 34242 14196 34244
rect 14140 34190 14142 34242
rect 14142 34190 14194 34242
rect 14194 34190 14196 34242
rect 14140 34188 14196 34190
rect 14028 32732 14084 32788
rect 14140 33404 14196 33460
rect 13916 32562 13972 32564
rect 13916 32510 13918 32562
rect 13918 32510 13970 32562
rect 13970 32510 13972 32562
rect 13916 32508 13972 32510
rect 13244 32450 13300 32452
rect 13244 32398 13246 32450
rect 13246 32398 13298 32450
rect 13298 32398 13300 32450
rect 13244 32396 13300 32398
rect 13356 31836 13412 31892
rect 11788 31666 11844 31668
rect 11788 31614 11790 31666
rect 11790 31614 11842 31666
rect 11842 31614 11844 31666
rect 11788 31612 11844 31614
rect 12124 31612 12180 31668
rect 12124 30994 12180 30996
rect 12124 30942 12126 30994
rect 12126 30942 12178 30994
rect 12178 30942 12180 30994
rect 12124 30940 12180 30942
rect 12572 30882 12628 30884
rect 12572 30830 12574 30882
rect 12574 30830 12626 30882
rect 12626 30830 12628 30882
rect 12572 30828 12628 30830
rect 12124 30156 12180 30212
rect 12460 30268 12516 30324
rect 11340 28140 11396 28196
rect 10556 26514 10612 26516
rect 10556 26462 10558 26514
rect 10558 26462 10610 26514
rect 10610 26462 10612 26514
rect 10556 26460 10612 26462
rect 9324 25228 9380 25284
rect 9884 25282 9940 25284
rect 9884 25230 9886 25282
rect 9886 25230 9938 25282
rect 9938 25230 9940 25282
rect 9884 25228 9940 25230
rect 9436 25116 9492 25172
rect 9772 25116 9828 25172
rect 9884 24834 9940 24836
rect 9884 24782 9886 24834
rect 9886 24782 9938 24834
rect 9938 24782 9940 24834
rect 9884 24780 9940 24782
rect 10444 25452 10500 25508
rect 9996 24668 10052 24724
rect 11676 29314 11732 29316
rect 11676 29262 11678 29314
rect 11678 29262 11730 29314
rect 11730 29262 11732 29314
rect 11676 29260 11732 29262
rect 12012 28812 12068 28868
rect 11676 28754 11732 28756
rect 11676 28702 11678 28754
rect 11678 28702 11730 28754
rect 11730 28702 11732 28754
rect 11676 28700 11732 28702
rect 12908 29820 12964 29876
rect 12460 29426 12516 29428
rect 12460 29374 12462 29426
rect 12462 29374 12514 29426
rect 12514 29374 12516 29426
rect 12460 29372 12516 29374
rect 12684 28812 12740 28868
rect 12796 29260 12852 29316
rect 12460 28476 12516 28532
rect 13020 29932 13076 29988
rect 13132 28700 13188 28756
rect 11452 26460 11508 26516
rect 10332 25116 10388 25172
rect 11228 25282 11284 25284
rect 11228 25230 11230 25282
rect 11230 25230 11282 25282
rect 11282 25230 11284 25282
rect 11228 25228 11284 25230
rect 11116 25116 11172 25172
rect 10556 23996 10612 24052
rect 10892 23212 10948 23268
rect 10780 21586 10836 21588
rect 10780 21534 10782 21586
rect 10782 21534 10834 21586
rect 10834 21534 10836 21586
rect 10780 21532 10836 21534
rect 11452 21474 11508 21476
rect 11452 21422 11454 21474
rect 11454 21422 11506 21474
rect 11506 21422 11508 21474
rect 11452 21420 11508 21422
rect 9660 21308 9716 21364
rect 8204 19852 8260 19908
rect 8764 19794 8820 19796
rect 8764 19742 8766 19794
rect 8766 19742 8818 19794
rect 8818 19742 8820 19794
rect 8764 19740 8820 19742
rect 7644 18956 7700 19012
rect 8204 18956 8260 19012
rect 6972 18284 7028 18340
rect 6860 17388 6916 17444
rect 8988 19852 9044 19908
rect 10780 21026 10836 21028
rect 10780 20974 10782 21026
rect 10782 20974 10834 21026
rect 10834 20974 10836 21026
rect 10780 20972 10836 20974
rect 9772 20578 9828 20580
rect 9772 20526 9774 20578
rect 9774 20526 9826 20578
rect 9826 20526 9828 20578
rect 9772 20524 9828 20526
rect 10444 20578 10500 20580
rect 10444 20526 10446 20578
rect 10446 20526 10498 20578
rect 10498 20526 10500 20578
rect 10444 20524 10500 20526
rect 9772 20130 9828 20132
rect 9772 20078 9774 20130
rect 9774 20078 9826 20130
rect 9826 20078 9828 20130
rect 9772 20076 9828 20078
rect 12236 26236 12292 26292
rect 12908 26290 12964 26292
rect 12908 26238 12910 26290
rect 12910 26238 12962 26290
rect 12962 26238 12964 26290
rect 12908 26236 12964 26238
rect 11788 25340 11844 25396
rect 12236 25004 12292 25060
rect 12124 24050 12180 24052
rect 12124 23998 12126 24050
rect 12126 23998 12178 24050
rect 12178 23998 12180 24050
rect 12124 23996 12180 23998
rect 12460 23884 12516 23940
rect 12460 23100 12516 23156
rect 12796 21532 12852 21588
rect 10780 20076 10836 20132
rect 9996 20018 10052 20020
rect 9996 19966 9998 20018
rect 9998 19966 10050 20018
rect 10050 19966 10052 20018
rect 9996 19964 10052 19966
rect 11004 19964 11060 20020
rect 10444 19740 10500 19796
rect 10892 19852 10948 19908
rect 8876 18956 8932 19012
rect 10556 19628 10612 19684
rect 8316 18396 8372 18452
rect 8652 18338 8708 18340
rect 8652 18286 8654 18338
rect 8654 18286 8706 18338
rect 8706 18286 8708 18338
rect 8652 18284 8708 18286
rect 6412 16098 6468 16100
rect 6412 16046 6414 16098
rect 6414 16046 6466 16098
rect 6466 16046 6468 16098
rect 6412 16044 6468 16046
rect 6076 15148 6132 15204
rect 6412 15260 6468 15316
rect 6860 15314 6916 15316
rect 6860 15262 6862 15314
rect 6862 15262 6914 15314
rect 6914 15262 6916 15314
rect 6860 15260 6916 15262
rect 4956 14476 5012 14532
rect 3724 13186 3780 13188
rect 3724 13134 3726 13186
rect 3726 13134 3778 13186
rect 3778 13134 3780 13186
rect 3724 13132 3780 13134
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 3836 12850 3892 12852
rect 3836 12798 3838 12850
rect 3838 12798 3890 12850
rect 3890 12798 3892 12850
rect 3836 12796 3892 12798
rect 4284 12796 4340 12852
rect 2492 11452 2548 11508
rect 1708 10498 1764 10500
rect 1708 10446 1710 10498
rect 1710 10446 1762 10498
rect 1762 10446 1764 10498
rect 1708 10444 1764 10446
rect 3612 10444 3668 10500
rect 3500 10332 3556 10388
rect 3388 9826 3444 9828
rect 3388 9774 3390 9826
rect 3390 9774 3442 9826
rect 3442 9774 3444 9826
rect 3388 9772 3444 9774
rect 4732 12850 4788 12852
rect 4732 12798 4734 12850
rect 4734 12798 4786 12850
rect 4786 12798 4788 12850
rect 4732 12796 4788 12798
rect 4844 12684 4900 12740
rect 4620 12066 4676 12068
rect 4620 12014 4622 12066
rect 4622 12014 4674 12066
rect 4674 12014 4676 12066
rect 4620 12012 4676 12014
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4396 11506 4452 11508
rect 4396 11454 4398 11506
rect 4398 11454 4450 11506
rect 4450 11454 4452 11506
rect 4396 11452 4452 11454
rect 4620 11394 4676 11396
rect 4620 11342 4622 11394
rect 4622 11342 4674 11394
rect 4674 11342 4676 11394
rect 4620 11340 4676 11342
rect 5292 12908 5348 12964
rect 5628 12850 5684 12852
rect 5628 12798 5630 12850
rect 5630 12798 5682 12850
rect 5682 12798 5684 12850
rect 5628 12796 5684 12798
rect 5740 12738 5796 12740
rect 5740 12686 5742 12738
rect 5742 12686 5794 12738
rect 5794 12686 5796 12738
rect 5740 12684 5796 12686
rect 5068 11788 5124 11844
rect 5516 12012 5572 12068
rect 5516 11340 5572 11396
rect 5964 11788 6020 11844
rect 9884 18396 9940 18452
rect 9100 17442 9156 17444
rect 9100 17390 9102 17442
rect 9102 17390 9154 17442
rect 9154 17390 9156 17442
rect 9100 17388 9156 17390
rect 8876 16268 8932 16324
rect 9212 16828 9268 16884
rect 9212 16210 9268 16212
rect 9212 16158 9214 16210
rect 9214 16158 9266 16210
rect 9266 16158 9268 16210
rect 9212 16156 9268 16158
rect 9212 15484 9268 15540
rect 7308 15148 7364 15204
rect 7084 13746 7140 13748
rect 7084 13694 7086 13746
rect 7086 13694 7138 13746
rect 7138 13694 7140 13746
rect 7084 13692 7140 13694
rect 6300 12348 6356 12404
rect 6860 12962 6916 12964
rect 6860 12910 6862 12962
rect 6862 12910 6914 12962
rect 6914 12910 6916 12962
rect 6860 12908 6916 12910
rect 7084 13074 7140 13076
rect 7084 13022 7086 13074
rect 7086 13022 7138 13074
rect 7138 13022 7140 13074
rect 7084 13020 7140 13022
rect 9548 16322 9604 16324
rect 9548 16270 9550 16322
rect 9550 16270 9602 16322
rect 9602 16270 9604 16322
rect 9548 16268 9604 16270
rect 9772 16882 9828 16884
rect 9772 16830 9774 16882
rect 9774 16830 9826 16882
rect 9826 16830 9828 16882
rect 9772 16828 9828 16830
rect 10220 16882 10276 16884
rect 10220 16830 10222 16882
rect 10222 16830 10274 16882
rect 10274 16830 10276 16882
rect 10220 16828 10276 16830
rect 10108 16322 10164 16324
rect 10108 16270 10110 16322
rect 10110 16270 10162 16322
rect 10162 16270 10164 16322
rect 10108 16268 10164 16270
rect 9660 16156 9716 16212
rect 9772 15538 9828 15540
rect 9772 15486 9774 15538
rect 9774 15486 9826 15538
rect 9826 15486 9828 15538
rect 9772 15484 9828 15486
rect 12124 20076 12180 20132
rect 11452 19740 11508 19796
rect 12012 19740 12068 19796
rect 11452 18450 11508 18452
rect 11452 18398 11454 18450
rect 11454 18398 11506 18450
rect 11506 18398 11508 18450
rect 11452 18396 11508 18398
rect 12348 18396 12404 18452
rect 12012 17612 12068 17668
rect 11900 16940 11956 16996
rect 11228 16716 11284 16772
rect 11340 16882 11396 16884
rect 11340 16830 11342 16882
rect 11342 16830 11394 16882
rect 11394 16830 11396 16882
rect 11340 16828 11396 16830
rect 10780 16156 10836 16212
rect 10668 15538 10724 15540
rect 10668 15486 10670 15538
rect 10670 15486 10722 15538
rect 10722 15486 10724 15538
rect 10668 15484 10724 15486
rect 10556 15314 10612 15316
rect 10556 15262 10558 15314
rect 10558 15262 10610 15314
rect 10610 15262 10612 15314
rect 10556 15260 10612 15262
rect 9660 15202 9716 15204
rect 9660 15150 9662 15202
rect 9662 15150 9714 15202
rect 9714 15150 9716 15202
rect 9660 15148 9716 15150
rect 10444 15202 10500 15204
rect 10444 15150 10446 15202
rect 10446 15150 10498 15202
rect 10498 15150 10500 15202
rect 10444 15148 10500 15150
rect 7532 13746 7588 13748
rect 7532 13694 7534 13746
rect 7534 13694 7586 13746
rect 7586 13694 7588 13746
rect 7532 13692 7588 13694
rect 9100 13580 9156 13636
rect 7756 13074 7812 13076
rect 7756 13022 7758 13074
rect 7758 13022 7810 13074
rect 7810 13022 7812 13074
rect 7756 13020 7812 13022
rect 7308 12908 7364 12964
rect 7196 12684 7252 12740
rect 6972 12236 7028 12292
rect 3948 10556 4004 10612
rect 3836 10498 3892 10500
rect 3836 10446 3838 10498
rect 3838 10446 3890 10498
rect 3890 10446 3892 10498
rect 3836 10444 3892 10446
rect 3724 9772 3780 9828
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4396 9996 4452 10052
rect 5180 10556 5236 10612
rect 5068 10498 5124 10500
rect 5068 10446 5070 10498
rect 5070 10446 5122 10498
rect 5122 10446 5124 10498
rect 5068 10444 5124 10446
rect 4956 10386 5012 10388
rect 4956 10334 4958 10386
rect 4958 10334 5010 10386
rect 5010 10334 5012 10386
rect 4956 10332 5012 10334
rect 4844 9884 4900 9940
rect 5068 9996 5124 10052
rect 1820 8258 1876 8260
rect 1820 8206 1822 8258
rect 1822 8206 1874 8258
rect 1874 8206 1876 8258
rect 1820 8204 1876 8206
rect 2940 7420 2996 7476
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 5964 9996 6020 10052
rect 5628 9884 5684 9940
rect 6076 9212 6132 9268
rect 6412 9154 6468 9156
rect 6412 9102 6414 9154
rect 6414 9102 6466 9154
rect 6466 9102 6468 9154
rect 6412 9100 6468 9102
rect 6748 9884 6804 9940
rect 8316 12962 8372 12964
rect 8316 12910 8318 12962
rect 8318 12910 8370 12962
rect 8370 12910 8372 12962
rect 8316 12908 8372 12910
rect 8764 12908 8820 12964
rect 8092 12684 8148 12740
rect 8092 11282 8148 11284
rect 8092 11230 8094 11282
rect 8094 11230 8146 11282
rect 8146 11230 8148 11282
rect 8092 11228 8148 11230
rect 7196 10610 7252 10612
rect 7196 10558 7198 10610
rect 7198 10558 7250 10610
rect 7250 10558 7252 10610
rect 7196 10556 7252 10558
rect 9884 12402 9940 12404
rect 9884 12350 9886 12402
rect 9886 12350 9938 12402
rect 9938 12350 9940 12402
rect 9884 12348 9940 12350
rect 9548 12290 9604 12292
rect 9548 12238 9550 12290
rect 9550 12238 9602 12290
rect 9602 12238 9604 12290
rect 9548 12236 9604 12238
rect 9884 11564 9940 11620
rect 9548 11116 9604 11172
rect 9660 11228 9716 11284
rect 9548 10722 9604 10724
rect 9548 10670 9550 10722
rect 9550 10670 9602 10722
rect 9602 10670 9604 10722
rect 9548 10668 9604 10670
rect 10332 12348 10388 12404
rect 10444 11564 10500 11620
rect 11900 16770 11956 16772
rect 11900 16718 11902 16770
rect 11902 16718 11954 16770
rect 11954 16718 11956 16770
rect 11900 16716 11956 16718
rect 11788 16268 11844 16324
rect 12012 16044 12068 16100
rect 11788 15538 11844 15540
rect 11788 15486 11790 15538
rect 11790 15486 11842 15538
rect 11842 15486 11844 15538
rect 11788 15484 11844 15486
rect 11228 13244 11284 13300
rect 13580 31724 13636 31780
rect 14700 33964 14756 34020
rect 14588 33516 14644 33572
rect 15036 34018 15092 34020
rect 15036 33966 15038 34018
rect 15038 33966 15090 34018
rect 15090 33966 15092 34018
rect 15036 33964 15092 33966
rect 14812 33852 14868 33908
rect 16492 34636 16548 34692
rect 15148 33404 15204 33460
rect 15708 33516 15764 33572
rect 14812 32732 14868 32788
rect 13804 31666 13860 31668
rect 13804 31614 13806 31666
rect 13806 31614 13858 31666
rect 13858 31614 13860 31666
rect 13804 31612 13860 31614
rect 13692 31052 13748 31108
rect 15148 32786 15204 32788
rect 15148 32734 15150 32786
rect 15150 32734 15202 32786
rect 15202 32734 15204 32786
rect 15148 32732 15204 32734
rect 16156 33740 16212 33796
rect 14588 31778 14644 31780
rect 14588 31726 14590 31778
rect 14590 31726 14642 31778
rect 14642 31726 14644 31778
rect 14588 31724 14644 31726
rect 14364 31052 14420 31108
rect 14924 31106 14980 31108
rect 14924 31054 14926 31106
rect 14926 31054 14978 31106
rect 14978 31054 14980 31106
rect 14924 31052 14980 31054
rect 14140 30882 14196 30884
rect 14140 30830 14142 30882
rect 14142 30830 14194 30882
rect 14194 30830 14196 30882
rect 14140 30828 14196 30830
rect 14588 30882 14644 30884
rect 14588 30830 14590 30882
rect 14590 30830 14642 30882
rect 14642 30830 14644 30882
rect 14588 30828 14644 30830
rect 15372 32284 15428 32340
rect 15148 30882 15204 30884
rect 15148 30830 15150 30882
rect 15150 30830 15202 30882
rect 15202 30830 15204 30882
rect 15148 30828 15204 30830
rect 15596 30828 15652 30884
rect 13804 30322 13860 30324
rect 13804 30270 13806 30322
rect 13806 30270 13858 30322
rect 13858 30270 13860 30322
rect 13804 30268 13860 30270
rect 13692 29986 13748 29988
rect 13692 29934 13694 29986
rect 13694 29934 13746 29986
rect 13746 29934 13748 29986
rect 13692 29932 13748 29934
rect 13580 29426 13636 29428
rect 13580 29374 13582 29426
rect 13582 29374 13634 29426
rect 13634 29374 13636 29426
rect 13580 29372 13636 29374
rect 14588 29986 14644 29988
rect 14588 29934 14590 29986
rect 14590 29934 14642 29986
rect 14642 29934 14644 29986
rect 14588 29932 14644 29934
rect 14140 29820 14196 29876
rect 14252 29314 14308 29316
rect 14252 29262 14254 29314
rect 14254 29262 14306 29314
rect 14306 29262 14308 29314
rect 14252 29260 14308 29262
rect 13580 28812 13636 28868
rect 13804 28700 13860 28756
rect 13580 26908 13636 26964
rect 13692 28028 13748 28084
rect 14924 29260 14980 29316
rect 14924 28642 14980 28644
rect 14924 28590 14926 28642
rect 14926 28590 14978 28642
rect 14978 28590 14980 28642
rect 14924 28588 14980 28590
rect 14364 27580 14420 27636
rect 14924 27970 14980 27972
rect 14924 27918 14926 27970
rect 14926 27918 14978 27970
rect 14978 27918 14980 27970
rect 14924 27916 14980 27918
rect 16380 33404 16436 33460
rect 18060 37826 18116 37828
rect 18060 37774 18062 37826
rect 18062 37774 18114 37826
rect 18114 37774 18116 37826
rect 18060 37772 18116 37774
rect 17836 37490 17892 37492
rect 17836 37438 17838 37490
rect 17838 37438 17890 37490
rect 17890 37438 17892 37490
rect 17836 37436 17892 37438
rect 18396 37772 18452 37828
rect 18396 37212 18452 37268
rect 18172 37154 18228 37156
rect 18172 37102 18174 37154
rect 18174 37102 18226 37154
rect 18226 37102 18228 37154
rect 18172 37100 18228 37102
rect 17836 36876 17892 36932
rect 19068 40908 19124 40964
rect 18732 39788 18788 39844
rect 18844 39564 18900 39620
rect 18620 39452 18676 39508
rect 18844 39228 18900 39284
rect 21308 42866 21364 42868
rect 21308 42814 21310 42866
rect 21310 42814 21362 42866
rect 21362 42814 21364 42866
rect 21308 42812 21364 42814
rect 21084 41970 21140 41972
rect 21084 41918 21086 41970
rect 21086 41918 21138 41970
rect 21138 41918 21140 41970
rect 21084 41916 21140 41918
rect 20636 41244 20692 41300
rect 21420 41186 21476 41188
rect 21420 41134 21422 41186
rect 21422 41134 21474 41186
rect 21474 41134 21476 41186
rect 21420 41132 21476 41134
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 20524 40684 20580 40740
rect 19516 39788 19572 39844
rect 20188 40572 20244 40628
rect 20748 40236 20804 40292
rect 19740 39564 19796 39620
rect 20076 39618 20132 39620
rect 20076 39566 20078 39618
rect 20078 39566 20130 39618
rect 20130 39566 20132 39618
rect 20076 39564 20132 39566
rect 19628 39506 19684 39508
rect 19628 39454 19630 39506
rect 19630 39454 19682 39506
rect 19682 39454 19684 39506
rect 19628 39452 19684 39454
rect 19852 39340 19908 39396
rect 19836 39226 19892 39228
rect 18956 39116 19012 39172
rect 19516 39116 19572 39172
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 18844 38610 18900 38612
rect 18844 38558 18846 38610
rect 18846 38558 18898 38610
rect 18898 38558 18900 38610
rect 18844 38556 18900 38558
rect 18844 38050 18900 38052
rect 18844 37998 18846 38050
rect 18846 37998 18898 38050
rect 18898 37998 18900 38050
rect 18844 37996 18900 37998
rect 18620 37436 18676 37492
rect 18844 36876 18900 36932
rect 17836 36204 17892 36260
rect 17724 35586 17780 35588
rect 17724 35534 17726 35586
rect 17726 35534 17778 35586
rect 17778 35534 17780 35586
rect 17724 35532 17780 35534
rect 16940 32620 16996 32676
rect 17276 35308 17332 35364
rect 16828 32562 16884 32564
rect 16828 32510 16830 32562
rect 16830 32510 16882 32562
rect 16882 32510 16884 32562
rect 16828 32508 16884 32510
rect 16268 31218 16324 31220
rect 16268 31166 16270 31218
rect 16270 31166 16322 31218
rect 16322 31166 16324 31218
rect 16268 31164 16324 31166
rect 16044 30828 16100 30884
rect 18396 34972 18452 35028
rect 17724 33852 17780 33908
rect 17500 33404 17556 33460
rect 18060 33964 18116 34020
rect 17388 32338 17444 32340
rect 17388 32286 17390 32338
rect 17390 32286 17442 32338
rect 17442 32286 17444 32338
rect 17388 32284 17444 32286
rect 17836 32620 17892 32676
rect 18172 34130 18228 34132
rect 18172 34078 18174 34130
rect 18174 34078 18226 34130
rect 18226 34078 18228 34130
rect 18172 34076 18228 34078
rect 18620 34690 18676 34692
rect 18620 34638 18622 34690
rect 18622 34638 18674 34690
rect 18674 34638 18676 34690
rect 18620 34636 18676 34638
rect 18508 34076 18564 34132
rect 18284 33852 18340 33908
rect 18508 33740 18564 33796
rect 18732 34076 18788 34132
rect 19404 38444 19460 38500
rect 19404 38274 19460 38276
rect 19404 38222 19406 38274
rect 19406 38222 19458 38274
rect 19458 38222 19460 38274
rect 19404 38220 19460 38222
rect 19292 37938 19348 37940
rect 19292 37886 19294 37938
rect 19294 37886 19346 37938
rect 19346 37886 19348 37938
rect 19292 37884 19348 37886
rect 19852 39004 19908 39060
rect 20076 38780 20132 38836
rect 19628 38556 19684 38612
rect 19740 38050 19796 38052
rect 19740 37998 19742 38050
rect 19742 37998 19794 38050
rect 19794 37998 19796 38050
rect 19740 37996 19796 37998
rect 19628 37772 19684 37828
rect 20076 38556 20132 38612
rect 20300 38332 20356 38388
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19068 37266 19124 37268
rect 19068 37214 19070 37266
rect 19070 37214 19122 37266
rect 19122 37214 19124 37266
rect 19068 37212 19124 37214
rect 20076 37154 20132 37156
rect 20076 37102 20078 37154
rect 20078 37102 20130 37154
rect 20130 37102 20132 37154
rect 20076 37100 20132 37102
rect 19180 36428 19236 36484
rect 21196 40124 21252 40180
rect 20524 36482 20580 36484
rect 20524 36430 20526 36482
rect 20526 36430 20578 36482
rect 20578 36430 20580 36482
rect 20524 36428 20580 36430
rect 19964 36204 20020 36260
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 20300 35532 20356 35588
rect 19964 35026 20020 35028
rect 19964 34974 19966 35026
rect 19966 34974 20018 35026
rect 20018 34974 20020 35026
rect 19964 34972 20020 34974
rect 20860 36482 20916 36484
rect 20860 36430 20862 36482
rect 20862 36430 20914 36482
rect 20914 36430 20916 36482
rect 20860 36428 20916 36430
rect 20748 35196 20804 35252
rect 20300 35026 20356 35028
rect 20300 34974 20302 35026
rect 20302 34974 20354 35026
rect 20354 34974 20356 35026
rect 20300 34972 20356 34974
rect 18956 33852 19012 33908
rect 20860 34690 20916 34692
rect 20860 34638 20862 34690
rect 20862 34638 20914 34690
rect 20914 34638 20916 34690
rect 20860 34636 20916 34638
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19068 33740 19124 33796
rect 18396 32562 18452 32564
rect 18396 32510 18398 32562
rect 18398 32510 18450 32562
rect 18450 32510 18452 32562
rect 18396 32508 18452 32510
rect 16828 31164 16884 31220
rect 16380 30044 16436 30100
rect 16604 30828 16660 30884
rect 16044 29372 16100 29428
rect 15820 28082 15876 28084
rect 15820 28030 15822 28082
rect 15822 28030 15874 28082
rect 15874 28030 15876 28082
rect 15820 28028 15876 28030
rect 15932 27916 15988 27972
rect 15148 27356 15204 27412
rect 15148 27020 15204 27076
rect 14588 26962 14644 26964
rect 14588 26910 14590 26962
rect 14590 26910 14642 26962
rect 14642 26910 14644 26962
rect 14588 26908 14644 26910
rect 13468 26236 13524 26292
rect 14252 25394 14308 25396
rect 14252 25342 14254 25394
rect 14254 25342 14306 25394
rect 14306 25342 14308 25394
rect 14252 25340 14308 25342
rect 13356 24668 13412 24724
rect 13580 23938 13636 23940
rect 13580 23886 13582 23938
rect 13582 23886 13634 23938
rect 13634 23886 13636 23938
rect 13580 23884 13636 23886
rect 14364 23436 14420 23492
rect 14588 23378 14644 23380
rect 14588 23326 14590 23378
rect 14590 23326 14642 23378
rect 14642 23326 14644 23378
rect 14588 23324 14644 23326
rect 15932 27634 15988 27636
rect 15932 27582 15934 27634
rect 15934 27582 15986 27634
rect 15986 27582 15988 27634
rect 15932 27580 15988 27582
rect 15820 27020 15876 27076
rect 16380 29314 16436 29316
rect 16380 29262 16382 29314
rect 16382 29262 16434 29314
rect 16434 29262 16436 29314
rect 16380 29260 16436 29262
rect 16156 27746 16212 27748
rect 16156 27694 16158 27746
rect 16158 27694 16210 27746
rect 16210 27694 16212 27746
rect 16156 27692 16212 27694
rect 16828 29484 16884 29540
rect 17388 29372 17444 29428
rect 17724 29260 17780 29316
rect 17500 27916 17556 27972
rect 16828 27746 16884 27748
rect 16828 27694 16830 27746
rect 16830 27694 16882 27746
rect 16882 27694 16884 27746
rect 16828 27692 16884 27694
rect 16716 27580 16772 27636
rect 17500 27746 17556 27748
rect 17500 27694 17502 27746
rect 17502 27694 17554 27746
rect 17554 27694 17556 27746
rect 17500 27692 17556 27694
rect 17388 27634 17444 27636
rect 17388 27582 17390 27634
rect 17390 27582 17442 27634
rect 17442 27582 17444 27634
rect 17388 27580 17444 27582
rect 16268 26572 16324 26628
rect 16604 26514 16660 26516
rect 16604 26462 16606 26514
rect 16606 26462 16658 26514
rect 16658 26462 16660 26514
rect 16604 26460 16660 26462
rect 16380 26402 16436 26404
rect 16380 26350 16382 26402
rect 16382 26350 16434 26402
rect 16434 26350 16436 26402
rect 16380 26348 16436 26350
rect 16828 26290 16884 26292
rect 16828 26238 16830 26290
rect 16830 26238 16882 26290
rect 16882 26238 16884 26290
rect 16828 26236 16884 26238
rect 16380 25788 16436 25844
rect 16380 24946 16436 24948
rect 16380 24894 16382 24946
rect 16382 24894 16434 24946
rect 16434 24894 16436 24946
rect 16380 24892 16436 24894
rect 15260 23324 15316 23380
rect 13468 23266 13524 23268
rect 13468 23214 13470 23266
rect 13470 23214 13522 23266
rect 13522 23214 13524 23266
rect 13468 23212 13524 23214
rect 13692 22930 13748 22932
rect 13692 22878 13694 22930
rect 13694 22878 13746 22930
rect 13746 22878 13748 22930
rect 13692 22876 13748 22878
rect 13916 21474 13972 21476
rect 13916 21422 13918 21474
rect 13918 21422 13970 21474
rect 13970 21422 13972 21474
rect 13916 21420 13972 21422
rect 13580 20860 13636 20916
rect 14028 20748 14084 20804
rect 14924 23266 14980 23268
rect 14924 23214 14926 23266
rect 14926 23214 14978 23266
rect 14978 23214 14980 23266
rect 14924 23212 14980 23214
rect 14476 22876 14532 22932
rect 15484 23436 15540 23492
rect 16828 24610 16884 24612
rect 16828 24558 16830 24610
rect 16830 24558 16882 24610
rect 16882 24558 16884 24610
rect 16828 24556 16884 24558
rect 15484 22764 15540 22820
rect 15708 22482 15764 22484
rect 15708 22430 15710 22482
rect 15710 22430 15762 22482
rect 15762 22430 15764 22482
rect 15708 22428 15764 22430
rect 14140 21084 14196 21140
rect 14588 20860 14644 20916
rect 14700 21308 14756 21364
rect 14812 21084 14868 21140
rect 15484 21362 15540 21364
rect 15484 21310 15486 21362
rect 15486 21310 15538 21362
rect 15538 21310 15540 21362
rect 15484 21308 15540 21310
rect 14812 20802 14868 20804
rect 14812 20750 14814 20802
rect 14814 20750 14866 20802
rect 14866 20750 14868 20802
rect 14812 20748 14868 20750
rect 15148 20802 15204 20804
rect 15148 20750 15150 20802
rect 15150 20750 15202 20802
rect 15202 20750 15204 20802
rect 15148 20748 15204 20750
rect 13020 19628 13076 19684
rect 14588 20188 14644 20244
rect 12796 18396 12852 18452
rect 12908 16940 12964 16996
rect 12572 16268 12628 16324
rect 12348 16210 12404 16212
rect 12348 16158 12350 16210
rect 12350 16158 12402 16210
rect 12402 16158 12404 16210
rect 12348 16156 12404 16158
rect 13020 17612 13076 17668
rect 13804 19122 13860 19124
rect 13804 19070 13806 19122
rect 13806 19070 13858 19122
rect 13858 19070 13860 19122
rect 13804 19068 13860 19070
rect 13580 19010 13636 19012
rect 13580 18958 13582 19010
rect 13582 18958 13634 19010
rect 13634 18958 13636 19010
rect 13580 18956 13636 18958
rect 14364 19010 14420 19012
rect 14364 18958 14366 19010
rect 14366 18958 14418 19010
rect 14418 18958 14420 19010
rect 14364 18956 14420 18958
rect 16828 23938 16884 23940
rect 16828 23886 16830 23938
rect 16830 23886 16882 23938
rect 16882 23886 16884 23938
rect 16828 23884 16884 23886
rect 16380 22764 16436 22820
rect 16828 23212 16884 23268
rect 19180 33964 19236 34020
rect 19404 33628 19460 33684
rect 19516 34076 19572 34132
rect 19180 33180 19236 33236
rect 18620 31612 18676 31668
rect 18284 31052 18340 31108
rect 18732 30098 18788 30100
rect 18732 30046 18734 30098
rect 18734 30046 18786 30098
rect 18786 30046 18788 30098
rect 18732 30044 18788 30046
rect 18172 29596 18228 29652
rect 18508 29484 18564 29540
rect 17948 28812 18004 28868
rect 18060 28700 18116 28756
rect 17836 26348 17892 26404
rect 17388 26236 17444 26292
rect 17948 25788 18004 25844
rect 17500 25506 17556 25508
rect 17500 25454 17502 25506
rect 17502 25454 17554 25506
rect 17554 25454 17556 25506
rect 17500 25452 17556 25454
rect 17612 23826 17668 23828
rect 17612 23774 17614 23826
rect 17614 23774 17666 23826
rect 17666 23774 17668 23826
rect 17612 23772 17668 23774
rect 18172 23996 18228 24052
rect 18060 23884 18116 23940
rect 17500 23100 17556 23156
rect 17276 22428 17332 22484
rect 16716 22146 16772 22148
rect 16716 22094 16718 22146
rect 16718 22094 16770 22146
rect 16770 22094 16772 22146
rect 16716 22092 16772 22094
rect 16604 21644 16660 21700
rect 16380 21586 16436 21588
rect 16380 21534 16382 21586
rect 16382 21534 16434 21586
rect 16434 21534 16436 21586
rect 16380 21532 16436 21534
rect 16156 21420 16212 21476
rect 16492 21308 16548 21364
rect 15596 20076 15652 20132
rect 15932 19852 15988 19908
rect 16380 19852 16436 19908
rect 14812 19122 14868 19124
rect 14812 19070 14814 19122
rect 14814 19070 14866 19122
rect 14866 19070 14868 19122
rect 14812 19068 14868 19070
rect 14140 17778 14196 17780
rect 14140 17726 14142 17778
rect 14142 17726 14194 17778
rect 14194 17726 14196 17778
rect 14140 17724 14196 17726
rect 13916 16828 13972 16884
rect 13580 16098 13636 16100
rect 13580 16046 13582 16098
rect 13582 16046 13634 16098
rect 13634 16046 13636 16098
rect 13580 16044 13636 16046
rect 15484 18956 15540 19012
rect 15708 17724 15764 17780
rect 15932 18226 15988 18228
rect 15932 18174 15934 18226
rect 15934 18174 15986 18226
rect 15986 18174 15988 18226
rect 15932 18172 15988 18174
rect 16156 17612 16212 17668
rect 16268 17554 16324 17556
rect 16268 17502 16270 17554
rect 16270 17502 16322 17554
rect 16322 17502 16324 17554
rect 16268 17500 16324 17502
rect 16156 17052 16212 17108
rect 15596 16882 15652 16884
rect 15596 16830 15598 16882
rect 15598 16830 15650 16882
rect 15650 16830 15652 16882
rect 15596 16828 15652 16830
rect 15148 16098 15204 16100
rect 15148 16046 15150 16098
rect 15150 16046 15202 16098
rect 15202 16046 15204 16098
rect 15148 16044 15204 16046
rect 14476 15874 14532 15876
rect 14476 15822 14478 15874
rect 14478 15822 14530 15874
rect 14530 15822 14532 15874
rect 14476 15820 14532 15822
rect 12572 14418 12628 14420
rect 12572 14366 12574 14418
rect 12574 14366 12626 14418
rect 12626 14366 12628 14418
rect 12572 14364 12628 14366
rect 12012 13634 12068 13636
rect 12012 13582 12014 13634
rect 12014 13582 12066 13634
rect 12066 13582 12068 13634
rect 12012 13580 12068 13582
rect 11676 13244 11732 13300
rect 12236 14140 12292 14196
rect 12124 13074 12180 13076
rect 12124 13022 12126 13074
rect 12126 13022 12178 13074
rect 12178 13022 12180 13074
rect 12124 13020 12180 13022
rect 9996 11116 10052 11172
rect 10668 11170 10724 11172
rect 10668 11118 10670 11170
rect 10670 11118 10722 11170
rect 10722 11118 10724 11170
rect 10668 11116 10724 11118
rect 10892 11564 10948 11620
rect 10108 10780 10164 10836
rect 9996 10556 10052 10612
rect 7196 9884 7252 9940
rect 8540 9938 8596 9940
rect 8540 9886 8542 9938
rect 8542 9886 8594 9938
rect 8594 9886 8596 9938
rect 8540 9884 8596 9886
rect 7196 9154 7252 9156
rect 7196 9102 7198 9154
rect 7198 9102 7250 9154
rect 7250 9102 7252 9154
rect 7196 9100 7252 9102
rect 7308 9212 7364 9268
rect 7756 8818 7812 8820
rect 7756 8766 7758 8818
rect 7758 8766 7810 8818
rect 7810 8766 7812 8818
rect 7756 8764 7812 8766
rect 8540 8764 8596 8820
rect 4172 7532 4228 7588
rect 3388 7420 3444 7476
rect 4060 7420 4116 7476
rect 2492 6076 2548 6132
rect 5068 7532 5124 7588
rect 4396 7474 4452 7476
rect 4396 7422 4398 7474
rect 4398 7422 4450 7474
rect 4450 7422 4452 7474
rect 4396 7420 4452 7422
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4732 6524 4788 6580
rect 5516 8204 5572 8260
rect 6748 6748 6804 6804
rect 5628 6578 5684 6580
rect 5628 6526 5630 6578
rect 5630 6526 5682 6578
rect 5682 6526 5684 6578
rect 5628 6524 5684 6526
rect 5404 6412 5460 6468
rect 5180 6130 5236 6132
rect 5180 6078 5182 6130
rect 5182 6078 5234 6130
rect 5234 6078 5236 6130
rect 5180 6076 5236 6078
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 6300 6412 6356 6468
rect 5964 6188 6020 6244
rect 1820 4956 1876 5012
rect 4172 4956 4228 5012
rect 6636 6188 6692 6244
rect 6524 5906 6580 5908
rect 6524 5854 6526 5906
rect 6526 5854 6578 5906
rect 6578 5854 6580 5906
rect 6524 5852 6580 5854
rect 7196 6466 7252 6468
rect 7196 6414 7198 6466
rect 7198 6414 7250 6466
rect 7250 6414 7252 6466
rect 7196 6412 7252 6414
rect 7084 5852 7140 5908
rect 7420 6188 7476 6244
rect 7868 6076 7924 6132
rect 7980 6188 8036 6244
rect 4956 4226 5012 4228
rect 4956 4174 4958 4226
rect 4958 4174 5010 4226
rect 5010 4174 5012 4226
rect 4956 4172 5012 4174
rect 7868 5906 7924 5908
rect 7868 5854 7870 5906
rect 7870 5854 7922 5906
rect 7922 5854 7924 5906
rect 7868 5852 7924 5854
rect 8204 7420 8260 7476
rect 8204 6748 8260 6804
rect 8316 6188 8372 6244
rect 8988 8092 9044 8148
rect 9660 7474 9716 7476
rect 9660 7422 9662 7474
rect 9662 7422 9714 7474
rect 9714 7422 9716 7474
rect 9660 7420 9716 7422
rect 8876 7362 8932 7364
rect 8876 7310 8878 7362
rect 8878 7310 8930 7362
rect 8930 7310 8932 7362
rect 8876 7308 8932 7310
rect 8988 6748 9044 6804
rect 8764 6130 8820 6132
rect 8764 6078 8766 6130
rect 8766 6078 8818 6130
rect 8818 6078 8820 6130
rect 8764 6076 8820 6078
rect 9660 5852 9716 5908
rect 8764 5740 8820 5796
rect 10332 10556 10388 10612
rect 11116 11394 11172 11396
rect 11116 11342 11118 11394
rect 11118 11342 11170 11394
rect 11170 11342 11172 11394
rect 11116 11340 11172 11342
rect 11004 10780 11060 10836
rect 11116 10668 11172 10724
rect 10892 10556 10948 10612
rect 10444 9548 10500 9604
rect 10332 7362 10388 7364
rect 10332 7310 10334 7362
rect 10334 7310 10386 7362
rect 10386 7310 10388 7362
rect 10332 7308 10388 7310
rect 11004 9660 11060 9716
rect 10780 9602 10836 9604
rect 10780 9550 10782 9602
rect 10782 9550 10834 9602
rect 10834 9550 10836 9602
rect 10780 9548 10836 9550
rect 13468 14418 13524 14420
rect 13468 14366 13470 14418
rect 13470 14366 13522 14418
rect 13522 14366 13524 14418
rect 13468 14364 13524 14366
rect 14028 14364 14084 14420
rect 12908 14306 12964 14308
rect 12908 14254 12910 14306
rect 12910 14254 12962 14306
rect 12962 14254 12964 14306
rect 12908 14252 12964 14254
rect 14924 14364 14980 14420
rect 14700 14252 14756 14308
rect 13804 13634 13860 13636
rect 13804 13582 13806 13634
rect 13806 13582 13858 13634
rect 13858 13582 13860 13634
rect 13804 13580 13860 13582
rect 11340 12402 11396 12404
rect 11340 12350 11342 12402
rect 11342 12350 11394 12402
rect 11394 12350 11396 12402
rect 11340 12348 11396 12350
rect 11676 12290 11732 12292
rect 11676 12238 11678 12290
rect 11678 12238 11730 12290
rect 11730 12238 11732 12290
rect 11676 12236 11732 12238
rect 12012 12124 12068 12180
rect 11676 11676 11732 11732
rect 11564 11282 11620 11284
rect 11564 11230 11566 11282
rect 11566 11230 11618 11282
rect 11618 11230 11620 11282
rect 11564 11228 11620 11230
rect 10444 6748 10500 6804
rect 10780 7532 10836 7588
rect 10220 6076 10276 6132
rect 11228 8146 11284 8148
rect 11228 8094 11230 8146
rect 11230 8094 11282 8146
rect 11282 8094 11284 8146
rect 11228 8092 11284 8094
rect 12684 12236 12740 12292
rect 13356 12066 13412 12068
rect 13356 12014 13358 12066
rect 13358 12014 13410 12066
rect 13410 12014 13412 12066
rect 13356 12012 13412 12014
rect 15484 14588 15540 14644
rect 15260 13692 15316 13748
rect 14028 12012 14084 12068
rect 15260 12796 15316 12852
rect 15708 15820 15764 15876
rect 15708 14588 15764 14644
rect 15596 12796 15652 12852
rect 12124 11394 12180 11396
rect 12124 11342 12126 11394
rect 12126 11342 12178 11394
rect 12178 11342 12180 11394
rect 12124 11340 12180 11342
rect 12236 11282 12292 11284
rect 12236 11230 12238 11282
rect 12238 11230 12290 11282
rect 12290 11230 12292 11282
rect 12236 11228 12292 11230
rect 12236 10610 12292 10612
rect 12236 10558 12238 10610
rect 12238 10558 12290 10610
rect 12290 10558 12292 10610
rect 12236 10556 12292 10558
rect 12684 10610 12740 10612
rect 12684 10558 12686 10610
rect 12686 10558 12738 10610
rect 12738 10558 12740 10610
rect 12684 10556 12740 10558
rect 12460 9996 12516 10052
rect 12572 9660 12628 9716
rect 12124 8428 12180 8484
rect 11900 8258 11956 8260
rect 11900 8206 11902 8258
rect 11902 8206 11954 8258
rect 11954 8206 11956 8258
rect 11900 8204 11956 8206
rect 11564 7420 11620 7476
rect 11116 6802 11172 6804
rect 11116 6750 11118 6802
rect 11118 6750 11170 6802
rect 11170 6750 11172 6802
rect 11116 6748 11172 6750
rect 12460 8204 12516 8260
rect 12124 6748 12180 6804
rect 11228 6636 11284 6692
rect 13804 11676 13860 11732
rect 13132 10108 13188 10164
rect 13580 10050 13636 10052
rect 13580 9998 13582 10050
rect 13582 9998 13634 10050
rect 13634 9998 13636 10050
rect 13580 9996 13636 9998
rect 13580 8482 13636 8484
rect 13580 8430 13582 8482
rect 13582 8430 13634 8482
rect 13634 8430 13636 8482
rect 13580 8428 13636 8430
rect 13804 8428 13860 8484
rect 12908 8258 12964 8260
rect 12908 8206 12910 8258
rect 12910 8206 12962 8258
rect 12962 8206 12964 8258
rect 12908 8204 12964 8206
rect 13692 8258 13748 8260
rect 13692 8206 13694 8258
rect 13694 8206 13746 8258
rect 13746 8206 13748 8258
rect 13692 8204 13748 8206
rect 12796 7586 12852 7588
rect 12796 7534 12798 7586
rect 12798 7534 12850 7586
rect 12850 7534 12852 7586
rect 12796 7532 12852 7534
rect 13356 6748 13412 6804
rect 16268 13074 16324 13076
rect 16268 13022 16270 13074
rect 16270 13022 16322 13074
rect 16322 13022 16324 13074
rect 16268 13020 16324 13022
rect 15596 11900 15652 11956
rect 16268 11676 16324 11732
rect 15372 11394 15428 11396
rect 15372 11342 15374 11394
rect 15374 11342 15426 11394
rect 15426 11342 15428 11394
rect 15372 11340 15428 11342
rect 15596 11282 15652 11284
rect 15596 11230 15598 11282
rect 15598 11230 15650 11282
rect 15650 11230 15652 11282
rect 15596 11228 15652 11230
rect 15372 10556 15428 10612
rect 14140 8428 14196 8484
rect 14588 7980 14644 8036
rect 15596 6636 15652 6692
rect 8988 4450 9044 4452
rect 8988 4398 8990 4450
rect 8990 4398 9042 4450
rect 9042 4398 9044 4450
rect 8988 4396 9044 4398
rect 11004 4450 11060 4452
rect 11004 4398 11006 4450
rect 11006 4398 11058 4450
rect 11058 4398 11060 4450
rect 11004 4396 11060 4398
rect 12908 4284 12964 4340
rect 14252 6578 14308 6580
rect 14252 6526 14254 6578
rect 14254 6526 14306 6578
rect 14306 6526 14308 6578
rect 14252 6524 14308 6526
rect 15036 5964 15092 6020
rect 16940 21084 16996 21140
rect 17836 22482 17892 22484
rect 17836 22430 17838 22482
rect 17838 22430 17890 22482
rect 17890 22430 17892 22482
rect 17836 22428 17892 22430
rect 17164 20972 17220 21028
rect 17500 21196 17556 21252
rect 16604 20524 16660 20580
rect 16828 20188 16884 20244
rect 16940 18338 16996 18340
rect 16940 18286 16942 18338
rect 16942 18286 16994 18338
rect 16994 18286 16996 18338
rect 16940 18284 16996 18286
rect 17500 18172 17556 18228
rect 17612 17612 17668 17668
rect 17500 17554 17556 17556
rect 17500 17502 17502 17554
rect 17502 17502 17554 17554
rect 17554 17502 17556 17554
rect 17500 17500 17556 17502
rect 17388 17052 17444 17108
rect 18060 21196 18116 21252
rect 18284 22764 18340 22820
rect 18396 21308 18452 21364
rect 19180 30044 19236 30100
rect 18956 29650 19012 29652
rect 18956 29598 18958 29650
rect 18958 29598 19010 29650
rect 19010 29598 19012 29650
rect 18956 29596 19012 29598
rect 18844 29484 18900 29540
rect 20076 33628 20132 33684
rect 20188 33404 20244 33460
rect 20412 33852 20468 33908
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 20860 33628 20916 33684
rect 20636 31778 20692 31780
rect 20636 31726 20638 31778
rect 20638 31726 20690 31778
rect 20690 31726 20692 31778
rect 20636 31724 20692 31726
rect 19628 31612 19684 31668
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 20748 31106 20804 31108
rect 20748 31054 20750 31106
rect 20750 31054 20802 31106
rect 20802 31054 20804 31106
rect 20748 31052 20804 31054
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19180 28754 19236 28756
rect 19180 28702 19182 28754
rect 19182 28702 19234 28754
rect 19234 28702 19236 28754
rect 19180 28700 19236 28702
rect 19740 28812 19796 28868
rect 18844 28588 18900 28644
rect 18620 28364 18676 28420
rect 19292 28588 19348 28644
rect 19068 28476 19124 28532
rect 20748 30210 20804 30212
rect 20748 30158 20750 30210
rect 20750 30158 20802 30210
rect 20802 30158 20804 30210
rect 20748 30156 20804 30158
rect 19964 28530 20020 28532
rect 19964 28478 19966 28530
rect 19966 28478 20018 28530
rect 20018 28478 20020 28530
rect 19964 28476 20020 28478
rect 19516 28364 19572 28420
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 18956 27746 19012 27748
rect 18956 27694 18958 27746
rect 18958 27694 19010 27746
rect 19010 27694 19012 27746
rect 18956 27692 19012 27694
rect 18620 26908 18676 26964
rect 18732 27020 18788 27076
rect 20636 28812 20692 28868
rect 20300 28476 20356 28532
rect 20412 27804 20468 27860
rect 20412 27186 20468 27188
rect 20412 27134 20414 27186
rect 20414 27134 20466 27186
rect 20466 27134 20468 27186
rect 20412 27132 20468 27134
rect 18620 26572 18676 26628
rect 19964 26850 20020 26852
rect 19964 26798 19966 26850
rect 19966 26798 20018 26850
rect 20018 26798 20020 26850
rect 19964 26796 20020 26798
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19068 26460 19124 26516
rect 18620 26290 18676 26292
rect 18620 26238 18622 26290
rect 18622 26238 18674 26290
rect 18674 26238 18676 26290
rect 18620 26236 18676 26238
rect 19068 26124 19124 26180
rect 19516 24780 19572 24836
rect 19516 24610 19572 24612
rect 19516 24558 19518 24610
rect 19518 24558 19570 24610
rect 19570 24558 19572 24610
rect 19516 24556 19572 24558
rect 21084 39452 21140 39508
rect 21420 40684 21476 40740
rect 21644 42924 21700 42980
rect 23212 45106 23268 45108
rect 23212 45054 23214 45106
rect 23214 45054 23266 45106
rect 23266 45054 23268 45106
rect 23212 45052 23268 45054
rect 22316 43260 22372 43316
rect 22204 42812 22260 42868
rect 22092 42588 22148 42644
rect 21756 41020 21812 41076
rect 21532 40348 21588 40404
rect 21308 38834 21364 38836
rect 21308 38782 21310 38834
rect 21310 38782 21362 38834
rect 21362 38782 21364 38834
rect 21308 38780 21364 38782
rect 21196 38668 21252 38724
rect 21084 38444 21140 38500
rect 21420 38444 21476 38500
rect 21644 40124 21700 40180
rect 22540 44380 22596 44436
rect 24668 45724 24724 45780
rect 24556 44994 24612 44996
rect 24556 44942 24558 44994
rect 24558 44942 24610 44994
rect 24610 44942 24612 44994
rect 24556 44940 24612 44942
rect 24556 44210 24612 44212
rect 24556 44158 24558 44210
rect 24558 44158 24610 44210
rect 24610 44158 24612 44210
rect 24556 44156 24612 44158
rect 22764 41244 22820 41300
rect 22764 40684 22820 40740
rect 23548 43036 23604 43092
rect 24332 43650 24388 43652
rect 24332 43598 24334 43650
rect 24334 43598 24386 43650
rect 24386 43598 24388 43650
rect 24332 43596 24388 43598
rect 23884 42812 23940 42868
rect 24220 43426 24276 43428
rect 24220 43374 24222 43426
rect 24222 43374 24274 43426
rect 24274 43374 24276 43426
rect 24220 43372 24276 43374
rect 25228 45106 25284 45108
rect 25228 45054 25230 45106
rect 25230 45054 25282 45106
rect 25282 45054 25284 45106
rect 25228 45052 25284 45054
rect 24332 43260 24388 43316
rect 24108 43148 24164 43204
rect 23996 42754 24052 42756
rect 23996 42702 23998 42754
rect 23998 42702 24050 42754
rect 24050 42702 24052 42754
rect 23996 42700 24052 42702
rect 23548 42588 23604 42644
rect 23996 41020 24052 41076
rect 24556 42978 24612 42980
rect 24556 42926 24558 42978
rect 24558 42926 24610 42978
rect 24610 42926 24612 42978
rect 24556 42924 24612 42926
rect 25676 45106 25732 45108
rect 25676 45054 25678 45106
rect 25678 45054 25730 45106
rect 25730 45054 25732 45106
rect 25676 45052 25732 45054
rect 25564 44994 25620 44996
rect 25564 44942 25566 44994
rect 25566 44942 25618 44994
rect 25618 44942 25620 44994
rect 25564 44940 25620 44942
rect 26348 45106 26404 45108
rect 26348 45054 26350 45106
rect 26350 45054 26402 45106
rect 26402 45054 26404 45106
rect 26348 45052 26404 45054
rect 24668 42754 24724 42756
rect 24668 42702 24670 42754
rect 24670 42702 24722 42754
rect 24722 42702 24724 42754
rect 24668 42700 24724 42702
rect 24780 43260 24836 43316
rect 24556 42642 24612 42644
rect 24556 42590 24558 42642
rect 24558 42590 24610 42642
rect 24610 42590 24612 42642
rect 24556 42588 24612 42590
rect 24668 42140 24724 42196
rect 24556 42028 24612 42084
rect 24444 40626 24500 40628
rect 24444 40574 24446 40626
rect 24446 40574 24498 40626
rect 24498 40574 24500 40626
rect 24444 40572 24500 40574
rect 25676 43538 25732 43540
rect 25676 43486 25678 43538
rect 25678 43486 25730 43538
rect 25730 43486 25732 43538
rect 25676 43484 25732 43486
rect 25452 43148 25508 43204
rect 24892 42812 24948 42868
rect 25004 42530 25060 42532
rect 25004 42478 25006 42530
rect 25006 42478 25058 42530
rect 25058 42478 25060 42530
rect 25004 42476 25060 42478
rect 26348 43538 26404 43540
rect 26348 43486 26350 43538
rect 26350 43486 26402 43538
rect 26402 43486 26404 43538
rect 26348 43484 26404 43486
rect 25788 43260 25844 43316
rect 25564 42028 25620 42084
rect 26460 42642 26516 42644
rect 26460 42590 26462 42642
rect 26462 42590 26514 42642
rect 26514 42590 26516 42642
rect 26460 42588 26516 42590
rect 25788 41916 25844 41972
rect 24780 40460 24836 40516
rect 24220 40402 24276 40404
rect 24220 40350 24222 40402
rect 24222 40350 24274 40402
rect 24274 40350 24276 40402
rect 24220 40348 24276 40350
rect 21756 39116 21812 39172
rect 22540 39116 22596 39172
rect 22316 39004 22372 39060
rect 22204 38780 22260 38836
rect 20972 31836 21028 31892
rect 21644 36988 21700 37044
rect 23212 38834 23268 38836
rect 23212 38782 23214 38834
rect 23214 38782 23266 38834
rect 23266 38782 23268 38834
rect 23212 38780 23268 38782
rect 24444 39004 24500 39060
rect 23996 38668 24052 38724
rect 23884 37378 23940 37380
rect 23884 37326 23886 37378
rect 23886 37326 23938 37378
rect 23938 37326 23940 37378
rect 23884 37324 23940 37326
rect 24780 37996 24836 38052
rect 21868 37100 21924 37156
rect 21532 36482 21588 36484
rect 21532 36430 21534 36482
rect 21534 36430 21586 36482
rect 21586 36430 21588 36482
rect 21532 36428 21588 36430
rect 21756 35532 21812 35588
rect 21532 35196 21588 35252
rect 21308 33404 21364 33460
rect 22540 36876 22596 36932
rect 22764 36988 22820 37044
rect 21980 35084 22036 35140
rect 22316 35532 22372 35588
rect 22204 34972 22260 35028
rect 21868 33516 21924 33572
rect 21980 34636 22036 34692
rect 21308 33234 21364 33236
rect 21308 33182 21310 33234
rect 21310 33182 21362 33234
rect 21362 33182 21364 33234
rect 21308 33180 21364 33182
rect 21420 31836 21476 31892
rect 21308 31666 21364 31668
rect 21308 31614 21310 31666
rect 21310 31614 21362 31666
rect 21362 31614 21364 31666
rect 21308 31612 21364 31614
rect 21196 31164 21252 31220
rect 21644 31666 21700 31668
rect 21644 31614 21646 31666
rect 21646 31614 21698 31666
rect 21698 31614 21700 31666
rect 21644 31612 21700 31614
rect 21420 31276 21476 31332
rect 21868 31164 21924 31220
rect 21308 30156 21364 30212
rect 21532 29260 21588 29316
rect 21420 28700 21476 28756
rect 21644 28530 21700 28532
rect 21644 28478 21646 28530
rect 21646 28478 21698 28530
rect 21698 28478 21700 28530
rect 21644 28476 21700 28478
rect 21420 27804 21476 27860
rect 20972 27244 21028 27300
rect 21084 27132 21140 27188
rect 21756 27858 21812 27860
rect 21756 27806 21758 27858
rect 21758 27806 21810 27858
rect 21810 27806 21812 27858
rect 21756 27804 21812 27806
rect 20748 26236 20804 26292
rect 20188 25452 20244 25508
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20300 24780 20356 24836
rect 19740 24444 19796 24500
rect 18620 23266 18676 23268
rect 18620 23214 18622 23266
rect 18622 23214 18674 23266
rect 18674 23214 18676 23266
rect 18620 23212 18676 23214
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19964 22258 20020 22260
rect 19964 22206 19966 22258
rect 19966 22206 20018 22258
rect 20018 22206 20020 22258
rect 19964 22204 20020 22206
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20636 24444 20692 24500
rect 20412 23212 20468 23268
rect 20412 22428 20468 22484
rect 19852 21644 19908 21700
rect 19740 21084 19796 21140
rect 19292 21026 19348 21028
rect 19292 20974 19294 21026
rect 19294 20974 19346 21026
rect 19346 20974 19348 21026
rect 19292 20972 19348 20974
rect 18956 20636 19012 20692
rect 19740 20524 19796 20580
rect 19964 21532 20020 21588
rect 18844 20018 18900 20020
rect 18844 19966 18846 20018
rect 18846 19966 18898 20018
rect 18898 19966 18900 20018
rect 18844 19964 18900 19966
rect 18508 18620 18564 18676
rect 17836 18450 17892 18452
rect 17836 18398 17838 18450
rect 17838 18398 17890 18450
rect 17890 18398 17892 18450
rect 17836 18396 17892 18398
rect 18060 16882 18116 16884
rect 18060 16830 18062 16882
rect 18062 16830 18114 16882
rect 18114 16830 18116 16882
rect 18060 16828 18116 16830
rect 18396 16882 18452 16884
rect 18396 16830 18398 16882
rect 18398 16830 18450 16882
rect 18450 16830 18452 16882
rect 18396 16828 18452 16830
rect 18620 18172 18676 18228
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19964 18396 20020 18452
rect 19068 17666 19124 17668
rect 19068 17614 19070 17666
rect 19070 17614 19122 17666
rect 19122 17614 19124 17666
rect 19068 17612 19124 17614
rect 18284 16492 18340 16548
rect 19068 16658 19124 16660
rect 19068 16606 19070 16658
rect 19070 16606 19122 16658
rect 19122 16606 19124 16658
rect 19068 16604 19124 16606
rect 18060 16380 18116 16436
rect 18396 16156 18452 16212
rect 18172 16098 18228 16100
rect 18172 16046 18174 16098
rect 18174 16046 18226 16098
rect 18226 16046 18228 16098
rect 18172 16044 18228 16046
rect 19068 16098 19124 16100
rect 19068 16046 19070 16098
rect 19070 16046 19122 16098
rect 19122 16046 19124 16098
rect 19068 16044 19124 16046
rect 19964 17554 20020 17556
rect 19964 17502 19966 17554
rect 19966 17502 20018 17554
rect 20018 17502 20020 17554
rect 19964 17500 20020 17502
rect 21532 25676 21588 25732
rect 22764 35532 22820 35588
rect 22988 36988 23044 37044
rect 23212 36370 23268 36372
rect 23212 36318 23214 36370
rect 23214 36318 23266 36370
rect 23266 36318 23268 36370
rect 23212 36316 23268 36318
rect 23996 35922 24052 35924
rect 23996 35870 23998 35922
rect 23998 35870 24050 35922
rect 24050 35870 24052 35922
rect 23996 35868 24052 35870
rect 24556 36428 24612 36484
rect 26460 41580 26516 41636
rect 25452 40572 25508 40628
rect 25900 40684 25956 40740
rect 25564 40514 25620 40516
rect 25564 40462 25566 40514
rect 25566 40462 25618 40514
rect 25618 40462 25620 40514
rect 25564 40460 25620 40462
rect 25340 39004 25396 39060
rect 26124 40348 26180 40404
rect 25340 38722 25396 38724
rect 25340 38670 25342 38722
rect 25342 38670 25394 38722
rect 25394 38670 25396 38722
rect 25340 38668 25396 38670
rect 25676 38444 25732 38500
rect 25676 36594 25732 36596
rect 25676 36542 25678 36594
rect 25678 36542 25730 36594
rect 25730 36542 25732 36594
rect 25676 36540 25732 36542
rect 25564 36316 25620 36372
rect 23212 35698 23268 35700
rect 23212 35646 23214 35698
rect 23214 35646 23266 35698
rect 23266 35646 23268 35698
rect 23212 35644 23268 35646
rect 23772 35698 23828 35700
rect 23772 35646 23774 35698
rect 23774 35646 23826 35698
rect 23826 35646 23828 35698
rect 23772 35644 23828 35646
rect 23548 35196 23604 35252
rect 23772 35196 23828 35252
rect 23100 34300 23156 34356
rect 22540 33516 22596 33572
rect 22428 33458 22484 33460
rect 22428 33406 22430 33458
rect 22430 33406 22482 33458
rect 22482 33406 22484 33458
rect 22428 33404 22484 33406
rect 22316 33346 22372 33348
rect 22316 33294 22318 33346
rect 22318 33294 22370 33346
rect 22370 33294 22372 33346
rect 22316 33292 22372 33294
rect 22652 32620 22708 32676
rect 22092 31778 22148 31780
rect 22092 31726 22094 31778
rect 22094 31726 22146 31778
rect 22146 31726 22148 31778
rect 22092 31724 22148 31726
rect 22652 31276 22708 31332
rect 22540 31164 22596 31220
rect 22316 30716 22372 30772
rect 22428 29314 22484 29316
rect 22428 29262 22430 29314
rect 22430 29262 22482 29314
rect 22482 29262 22484 29314
rect 22428 29260 22484 29262
rect 23436 34636 23492 34692
rect 23772 34242 23828 34244
rect 23772 34190 23774 34242
rect 23774 34190 23826 34242
rect 23826 34190 23828 34242
rect 23772 34188 23828 34190
rect 23996 34354 24052 34356
rect 23996 34302 23998 34354
rect 23998 34302 24050 34354
rect 24050 34302 24052 34354
rect 23996 34300 24052 34302
rect 25340 35698 25396 35700
rect 25340 35646 25342 35698
rect 25342 35646 25394 35698
rect 25394 35646 25396 35698
rect 25340 35644 25396 35646
rect 25004 35138 25060 35140
rect 25004 35086 25006 35138
rect 25006 35086 25058 35138
rect 25058 35086 25060 35138
rect 25004 35084 25060 35086
rect 24668 34972 24724 35028
rect 25452 35196 25508 35252
rect 24220 34636 24276 34692
rect 23212 33740 23268 33796
rect 22876 33068 22932 33124
rect 23548 33122 23604 33124
rect 23548 33070 23550 33122
rect 23550 33070 23602 33122
rect 23602 33070 23604 33122
rect 23548 33068 23604 33070
rect 23548 32562 23604 32564
rect 23548 32510 23550 32562
rect 23550 32510 23602 32562
rect 23602 32510 23604 32562
rect 23548 32508 23604 32510
rect 22988 30940 23044 30996
rect 23100 31164 23156 31220
rect 23100 30604 23156 30660
rect 23660 31164 23716 31220
rect 23772 31612 23828 31668
rect 23772 30716 23828 30772
rect 23660 30044 23716 30100
rect 23996 31052 24052 31108
rect 24332 33852 24388 33908
rect 24892 33740 24948 33796
rect 23884 30492 23940 30548
rect 23996 30268 24052 30324
rect 24220 30268 24276 30324
rect 22764 28700 22820 28756
rect 22540 28642 22596 28644
rect 22540 28590 22542 28642
rect 22542 28590 22594 28642
rect 22594 28590 22596 28642
rect 22540 28588 22596 28590
rect 24556 33292 24612 33348
rect 25788 34802 25844 34804
rect 25788 34750 25790 34802
rect 25790 34750 25842 34802
rect 25842 34750 25844 34802
rect 25788 34748 25844 34750
rect 25004 33628 25060 33684
rect 24556 32844 24612 32900
rect 24668 32562 24724 32564
rect 24668 32510 24670 32562
rect 24670 32510 24722 32562
rect 24722 32510 24724 32562
rect 24668 32508 24724 32510
rect 24780 31052 24836 31108
rect 24668 30882 24724 30884
rect 24668 30830 24670 30882
rect 24670 30830 24722 30882
rect 24722 30830 24724 30882
rect 24668 30828 24724 30830
rect 24556 29986 24612 29988
rect 24556 29934 24558 29986
rect 24558 29934 24610 29986
rect 24610 29934 24612 29986
rect 24556 29932 24612 29934
rect 24444 29314 24500 29316
rect 24444 29262 24446 29314
rect 24446 29262 24498 29314
rect 24498 29262 24500 29314
rect 24444 29260 24500 29262
rect 23996 28754 24052 28756
rect 23996 28702 23998 28754
rect 23998 28702 24050 28754
rect 24050 28702 24052 28754
rect 23996 28700 24052 28702
rect 21868 26348 21924 26404
rect 22204 26290 22260 26292
rect 22204 26238 22206 26290
rect 22206 26238 22258 26290
rect 22258 26238 22260 26290
rect 22204 26236 22260 26238
rect 21980 25452 22036 25508
rect 21756 25228 21812 25284
rect 22204 24556 22260 24612
rect 21980 24444 22036 24500
rect 21756 23996 21812 24052
rect 20748 23324 20804 23380
rect 21308 23154 21364 23156
rect 21308 23102 21310 23154
rect 21310 23102 21362 23154
rect 21362 23102 21364 23154
rect 21308 23100 21364 23102
rect 20748 20748 20804 20804
rect 20636 20636 20692 20692
rect 20748 20300 20804 20356
rect 21420 20690 21476 20692
rect 21420 20638 21422 20690
rect 21422 20638 21474 20690
rect 21474 20638 21476 20690
rect 21420 20636 21476 20638
rect 21756 23714 21812 23716
rect 21756 23662 21758 23714
rect 21758 23662 21810 23714
rect 21810 23662 21812 23714
rect 21756 23660 21812 23662
rect 21644 23548 21700 23604
rect 21868 22876 21924 22932
rect 22204 23324 22260 23380
rect 21868 22146 21924 22148
rect 21868 22094 21870 22146
rect 21870 22094 21922 22146
rect 21922 22094 21924 22146
rect 21868 22092 21924 22094
rect 21980 21868 22036 21924
rect 20860 18284 20916 18340
rect 20860 17836 20916 17892
rect 20524 17612 20580 17668
rect 20300 17500 20356 17556
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19292 16044 19348 16100
rect 17724 15820 17780 15876
rect 17948 15484 18004 15540
rect 18284 15372 18340 15428
rect 18396 15820 18452 15876
rect 18844 15538 18900 15540
rect 18844 15486 18846 15538
rect 18846 15486 18898 15538
rect 18898 15486 18900 15538
rect 18844 15484 18900 15486
rect 16604 14252 16660 14308
rect 18396 14364 18452 14420
rect 16716 13020 16772 13076
rect 17724 12962 17780 12964
rect 17724 12910 17726 12962
rect 17726 12910 17778 12962
rect 17778 12910 17780 12962
rect 17724 12908 17780 12910
rect 17948 13692 18004 13748
rect 17948 13522 18004 13524
rect 17948 13470 17950 13522
rect 17950 13470 18002 13522
rect 18002 13470 18004 13522
rect 17948 13468 18004 13470
rect 18508 13132 18564 13188
rect 19404 15484 19460 15540
rect 19516 16492 19572 16548
rect 19740 16658 19796 16660
rect 19740 16606 19742 16658
rect 19742 16606 19794 16658
rect 19794 16606 19796 16658
rect 19740 16604 19796 16606
rect 19628 16210 19684 16212
rect 19628 16158 19630 16210
rect 19630 16158 19682 16210
rect 19682 16158 19684 16210
rect 19628 16156 19684 16158
rect 21868 18674 21924 18676
rect 21868 18622 21870 18674
rect 21870 18622 21922 18674
rect 21922 18622 21924 18674
rect 21868 18620 21924 18622
rect 22204 18508 22260 18564
rect 22652 25676 22708 25732
rect 22876 24610 22932 24612
rect 22876 24558 22878 24610
rect 22878 24558 22930 24610
rect 22930 24558 22932 24610
rect 22876 24556 22932 24558
rect 22988 24444 23044 24500
rect 22428 21980 22484 22036
rect 22540 20300 22596 20356
rect 22764 23548 22820 23604
rect 22988 23938 23044 23940
rect 22988 23886 22990 23938
rect 22990 23886 23042 23938
rect 23042 23886 23044 23938
rect 22988 23884 23044 23886
rect 23100 23826 23156 23828
rect 23100 23774 23102 23826
rect 23102 23774 23154 23826
rect 23154 23774 23156 23826
rect 23100 23772 23156 23774
rect 22988 23660 23044 23716
rect 22764 23154 22820 23156
rect 22764 23102 22766 23154
rect 22766 23102 22818 23154
rect 22818 23102 22820 23154
rect 22764 23100 22820 23102
rect 23548 27020 23604 27076
rect 23436 26460 23492 26516
rect 23996 26796 24052 26852
rect 23548 25452 23604 25508
rect 24556 28028 24612 28084
rect 24220 27074 24276 27076
rect 24220 27022 24222 27074
rect 24222 27022 24274 27074
rect 24274 27022 24276 27074
rect 24220 27020 24276 27022
rect 24332 26796 24388 26852
rect 24668 26684 24724 26740
rect 24556 26236 24612 26292
rect 24556 25788 24612 25844
rect 24332 25004 24388 25060
rect 24444 24946 24500 24948
rect 24444 24894 24446 24946
rect 24446 24894 24498 24946
rect 24498 24894 24500 24946
rect 24444 24892 24500 24894
rect 24444 24498 24500 24500
rect 24444 24446 24446 24498
rect 24446 24446 24498 24498
rect 24498 24446 24500 24498
rect 24444 24444 24500 24446
rect 23436 23436 23492 23492
rect 23212 23324 23268 23380
rect 23100 23266 23156 23268
rect 23100 23214 23102 23266
rect 23102 23214 23154 23266
rect 23154 23214 23156 23266
rect 23100 23212 23156 23214
rect 22876 22258 22932 22260
rect 22876 22206 22878 22258
rect 22878 22206 22930 22258
rect 22930 22206 22932 22258
rect 22876 22204 22932 22206
rect 22652 21868 22708 21924
rect 22428 19906 22484 19908
rect 22428 19854 22430 19906
rect 22430 19854 22482 19906
rect 22482 19854 22484 19906
rect 22428 19852 22484 19854
rect 22764 21644 22820 21700
rect 22876 21980 22932 22036
rect 22876 20578 22932 20580
rect 22876 20526 22878 20578
rect 22878 20526 22930 20578
rect 22930 20526 22932 20578
rect 22876 20524 22932 20526
rect 23100 21810 23156 21812
rect 23100 21758 23102 21810
rect 23102 21758 23154 21810
rect 23154 21758 23156 21810
rect 23100 21756 23156 21758
rect 23884 23324 23940 23380
rect 23996 23266 24052 23268
rect 23996 23214 23998 23266
rect 23998 23214 24050 23266
rect 24050 23214 24052 23266
rect 23996 23212 24052 23214
rect 24556 23378 24612 23380
rect 24556 23326 24558 23378
rect 24558 23326 24610 23378
rect 24610 23326 24612 23378
rect 24556 23324 24612 23326
rect 23324 21868 23380 21924
rect 23436 21698 23492 21700
rect 23436 21646 23438 21698
rect 23438 21646 23490 21698
rect 23490 21646 23492 21698
rect 23436 21644 23492 21646
rect 23548 20690 23604 20692
rect 23548 20638 23550 20690
rect 23550 20638 23602 20690
rect 23602 20638 23604 20690
rect 23548 20636 23604 20638
rect 23772 20636 23828 20692
rect 23996 21756 24052 21812
rect 23100 19740 23156 19796
rect 22316 18396 22372 18452
rect 22652 18450 22708 18452
rect 22652 18398 22654 18450
rect 22654 18398 22706 18450
rect 22706 18398 22708 18450
rect 22652 18396 22708 18398
rect 21420 17500 21476 17556
rect 20188 16268 20244 16324
rect 20300 16604 20356 16660
rect 20412 15874 20468 15876
rect 20412 15822 20414 15874
rect 20414 15822 20466 15874
rect 20466 15822 20468 15874
rect 20412 15820 20468 15822
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19628 15484 19684 15540
rect 19964 15484 20020 15540
rect 19740 15426 19796 15428
rect 19740 15374 19742 15426
rect 19742 15374 19794 15426
rect 19794 15374 19796 15426
rect 19740 15372 19796 15374
rect 20188 15484 20244 15540
rect 19516 15314 19572 15316
rect 19516 15262 19518 15314
rect 19518 15262 19570 15314
rect 19570 15262 19572 15314
rect 19516 15260 19572 15262
rect 21084 16828 21140 16884
rect 20860 16156 20916 16212
rect 20972 16716 21028 16772
rect 21308 16492 21364 16548
rect 21196 16268 21252 16324
rect 20972 15538 21028 15540
rect 20972 15486 20974 15538
rect 20974 15486 21026 15538
rect 21026 15486 21028 15538
rect 20972 15484 21028 15486
rect 20748 15426 20804 15428
rect 20748 15374 20750 15426
rect 20750 15374 20802 15426
rect 20802 15374 20804 15426
rect 20748 15372 20804 15374
rect 20636 15314 20692 15316
rect 20636 15262 20638 15314
rect 20638 15262 20690 15314
rect 20690 15262 20692 15314
rect 20636 15260 20692 15262
rect 21868 17052 21924 17108
rect 21532 16770 21588 16772
rect 21532 16718 21534 16770
rect 21534 16718 21586 16770
rect 21586 16718 21588 16770
rect 21532 16716 21588 16718
rect 21868 16156 21924 16212
rect 21532 16098 21588 16100
rect 21532 16046 21534 16098
rect 21534 16046 21586 16098
rect 21586 16046 21588 16098
rect 21532 16044 21588 16046
rect 19628 15148 19684 15204
rect 20860 15202 20916 15204
rect 20860 15150 20862 15202
rect 20862 15150 20914 15202
rect 20914 15150 20916 15202
rect 20860 15148 20916 15150
rect 22876 18396 22932 18452
rect 23884 20130 23940 20132
rect 23884 20078 23886 20130
rect 23886 20078 23938 20130
rect 23938 20078 23940 20130
rect 23884 20076 23940 20078
rect 24556 22482 24612 22484
rect 24556 22430 24558 22482
rect 24558 22430 24610 22482
rect 24610 22430 24612 22482
rect 24556 22428 24612 22430
rect 24444 21644 24500 21700
rect 24220 20972 24276 21028
rect 24332 19740 24388 19796
rect 25228 32562 25284 32564
rect 25228 32510 25230 32562
rect 25230 32510 25282 32562
rect 25282 32510 25284 32562
rect 25228 32508 25284 32510
rect 25004 31890 25060 31892
rect 25004 31838 25006 31890
rect 25006 31838 25058 31890
rect 25058 31838 25060 31890
rect 25004 31836 25060 31838
rect 25676 34690 25732 34692
rect 25676 34638 25678 34690
rect 25678 34638 25730 34690
rect 25730 34638 25732 34690
rect 25676 34636 25732 34638
rect 26236 39340 26292 39396
rect 26236 38834 26292 38836
rect 26236 38782 26238 38834
rect 26238 38782 26290 38834
rect 26290 38782 26292 38834
rect 26236 38780 26292 38782
rect 26124 38668 26180 38724
rect 26684 42140 26740 42196
rect 27020 45052 27076 45108
rect 29148 45778 29204 45780
rect 29148 45726 29150 45778
rect 29150 45726 29202 45778
rect 29202 45726 29204 45778
rect 29148 45724 29204 45726
rect 30604 45724 30660 45780
rect 26684 41746 26740 41748
rect 26684 41694 26686 41746
rect 26686 41694 26738 41746
rect 26738 41694 26740 41746
rect 26684 41692 26740 41694
rect 26796 41020 26852 41076
rect 26684 40402 26740 40404
rect 26684 40350 26686 40402
rect 26686 40350 26738 40402
rect 26738 40350 26740 40402
rect 26684 40348 26740 40350
rect 26908 39788 26964 39844
rect 26684 39394 26740 39396
rect 26684 39342 26686 39394
rect 26686 39342 26738 39394
rect 26738 39342 26740 39394
rect 26684 39340 26740 39342
rect 26572 38050 26628 38052
rect 26572 37998 26574 38050
rect 26574 37998 26626 38050
rect 26626 37998 26628 38050
rect 26572 37996 26628 37998
rect 27132 43596 27188 43652
rect 28476 44994 28532 44996
rect 28476 44942 28478 44994
rect 28478 44942 28530 44994
rect 28530 44942 28532 44994
rect 28476 44940 28532 44942
rect 31388 45276 31444 45332
rect 31612 45612 31668 45668
rect 31948 45330 32004 45332
rect 31948 45278 31950 45330
rect 31950 45278 32002 45330
rect 32002 45278 32004 45330
rect 31948 45276 32004 45278
rect 31724 45052 31780 45108
rect 31052 44994 31108 44996
rect 31052 44942 31054 44994
rect 31054 44942 31106 44994
rect 31106 44942 31108 44994
rect 31052 44940 31108 44942
rect 30940 44434 30996 44436
rect 30940 44382 30942 44434
rect 30942 44382 30994 44434
rect 30994 44382 30996 44434
rect 30940 44380 30996 44382
rect 28476 43596 28532 43652
rect 31164 44492 31220 44548
rect 30268 43596 30324 43652
rect 29596 43372 29652 43428
rect 28476 42812 28532 42868
rect 27244 41970 27300 41972
rect 27244 41918 27246 41970
rect 27246 41918 27298 41970
rect 27298 41918 27300 41970
rect 27244 41916 27300 41918
rect 29148 41916 29204 41972
rect 28028 41858 28084 41860
rect 28028 41806 28030 41858
rect 28030 41806 28082 41858
rect 28082 41806 28084 41858
rect 28028 41804 28084 41806
rect 27692 41692 27748 41748
rect 28028 40460 28084 40516
rect 27020 37548 27076 37604
rect 27804 40402 27860 40404
rect 27804 40350 27806 40402
rect 27806 40350 27858 40402
rect 27858 40350 27860 40402
rect 27804 40348 27860 40350
rect 28364 40460 28420 40516
rect 28252 39788 28308 39844
rect 27356 39452 27412 39508
rect 26572 36988 26628 37044
rect 26348 35868 26404 35924
rect 26012 35586 26068 35588
rect 26012 35534 26014 35586
rect 26014 35534 26066 35586
rect 26066 35534 26068 35586
rect 26012 35532 26068 35534
rect 27244 37660 27300 37716
rect 28924 40460 28980 40516
rect 29484 42700 29540 42756
rect 29372 41074 29428 41076
rect 29372 41022 29374 41074
rect 29374 41022 29426 41074
rect 29426 41022 29428 41074
rect 29372 41020 29428 41022
rect 28476 40402 28532 40404
rect 28476 40350 28478 40402
rect 28478 40350 28530 40402
rect 28530 40350 28532 40402
rect 28476 40348 28532 40350
rect 28924 40290 28980 40292
rect 28924 40238 28926 40290
rect 28926 40238 28978 40290
rect 28978 40238 28980 40290
rect 28924 40236 28980 40238
rect 29148 40124 29204 40180
rect 29260 39618 29316 39620
rect 29260 39566 29262 39618
rect 29262 39566 29314 39618
rect 29314 39566 29316 39618
rect 29260 39564 29316 39566
rect 29148 39452 29204 39508
rect 27804 37660 27860 37716
rect 26348 35420 26404 35476
rect 27692 35698 27748 35700
rect 27692 35646 27694 35698
rect 27694 35646 27746 35698
rect 27746 35646 27748 35698
rect 27692 35644 27748 35646
rect 26684 35308 26740 35364
rect 25900 34188 25956 34244
rect 25788 32956 25844 33012
rect 25676 31836 25732 31892
rect 25676 31554 25732 31556
rect 25676 31502 25678 31554
rect 25678 31502 25730 31554
rect 25730 31502 25732 31554
rect 25676 31500 25732 31502
rect 25564 31218 25620 31220
rect 25564 31166 25566 31218
rect 25566 31166 25618 31218
rect 25618 31166 25620 31218
rect 25564 31164 25620 31166
rect 25676 30940 25732 30996
rect 25340 30492 25396 30548
rect 25004 30044 25060 30100
rect 26796 33628 26852 33684
rect 26012 33346 26068 33348
rect 26012 33294 26014 33346
rect 26014 33294 26066 33346
rect 26066 33294 26068 33346
rect 26012 33292 26068 33294
rect 26012 32508 26068 32564
rect 26236 32396 26292 32452
rect 26684 31836 26740 31892
rect 27020 33404 27076 33460
rect 27468 34690 27524 34692
rect 27468 34638 27470 34690
rect 27470 34638 27522 34690
rect 27522 34638 27524 34690
rect 27468 34636 27524 34638
rect 26908 31948 26964 32004
rect 27356 32844 27412 32900
rect 26572 31554 26628 31556
rect 26572 31502 26574 31554
rect 26574 31502 26626 31554
rect 26626 31502 26628 31554
rect 26572 31500 26628 31502
rect 27132 31724 27188 31780
rect 26796 31388 26852 31444
rect 26572 31276 26628 31332
rect 26796 31218 26852 31220
rect 26796 31166 26798 31218
rect 26798 31166 26850 31218
rect 26850 31166 26852 31218
rect 26796 31164 26852 31166
rect 27020 31164 27076 31220
rect 27580 33346 27636 33348
rect 27580 33294 27582 33346
rect 27582 33294 27634 33346
rect 27634 33294 27636 33346
rect 27580 33292 27636 33294
rect 27692 33122 27748 33124
rect 27692 33070 27694 33122
rect 27694 33070 27746 33122
rect 27746 33070 27748 33122
rect 27692 33068 27748 33070
rect 27468 32732 27524 32788
rect 27468 32172 27524 32228
rect 27356 31778 27412 31780
rect 27356 31726 27358 31778
rect 27358 31726 27410 31778
rect 27410 31726 27412 31778
rect 27356 31724 27412 31726
rect 26124 30828 26180 30884
rect 26460 30210 26516 30212
rect 26460 30158 26462 30210
rect 26462 30158 26514 30210
rect 26514 30158 26516 30210
rect 26460 30156 26516 30158
rect 25900 30098 25956 30100
rect 25900 30046 25902 30098
rect 25902 30046 25954 30098
rect 25954 30046 25956 30098
rect 25900 30044 25956 30046
rect 26236 30098 26292 30100
rect 26236 30046 26238 30098
rect 26238 30046 26290 30098
rect 26290 30046 26292 30098
rect 26236 30044 26292 30046
rect 24892 28028 24948 28084
rect 24892 26796 24948 26852
rect 24892 25564 24948 25620
rect 26012 28700 26068 28756
rect 26124 28588 26180 28644
rect 26236 28082 26292 28084
rect 26236 28030 26238 28082
rect 26238 28030 26290 28082
rect 26290 28030 26292 28082
rect 26236 28028 26292 28030
rect 26124 27804 26180 27860
rect 25228 26684 25284 26740
rect 25452 27468 25508 27524
rect 25228 26348 25284 26404
rect 25788 27244 25844 27300
rect 25676 26962 25732 26964
rect 25676 26910 25678 26962
rect 25678 26910 25730 26962
rect 25730 26910 25732 26962
rect 25676 26908 25732 26910
rect 26012 27132 26068 27188
rect 25788 26514 25844 26516
rect 25788 26462 25790 26514
rect 25790 26462 25842 26514
rect 25842 26462 25844 26514
rect 25788 26460 25844 26462
rect 25452 25676 25508 25732
rect 25116 25228 25172 25284
rect 24892 20748 24948 20804
rect 23212 18508 23268 18564
rect 23436 17836 23492 17892
rect 22764 17724 22820 17780
rect 22428 17052 22484 17108
rect 22316 16098 22372 16100
rect 22316 16046 22318 16098
rect 22318 16046 22370 16098
rect 22370 16046 22372 16098
rect 22316 16044 22372 16046
rect 22652 17442 22708 17444
rect 22652 17390 22654 17442
rect 22654 17390 22706 17442
rect 22706 17390 22708 17442
rect 22652 17388 22708 17390
rect 22764 16716 22820 16772
rect 23100 17052 23156 17108
rect 23660 17388 23716 17444
rect 23324 16716 23380 16772
rect 25452 25228 25508 25284
rect 25452 24780 25508 24836
rect 25340 24722 25396 24724
rect 25340 24670 25342 24722
rect 25342 24670 25394 24722
rect 25394 24670 25396 24722
rect 25340 24668 25396 24670
rect 25228 23772 25284 23828
rect 25116 22988 25172 23044
rect 25228 21474 25284 21476
rect 25228 21422 25230 21474
rect 25230 21422 25282 21474
rect 25282 21422 25284 21474
rect 25228 21420 25284 21422
rect 25788 24722 25844 24724
rect 25788 24670 25790 24722
rect 25790 24670 25842 24722
rect 25842 24670 25844 24722
rect 25788 24668 25844 24670
rect 25900 24444 25956 24500
rect 26012 26236 26068 26292
rect 25788 23660 25844 23716
rect 25564 22876 25620 22932
rect 25676 22428 25732 22484
rect 26796 29484 26852 29540
rect 26684 28588 26740 28644
rect 26236 27468 26292 27524
rect 27244 30156 27300 30212
rect 28252 36204 28308 36260
rect 27916 35644 27972 35700
rect 27916 34690 27972 34692
rect 27916 34638 27918 34690
rect 27918 34638 27970 34690
rect 27970 34638 27972 34690
rect 27916 34636 27972 34638
rect 28588 38556 28644 38612
rect 29148 38834 29204 38836
rect 29148 38782 29150 38834
rect 29150 38782 29202 38834
rect 29202 38782 29204 38834
rect 29148 38780 29204 38782
rect 29708 43260 29764 43316
rect 30044 42642 30100 42644
rect 30044 42590 30046 42642
rect 30046 42590 30098 42642
rect 30098 42590 30100 42642
rect 30044 42588 30100 42590
rect 31276 43596 31332 43652
rect 30604 43484 30660 43540
rect 31164 43484 31220 43540
rect 30604 43260 30660 43316
rect 30380 42754 30436 42756
rect 30380 42702 30382 42754
rect 30382 42702 30434 42754
rect 30434 42702 30436 42754
rect 30380 42700 30436 42702
rect 31388 43260 31444 43316
rect 31948 44322 32004 44324
rect 31948 44270 31950 44322
rect 31950 44270 32002 44322
rect 32002 44270 32004 44322
rect 31948 44268 32004 44270
rect 33068 45778 33124 45780
rect 33068 45726 33070 45778
rect 33070 45726 33122 45778
rect 33122 45726 33124 45778
rect 33068 45724 33124 45726
rect 32508 45388 32564 45444
rect 32284 45106 32340 45108
rect 32284 45054 32286 45106
rect 32286 45054 32338 45106
rect 32338 45054 32340 45106
rect 32284 45052 32340 45054
rect 32284 44546 32340 44548
rect 32284 44494 32286 44546
rect 32286 44494 32338 44546
rect 32338 44494 32340 44546
rect 32284 44492 32340 44494
rect 30492 41970 30548 41972
rect 30492 41918 30494 41970
rect 30494 41918 30546 41970
rect 30546 41918 30548 41970
rect 30492 41916 30548 41918
rect 29932 41580 29988 41636
rect 32620 45052 32676 45108
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 33404 45388 33460 45444
rect 33852 45666 33908 45668
rect 33852 45614 33854 45666
rect 33854 45614 33906 45666
rect 33906 45614 33908 45666
rect 33852 45612 33908 45614
rect 33964 45388 34020 45444
rect 34412 45276 34468 45332
rect 33740 45052 33796 45108
rect 33404 44994 33460 44996
rect 33404 44942 33406 44994
rect 33406 44942 33458 44994
rect 33458 44942 33460 44994
rect 33404 44940 33460 44942
rect 34636 44940 34692 44996
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 33964 44492 34020 44548
rect 33292 44380 33348 44436
rect 31948 42028 32004 42084
rect 31276 41580 31332 41636
rect 29708 40908 29764 40964
rect 30604 40908 30660 40964
rect 30492 40684 30548 40740
rect 30044 39618 30100 39620
rect 30044 39566 30046 39618
rect 30046 39566 30098 39618
rect 30098 39566 30100 39618
rect 30044 39564 30100 39566
rect 29708 39452 29764 39508
rect 28588 37660 28644 37716
rect 29260 36540 29316 36596
rect 30268 39842 30324 39844
rect 30268 39790 30270 39842
rect 30270 39790 30322 39842
rect 30322 39790 30324 39842
rect 30268 39788 30324 39790
rect 29596 38556 29652 38612
rect 30716 40402 30772 40404
rect 30716 40350 30718 40402
rect 30718 40350 30770 40402
rect 30770 40350 30772 40402
rect 30716 40348 30772 40350
rect 32396 42028 32452 42084
rect 33068 43314 33124 43316
rect 33068 43262 33070 43314
rect 33070 43262 33122 43314
rect 33122 43262 33124 43314
rect 33068 43260 33124 43262
rect 34188 44546 34244 44548
rect 34188 44494 34190 44546
rect 34190 44494 34242 44546
rect 34242 44494 34244 44546
rect 34188 44492 34244 44494
rect 35532 44492 35588 44548
rect 33628 44322 33684 44324
rect 33628 44270 33630 44322
rect 33630 44270 33682 44322
rect 33682 44270 33684 44322
rect 33628 44268 33684 44270
rect 33628 43708 33684 43764
rect 33404 43538 33460 43540
rect 33404 43486 33406 43538
rect 33406 43486 33458 43538
rect 33458 43486 33460 43538
rect 33404 43484 33460 43486
rect 33628 42754 33684 42756
rect 33628 42702 33630 42754
rect 33630 42702 33682 42754
rect 33682 42702 33684 42754
rect 33628 42700 33684 42702
rect 33404 42252 33460 42308
rect 32732 41804 32788 41860
rect 31388 40962 31444 40964
rect 31388 40910 31390 40962
rect 31390 40910 31442 40962
rect 31442 40910 31444 40962
rect 31388 40908 31444 40910
rect 31388 40514 31444 40516
rect 31388 40462 31390 40514
rect 31390 40462 31442 40514
rect 31442 40462 31444 40514
rect 31388 40460 31444 40462
rect 31164 40348 31220 40404
rect 30380 38780 30436 38836
rect 30492 39618 30548 39620
rect 30492 39566 30494 39618
rect 30494 39566 30546 39618
rect 30546 39566 30548 39618
rect 30492 39564 30548 39566
rect 31052 39564 31108 39620
rect 31500 40402 31556 40404
rect 31500 40350 31502 40402
rect 31502 40350 31554 40402
rect 31554 40350 31556 40402
rect 31500 40348 31556 40350
rect 31276 40124 31332 40180
rect 31500 40124 31556 40180
rect 29596 38050 29652 38052
rect 29596 37998 29598 38050
rect 29598 37998 29650 38050
rect 29650 37998 29652 38050
rect 29596 37996 29652 37998
rect 30380 37996 30436 38052
rect 30268 37938 30324 37940
rect 30268 37886 30270 37938
rect 30270 37886 30322 37938
rect 30322 37886 30324 37938
rect 30268 37884 30324 37886
rect 29484 37436 29540 37492
rect 29820 36540 29876 36596
rect 29708 36370 29764 36372
rect 29708 36318 29710 36370
rect 29710 36318 29762 36370
rect 29762 36318 29764 36370
rect 29708 36316 29764 36318
rect 28588 34748 28644 34804
rect 29148 35980 29204 36036
rect 29596 36258 29652 36260
rect 29596 36206 29598 36258
rect 29598 36206 29650 36258
rect 29650 36206 29652 36258
rect 29596 36204 29652 36206
rect 29596 35980 29652 36036
rect 29484 35756 29540 35812
rect 29148 35644 29204 35700
rect 29372 35644 29428 35700
rect 29484 34860 29540 34916
rect 30940 37100 30996 37156
rect 31164 37212 31220 37268
rect 30716 36092 30772 36148
rect 30940 35756 30996 35812
rect 29372 34690 29428 34692
rect 29372 34638 29374 34690
rect 29374 34638 29426 34690
rect 29426 34638 29428 34690
rect 29372 34636 29428 34638
rect 29708 34636 29764 34692
rect 29036 34130 29092 34132
rect 29036 34078 29038 34130
rect 29038 34078 29090 34130
rect 29090 34078 29092 34130
rect 29036 34076 29092 34078
rect 28252 33180 28308 33236
rect 28588 33122 28644 33124
rect 28588 33070 28590 33122
rect 28590 33070 28642 33122
rect 28642 33070 28644 33122
rect 28588 33068 28644 33070
rect 28028 32732 28084 32788
rect 28140 32956 28196 33012
rect 27916 32674 27972 32676
rect 27916 32622 27918 32674
rect 27918 32622 27970 32674
rect 27970 32622 27972 32674
rect 27916 32620 27972 32622
rect 27804 31724 27860 31780
rect 27916 32172 27972 32228
rect 27692 31612 27748 31668
rect 27804 31554 27860 31556
rect 27804 31502 27806 31554
rect 27806 31502 27858 31554
rect 27858 31502 27860 31554
rect 27804 31500 27860 31502
rect 27916 31276 27972 31332
rect 27580 31106 27636 31108
rect 27580 31054 27582 31106
rect 27582 31054 27634 31106
rect 27634 31054 27636 31106
rect 27580 31052 27636 31054
rect 27916 31052 27972 31108
rect 28476 32956 28532 33012
rect 28476 32732 28532 32788
rect 28588 31724 28644 31780
rect 28476 31276 28532 31332
rect 27468 29932 27524 29988
rect 27692 30098 27748 30100
rect 27692 30046 27694 30098
rect 27694 30046 27746 30098
rect 27746 30046 27748 30098
rect 27692 30044 27748 30046
rect 28028 29708 28084 29764
rect 27356 29538 27412 29540
rect 27356 29486 27358 29538
rect 27358 29486 27410 29538
rect 27410 29486 27412 29538
rect 27356 29484 27412 29486
rect 27580 28642 27636 28644
rect 27580 28590 27582 28642
rect 27582 28590 27634 28642
rect 27634 28590 27636 28642
rect 27580 28588 27636 28590
rect 27132 28028 27188 28084
rect 27356 28140 27412 28196
rect 26796 27020 26852 27076
rect 26572 26962 26628 26964
rect 26572 26910 26574 26962
rect 26574 26910 26626 26962
rect 26626 26910 26628 26962
rect 26572 26908 26628 26910
rect 27020 27132 27076 27188
rect 26908 26850 26964 26852
rect 26908 26798 26910 26850
rect 26910 26798 26962 26850
rect 26962 26798 26964 26850
rect 26908 26796 26964 26798
rect 27356 27244 27412 27300
rect 26796 25116 26852 25172
rect 26124 23884 26180 23940
rect 26684 23772 26740 23828
rect 26348 23042 26404 23044
rect 26348 22990 26350 23042
rect 26350 22990 26402 23042
rect 26402 22990 26404 23042
rect 26348 22988 26404 22990
rect 26460 21420 26516 21476
rect 25004 20076 25060 20132
rect 24108 18338 24164 18340
rect 24108 18286 24110 18338
rect 24110 18286 24162 18338
rect 24162 18286 24164 18338
rect 24108 18284 24164 18286
rect 23884 17778 23940 17780
rect 23884 17726 23886 17778
rect 23886 17726 23938 17778
rect 23938 17726 23940 17778
rect 23884 17724 23940 17726
rect 23996 15874 24052 15876
rect 23996 15822 23998 15874
rect 23998 15822 24050 15874
rect 24050 15822 24052 15874
rect 23996 15820 24052 15822
rect 23436 15538 23492 15540
rect 23436 15486 23438 15538
rect 23438 15486 23490 15538
rect 23490 15486 23492 15538
rect 23436 15484 23492 15486
rect 22540 15260 22596 15316
rect 20300 14418 20356 14420
rect 20300 14366 20302 14418
rect 20302 14366 20354 14418
rect 20354 14366 20356 14418
rect 20300 14364 20356 14366
rect 19516 14306 19572 14308
rect 19516 14254 19518 14306
rect 19518 14254 19570 14306
rect 19570 14254 19572 14306
rect 19516 14252 19572 14254
rect 18844 12908 18900 12964
rect 18172 12850 18228 12852
rect 18172 12798 18174 12850
rect 18174 12798 18226 12850
rect 18226 12798 18228 12850
rect 18172 12796 18228 12798
rect 18508 12796 18564 12852
rect 16716 12012 16772 12068
rect 17836 12066 17892 12068
rect 17836 12014 17838 12066
rect 17838 12014 17890 12066
rect 17890 12014 17892 12066
rect 17836 12012 17892 12014
rect 18172 11676 18228 11732
rect 16604 11228 16660 11284
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19516 13132 19572 13188
rect 19852 12962 19908 12964
rect 19852 12910 19854 12962
rect 19854 12910 19906 12962
rect 19906 12910 19908 12962
rect 19852 12908 19908 12910
rect 20300 12962 20356 12964
rect 20300 12910 20302 12962
rect 20302 12910 20354 12962
rect 20354 12910 20356 12962
rect 20300 12908 20356 12910
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19068 11340 19124 11396
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 21308 13804 21364 13860
rect 21756 14476 21812 14532
rect 21084 13468 21140 13524
rect 20524 12908 20580 12964
rect 20860 12738 20916 12740
rect 20860 12686 20862 12738
rect 20862 12686 20914 12738
rect 20914 12686 20916 12738
rect 20860 12684 20916 12686
rect 20412 10780 20468 10836
rect 16828 9266 16884 9268
rect 16828 9214 16830 9266
rect 16830 9214 16882 9266
rect 16882 9214 16884 9266
rect 16828 9212 16884 9214
rect 16044 9100 16100 9156
rect 16044 8428 16100 8484
rect 16604 8428 16660 8484
rect 16268 8258 16324 8260
rect 16268 8206 16270 8258
rect 16270 8206 16322 8258
rect 16322 8206 16324 8258
rect 16268 8204 16324 8206
rect 16156 8034 16212 8036
rect 16156 7982 16158 8034
rect 16158 7982 16210 8034
rect 16210 7982 16212 8034
rect 16156 7980 16212 7982
rect 16044 7868 16100 7924
rect 15932 5964 15988 6020
rect 16492 6748 16548 6804
rect 16044 6412 16100 6468
rect 15148 5516 15204 5572
rect 7532 4172 7588 4228
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 13132 3500 13188 3556
rect 7756 3388 7812 3444
rect 8204 3442 8260 3444
rect 8204 3390 8206 3442
rect 8206 3390 8258 3442
rect 8258 3390 8260 3442
rect 8204 3388 8260 3390
rect 16268 6524 16324 6580
rect 16156 6018 16212 6020
rect 16156 5966 16158 6018
rect 16158 5966 16210 6018
rect 16210 5966 16212 6018
rect 16156 5964 16212 5966
rect 16716 8204 16772 8260
rect 16716 8034 16772 8036
rect 16716 7982 16718 8034
rect 16718 7982 16770 8034
rect 16770 7982 16772 8034
rect 16716 7980 16772 7982
rect 17276 9660 17332 9716
rect 21308 13132 21364 13188
rect 22428 13804 22484 13860
rect 23212 13692 23268 13748
rect 21868 12738 21924 12740
rect 21868 12686 21870 12738
rect 21870 12686 21922 12738
rect 21922 12686 21924 12738
rect 21868 12684 21924 12686
rect 21420 11788 21476 11844
rect 22540 12684 22596 12740
rect 21868 11004 21924 11060
rect 22204 11900 22260 11956
rect 21532 10834 21588 10836
rect 21532 10782 21534 10834
rect 21534 10782 21586 10834
rect 21586 10782 21588 10834
rect 21532 10780 21588 10782
rect 20972 9772 21028 9828
rect 18844 9660 18900 9716
rect 17500 9212 17556 9268
rect 18732 9548 18788 9604
rect 17388 9100 17444 9156
rect 17276 8146 17332 8148
rect 17276 8094 17278 8146
rect 17278 8094 17330 8146
rect 17330 8094 17332 8146
rect 17276 8092 17332 8094
rect 17388 7980 17444 8036
rect 17276 7868 17332 7924
rect 17052 6802 17108 6804
rect 17052 6750 17054 6802
rect 17054 6750 17106 6802
rect 17106 6750 17108 6802
rect 17052 6748 17108 6750
rect 16604 5122 16660 5124
rect 16604 5070 16606 5122
rect 16606 5070 16658 5122
rect 16658 5070 16660 5122
rect 16604 5068 16660 5070
rect 15708 5010 15764 5012
rect 15708 4958 15710 5010
rect 15710 4958 15762 5010
rect 15762 4958 15764 5010
rect 15708 4956 15764 4958
rect 16044 4898 16100 4900
rect 16044 4846 16046 4898
rect 16046 4846 16098 4898
rect 16098 4846 16100 4898
rect 16044 4844 16100 4846
rect 16380 4396 16436 4452
rect 17164 6466 17220 6468
rect 17164 6414 17166 6466
rect 17166 6414 17218 6466
rect 17218 6414 17220 6466
rect 17164 6412 17220 6414
rect 16940 6076 16996 6132
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 20524 9436 20580 9492
rect 19180 8316 19236 8372
rect 18060 8258 18116 8260
rect 18060 8206 18062 8258
rect 18062 8206 18114 8258
rect 18114 8206 18116 8258
rect 18060 8204 18116 8206
rect 17724 8092 17780 8148
rect 17836 7868 17892 7924
rect 17612 6076 17668 6132
rect 17052 5964 17108 6020
rect 15148 3388 15204 3444
rect 17612 5794 17668 5796
rect 17612 5742 17614 5794
rect 17614 5742 17666 5794
rect 17666 5742 17668 5794
rect 17612 5740 17668 5742
rect 19404 8034 19460 8036
rect 19404 7982 19406 8034
rect 19406 7982 19458 8034
rect 19458 7982 19460 8034
rect 19404 7980 19460 7982
rect 18396 7868 18452 7924
rect 20188 8204 20244 8260
rect 21196 8930 21252 8932
rect 21196 8878 21198 8930
rect 21198 8878 21250 8930
rect 21250 8878 21252 8930
rect 21196 8876 21252 8878
rect 20860 8428 20916 8484
rect 20300 8146 20356 8148
rect 20300 8094 20302 8146
rect 20302 8094 20354 8146
rect 20354 8094 20356 8146
rect 20300 8092 20356 8094
rect 21532 9772 21588 9828
rect 21868 9826 21924 9828
rect 21868 9774 21870 9826
rect 21870 9774 21922 9826
rect 21922 9774 21924 9826
rect 21868 9772 21924 9774
rect 21644 9602 21700 9604
rect 21644 9550 21646 9602
rect 21646 9550 21698 9602
rect 21698 9550 21700 9602
rect 21644 9548 21700 9550
rect 21532 9436 21588 9492
rect 21420 8370 21476 8372
rect 21420 8318 21422 8370
rect 21422 8318 21474 8370
rect 21474 8318 21476 8370
rect 21420 8316 21476 8318
rect 21420 8146 21476 8148
rect 21420 8094 21422 8146
rect 21422 8094 21474 8146
rect 21474 8094 21476 8146
rect 21420 8092 21476 8094
rect 20188 8034 20244 8036
rect 20188 7982 20190 8034
rect 20190 7982 20242 8034
rect 20242 7982 20244 8034
rect 20188 7980 20244 7982
rect 21980 8876 22036 8932
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19740 7644 19796 7700
rect 20300 7644 20356 7700
rect 17948 6524 18004 6580
rect 19964 6578 20020 6580
rect 19964 6526 19966 6578
rect 19966 6526 20018 6578
rect 20018 6526 20020 6578
rect 19964 6524 20020 6526
rect 19292 6412 19348 6468
rect 17948 5906 18004 5908
rect 17948 5854 17950 5906
rect 17950 5854 18002 5906
rect 18002 5854 18004 5906
rect 17948 5852 18004 5854
rect 17948 5292 18004 5348
rect 17500 4844 17556 4900
rect 17836 5180 17892 5236
rect 18172 5628 18228 5684
rect 17388 4450 17444 4452
rect 17388 4398 17390 4450
rect 17390 4398 17442 4450
rect 17442 4398 17444 4450
rect 17388 4396 17444 4398
rect 17612 3554 17668 3556
rect 17612 3502 17614 3554
rect 17614 3502 17666 3554
rect 17666 3502 17668 3554
rect 17612 3500 17668 3502
rect 18956 5682 19012 5684
rect 18956 5630 18958 5682
rect 18958 5630 19010 5682
rect 19010 5630 19012 5682
rect 18956 5628 19012 5630
rect 18508 5068 18564 5124
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 20076 5852 20132 5908
rect 19516 5234 19572 5236
rect 19516 5182 19518 5234
rect 19518 5182 19570 5234
rect 19570 5182 19572 5234
rect 19516 5180 19572 5182
rect 20748 6524 20804 6580
rect 20860 6130 20916 6132
rect 20860 6078 20862 6130
rect 20862 6078 20914 6130
rect 20914 6078 20916 6130
rect 20860 6076 20916 6078
rect 21756 6524 21812 6580
rect 21420 6466 21476 6468
rect 21420 6414 21422 6466
rect 21422 6414 21474 6466
rect 21474 6414 21476 6466
rect 21420 6412 21476 6414
rect 21532 5964 21588 6020
rect 21196 5906 21252 5908
rect 21196 5854 21198 5906
rect 21198 5854 21250 5906
rect 21250 5854 21252 5906
rect 21196 5852 21252 5854
rect 21980 5964 22036 6020
rect 20300 5292 20356 5348
rect 21308 5740 21364 5796
rect 20524 5292 20580 5348
rect 21532 5740 21588 5796
rect 21644 5122 21700 5124
rect 21644 5070 21646 5122
rect 21646 5070 21698 5122
rect 21698 5070 21700 5122
rect 21644 5068 21700 5070
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 20300 4172 20356 4228
rect 21084 4284 21140 4340
rect 20860 3612 20916 3668
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 24332 17778 24388 17780
rect 24332 17726 24334 17778
rect 24334 17726 24386 17778
rect 24386 17726 24388 17778
rect 24332 17724 24388 17726
rect 25004 19740 25060 19796
rect 25228 18450 25284 18452
rect 25228 18398 25230 18450
rect 25230 18398 25282 18450
rect 25282 18398 25284 18450
rect 25228 18396 25284 18398
rect 24444 16882 24500 16884
rect 24444 16830 24446 16882
rect 24446 16830 24498 16882
rect 24498 16830 24500 16882
rect 24444 16828 24500 16830
rect 24556 18284 24612 18340
rect 24220 14588 24276 14644
rect 25452 17388 25508 17444
rect 24444 15538 24500 15540
rect 24444 15486 24446 15538
rect 24446 15486 24498 15538
rect 24498 15486 24500 15538
rect 24444 15484 24500 15486
rect 24108 14530 24164 14532
rect 24108 14478 24110 14530
rect 24110 14478 24162 14530
rect 24162 14478 24164 14530
rect 24108 14476 24164 14478
rect 24444 13692 24500 13748
rect 23884 13580 23940 13636
rect 23324 12908 23380 12964
rect 23436 12012 23492 12068
rect 23772 11900 23828 11956
rect 22764 11004 22820 11060
rect 23436 9996 23492 10052
rect 22652 8876 22708 8932
rect 22428 8428 22484 8484
rect 22988 8258 23044 8260
rect 22988 8206 22990 8258
rect 22990 8206 23042 8258
rect 23042 8206 23044 8258
rect 22988 8204 23044 8206
rect 22540 8146 22596 8148
rect 22540 8094 22542 8146
rect 22542 8094 22594 8146
rect 22594 8094 22596 8146
rect 22540 8092 22596 8094
rect 24108 12738 24164 12740
rect 24108 12686 24110 12738
rect 24110 12686 24162 12738
rect 24162 12686 24164 12738
rect 24108 12684 24164 12686
rect 23772 8204 23828 8260
rect 23884 8316 23940 8372
rect 23660 8092 23716 8148
rect 23212 7532 23268 7588
rect 24108 7980 24164 8036
rect 24108 7586 24164 7588
rect 24108 7534 24110 7586
rect 24110 7534 24162 7586
rect 24162 7534 24164 7586
rect 24108 7532 24164 7534
rect 22652 7474 22708 7476
rect 22652 7422 22654 7474
rect 22654 7422 22706 7474
rect 22706 7422 22708 7474
rect 22652 7420 22708 7422
rect 22428 6860 22484 6916
rect 22428 5794 22484 5796
rect 22428 5742 22430 5794
rect 22430 5742 22482 5794
rect 22482 5742 22484 5794
rect 22428 5740 22484 5742
rect 22204 5516 22260 5572
rect 22316 5628 22372 5684
rect 22764 5516 22820 5572
rect 22428 4396 22484 4452
rect 21420 4226 21476 4228
rect 21420 4174 21422 4226
rect 21422 4174 21474 4226
rect 21474 4174 21476 4226
rect 21420 4172 21476 4174
rect 22092 3666 22148 3668
rect 22092 3614 22094 3666
rect 22094 3614 22146 3666
rect 22146 3614 22148 3666
rect 22092 3612 22148 3614
rect 23660 5292 23716 5348
rect 23436 5180 23492 5236
rect 23548 5068 23604 5124
rect 24668 16044 24724 16100
rect 24780 15260 24836 15316
rect 24668 12236 24724 12292
rect 25340 17052 25396 17108
rect 25228 16828 25284 16884
rect 27020 23826 27076 23828
rect 27020 23774 27022 23826
rect 27022 23774 27074 23826
rect 27074 23774 27076 23826
rect 27020 23772 27076 23774
rect 27804 28364 27860 28420
rect 27916 28140 27972 28196
rect 28476 29484 28532 29540
rect 28252 28476 28308 28532
rect 28028 26796 28084 26852
rect 27244 23996 27300 24052
rect 27580 23884 27636 23940
rect 27356 23714 27412 23716
rect 27356 23662 27358 23714
rect 27358 23662 27410 23714
rect 27410 23662 27412 23714
rect 27356 23660 27412 23662
rect 27468 23548 27524 23604
rect 27132 23324 27188 23380
rect 27804 25394 27860 25396
rect 27804 25342 27806 25394
rect 27806 25342 27858 25394
rect 27858 25342 27860 25394
rect 27804 25340 27860 25342
rect 27916 23996 27972 24052
rect 28140 23938 28196 23940
rect 28140 23886 28142 23938
rect 28142 23886 28194 23938
rect 28194 23886 28196 23938
rect 28140 23884 28196 23886
rect 28028 23100 28084 23156
rect 27580 21756 27636 21812
rect 27804 22146 27860 22148
rect 27804 22094 27806 22146
rect 27806 22094 27858 22146
rect 27858 22094 27860 22146
rect 27804 22092 27860 22094
rect 26796 20018 26852 20020
rect 26796 19966 26798 20018
rect 26798 19966 26850 20018
rect 26850 19966 26852 20018
rect 26796 19964 26852 19966
rect 26348 19906 26404 19908
rect 26348 19854 26350 19906
rect 26350 19854 26402 19906
rect 26402 19854 26404 19906
rect 26348 19852 26404 19854
rect 26348 18396 26404 18452
rect 27804 21420 27860 21476
rect 27580 20188 27636 20244
rect 27692 19964 27748 20020
rect 27468 18284 27524 18340
rect 25788 17724 25844 17780
rect 27692 17724 27748 17780
rect 26348 17500 26404 17556
rect 26908 17612 26964 17668
rect 26908 16492 26964 16548
rect 26012 15484 26068 15540
rect 25900 15260 25956 15316
rect 25788 15202 25844 15204
rect 25788 15150 25790 15202
rect 25790 15150 25842 15202
rect 25842 15150 25844 15202
rect 25788 15148 25844 15150
rect 25004 14642 25060 14644
rect 25004 14590 25006 14642
rect 25006 14590 25058 14642
rect 25058 14590 25060 14642
rect 25004 14588 25060 14590
rect 24892 13580 24948 13636
rect 27132 16156 27188 16212
rect 26236 15148 26292 15204
rect 25340 13634 25396 13636
rect 25340 13582 25342 13634
rect 25342 13582 25394 13634
rect 25394 13582 25396 13634
rect 25340 13580 25396 13582
rect 27020 15820 27076 15876
rect 27244 17554 27300 17556
rect 27244 17502 27246 17554
rect 27246 17502 27298 17554
rect 27298 17502 27300 17554
rect 27244 17500 27300 17502
rect 28588 28364 28644 28420
rect 28476 28028 28532 28084
rect 28812 32562 28868 32564
rect 28812 32510 28814 32562
rect 28814 32510 28866 32562
rect 28866 32510 28868 32562
rect 28812 32508 28868 32510
rect 29484 33458 29540 33460
rect 29484 33406 29486 33458
rect 29486 33406 29538 33458
rect 29538 33406 29540 33458
rect 29484 33404 29540 33406
rect 29372 33346 29428 33348
rect 29372 33294 29374 33346
rect 29374 33294 29426 33346
rect 29426 33294 29428 33346
rect 29372 33292 29428 33294
rect 30492 35420 30548 35476
rect 30716 35698 30772 35700
rect 30716 35646 30718 35698
rect 30718 35646 30770 35698
rect 30770 35646 30772 35698
rect 30716 35644 30772 35646
rect 31052 35698 31108 35700
rect 31052 35646 31054 35698
rect 31054 35646 31106 35698
rect 31106 35646 31108 35698
rect 31052 35644 31108 35646
rect 30604 35308 30660 35364
rect 29932 34802 29988 34804
rect 29932 34750 29934 34802
rect 29934 34750 29986 34802
rect 29986 34750 29988 34802
rect 29932 34748 29988 34750
rect 29932 34076 29988 34132
rect 29596 32844 29652 32900
rect 29372 32172 29428 32228
rect 30268 32956 30324 33012
rect 30380 33180 30436 33236
rect 30380 32732 30436 32788
rect 29820 32674 29876 32676
rect 29820 32622 29822 32674
rect 29822 32622 29874 32674
rect 29874 32622 29876 32674
rect 29820 32620 29876 32622
rect 29036 31500 29092 31556
rect 30268 31612 30324 31668
rect 28924 30044 28980 30100
rect 29372 29260 29428 29316
rect 29260 28530 29316 28532
rect 29260 28478 29262 28530
rect 29262 28478 29314 28530
rect 29314 28478 29316 28530
rect 29260 28476 29316 28478
rect 29148 28364 29204 28420
rect 29148 27692 29204 27748
rect 28812 26684 28868 26740
rect 28924 26124 28980 26180
rect 28476 25394 28532 25396
rect 28476 25342 28478 25394
rect 28478 25342 28530 25394
rect 28530 25342 28532 25394
rect 28476 25340 28532 25342
rect 28588 25116 28644 25172
rect 28476 23826 28532 23828
rect 28476 23774 28478 23826
rect 28478 23774 28530 23826
rect 28530 23774 28532 23826
rect 28476 23772 28532 23774
rect 28588 23714 28644 23716
rect 28588 23662 28590 23714
rect 28590 23662 28642 23714
rect 28642 23662 28644 23714
rect 28588 23660 28644 23662
rect 29148 23938 29204 23940
rect 29148 23886 29150 23938
rect 29150 23886 29202 23938
rect 29202 23886 29204 23938
rect 29148 23884 29204 23886
rect 29484 28476 29540 28532
rect 29596 27692 29652 27748
rect 29708 27580 29764 27636
rect 29372 23996 29428 24052
rect 29820 26962 29876 26964
rect 29820 26910 29822 26962
rect 29822 26910 29874 26962
rect 29874 26910 29876 26962
rect 29820 26908 29876 26910
rect 31164 34524 31220 34580
rect 32060 40962 32116 40964
rect 32060 40910 32062 40962
rect 32062 40910 32114 40962
rect 32114 40910 32116 40962
rect 32060 40908 32116 40910
rect 32508 40908 32564 40964
rect 32396 40626 32452 40628
rect 32396 40574 32398 40626
rect 32398 40574 32450 40626
rect 32450 40574 32452 40626
rect 32396 40572 32452 40574
rect 31836 40124 31892 40180
rect 31948 40236 32004 40292
rect 32172 38946 32228 38948
rect 32172 38894 32174 38946
rect 32174 38894 32226 38946
rect 32226 38894 32228 38946
rect 32172 38892 32228 38894
rect 31612 38780 31668 38836
rect 31948 38780 32004 38836
rect 31388 37884 31444 37940
rect 31500 36204 31556 36260
rect 31388 35810 31444 35812
rect 31388 35758 31390 35810
rect 31390 35758 31442 35810
rect 31442 35758 31444 35810
rect 31388 35756 31444 35758
rect 31500 35532 31556 35588
rect 31500 35308 31556 35364
rect 32396 39340 32452 39396
rect 32732 40908 32788 40964
rect 34748 43538 34804 43540
rect 34748 43486 34750 43538
rect 34750 43486 34802 43538
rect 34802 43486 34804 43538
rect 34748 43484 34804 43486
rect 34524 43260 34580 43316
rect 33964 42252 34020 42308
rect 33964 42028 34020 42084
rect 33740 41186 33796 41188
rect 33740 41134 33742 41186
rect 33742 41134 33794 41186
rect 33794 41134 33796 41186
rect 33740 41132 33796 41134
rect 33404 41020 33460 41076
rect 33852 41074 33908 41076
rect 33852 41022 33854 41074
rect 33854 41022 33906 41074
rect 33906 41022 33908 41074
rect 33852 41020 33908 41022
rect 32620 39004 32676 39060
rect 32172 38108 32228 38164
rect 32060 37154 32116 37156
rect 32060 37102 32062 37154
rect 32062 37102 32114 37154
rect 32114 37102 32116 37154
rect 32060 37100 32116 37102
rect 31724 35308 31780 35364
rect 31836 35644 31892 35700
rect 33292 38780 33348 38836
rect 32732 38162 32788 38164
rect 32732 38110 32734 38162
rect 32734 38110 32786 38162
rect 32786 38110 32788 38162
rect 32732 38108 32788 38110
rect 33180 37154 33236 37156
rect 33180 37102 33182 37154
rect 33182 37102 33234 37154
rect 33234 37102 33236 37154
rect 33180 37100 33236 37102
rect 32172 35698 32228 35700
rect 32172 35646 32174 35698
rect 32174 35646 32226 35698
rect 32226 35646 32228 35698
rect 32172 35644 32228 35646
rect 32172 35420 32228 35476
rect 31836 34748 31892 34804
rect 32060 35308 32116 35364
rect 31276 33404 31332 33460
rect 32172 33852 32228 33908
rect 31164 33068 31220 33124
rect 32060 32060 32116 32116
rect 31164 31388 31220 31444
rect 31052 30268 31108 30324
rect 30380 29932 30436 29988
rect 30268 28364 30324 28420
rect 30044 28082 30100 28084
rect 30044 28030 30046 28082
rect 30046 28030 30098 28082
rect 30098 28030 30100 28082
rect 30044 28028 30100 28030
rect 30156 27804 30212 27860
rect 30716 28364 30772 28420
rect 30492 27468 30548 27524
rect 31388 30434 31444 30436
rect 31388 30382 31390 30434
rect 31390 30382 31442 30434
rect 31442 30382 31444 30434
rect 31388 30380 31444 30382
rect 31500 30268 31556 30324
rect 31164 29932 31220 29988
rect 31724 29932 31780 29988
rect 33180 36876 33236 36932
rect 33068 36316 33124 36372
rect 33068 35308 33124 35364
rect 33068 34748 33124 34804
rect 33068 33292 33124 33348
rect 32396 32508 32452 32564
rect 32060 30322 32116 30324
rect 32060 30270 32062 30322
rect 32062 30270 32114 30322
rect 32114 30270 32116 30322
rect 32060 30268 32116 30270
rect 31836 29708 31892 29764
rect 32172 30044 32228 30100
rect 31612 28812 31668 28868
rect 31164 28364 31220 28420
rect 31276 28082 31332 28084
rect 31276 28030 31278 28082
rect 31278 28030 31330 28082
rect 31330 28030 31332 28082
rect 31276 28028 31332 28030
rect 32172 28364 32228 28420
rect 31948 28028 32004 28084
rect 32060 28140 32116 28196
rect 31836 27804 31892 27860
rect 29484 23826 29540 23828
rect 29484 23774 29486 23826
rect 29486 23774 29538 23826
rect 29538 23774 29540 23826
rect 29484 23772 29540 23774
rect 29260 23212 29316 23268
rect 29372 23660 29428 23716
rect 29148 22482 29204 22484
rect 29148 22430 29150 22482
rect 29150 22430 29202 22482
rect 29202 22430 29204 22482
rect 29148 22428 29204 22430
rect 29596 22316 29652 22372
rect 28476 22146 28532 22148
rect 28476 22094 28478 22146
rect 28478 22094 28530 22146
rect 28530 22094 28532 22146
rect 28476 22092 28532 22094
rect 28812 21810 28868 21812
rect 28812 21758 28814 21810
rect 28814 21758 28866 21810
rect 28866 21758 28868 21810
rect 28812 21756 28868 21758
rect 31500 27186 31556 27188
rect 31500 27134 31502 27186
rect 31502 27134 31554 27186
rect 31554 27134 31556 27186
rect 31500 27132 31556 27134
rect 31500 26908 31556 26964
rect 32284 27356 32340 27412
rect 32844 27356 32900 27412
rect 32508 27132 32564 27188
rect 32396 27020 32452 27076
rect 32620 27074 32676 27076
rect 32620 27022 32622 27074
rect 32622 27022 32674 27074
rect 32674 27022 32676 27074
rect 32620 27020 32676 27022
rect 32060 26908 32116 26964
rect 32844 26852 32900 26908
rect 32732 26684 32788 26740
rect 31612 25004 31668 25060
rect 32508 25228 32564 25284
rect 31164 24220 31220 24276
rect 30492 24162 30548 24164
rect 30492 24110 30494 24162
rect 30494 24110 30546 24162
rect 30546 24110 30548 24162
rect 30492 24108 30548 24110
rect 30156 23772 30212 23828
rect 28476 21420 28532 21476
rect 28364 20188 28420 20244
rect 28364 20018 28420 20020
rect 28364 19966 28366 20018
rect 28366 19966 28418 20018
rect 28418 19966 28420 20018
rect 28364 19964 28420 19966
rect 28476 18844 28532 18900
rect 27804 17500 27860 17556
rect 27356 17442 27412 17444
rect 27356 17390 27358 17442
rect 27358 17390 27410 17442
rect 27410 17390 27412 17442
rect 27356 17388 27412 17390
rect 27356 16940 27412 16996
rect 28028 17778 28084 17780
rect 28028 17726 28030 17778
rect 28030 17726 28082 17778
rect 28082 17726 28084 17778
rect 28028 17724 28084 17726
rect 29484 21026 29540 21028
rect 29484 20974 29486 21026
rect 29486 20974 29538 21026
rect 29538 20974 29540 21026
rect 29484 20972 29540 20974
rect 30492 21698 30548 21700
rect 30492 21646 30494 21698
rect 30494 21646 30546 21698
rect 30546 21646 30548 21698
rect 30492 21644 30548 21646
rect 29596 20524 29652 20580
rect 30268 20578 30324 20580
rect 30268 20526 30270 20578
rect 30270 20526 30322 20578
rect 30322 20526 30324 20578
rect 30268 20524 30324 20526
rect 29036 20188 29092 20244
rect 29484 20188 29540 20244
rect 30380 20130 30436 20132
rect 30380 20078 30382 20130
rect 30382 20078 30434 20130
rect 30434 20078 30436 20130
rect 30380 20076 30436 20078
rect 29260 19180 29316 19236
rect 28812 17724 28868 17780
rect 29148 17778 29204 17780
rect 29148 17726 29150 17778
rect 29150 17726 29202 17778
rect 29202 17726 29204 17778
rect 29148 17724 29204 17726
rect 27916 16828 27972 16884
rect 27356 15820 27412 15876
rect 27692 15484 27748 15540
rect 26460 14588 26516 14644
rect 28028 16940 28084 16996
rect 27916 15314 27972 15316
rect 27916 15262 27918 15314
rect 27918 15262 27970 15314
rect 27970 15262 27972 15314
rect 27916 15260 27972 15262
rect 28140 16210 28196 16212
rect 28140 16158 28142 16210
rect 28142 16158 28194 16210
rect 28194 16158 28196 16210
rect 28140 16156 28196 16158
rect 28140 15314 28196 15316
rect 28140 15262 28142 15314
rect 28142 15262 28194 15314
rect 28194 15262 28196 15314
rect 28140 15260 28196 15262
rect 26460 13916 26516 13972
rect 28588 16604 28644 16660
rect 30828 22428 30884 22484
rect 30828 21756 30884 21812
rect 30716 20972 30772 21028
rect 30716 20578 30772 20580
rect 30716 20526 30718 20578
rect 30718 20526 30770 20578
rect 30770 20526 30772 20578
rect 30716 20524 30772 20526
rect 31052 21474 31108 21476
rect 31052 21422 31054 21474
rect 31054 21422 31106 21474
rect 31106 21422 31108 21474
rect 31052 21420 31108 21422
rect 31276 23436 31332 23492
rect 31276 22876 31332 22932
rect 31948 23826 32004 23828
rect 31948 23774 31950 23826
rect 31950 23774 32002 23826
rect 32002 23774 32004 23826
rect 31948 23772 32004 23774
rect 31836 23154 31892 23156
rect 31836 23102 31838 23154
rect 31838 23102 31890 23154
rect 31890 23102 31892 23154
rect 31836 23100 31892 23102
rect 32508 23100 32564 23156
rect 31276 22258 31332 22260
rect 31276 22206 31278 22258
rect 31278 22206 31330 22258
rect 31330 22206 31332 22258
rect 31276 22204 31332 22206
rect 31276 21586 31332 21588
rect 31276 21534 31278 21586
rect 31278 21534 31330 21586
rect 31330 21534 31332 21586
rect 31276 21532 31332 21534
rect 31164 21308 31220 21364
rect 31724 22092 31780 22148
rect 31836 21756 31892 21812
rect 30940 19964 30996 20020
rect 30492 19740 30548 19796
rect 30380 19628 30436 19684
rect 30044 19234 30100 19236
rect 30044 19182 30046 19234
rect 30046 19182 30098 19234
rect 30098 19182 30100 19234
rect 30044 19180 30100 19182
rect 31164 20578 31220 20580
rect 31164 20526 31166 20578
rect 31166 20526 31218 20578
rect 31218 20526 31220 20578
rect 31164 20524 31220 20526
rect 31500 19906 31556 19908
rect 31500 19854 31502 19906
rect 31502 19854 31554 19906
rect 31554 19854 31556 19906
rect 31500 19852 31556 19854
rect 30716 19234 30772 19236
rect 30716 19182 30718 19234
rect 30718 19182 30770 19234
rect 30770 19182 30772 19234
rect 30716 19180 30772 19182
rect 30156 19122 30212 19124
rect 30156 19070 30158 19122
rect 30158 19070 30210 19122
rect 30210 19070 30212 19122
rect 30156 19068 30212 19070
rect 29932 19010 29988 19012
rect 29932 18958 29934 19010
rect 29934 18958 29986 19010
rect 29986 18958 29988 19010
rect 29932 18956 29988 18958
rect 29708 16940 29764 16996
rect 30044 18844 30100 18900
rect 29708 16604 29764 16660
rect 28588 16098 28644 16100
rect 28588 16046 28590 16098
rect 28590 16046 28642 16098
rect 28642 16046 28644 16098
rect 28588 16044 28644 16046
rect 28476 15986 28532 15988
rect 28476 15934 28478 15986
rect 28478 15934 28530 15986
rect 28530 15934 28532 15986
rect 28476 15932 28532 15934
rect 29148 16210 29204 16212
rect 29148 16158 29150 16210
rect 29150 16158 29202 16210
rect 29202 16158 29204 16210
rect 29148 16156 29204 16158
rect 29260 16044 29316 16100
rect 28588 15314 28644 15316
rect 28588 15262 28590 15314
rect 28590 15262 28642 15314
rect 28642 15262 28644 15314
rect 28588 15260 28644 15262
rect 28476 15202 28532 15204
rect 28476 15150 28478 15202
rect 28478 15150 28530 15202
rect 28530 15150 28532 15202
rect 28476 15148 28532 15150
rect 28028 14364 28084 14420
rect 27356 13692 27412 13748
rect 25228 12460 25284 12516
rect 25452 12572 25508 12628
rect 25228 11954 25284 11956
rect 25228 11902 25230 11954
rect 25230 11902 25282 11954
rect 25282 11902 25284 11954
rect 25228 11900 25284 11902
rect 25900 12738 25956 12740
rect 25900 12686 25902 12738
rect 25902 12686 25954 12738
rect 25954 12686 25956 12738
rect 25900 12684 25956 12686
rect 26572 12962 26628 12964
rect 26572 12910 26574 12962
rect 26574 12910 26626 12962
rect 26626 12910 26628 12962
rect 26572 12908 26628 12910
rect 26908 12850 26964 12852
rect 26908 12798 26910 12850
rect 26910 12798 26962 12850
rect 26962 12798 26964 12850
rect 26908 12796 26964 12798
rect 27244 12796 27300 12852
rect 26460 12738 26516 12740
rect 26460 12686 26462 12738
rect 26462 12686 26514 12738
rect 26514 12686 26516 12738
rect 26460 12684 26516 12686
rect 26124 12460 26180 12516
rect 25788 12290 25844 12292
rect 25788 12238 25790 12290
rect 25790 12238 25842 12290
rect 25842 12238 25844 12290
rect 25788 12236 25844 12238
rect 25676 12012 25732 12068
rect 26236 12012 26292 12068
rect 25004 10444 25060 10500
rect 25116 9996 25172 10052
rect 25676 10498 25732 10500
rect 25676 10446 25678 10498
rect 25678 10446 25730 10498
rect 25730 10446 25732 10498
rect 25676 10444 25732 10446
rect 25452 9100 25508 9156
rect 24556 8370 24612 8372
rect 24556 8318 24558 8370
rect 24558 8318 24610 8370
rect 24610 8318 24612 8370
rect 24556 8316 24612 8318
rect 25228 8146 25284 8148
rect 25228 8094 25230 8146
rect 25230 8094 25282 8146
rect 25282 8094 25284 8146
rect 25228 8092 25284 8094
rect 25452 8092 25508 8148
rect 24556 7868 24612 7924
rect 25676 8204 25732 8260
rect 26124 9548 26180 9604
rect 26236 9772 26292 9828
rect 25900 9154 25956 9156
rect 25900 9102 25902 9154
rect 25902 9102 25954 9154
rect 25954 9102 25956 9154
rect 25900 9100 25956 9102
rect 26012 8876 26068 8932
rect 25788 8092 25844 8148
rect 25564 7980 25620 8036
rect 24556 6860 24612 6916
rect 24332 6636 24388 6692
rect 24220 6578 24276 6580
rect 24220 6526 24222 6578
rect 24222 6526 24274 6578
rect 24274 6526 24276 6578
rect 24220 6524 24276 6526
rect 23772 5068 23828 5124
rect 24668 5234 24724 5236
rect 24668 5182 24670 5234
rect 24670 5182 24722 5234
rect 24722 5182 24724 5234
rect 24668 5180 24724 5182
rect 24780 6636 24836 6692
rect 25228 6018 25284 6020
rect 25228 5966 25230 6018
rect 25230 5966 25282 6018
rect 25282 5966 25284 6018
rect 25228 5964 25284 5966
rect 25340 5852 25396 5908
rect 23548 4898 23604 4900
rect 23548 4846 23550 4898
rect 23550 4846 23602 4898
rect 23602 4846 23604 4898
rect 23548 4844 23604 4846
rect 22652 3724 22708 3780
rect 24556 3778 24612 3780
rect 24556 3726 24558 3778
rect 24558 3726 24610 3778
rect 24610 3726 24612 3778
rect 24556 3724 24612 3726
rect 26012 7420 26068 7476
rect 26236 7362 26292 7364
rect 26236 7310 26238 7362
rect 26238 7310 26290 7362
rect 26290 7310 26292 7362
rect 26236 7308 26292 7310
rect 26124 6636 26180 6692
rect 25900 5682 25956 5684
rect 25900 5630 25902 5682
rect 25902 5630 25954 5682
rect 25954 5630 25956 5682
rect 25900 5628 25956 5630
rect 25788 4956 25844 5012
rect 25228 4450 25284 4452
rect 25228 4398 25230 4450
rect 25230 4398 25282 4450
rect 25282 4398 25284 4450
rect 25228 4396 25284 4398
rect 24668 3500 24724 3556
rect 26124 5068 26180 5124
rect 26684 12290 26740 12292
rect 26684 12238 26686 12290
rect 26686 12238 26738 12290
rect 26738 12238 26740 12290
rect 26684 12236 26740 12238
rect 26460 6748 26516 6804
rect 26572 7308 26628 7364
rect 27132 9042 27188 9044
rect 27132 8990 27134 9042
rect 27134 8990 27186 9042
rect 27186 8990 27188 9042
rect 27132 8988 27188 8990
rect 27020 8876 27076 8932
rect 26684 6636 26740 6692
rect 27692 13020 27748 13076
rect 28364 14306 28420 14308
rect 28364 14254 28366 14306
rect 28366 14254 28418 14306
rect 28418 14254 28420 14306
rect 28364 14252 28420 14254
rect 29596 15874 29652 15876
rect 29596 15822 29598 15874
rect 29598 15822 29650 15874
rect 29650 15822 29652 15874
rect 29596 15820 29652 15822
rect 29820 15874 29876 15876
rect 29820 15822 29822 15874
rect 29822 15822 29874 15874
rect 29874 15822 29876 15874
rect 29820 15820 29876 15822
rect 28364 13970 28420 13972
rect 28364 13918 28366 13970
rect 28366 13918 28418 13970
rect 28418 13918 28420 13970
rect 28364 13916 28420 13918
rect 29484 13132 29540 13188
rect 29372 13074 29428 13076
rect 29372 13022 29374 13074
rect 29374 13022 29426 13074
rect 29426 13022 29428 13074
rect 29372 13020 29428 13022
rect 31388 19740 31444 19796
rect 30716 18620 30772 18676
rect 30940 19010 30996 19012
rect 30940 18958 30942 19010
rect 30942 18958 30994 19010
rect 30994 18958 30996 19010
rect 30940 18956 30996 18958
rect 30828 17724 30884 17780
rect 30268 16882 30324 16884
rect 30268 16830 30270 16882
rect 30270 16830 30322 16882
rect 30322 16830 30324 16882
rect 30268 16828 30324 16830
rect 30716 15932 30772 15988
rect 30268 15874 30324 15876
rect 30268 15822 30270 15874
rect 30270 15822 30322 15874
rect 30322 15822 30324 15874
rect 30268 15820 30324 15822
rect 30604 15314 30660 15316
rect 30604 15262 30606 15314
rect 30606 15262 30658 15314
rect 30658 15262 30660 15314
rect 30604 15260 30660 15262
rect 27804 12236 27860 12292
rect 30156 14418 30212 14420
rect 30156 14366 30158 14418
rect 30158 14366 30210 14418
rect 30210 14366 30212 14418
rect 30156 14364 30212 14366
rect 29932 14252 29988 14308
rect 30156 13746 30212 13748
rect 30156 13694 30158 13746
rect 30158 13694 30210 13746
rect 30210 13694 30212 13746
rect 30156 13692 30212 13694
rect 29036 12290 29092 12292
rect 29036 12238 29038 12290
rect 29038 12238 29090 12290
rect 29090 12238 29092 12290
rect 29036 12236 29092 12238
rect 29148 12684 29204 12740
rect 29708 12796 29764 12852
rect 29820 12738 29876 12740
rect 29820 12686 29822 12738
rect 29822 12686 29874 12738
rect 29874 12686 29876 12738
rect 29820 12684 29876 12686
rect 29820 12124 29876 12180
rect 30716 12796 30772 12852
rect 30604 12684 30660 12740
rect 31276 17276 31332 17332
rect 31164 16994 31220 16996
rect 31164 16942 31166 16994
rect 31166 16942 31218 16994
rect 31218 16942 31220 16994
rect 31164 16940 31220 16942
rect 31500 19010 31556 19012
rect 31500 18958 31502 19010
rect 31502 18958 31554 19010
rect 31554 18958 31556 19010
rect 31500 18956 31556 18958
rect 31500 18562 31556 18564
rect 31500 18510 31502 18562
rect 31502 18510 31554 18562
rect 31554 18510 31556 18562
rect 31500 18508 31556 18510
rect 31836 20130 31892 20132
rect 31836 20078 31838 20130
rect 31838 20078 31890 20130
rect 31890 20078 31892 20130
rect 31836 20076 31892 20078
rect 32060 21980 32116 22036
rect 31836 19852 31892 19908
rect 31948 19794 32004 19796
rect 31948 19742 31950 19794
rect 31950 19742 32002 19794
rect 32002 19742 32004 19794
rect 31948 19740 32004 19742
rect 31836 17276 31892 17332
rect 31500 17052 31556 17108
rect 31276 16716 31332 16772
rect 31276 15932 31332 15988
rect 31500 15484 31556 15540
rect 31724 17052 31780 17108
rect 31948 16994 32004 16996
rect 31948 16942 31950 16994
rect 31950 16942 32002 16994
rect 32002 16942 32004 16994
rect 31948 16940 32004 16942
rect 32060 16828 32116 16884
rect 31836 15538 31892 15540
rect 31836 15486 31838 15538
rect 31838 15486 31890 15538
rect 31890 15486 31892 15538
rect 31836 15484 31892 15486
rect 31724 15426 31780 15428
rect 31724 15374 31726 15426
rect 31726 15374 31778 15426
rect 31778 15374 31780 15426
rect 31724 15372 31780 15374
rect 31052 13692 31108 13748
rect 31388 13746 31444 13748
rect 31388 13694 31390 13746
rect 31390 13694 31442 13746
rect 31442 13694 31444 13746
rect 31388 13692 31444 13694
rect 31836 13746 31892 13748
rect 31836 13694 31838 13746
rect 31838 13694 31890 13746
rect 31890 13694 31892 13746
rect 31836 13692 31892 13694
rect 31724 13634 31780 13636
rect 31724 13582 31726 13634
rect 31726 13582 31778 13634
rect 31778 13582 31780 13634
rect 31724 13580 31780 13582
rect 32060 13244 32116 13300
rect 30492 12236 30548 12292
rect 30940 12178 30996 12180
rect 30940 12126 30942 12178
rect 30942 12126 30994 12178
rect 30994 12126 30996 12178
rect 30940 12124 30996 12126
rect 31388 12402 31444 12404
rect 31388 12350 31390 12402
rect 31390 12350 31442 12402
rect 31442 12350 31444 12402
rect 31388 12348 31444 12350
rect 31276 12290 31332 12292
rect 31276 12238 31278 12290
rect 31278 12238 31330 12290
rect 31330 12238 31332 12290
rect 31276 12236 31332 12238
rect 32060 12402 32116 12404
rect 32060 12350 32062 12402
rect 32062 12350 32114 12402
rect 32114 12350 32116 12402
rect 32060 12348 32116 12350
rect 30828 11170 30884 11172
rect 30828 11118 30830 11170
rect 30830 11118 30882 11170
rect 30882 11118 30884 11170
rect 30828 11116 30884 11118
rect 30492 10668 30548 10724
rect 27580 9826 27636 9828
rect 27580 9774 27582 9826
rect 27582 9774 27634 9826
rect 27634 9774 27636 9826
rect 27580 9772 27636 9774
rect 27468 9714 27524 9716
rect 27468 9662 27470 9714
rect 27470 9662 27522 9714
rect 27522 9662 27524 9714
rect 27468 9660 27524 9662
rect 28700 9660 28756 9716
rect 27916 9548 27972 9604
rect 30716 9548 30772 9604
rect 29596 8988 29652 9044
rect 27804 8316 27860 8372
rect 29148 8876 29204 8932
rect 28252 8034 28308 8036
rect 28252 7982 28254 8034
rect 28254 7982 28306 8034
rect 28306 7982 28308 8034
rect 28252 7980 28308 7982
rect 29260 8370 29316 8372
rect 29260 8318 29262 8370
rect 29262 8318 29314 8370
rect 29314 8318 29316 8370
rect 29260 8316 29316 8318
rect 30828 8988 30884 9044
rect 27468 6524 27524 6580
rect 28252 6860 28308 6916
rect 29484 8146 29540 8148
rect 29484 8094 29486 8146
rect 29486 8094 29538 8146
rect 29538 8094 29540 8146
rect 29484 8092 29540 8094
rect 29036 7084 29092 7140
rect 29596 7084 29652 7140
rect 28364 6636 28420 6692
rect 29372 6690 29428 6692
rect 29372 6638 29374 6690
rect 29374 6638 29426 6690
rect 29426 6638 29428 6690
rect 29372 6636 29428 6638
rect 30268 7084 30324 7140
rect 30380 6748 30436 6804
rect 30044 6690 30100 6692
rect 30044 6638 30046 6690
rect 30046 6638 30098 6690
rect 30098 6638 30100 6690
rect 30044 6636 30100 6638
rect 29148 6578 29204 6580
rect 29148 6526 29150 6578
rect 29150 6526 29202 6578
rect 29202 6526 29204 6578
rect 29148 6524 29204 6526
rect 28588 6466 28644 6468
rect 28588 6414 28590 6466
rect 28590 6414 28642 6466
rect 28642 6414 28644 6466
rect 28588 6412 28644 6414
rect 29596 6412 29652 6468
rect 27356 6300 27412 6356
rect 26348 5404 26404 5460
rect 26348 4844 26404 4900
rect 25900 4172 25956 4228
rect 26908 5516 26964 5572
rect 29148 5234 29204 5236
rect 29148 5182 29150 5234
rect 29150 5182 29202 5234
rect 29202 5182 29204 5234
rect 29148 5180 29204 5182
rect 27804 5068 27860 5124
rect 30044 5292 30100 5348
rect 29260 4956 29316 5012
rect 28700 3778 28756 3780
rect 28700 3726 28702 3778
rect 28702 3726 28754 3778
rect 28754 3726 28756 3778
rect 28700 3724 28756 3726
rect 23996 3276 24052 3332
rect 25228 3330 25284 3332
rect 25228 3278 25230 3330
rect 25230 3278 25282 3330
rect 25282 3278 25284 3330
rect 25228 3276 25284 3278
rect 29484 5122 29540 5124
rect 29484 5070 29486 5122
rect 29486 5070 29538 5122
rect 29538 5070 29540 5122
rect 29484 5068 29540 5070
rect 30940 6860 30996 6916
rect 30604 6466 30660 6468
rect 30604 6414 30606 6466
rect 30606 6414 30658 6466
rect 30658 6414 30660 6466
rect 30604 6412 30660 6414
rect 31052 6300 31108 6356
rect 31052 5628 31108 5684
rect 31276 5292 31332 5348
rect 30492 5068 30548 5124
rect 30380 4898 30436 4900
rect 30380 4846 30382 4898
rect 30382 4846 30434 4898
rect 30434 4846 30436 4898
rect 30380 4844 30436 4846
rect 29260 3724 29316 3780
rect 29036 3554 29092 3556
rect 29036 3502 29038 3554
rect 29038 3502 29090 3554
rect 29090 3502 29092 3554
rect 29036 3500 29092 3502
rect 31948 11788 32004 11844
rect 31500 10332 31556 10388
rect 31948 9548 32004 9604
rect 33740 40572 33796 40628
rect 33628 40402 33684 40404
rect 33628 40350 33630 40402
rect 33630 40350 33682 40402
rect 33682 40350 33684 40402
rect 33628 40348 33684 40350
rect 33740 38834 33796 38836
rect 33740 38782 33742 38834
rect 33742 38782 33794 38834
rect 33794 38782 33796 38834
rect 33740 38780 33796 38782
rect 34300 41186 34356 41188
rect 34300 41134 34302 41186
rect 34302 41134 34354 41186
rect 34354 41134 34356 41186
rect 34300 41132 34356 41134
rect 35644 43708 35700 43764
rect 35420 43260 35476 43316
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 37212 44940 37268 44996
rect 36988 44268 37044 44324
rect 36652 43708 36708 43764
rect 37996 45666 38052 45668
rect 37996 45614 37998 45666
rect 37998 45614 38050 45666
rect 38050 45614 38052 45666
rect 37996 45612 38052 45614
rect 38444 45500 38500 45556
rect 37212 43708 37268 43764
rect 37436 43932 37492 43988
rect 37100 43484 37156 43540
rect 36540 42700 36596 42756
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 36652 42252 36708 42308
rect 38556 45724 38612 45780
rect 39116 45612 39172 45668
rect 39340 45612 39396 45668
rect 38556 44322 38612 44324
rect 38556 44270 38558 44322
rect 38558 44270 38610 44322
rect 38610 44270 38612 44322
rect 38556 44268 38612 44270
rect 39676 44828 39732 44884
rect 38220 43762 38276 43764
rect 38220 43710 38222 43762
rect 38222 43710 38274 43762
rect 38274 43710 38276 43762
rect 38220 43708 38276 43710
rect 38108 43538 38164 43540
rect 38108 43486 38110 43538
rect 38110 43486 38162 43538
rect 38162 43486 38164 43538
rect 38108 43484 38164 43486
rect 37884 42924 37940 42980
rect 37548 42252 37604 42308
rect 39228 43708 39284 43764
rect 38556 43596 38612 43652
rect 38444 43538 38500 43540
rect 38444 43486 38446 43538
rect 38446 43486 38498 43538
rect 38498 43486 38500 43538
rect 38444 43484 38500 43486
rect 39004 43650 39060 43652
rect 39004 43598 39006 43650
rect 39006 43598 39058 43650
rect 39058 43598 39060 43650
rect 39004 43596 39060 43598
rect 39676 43932 39732 43988
rect 39004 42812 39060 42868
rect 36988 41692 37044 41748
rect 36540 41132 36596 41188
rect 34636 41074 34692 41076
rect 34636 41022 34638 41074
rect 34638 41022 34690 41074
rect 34690 41022 34692 41074
rect 34636 41020 34692 41022
rect 34412 40460 34468 40516
rect 34076 39788 34132 39844
rect 34412 39788 34468 39844
rect 34972 40460 35028 40516
rect 34636 39788 34692 39844
rect 34860 39506 34916 39508
rect 34860 39454 34862 39506
rect 34862 39454 34914 39506
rect 34914 39454 34916 39506
rect 34860 39452 34916 39454
rect 34972 39394 35028 39396
rect 34972 39342 34974 39394
rect 34974 39342 35026 39394
rect 35026 39342 35028 39394
rect 34972 39340 35028 39342
rect 34076 39004 34132 39060
rect 34188 39116 34244 39172
rect 33628 38050 33684 38052
rect 33628 37998 33630 38050
rect 33630 37998 33682 38050
rect 33682 37998 33684 38050
rect 33628 37996 33684 37998
rect 33740 37548 33796 37604
rect 33628 37266 33684 37268
rect 33628 37214 33630 37266
rect 33630 37214 33682 37266
rect 33682 37214 33684 37266
rect 33628 37212 33684 37214
rect 33852 37154 33908 37156
rect 33852 37102 33854 37154
rect 33854 37102 33906 37154
rect 33906 37102 33908 37154
rect 33852 37100 33908 37102
rect 33628 36988 33684 37044
rect 33516 36316 33572 36372
rect 33964 36876 34020 36932
rect 35532 41020 35588 41076
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35420 39676 35476 39732
rect 35308 39618 35364 39620
rect 35308 39566 35310 39618
rect 35310 39566 35362 39618
rect 35362 39566 35364 39618
rect 35308 39564 35364 39566
rect 35420 39340 35476 39396
rect 35084 39116 35140 39172
rect 34300 38556 34356 38612
rect 35644 39618 35700 39620
rect 35644 39566 35646 39618
rect 35646 39566 35698 39618
rect 35698 39566 35700 39618
rect 35644 39564 35700 39566
rect 35756 39506 35812 39508
rect 35756 39454 35758 39506
rect 35758 39454 35810 39506
rect 35810 39454 35812 39506
rect 35756 39452 35812 39454
rect 36092 39676 36148 39732
rect 36092 39340 36148 39396
rect 35084 38610 35140 38612
rect 35084 38558 35086 38610
rect 35086 38558 35138 38610
rect 35138 38558 35140 38610
rect 35084 38556 35140 38558
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 34748 37490 34804 37492
rect 34748 37438 34750 37490
rect 34750 37438 34802 37490
rect 34802 37438 34804 37490
rect 34748 37436 34804 37438
rect 35644 37548 35700 37604
rect 35196 37378 35252 37380
rect 35196 37326 35198 37378
rect 35198 37326 35250 37378
rect 35250 37326 35252 37378
rect 35196 37324 35252 37326
rect 34636 37266 34692 37268
rect 34636 37214 34638 37266
rect 34638 37214 34690 37266
rect 34690 37214 34692 37266
rect 34636 37212 34692 37214
rect 35644 37100 35700 37156
rect 34972 36876 35028 36932
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 34188 34972 34244 35028
rect 34524 35586 34580 35588
rect 34524 35534 34526 35586
rect 34526 35534 34578 35586
rect 34578 35534 34580 35586
rect 34524 35532 34580 35534
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35420 35026 35476 35028
rect 35420 34974 35422 35026
rect 35422 34974 35474 35026
rect 35474 34974 35476 35026
rect 35420 34972 35476 34974
rect 34524 34748 34580 34804
rect 34076 34300 34132 34356
rect 33852 33964 33908 34020
rect 36316 39788 36372 39844
rect 37324 41186 37380 41188
rect 37324 41134 37326 41186
rect 37326 41134 37378 41186
rect 37378 41134 37380 41186
rect 37324 41132 37380 41134
rect 37324 39730 37380 39732
rect 37324 39678 37326 39730
rect 37326 39678 37378 39730
rect 37378 39678 37380 39730
rect 37324 39676 37380 39678
rect 37100 39564 37156 39620
rect 36988 38892 37044 38948
rect 38892 41916 38948 41972
rect 38668 40796 38724 40852
rect 37212 39116 37268 39172
rect 38444 39228 38500 39284
rect 36428 38722 36484 38724
rect 36428 38670 36430 38722
rect 36430 38670 36482 38722
rect 36482 38670 36484 38722
rect 36428 38668 36484 38670
rect 36204 37996 36260 38052
rect 36428 38162 36484 38164
rect 36428 38110 36430 38162
rect 36430 38110 36482 38162
rect 36482 38110 36484 38162
rect 36428 38108 36484 38110
rect 36092 37490 36148 37492
rect 36092 37438 36094 37490
rect 36094 37438 36146 37490
rect 36146 37438 36148 37490
rect 36092 37436 36148 37438
rect 37996 38834 38052 38836
rect 37996 38782 37998 38834
rect 37998 38782 38050 38834
rect 38050 38782 38052 38834
rect 37996 38780 38052 38782
rect 38108 38668 38164 38724
rect 38892 40402 38948 40404
rect 38892 40350 38894 40402
rect 38894 40350 38946 40402
rect 38946 40350 38948 40402
rect 38892 40348 38948 40350
rect 37436 38108 37492 38164
rect 36428 37324 36484 37380
rect 36540 37996 36596 38052
rect 36428 36258 36484 36260
rect 36428 36206 36430 36258
rect 36430 36206 36482 36258
rect 36482 36206 36484 36258
rect 36428 36204 36484 36206
rect 36092 36092 36148 36148
rect 35980 35698 36036 35700
rect 35980 35646 35982 35698
rect 35982 35646 36034 35698
rect 36034 35646 36036 35698
rect 35980 35644 36036 35646
rect 36316 35084 36372 35140
rect 37100 37996 37156 38052
rect 38108 37996 38164 38052
rect 38780 37660 38836 37716
rect 38780 37100 38836 37156
rect 37100 36258 37156 36260
rect 37100 36206 37102 36258
rect 37102 36206 37154 36258
rect 37154 36206 37156 36258
rect 37100 36204 37156 36206
rect 36988 35644 37044 35700
rect 37100 35868 37156 35924
rect 36988 35138 37044 35140
rect 36988 35086 36990 35138
rect 36990 35086 37042 35138
rect 37042 35086 37044 35138
rect 36988 35084 37044 35086
rect 36092 34412 36148 34468
rect 33740 33292 33796 33348
rect 33180 32620 33236 32676
rect 33404 32674 33460 32676
rect 33404 32622 33406 32674
rect 33406 32622 33458 32674
rect 33458 32622 33460 32674
rect 33404 32620 33460 32622
rect 36652 34354 36708 34356
rect 36652 34302 36654 34354
rect 36654 34302 36706 34354
rect 36706 34302 36708 34354
rect 36652 34300 36708 34302
rect 36764 34130 36820 34132
rect 36764 34078 36766 34130
rect 36766 34078 36818 34130
rect 36818 34078 36820 34130
rect 36764 34076 36820 34078
rect 36540 33964 36596 34020
rect 36428 33852 36484 33908
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35868 33404 35924 33460
rect 35420 33068 35476 33124
rect 33068 32562 33124 32564
rect 33068 32510 33070 32562
rect 33070 32510 33122 32562
rect 33122 32510 33124 32562
rect 33068 32508 33124 32510
rect 34300 32562 34356 32564
rect 34300 32510 34302 32562
rect 34302 32510 34354 32562
rect 34354 32510 34356 32562
rect 34300 32508 34356 32510
rect 34188 32396 34244 32452
rect 33404 32060 33460 32116
rect 33180 31554 33236 31556
rect 33180 31502 33182 31554
rect 33182 31502 33234 31554
rect 33234 31502 33236 31554
rect 33180 31500 33236 31502
rect 33964 31612 34020 31668
rect 33516 31554 33572 31556
rect 33516 31502 33518 31554
rect 33518 31502 33570 31554
rect 33570 31502 33572 31554
rect 33516 31500 33572 31502
rect 35420 32396 35476 32452
rect 36428 33122 36484 33124
rect 36428 33070 36430 33122
rect 36430 33070 36482 33122
rect 36482 33070 36484 33122
rect 36428 33068 36484 33070
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 33964 31164 34020 31220
rect 33180 30604 33236 30660
rect 34076 30434 34132 30436
rect 34076 30382 34078 30434
rect 34078 30382 34130 30434
rect 34130 30382 34132 30434
rect 34076 30380 34132 30382
rect 33516 30268 33572 30324
rect 34188 30268 34244 30324
rect 34636 30492 34692 30548
rect 34748 31500 34804 31556
rect 34748 30380 34804 30436
rect 34300 30156 34356 30212
rect 34636 30268 34692 30324
rect 33740 30098 33796 30100
rect 33740 30046 33742 30098
rect 33742 30046 33794 30098
rect 33794 30046 33796 30098
rect 33740 30044 33796 30046
rect 33628 29650 33684 29652
rect 33628 29598 33630 29650
rect 33630 29598 33682 29650
rect 33682 29598 33684 29650
rect 33628 29596 33684 29598
rect 33740 29538 33796 29540
rect 33740 29486 33742 29538
rect 33742 29486 33794 29538
rect 33794 29486 33796 29538
rect 33740 29484 33796 29486
rect 33292 28140 33348 28196
rect 33292 27746 33348 27748
rect 33292 27694 33294 27746
rect 33294 27694 33346 27746
rect 33346 27694 33348 27746
rect 33292 27692 33348 27694
rect 33180 27244 33236 27300
rect 33068 26850 33124 26852
rect 33068 26798 33070 26850
rect 33070 26798 33122 26850
rect 33122 26798 33124 26850
rect 33068 26796 33124 26798
rect 32956 25618 33012 25620
rect 32956 25566 32958 25618
rect 32958 25566 33010 25618
rect 33010 25566 33012 25618
rect 32956 25564 33012 25566
rect 33516 28866 33572 28868
rect 33516 28814 33518 28866
rect 33518 28814 33570 28866
rect 33570 28814 33572 28866
rect 33516 28812 33572 28814
rect 33852 28866 33908 28868
rect 33852 28814 33854 28866
rect 33854 28814 33906 28866
rect 33906 28814 33908 28866
rect 33852 28812 33908 28814
rect 34076 29426 34132 29428
rect 34076 29374 34078 29426
rect 34078 29374 34130 29426
rect 34130 29374 34132 29426
rect 34076 29372 34132 29374
rect 33852 28364 33908 28420
rect 33740 27858 33796 27860
rect 33740 27806 33742 27858
rect 33742 27806 33794 27858
rect 33794 27806 33796 27858
rect 33740 27804 33796 27806
rect 33964 27244 34020 27300
rect 34076 27132 34132 27188
rect 33404 27020 33460 27076
rect 33852 27074 33908 27076
rect 33852 27022 33854 27074
rect 33854 27022 33906 27074
rect 33906 27022 33908 27074
rect 33852 27020 33908 27022
rect 35980 31388 36036 31444
rect 35084 30940 35140 30996
rect 34748 28642 34804 28644
rect 34748 28590 34750 28642
rect 34750 28590 34802 28642
rect 34802 28590 34804 28642
rect 34748 28588 34804 28590
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35420 30380 35476 30436
rect 35084 30098 35140 30100
rect 35084 30046 35086 30098
rect 35086 30046 35138 30098
rect 35138 30046 35140 30098
rect 35084 30044 35140 30046
rect 34972 29484 35028 29540
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 34524 27804 34580 27860
rect 34412 27746 34468 27748
rect 34412 27694 34414 27746
rect 34414 27694 34466 27746
rect 34466 27694 34468 27746
rect 34412 27692 34468 27694
rect 34524 27074 34580 27076
rect 34524 27022 34526 27074
rect 34526 27022 34578 27074
rect 34578 27022 34580 27074
rect 34524 27020 34580 27022
rect 33852 26796 33908 26852
rect 33740 26572 33796 26628
rect 34636 26572 34692 26628
rect 33180 25564 33236 25620
rect 33740 25618 33796 25620
rect 33740 25566 33742 25618
rect 33742 25566 33794 25618
rect 33794 25566 33796 25618
rect 33740 25564 33796 25566
rect 33852 25282 33908 25284
rect 33852 25230 33854 25282
rect 33854 25230 33906 25282
rect 33906 25230 33908 25282
rect 33852 25228 33908 25230
rect 33068 23772 33124 23828
rect 32284 22258 32340 22260
rect 32284 22206 32286 22258
rect 32286 22206 32338 22258
rect 32338 22206 32340 22258
rect 32284 22204 32340 22206
rect 32620 22146 32676 22148
rect 32620 22094 32622 22146
rect 32622 22094 32674 22146
rect 32674 22094 32676 22146
rect 32620 22092 32676 22094
rect 32284 21980 32340 22036
rect 32844 21980 32900 22036
rect 32508 21586 32564 21588
rect 32508 21534 32510 21586
rect 32510 21534 32562 21586
rect 32562 21534 32564 21586
rect 32508 21532 32564 21534
rect 32284 21420 32340 21476
rect 33292 23154 33348 23156
rect 33292 23102 33294 23154
rect 33294 23102 33346 23154
rect 33346 23102 33348 23154
rect 33292 23100 33348 23102
rect 34076 24556 34132 24612
rect 34636 23660 34692 23716
rect 34300 23154 34356 23156
rect 34300 23102 34302 23154
rect 34302 23102 34354 23154
rect 34354 23102 34356 23154
rect 34300 23100 34356 23102
rect 33292 20242 33348 20244
rect 33292 20190 33294 20242
rect 33294 20190 33346 20242
rect 33346 20190 33348 20242
rect 33292 20188 33348 20190
rect 33628 21532 33684 21588
rect 33740 22764 33796 22820
rect 33964 22258 34020 22260
rect 33964 22206 33966 22258
rect 33966 22206 34018 22258
rect 34018 22206 34020 22258
rect 33964 22204 34020 22206
rect 34860 27692 34916 27748
rect 34972 23660 35028 23716
rect 34748 23324 34804 23380
rect 34748 23042 34804 23044
rect 34748 22990 34750 23042
rect 34750 22990 34802 23042
rect 34802 22990 34804 23042
rect 34748 22988 34804 22990
rect 34972 22876 35028 22932
rect 34748 21980 34804 22036
rect 34412 21868 34468 21924
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35420 27186 35476 27188
rect 35420 27134 35422 27186
rect 35422 27134 35474 27186
rect 35474 27134 35476 27186
rect 35420 27132 35476 27134
rect 35868 29596 35924 29652
rect 35980 30828 36036 30884
rect 36540 31724 36596 31780
rect 36204 31276 36260 31332
rect 36540 30994 36596 30996
rect 36540 30942 36542 30994
rect 36542 30942 36594 30994
rect 36594 30942 36596 30994
rect 36540 30940 36596 30942
rect 37660 35868 37716 35924
rect 37548 35420 37604 35476
rect 37324 33346 37380 33348
rect 37324 33294 37326 33346
rect 37326 33294 37378 33346
rect 37378 33294 37380 33346
rect 37324 33292 37380 33294
rect 38556 36316 38612 36372
rect 38220 34412 38276 34468
rect 38332 34802 38388 34804
rect 38332 34750 38334 34802
rect 38334 34750 38386 34802
rect 38386 34750 38388 34802
rect 38332 34748 38388 34750
rect 37996 33292 38052 33348
rect 38220 34188 38276 34244
rect 38220 33852 38276 33908
rect 37548 33180 37604 33236
rect 37884 33234 37940 33236
rect 37884 33182 37886 33234
rect 37886 33182 37938 33234
rect 37938 33182 37940 33234
rect 37884 33180 37940 33182
rect 36988 32508 37044 32564
rect 37772 31836 37828 31892
rect 37548 31724 37604 31780
rect 37100 31554 37156 31556
rect 37100 31502 37102 31554
rect 37102 31502 37154 31554
rect 37154 31502 37156 31554
rect 37100 31500 37156 31502
rect 37436 31554 37492 31556
rect 37436 31502 37438 31554
rect 37438 31502 37490 31554
rect 37490 31502 37492 31554
rect 37436 31500 37492 31502
rect 38556 33292 38612 33348
rect 38892 34690 38948 34692
rect 38892 34638 38894 34690
rect 38894 34638 38946 34690
rect 38946 34638 38948 34690
rect 38892 34636 38948 34638
rect 39900 44268 39956 44324
rect 39788 43820 39844 43876
rect 40684 45388 40740 45444
rect 40348 43820 40404 43876
rect 40460 43708 40516 43764
rect 40124 43596 40180 43652
rect 40012 43314 40068 43316
rect 40012 43262 40014 43314
rect 40014 43262 40066 43314
rect 40066 43262 40068 43314
rect 40012 43260 40068 43262
rect 39788 42978 39844 42980
rect 39788 42926 39790 42978
rect 39790 42926 39842 42978
rect 39842 42926 39844 42978
rect 39788 42924 39844 42926
rect 39452 41580 39508 41636
rect 39900 42642 39956 42644
rect 39900 42590 39902 42642
rect 39902 42590 39954 42642
rect 39954 42590 39956 42642
rect 39900 42588 39956 42590
rect 39900 41858 39956 41860
rect 39900 41806 39902 41858
rect 39902 41806 39954 41858
rect 39954 41806 39956 41858
rect 39900 41804 39956 41806
rect 40236 43036 40292 43092
rect 40236 42476 40292 42532
rect 40124 41804 40180 41860
rect 40348 41692 40404 41748
rect 40012 41580 40068 41636
rect 40236 41298 40292 41300
rect 40236 41246 40238 41298
rect 40238 41246 40290 41298
rect 40290 41246 40292 41298
rect 40236 41244 40292 41246
rect 39676 40908 39732 40964
rect 41020 45106 41076 45108
rect 41020 45054 41022 45106
rect 41022 45054 41074 45106
rect 41074 45054 41076 45106
rect 41020 45052 41076 45054
rect 40908 44882 40964 44884
rect 40908 44830 40910 44882
rect 40910 44830 40962 44882
rect 40962 44830 40964 44882
rect 40908 44828 40964 44830
rect 41692 45778 41748 45780
rect 41692 45726 41694 45778
rect 41694 45726 41746 45778
rect 41746 45726 41748 45778
rect 41692 45724 41748 45726
rect 45276 47068 45332 47124
rect 43260 45948 43316 46004
rect 43820 45890 43876 45892
rect 43820 45838 43822 45890
rect 43822 45838 43874 45890
rect 43874 45838 43876 45890
rect 43820 45836 43876 45838
rect 46620 45724 46676 45780
rect 41692 44994 41748 44996
rect 41692 44942 41694 44994
rect 41694 44942 41746 44994
rect 41746 44942 41748 44994
rect 41692 44940 41748 44942
rect 41580 44492 41636 44548
rect 41020 44322 41076 44324
rect 41020 44270 41022 44322
rect 41022 44270 41074 44322
rect 41074 44270 41076 44322
rect 41020 44268 41076 44270
rect 41468 44268 41524 44324
rect 40908 43260 40964 43316
rect 40572 43036 40628 43092
rect 40572 42754 40628 42756
rect 40572 42702 40574 42754
rect 40574 42702 40626 42754
rect 40626 42702 40628 42754
rect 40572 42700 40628 42702
rect 41356 42700 41412 42756
rect 40684 42476 40740 42532
rect 42028 43820 42084 43876
rect 40572 41804 40628 41860
rect 41020 41692 41076 41748
rect 40908 41580 40964 41636
rect 40908 41244 40964 41300
rect 40572 40908 40628 40964
rect 40348 40572 40404 40628
rect 39900 40460 39956 40516
rect 39788 39452 39844 39508
rect 39788 38780 39844 38836
rect 39788 38444 39844 38500
rect 40684 40460 40740 40516
rect 40460 38780 40516 38836
rect 41692 41746 41748 41748
rect 41692 41694 41694 41746
rect 41694 41694 41746 41746
rect 41746 41694 41748 41746
rect 41692 41692 41748 41694
rect 41468 40460 41524 40516
rect 43596 45666 43652 45668
rect 43596 45614 43598 45666
rect 43598 45614 43650 45666
rect 43650 45614 43652 45666
rect 43596 45612 43652 45614
rect 42924 44940 42980 44996
rect 43708 44940 43764 44996
rect 42476 43650 42532 43652
rect 42476 43598 42478 43650
rect 42478 43598 42530 43650
rect 42530 43598 42532 43650
rect 42476 43596 42532 43598
rect 42588 43372 42644 43428
rect 42252 42924 42308 42980
rect 42140 42642 42196 42644
rect 42140 42590 42142 42642
rect 42142 42590 42194 42642
rect 42194 42590 42196 42642
rect 42140 42588 42196 42590
rect 43372 43426 43428 43428
rect 43372 43374 43374 43426
rect 43374 43374 43426 43426
rect 43426 43374 43428 43426
rect 43372 43372 43428 43374
rect 42364 41746 42420 41748
rect 42364 41694 42366 41746
rect 42366 41694 42418 41746
rect 42418 41694 42420 41746
rect 42364 41692 42420 41694
rect 41916 40402 41972 40404
rect 41916 40350 41918 40402
rect 41918 40350 41970 40402
rect 41970 40350 41972 40402
rect 41916 40348 41972 40350
rect 43484 41804 43540 41860
rect 42588 40402 42644 40404
rect 42588 40350 42590 40402
rect 42590 40350 42642 40402
rect 42642 40350 42644 40402
rect 42588 40348 42644 40350
rect 43036 40348 43092 40404
rect 40124 38444 40180 38500
rect 40236 38332 40292 38388
rect 40124 38050 40180 38052
rect 40124 37998 40126 38050
rect 40126 37998 40178 38050
rect 40178 37998 40180 38050
rect 40124 37996 40180 37998
rect 40348 37996 40404 38052
rect 40124 37436 40180 37492
rect 41020 37490 41076 37492
rect 41020 37438 41022 37490
rect 41022 37438 41074 37490
rect 41074 37438 41076 37490
rect 41020 37436 41076 37438
rect 40012 37154 40068 37156
rect 40012 37102 40014 37154
rect 40014 37102 40066 37154
rect 40066 37102 40068 37154
rect 40012 37100 40068 37102
rect 40908 37154 40964 37156
rect 40908 37102 40910 37154
rect 40910 37102 40962 37154
rect 40962 37102 40964 37154
rect 40908 37100 40964 37102
rect 40348 36988 40404 37044
rect 39900 36428 39956 36484
rect 39788 36370 39844 36372
rect 39788 36318 39790 36370
rect 39790 36318 39842 36370
rect 39842 36318 39844 36370
rect 39788 36316 39844 36318
rect 40012 35868 40068 35924
rect 39900 35420 39956 35476
rect 42476 39506 42532 39508
rect 42476 39454 42478 39506
rect 42478 39454 42530 39506
rect 42530 39454 42532 39506
rect 42476 39452 42532 39454
rect 42364 39394 42420 39396
rect 42364 39342 42366 39394
rect 42366 39342 42418 39394
rect 42418 39342 42420 39394
rect 42364 39340 42420 39342
rect 42140 39004 42196 39060
rect 41916 38556 41972 38612
rect 41580 38332 41636 38388
rect 41580 37212 41636 37268
rect 41132 36428 41188 36484
rect 40572 35420 40628 35476
rect 39788 34914 39844 34916
rect 39788 34862 39790 34914
rect 39790 34862 39842 34914
rect 39842 34862 39844 34914
rect 39788 34860 39844 34862
rect 39228 34524 39284 34580
rect 39004 34300 39060 34356
rect 38780 33516 38836 33572
rect 39788 33964 39844 34020
rect 38780 33346 38836 33348
rect 38780 33294 38782 33346
rect 38782 33294 38834 33346
rect 38834 33294 38836 33346
rect 38780 33292 38836 33294
rect 38668 31948 38724 32004
rect 40012 34242 40068 34244
rect 40012 34190 40014 34242
rect 40014 34190 40066 34242
rect 40066 34190 40068 34242
rect 40012 34188 40068 34190
rect 38780 33068 38836 33124
rect 39116 33292 39172 33348
rect 39228 33068 39284 33124
rect 37772 31388 37828 31444
rect 38668 31388 38724 31444
rect 39900 33234 39956 33236
rect 39900 33182 39902 33234
rect 39902 33182 39954 33234
rect 39954 33182 39956 33234
rect 39900 33180 39956 33182
rect 39676 32562 39732 32564
rect 39676 32510 39678 32562
rect 39678 32510 39730 32562
rect 39730 32510 39732 32562
rect 39676 32508 39732 32510
rect 40908 34242 40964 34244
rect 40908 34190 40910 34242
rect 40910 34190 40962 34242
rect 40962 34190 40964 34242
rect 40908 34188 40964 34190
rect 41020 33964 41076 34020
rect 41244 35644 41300 35700
rect 41132 34860 41188 34916
rect 41244 35420 41300 35476
rect 42700 38892 42756 38948
rect 41916 38050 41972 38052
rect 41916 37998 41918 38050
rect 41918 37998 41970 38050
rect 41970 37998 41972 38050
rect 41916 37996 41972 37998
rect 41804 36988 41860 37044
rect 41692 35922 41748 35924
rect 41692 35870 41694 35922
rect 41694 35870 41746 35922
rect 41746 35870 41748 35922
rect 41692 35868 41748 35870
rect 42476 35698 42532 35700
rect 42476 35646 42478 35698
rect 42478 35646 42530 35698
rect 42530 35646 42532 35698
rect 42476 35644 42532 35646
rect 42700 35532 42756 35588
rect 42812 35420 42868 35476
rect 43820 44492 43876 44548
rect 44828 44322 44884 44324
rect 44828 44270 44830 44322
rect 44830 44270 44882 44322
rect 44882 44270 44884 44322
rect 44828 44268 44884 44270
rect 44828 43650 44884 43652
rect 44828 43598 44830 43650
rect 44830 43598 44882 43650
rect 44882 43598 44884 43650
rect 44828 43596 44884 43598
rect 45724 43484 45780 43540
rect 44940 42642 44996 42644
rect 44940 42590 44942 42642
rect 44942 42590 44994 42642
rect 44994 42590 44996 42642
rect 44940 42588 44996 42590
rect 44268 41186 44324 41188
rect 44268 41134 44270 41186
rect 44270 41134 44322 41186
rect 44322 41134 44324 41186
rect 44268 41132 44324 41134
rect 44604 40402 44660 40404
rect 44604 40350 44606 40402
rect 44606 40350 44658 40402
rect 44658 40350 44660 40402
rect 44604 40348 44660 40350
rect 43484 39340 43540 39396
rect 43148 39058 43204 39060
rect 43148 39006 43150 39058
rect 43150 39006 43202 39058
rect 43202 39006 43204 39058
rect 43148 39004 43204 39006
rect 43036 38556 43092 38612
rect 43148 38332 43204 38388
rect 43148 38162 43204 38164
rect 43148 38110 43150 38162
rect 43150 38110 43202 38162
rect 43202 38110 43204 38162
rect 43148 38108 43204 38110
rect 43036 37378 43092 37380
rect 43036 37326 43038 37378
rect 43038 37326 43090 37378
rect 43090 37326 43092 37378
rect 43036 37324 43092 37326
rect 43820 39116 43876 39172
rect 43708 38834 43764 38836
rect 43708 38782 43710 38834
rect 43710 38782 43762 38834
rect 43762 38782 43764 38834
rect 43708 38780 43764 38782
rect 44156 38220 44212 38276
rect 43932 38108 43988 38164
rect 43708 37324 43764 37380
rect 43820 37772 43876 37828
rect 44156 37884 44212 37940
rect 44380 39394 44436 39396
rect 44380 39342 44382 39394
rect 44382 39342 44434 39394
rect 44434 39342 44436 39394
rect 44380 39340 44436 39342
rect 45612 43036 45668 43092
rect 45724 42754 45780 42756
rect 45724 42702 45726 42754
rect 45726 42702 45778 42754
rect 45778 42702 45780 42754
rect 45724 42700 45780 42702
rect 45612 42588 45668 42644
rect 45500 42028 45556 42084
rect 46508 45500 46564 45556
rect 46508 43596 46564 43652
rect 46396 42754 46452 42756
rect 46396 42702 46398 42754
rect 46398 42702 46450 42754
rect 46450 42702 46452 42754
rect 46396 42700 46452 42702
rect 46284 42476 46340 42532
rect 45948 40796 46004 40852
rect 44940 39842 44996 39844
rect 44940 39790 44942 39842
rect 44942 39790 44994 39842
rect 44994 39790 44996 39842
rect 44940 39788 44996 39790
rect 45276 39004 45332 39060
rect 44940 38892 44996 38948
rect 44268 36652 44324 36708
rect 43260 35308 43316 35364
rect 43596 35532 43652 35588
rect 44940 37996 44996 38052
rect 45164 37884 45220 37940
rect 45052 37826 45108 37828
rect 45052 37774 45054 37826
rect 45054 37774 45106 37826
rect 45106 37774 45108 37826
rect 45052 37772 45108 37774
rect 45724 40124 45780 40180
rect 45836 39058 45892 39060
rect 45836 39006 45838 39058
rect 45838 39006 45890 39058
rect 45890 39006 45892 39058
rect 45836 39004 45892 39006
rect 45724 38834 45780 38836
rect 45724 38782 45726 38834
rect 45726 38782 45778 38834
rect 45778 38782 45780 38834
rect 45724 38780 45780 38782
rect 45948 38834 46004 38836
rect 45948 38782 45950 38834
rect 45950 38782 46002 38834
rect 46002 38782 46004 38834
rect 45948 38780 46004 38782
rect 45612 38332 45668 38388
rect 45724 38050 45780 38052
rect 45724 37998 45726 38050
rect 45726 37998 45778 38050
rect 45778 37998 45780 38050
rect 45724 37996 45780 37998
rect 45836 37938 45892 37940
rect 45836 37886 45838 37938
rect 45838 37886 45890 37938
rect 45890 37886 45892 37938
rect 45836 37884 45892 37886
rect 45500 37436 45556 37492
rect 44828 36258 44884 36260
rect 44828 36206 44830 36258
rect 44830 36206 44882 36258
rect 44882 36206 44884 36258
rect 44828 36204 44884 36206
rect 44828 35308 44884 35364
rect 44940 35532 44996 35588
rect 43596 34802 43652 34804
rect 43596 34750 43598 34802
rect 43598 34750 43650 34802
rect 43650 34750 43652 34802
rect 43596 34748 43652 34750
rect 43148 34636 43204 34692
rect 42476 34300 42532 34356
rect 42140 34130 42196 34132
rect 42140 34078 42142 34130
rect 42142 34078 42194 34130
rect 42194 34078 42196 34130
rect 42140 34076 42196 34078
rect 41580 33628 41636 33684
rect 40348 32956 40404 33012
rect 41580 33346 41636 33348
rect 41580 33294 41582 33346
rect 41582 33294 41634 33346
rect 41634 33294 41636 33346
rect 41580 33292 41636 33294
rect 41692 33068 41748 33124
rect 43708 34636 43764 34692
rect 39564 31778 39620 31780
rect 39564 31726 39566 31778
rect 39566 31726 39618 31778
rect 39618 31726 39620 31778
rect 39564 31724 39620 31726
rect 36764 30828 36820 30884
rect 36092 30716 36148 30772
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35532 23154 35588 23156
rect 35532 23102 35534 23154
rect 35534 23102 35586 23154
rect 35586 23102 35588 23154
rect 35532 23100 35588 23102
rect 35420 22988 35476 23044
rect 35532 22876 35588 22932
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 34188 21698 34244 21700
rect 34188 21646 34190 21698
rect 34190 21646 34242 21698
rect 34242 21646 34244 21698
rect 34188 21644 34244 21646
rect 34636 21698 34692 21700
rect 34636 21646 34638 21698
rect 34638 21646 34690 21698
rect 34690 21646 34692 21698
rect 34636 21644 34692 21646
rect 34412 21586 34468 21588
rect 34412 21534 34414 21586
rect 34414 21534 34466 21586
rect 34466 21534 34468 21586
rect 34412 21532 34468 21534
rect 35644 22092 35700 22148
rect 34972 21196 35028 21252
rect 33180 20076 33236 20132
rect 32396 19906 32452 19908
rect 32396 19854 32398 19906
rect 32398 19854 32450 19906
rect 32450 19854 32452 19906
rect 32396 19852 32452 19854
rect 32284 19740 32340 19796
rect 32844 19740 32900 19796
rect 32732 17442 32788 17444
rect 32732 17390 32734 17442
rect 32734 17390 32786 17442
rect 32786 17390 32788 17442
rect 32732 17388 32788 17390
rect 32284 17052 32340 17108
rect 33180 19180 33236 19236
rect 33180 18172 33236 18228
rect 33180 17388 33236 17444
rect 32956 14476 33012 14532
rect 33292 16716 33348 16772
rect 33180 13746 33236 13748
rect 33180 13694 33182 13746
rect 33182 13694 33234 13746
rect 33234 13694 33236 13746
rect 33180 13692 33236 13694
rect 32396 13634 32452 13636
rect 32396 13582 32398 13634
rect 32398 13582 32450 13634
rect 32450 13582 32452 13634
rect 32396 13580 32452 13582
rect 33516 19906 33572 19908
rect 33516 19854 33518 19906
rect 33518 19854 33570 19906
rect 33570 19854 33572 19906
rect 33516 19852 33572 19854
rect 33516 19180 33572 19236
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 38108 29596 38164 29652
rect 37324 29372 37380 29428
rect 36428 29260 36484 29316
rect 37884 29314 37940 29316
rect 37884 29262 37886 29314
rect 37886 29262 37938 29314
rect 37938 29262 37940 29314
rect 37884 29260 37940 29262
rect 36428 28642 36484 28644
rect 36428 28590 36430 28642
rect 36430 28590 36482 28642
rect 36482 28590 36484 28642
rect 36428 28588 36484 28590
rect 36988 28476 37044 28532
rect 36988 27858 37044 27860
rect 36988 27806 36990 27858
rect 36990 27806 37042 27858
rect 37042 27806 37044 27858
rect 36988 27804 37044 27806
rect 36540 27020 36596 27076
rect 37772 28252 37828 28308
rect 41916 31836 41972 31892
rect 39900 31612 39956 31668
rect 40236 31666 40292 31668
rect 40236 31614 40238 31666
rect 40238 31614 40290 31666
rect 40290 31614 40292 31666
rect 40236 31612 40292 31614
rect 41916 31612 41972 31668
rect 41356 31500 41412 31556
rect 39900 29596 39956 29652
rect 39116 29260 39172 29316
rect 38668 28530 38724 28532
rect 38668 28478 38670 28530
rect 38670 28478 38722 28530
rect 38722 28478 38724 28530
rect 38668 28476 38724 28478
rect 38332 28252 38388 28308
rect 40908 30380 40964 30436
rect 41692 30940 41748 30996
rect 41244 30882 41300 30884
rect 41244 30830 41246 30882
rect 41246 30830 41298 30882
rect 41298 30830 41300 30882
rect 41244 30828 41300 30830
rect 41132 30716 41188 30772
rect 40012 29372 40068 29428
rect 39788 28700 39844 28756
rect 40012 29148 40068 29204
rect 39676 28476 39732 28532
rect 38668 27804 38724 27860
rect 38556 26908 38612 26964
rect 36204 25116 36260 25172
rect 36428 25506 36484 25508
rect 36428 25454 36430 25506
rect 36430 25454 36482 25506
rect 36482 25454 36484 25506
rect 36428 25452 36484 25454
rect 35980 24610 36036 24612
rect 35980 24558 35982 24610
rect 35982 24558 36034 24610
rect 36034 24558 36036 24610
rect 35980 24556 36036 24558
rect 36428 23772 36484 23828
rect 36316 23212 36372 23268
rect 36988 25340 37044 25396
rect 37324 25506 37380 25508
rect 37324 25454 37326 25506
rect 37326 25454 37378 25506
rect 37378 25454 37380 25506
rect 37324 25452 37380 25454
rect 37212 25116 37268 25172
rect 36876 23324 36932 23380
rect 36092 23042 36148 23044
rect 36092 22990 36094 23042
rect 36094 22990 36146 23042
rect 36146 22990 36148 23042
rect 36092 22988 36148 22990
rect 35980 22876 36036 22932
rect 35980 22316 36036 22372
rect 36092 21868 36148 21924
rect 36876 22988 36932 23044
rect 37100 23042 37156 23044
rect 37100 22990 37102 23042
rect 37102 22990 37154 23042
rect 37154 22990 37156 23042
rect 37100 22988 37156 22990
rect 37324 25004 37380 25060
rect 37324 23436 37380 23492
rect 37548 26684 37604 26740
rect 37548 26236 37604 26292
rect 37436 23324 37492 23380
rect 37660 25452 37716 25508
rect 36876 21474 36932 21476
rect 36876 21422 36878 21474
rect 36878 21422 36930 21474
rect 36930 21422 36932 21474
rect 36876 21420 36932 21422
rect 35980 21308 36036 21364
rect 34188 20188 34244 20244
rect 34524 20300 34580 20356
rect 33852 20130 33908 20132
rect 33852 20078 33854 20130
rect 33854 20078 33906 20130
rect 33906 20078 33908 20130
rect 33852 20076 33908 20078
rect 33628 19068 33684 19124
rect 33740 19964 33796 20020
rect 34300 20018 34356 20020
rect 34300 19966 34302 20018
rect 34302 19966 34354 20018
rect 34354 19966 34356 20018
rect 34300 19964 34356 19966
rect 33516 16492 33572 16548
rect 33628 16828 33684 16884
rect 33404 15372 33460 15428
rect 33516 15260 33572 15316
rect 34300 18508 34356 18564
rect 33852 18172 33908 18228
rect 33964 17612 34020 17668
rect 34188 17836 34244 17892
rect 33964 17442 34020 17444
rect 33964 17390 33966 17442
rect 33966 17390 34018 17442
rect 34018 17390 34020 17442
rect 33964 17388 34020 17390
rect 34188 15596 34244 15652
rect 34748 20076 34804 20132
rect 35084 20188 35140 20244
rect 34636 18396 34692 18452
rect 34524 17778 34580 17780
rect 34524 17726 34526 17778
rect 34526 17726 34578 17778
rect 34578 17726 34580 17778
rect 34524 17724 34580 17726
rect 35532 20300 35588 20356
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 36540 20188 36596 20244
rect 34972 18508 35028 18564
rect 35084 18620 35140 18676
rect 34860 18450 34916 18452
rect 34860 18398 34862 18450
rect 34862 18398 34914 18450
rect 34914 18398 34916 18450
rect 34860 18396 34916 18398
rect 35420 19234 35476 19236
rect 35420 19182 35422 19234
rect 35422 19182 35474 19234
rect 35474 19182 35476 19234
rect 35420 19180 35476 19182
rect 35532 19122 35588 19124
rect 35532 19070 35534 19122
rect 35534 19070 35586 19122
rect 35586 19070 35588 19122
rect 35532 19068 35588 19070
rect 35756 19122 35812 19124
rect 35756 19070 35758 19122
rect 35758 19070 35810 19122
rect 35810 19070 35812 19122
rect 35756 19068 35812 19070
rect 35420 18562 35476 18564
rect 35420 18510 35422 18562
rect 35422 18510 35474 18562
rect 35474 18510 35476 18562
rect 35420 18508 35476 18510
rect 35868 18562 35924 18564
rect 35868 18510 35870 18562
rect 35870 18510 35922 18562
rect 35922 18510 35924 18562
rect 35868 18508 35924 18510
rect 36092 19906 36148 19908
rect 36092 19854 36094 19906
rect 36094 19854 36146 19906
rect 36146 19854 36148 19906
rect 36092 19852 36148 19854
rect 36092 19180 36148 19236
rect 36316 18284 36372 18340
rect 37212 21474 37268 21476
rect 37212 21422 37214 21474
rect 37214 21422 37266 21474
rect 37266 21422 37268 21474
rect 37212 21420 37268 21422
rect 37212 20188 37268 20244
rect 34524 17500 34580 17556
rect 34860 17276 34916 17332
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35644 17724 35700 17780
rect 35420 17500 35476 17556
rect 35084 16828 35140 16884
rect 35644 16828 35700 16884
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 34524 15820 34580 15876
rect 34748 15148 34804 15204
rect 33740 14588 33796 14644
rect 33628 12684 33684 12740
rect 35420 15708 35476 15764
rect 35756 15484 35812 15540
rect 34748 14642 34804 14644
rect 34748 14590 34750 14642
rect 34750 14590 34802 14642
rect 34802 14590 34804 14642
rect 34748 14588 34804 14590
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35308 14588 35364 14644
rect 34412 13244 34468 13300
rect 34188 12796 34244 12852
rect 33964 12684 34020 12740
rect 33292 11788 33348 11844
rect 34524 12738 34580 12740
rect 34524 12686 34526 12738
rect 34526 12686 34578 12738
rect 34578 12686 34580 12738
rect 34524 12684 34580 12686
rect 34412 12572 34468 12628
rect 34300 12460 34356 12516
rect 34188 12236 34244 12292
rect 33852 11452 33908 11508
rect 33404 11004 33460 11060
rect 32284 10780 32340 10836
rect 32620 10780 32676 10836
rect 33628 10834 33684 10836
rect 33628 10782 33630 10834
rect 33630 10782 33682 10834
rect 33682 10782 33684 10834
rect 33628 10780 33684 10782
rect 33964 11340 34020 11396
rect 32396 10386 32452 10388
rect 32396 10334 32398 10386
rect 32398 10334 32450 10386
rect 32450 10334 32452 10386
rect 32396 10332 32452 10334
rect 32284 10108 32340 10164
rect 32508 9266 32564 9268
rect 32508 9214 32510 9266
rect 32510 9214 32562 9266
rect 32562 9214 32564 9266
rect 32508 9212 32564 9214
rect 33516 9212 33572 9268
rect 32172 8988 32228 9044
rect 33292 9042 33348 9044
rect 33292 8990 33294 9042
rect 33294 8990 33346 9042
rect 33346 8990 33348 9042
rect 33292 8988 33348 8990
rect 32508 7980 32564 8036
rect 32732 7868 32788 7924
rect 31948 7474 32004 7476
rect 31948 7422 31950 7474
rect 31950 7422 32002 7474
rect 32002 7422 32004 7474
rect 31948 7420 32004 7422
rect 32508 6748 32564 6804
rect 32172 6690 32228 6692
rect 32172 6638 32174 6690
rect 32174 6638 32226 6690
rect 32226 6638 32228 6690
rect 32172 6636 32228 6638
rect 31612 6300 31668 6356
rect 34412 11004 34468 11060
rect 33628 7868 33684 7924
rect 33628 7532 33684 7588
rect 32956 6860 33012 6916
rect 33292 6690 33348 6692
rect 33292 6638 33294 6690
rect 33294 6638 33346 6690
rect 33346 6638 33348 6690
rect 33292 6636 33348 6638
rect 32732 6300 32788 6356
rect 33404 5964 33460 6020
rect 33180 5794 33236 5796
rect 33180 5742 33182 5794
rect 33182 5742 33234 5794
rect 33234 5742 33236 5794
rect 33180 5740 33236 5742
rect 32956 4844 33012 4900
rect 32284 4284 32340 4340
rect 31836 3612 31892 3668
rect 31500 3388 31556 3444
rect 32172 3500 32228 3556
rect 33292 4562 33348 4564
rect 33292 4510 33294 4562
rect 33294 4510 33346 4562
rect 33346 4510 33348 4562
rect 33292 4508 33348 4510
rect 33740 6860 33796 6916
rect 34076 8930 34132 8932
rect 34076 8878 34078 8930
rect 34078 8878 34130 8930
rect 34130 8878 34132 8930
rect 34076 8876 34132 8878
rect 33852 5964 33908 6020
rect 34300 10498 34356 10500
rect 34300 10446 34302 10498
rect 34302 10446 34354 10498
rect 34354 10446 34356 10498
rect 34300 10444 34356 10446
rect 34748 11452 34804 11508
rect 34972 13244 35028 13300
rect 34972 12850 35028 12852
rect 34972 12798 34974 12850
rect 34974 12798 35026 12850
rect 35026 12798 35028 12850
rect 34972 12796 35028 12798
rect 36428 17276 36484 17332
rect 36428 16044 36484 16100
rect 36540 16828 36596 16884
rect 36092 15426 36148 15428
rect 36092 15374 36094 15426
rect 36094 15374 36146 15426
rect 36146 15374 36148 15426
rect 36092 15372 36148 15374
rect 36428 15260 36484 15316
rect 35756 14588 35812 14644
rect 35868 14530 35924 14532
rect 35868 14478 35870 14530
rect 35870 14478 35922 14530
rect 35922 14478 35924 14530
rect 35868 14476 35924 14478
rect 35980 14418 36036 14420
rect 35980 14366 35982 14418
rect 35982 14366 36034 14418
rect 36034 14366 36036 14418
rect 35980 14364 36036 14366
rect 36092 14306 36148 14308
rect 36092 14254 36094 14306
rect 36094 14254 36146 14306
rect 36146 14254 36148 14306
rect 36092 14252 36148 14254
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 37212 19906 37268 19908
rect 37212 19854 37214 19906
rect 37214 19854 37266 19906
rect 37266 19854 37268 19906
rect 37212 19852 37268 19854
rect 37100 18450 37156 18452
rect 37100 18398 37102 18450
rect 37102 18398 37154 18450
rect 37154 18398 37156 18450
rect 37100 18396 37156 18398
rect 36764 16156 36820 16212
rect 36652 14028 36708 14084
rect 36876 16044 36932 16100
rect 36540 13132 36596 13188
rect 35084 12572 35140 12628
rect 36204 12796 36260 12852
rect 36204 12066 36260 12068
rect 36204 12014 36206 12066
rect 36206 12014 36258 12066
rect 36258 12014 36260 12066
rect 36204 12012 36260 12014
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 34636 9884 34692 9940
rect 34972 11452 35028 11508
rect 34412 9602 34468 9604
rect 34412 9550 34414 9602
rect 34414 9550 34466 9602
rect 34466 9550 34468 9602
rect 34412 9548 34468 9550
rect 34860 10444 34916 10500
rect 35196 11116 35252 11172
rect 35532 11004 35588 11060
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35756 10556 35812 10612
rect 34972 9826 35028 9828
rect 34972 9774 34974 9826
rect 34974 9774 35026 9826
rect 35026 9774 35028 9826
rect 34972 9772 35028 9774
rect 35420 9660 35476 9716
rect 35196 9602 35252 9604
rect 35196 9550 35198 9602
rect 35198 9550 35250 9602
rect 35250 9550 35252 9602
rect 35196 9548 35252 9550
rect 35196 9212 35252 9268
rect 35308 9154 35364 9156
rect 35308 9102 35310 9154
rect 35310 9102 35362 9154
rect 35362 9102 35364 9154
rect 35308 9100 35364 9102
rect 35980 9884 36036 9940
rect 36204 9826 36260 9828
rect 36204 9774 36206 9826
rect 36206 9774 36258 9826
rect 36258 9774 36260 9826
rect 36204 9772 36260 9774
rect 35756 9660 35812 9716
rect 35868 9548 35924 9604
rect 34300 8370 34356 8372
rect 34300 8318 34302 8370
rect 34302 8318 34354 8370
rect 34354 8318 34356 8370
rect 34300 8316 34356 8318
rect 34188 6860 34244 6916
rect 34188 6636 34244 6692
rect 34972 8876 35028 8932
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 34972 8034 35028 8036
rect 34972 7982 34974 8034
rect 34974 7982 35026 8034
rect 35026 7982 35028 8034
rect 34972 7980 35028 7982
rect 34860 7868 34916 7924
rect 34748 7532 34804 7588
rect 34636 6524 34692 6580
rect 34524 6412 34580 6468
rect 33516 5180 33572 5236
rect 33852 5794 33908 5796
rect 33852 5742 33854 5794
rect 33854 5742 33906 5794
rect 33906 5742 33908 5794
rect 33852 5740 33908 5742
rect 33628 5068 33684 5124
rect 34972 6018 35028 6020
rect 34972 5966 34974 6018
rect 34974 5966 35026 6018
rect 35026 5966 35028 6018
rect 34972 5964 35028 5966
rect 34188 5906 34244 5908
rect 34188 5854 34190 5906
rect 34190 5854 34242 5906
rect 34242 5854 34244 5906
rect 34188 5852 34244 5854
rect 34860 5906 34916 5908
rect 34860 5854 34862 5906
rect 34862 5854 34914 5906
rect 34914 5854 34916 5906
rect 34860 5852 34916 5854
rect 34748 5234 34804 5236
rect 34748 5182 34750 5234
rect 34750 5182 34802 5234
rect 34802 5182 34804 5234
rect 34748 5180 34804 5182
rect 34636 5122 34692 5124
rect 34636 5070 34638 5122
rect 34638 5070 34690 5122
rect 34690 5070 34692 5122
rect 34636 5068 34692 5070
rect 35196 8316 35252 8372
rect 35644 8370 35700 8372
rect 35644 8318 35646 8370
rect 35646 8318 35698 8370
rect 35698 8318 35700 8370
rect 35644 8316 35700 8318
rect 35756 7644 35812 7700
rect 35532 7420 35588 7476
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35532 6636 35588 6692
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35420 5292 35476 5348
rect 35308 5180 35364 5236
rect 33964 4732 34020 4788
rect 34076 4956 34132 5012
rect 34860 4508 34916 4564
rect 35756 5180 35812 5236
rect 35868 6412 35924 6468
rect 35644 5122 35700 5124
rect 35644 5070 35646 5122
rect 35646 5070 35698 5122
rect 35698 5070 35700 5122
rect 35644 5068 35700 5070
rect 35532 4956 35588 5012
rect 37548 21980 37604 22036
rect 37436 21756 37492 21812
rect 37436 17052 37492 17108
rect 37100 15596 37156 15652
rect 36876 12796 36932 12852
rect 37212 15372 37268 15428
rect 37212 14530 37268 14532
rect 37212 14478 37214 14530
rect 37214 14478 37266 14530
rect 37266 14478 37268 14530
rect 37212 14476 37268 14478
rect 37324 14418 37380 14420
rect 37324 14366 37326 14418
rect 37326 14366 37378 14418
rect 37378 14366 37380 14418
rect 37324 14364 37380 14366
rect 37436 14252 37492 14308
rect 37436 13580 37492 13636
rect 37100 13468 37156 13524
rect 37324 13132 37380 13188
rect 37100 12124 37156 12180
rect 36428 10780 36484 10836
rect 36988 12012 37044 12068
rect 37100 11452 37156 11508
rect 36652 11116 36708 11172
rect 36652 10668 36708 10724
rect 36428 9826 36484 9828
rect 36428 9774 36430 9826
rect 36430 9774 36482 9826
rect 36482 9774 36484 9826
rect 36428 9772 36484 9774
rect 36092 9212 36148 9268
rect 36204 9100 36260 9156
rect 36540 8428 36596 8484
rect 37100 10610 37156 10612
rect 37100 10558 37102 10610
rect 37102 10558 37154 10610
rect 37154 10558 37156 10610
rect 37100 10556 37156 10558
rect 39340 27074 39396 27076
rect 39340 27022 39342 27074
rect 39342 27022 39394 27074
rect 39394 27022 39396 27074
rect 39340 27020 39396 27022
rect 40236 29314 40292 29316
rect 40236 29262 40238 29314
rect 40238 29262 40290 29314
rect 40290 29262 40292 29314
rect 40236 29260 40292 29262
rect 40348 28364 40404 28420
rect 41244 29538 41300 29540
rect 41244 29486 41246 29538
rect 41246 29486 41298 29538
rect 41298 29486 41300 29538
rect 41244 29484 41300 29486
rect 41244 28364 41300 28420
rect 39228 26908 39284 26964
rect 40348 27074 40404 27076
rect 40348 27022 40350 27074
rect 40350 27022 40402 27074
rect 40402 27022 40404 27074
rect 40348 27020 40404 27022
rect 40124 26962 40180 26964
rect 40124 26910 40126 26962
rect 40126 26910 40178 26962
rect 40178 26910 40180 26962
rect 40124 26908 40180 26910
rect 41020 27804 41076 27860
rect 42476 31724 42532 31780
rect 42924 33628 42980 33684
rect 44044 34412 44100 34468
rect 43932 34076 43988 34132
rect 43708 33458 43764 33460
rect 43708 33406 43710 33458
rect 43710 33406 43762 33458
rect 43762 33406 43764 33458
rect 43708 33404 43764 33406
rect 43708 32508 43764 32564
rect 43036 31890 43092 31892
rect 43036 31838 43038 31890
rect 43038 31838 43090 31890
rect 43090 31838 43092 31890
rect 43036 31836 43092 31838
rect 42924 31612 42980 31668
rect 43260 31500 43316 31556
rect 43260 31052 43316 31108
rect 42364 30940 42420 30996
rect 42812 30994 42868 30996
rect 42812 30942 42814 30994
rect 42814 30942 42866 30994
rect 42866 30942 42868 30994
rect 42812 30940 42868 30942
rect 42028 30882 42084 30884
rect 42028 30830 42030 30882
rect 42030 30830 42082 30882
rect 42082 30830 42084 30882
rect 42028 30828 42084 30830
rect 42476 30716 42532 30772
rect 42812 30380 42868 30436
rect 43708 31836 43764 31892
rect 42364 30268 42420 30324
rect 41468 28082 41524 28084
rect 41468 28030 41470 28082
rect 41470 28030 41522 28082
rect 41522 28030 41524 28082
rect 41468 28028 41524 28030
rect 41804 30156 41860 30212
rect 42140 28082 42196 28084
rect 42140 28030 42142 28082
rect 42142 28030 42194 28082
rect 42194 28030 42196 28082
rect 42140 28028 42196 28030
rect 41356 27074 41412 27076
rect 41356 27022 41358 27074
rect 41358 27022 41410 27074
rect 41410 27022 41412 27074
rect 41356 27020 41412 27022
rect 39452 26460 39508 26516
rect 40124 26684 40180 26740
rect 38892 26236 38948 26292
rect 37996 25676 38052 25732
rect 38780 25730 38836 25732
rect 38780 25678 38782 25730
rect 38782 25678 38834 25730
rect 38834 25678 38836 25730
rect 38780 25676 38836 25678
rect 38108 25394 38164 25396
rect 38108 25342 38110 25394
rect 38110 25342 38162 25394
rect 38162 25342 38164 25394
rect 38108 25340 38164 25342
rect 38332 24668 38388 24724
rect 37884 24556 37940 24612
rect 37884 23938 37940 23940
rect 37884 23886 37886 23938
rect 37886 23886 37938 23938
rect 37938 23886 37940 23938
rect 37884 23884 37940 23886
rect 38444 23884 38500 23940
rect 38668 23660 38724 23716
rect 39340 26290 39396 26292
rect 39340 26238 39342 26290
rect 39342 26238 39394 26290
rect 39394 26238 39396 26290
rect 39340 26236 39396 26238
rect 39004 25394 39060 25396
rect 39004 25342 39006 25394
rect 39006 25342 39058 25394
rect 39058 25342 39060 25394
rect 39004 25340 39060 25342
rect 39676 25394 39732 25396
rect 39676 25342 39678 25394
rect 39678 25342 39730 25394
rect 39730 25342 39732 25394
rect 39676 25340 39732 25342
rect 39452 25228 39508 25284
rect 39228 23884 39284 23940
rect 39788 23884 39844 23940
rect 38444 23378 38500 23380
rect 38444 23326 38446 23378
rect 38446 23326 38498 23378
rect 38498 23326 38500 23378
rect 38444 23324 38500 23326
rect 37772 22988 37828 23044
rect 37884 22876 37940 22932
rect 38444 22652 38500 22708
rect 38780 23154 38836 23156
rect 38780 23102 38782 23154
rect 38782 23102 38834 23154
rect 38834 23102 38836 23154
rect 38780 23100 38836 23102
rect 38780 21810 38836 21812
rect 38780 21758 38782 21810
rect 38782 21758 38834 21810
rect 38834 21758 38836 21810
rect 38780 21756 38836 21758
rect 39452 23436 39508 23492
rect 39564 23714 39620 23716
rect 39564 23662 39566 23714
rect 39566 23662 39618 23714
rect 39618 23662 39620 23714
rect 39564 23660 39620 23662
rect 39564 23212 39620 23268
rect 39452 23100 39508 23156
rect 39340 19740 39396 19796
rect 39340 18508 39396 18564
rect 37772 18338 37828 18340
rect 37772 18286 37774 18338
rect 37774 18286 37826 18338
rect 37826 18286 37828 18338
rect 37772 18284 37828 18286
rect 37884 16882 37940 16884
rect 37884 16830 37886 16882
rect 37886 16830 37938 16882
rect 37938 16830 37940 16882
rect 37884 16828 37940 16830
rect 38668 17052 38724 17108
rect 38556 16828 38612 16884
rect 37772 16210 37828 16212
rect 37772 16158 37774 16210
rect 37774 16158 37826 16210
rect 37826 16158 37828 16210
rect 37772 16156 37828 16158
rect 38892 16156 38948 16212
rect 37772 15820 37828 15876
rect 37660 15148 37716 15204
rect 38332 15260 38388 15316
rect 39116 15820 39172 15876
rect 39564 15708 39620 15764
rect 39564 15202 39620 15204
rect 39564 15150 39566 15202
rect 39566 15150 39618 15202
rect 39618 15150 39620 15202
rect 39564 15148 39620 15150
rect 38220 14476 38276 14532
rect 39004 14530 39060 14532
rect 39004 14478 39006 14530
rect 39006 14478 39058 14530
rect 39058 14478 39060 14530
rect 39004 14476 39060 14478
rect 38780 14252 38836 14308
rect 38556 13804 38612 13860
rect 37324 12178 37380 12180
rect 37324 12126 37326 12178
rect 37326 12126 37378 12178
rect 37378 12126 37380 12178
rect 37324 12124 37380 12126
rect 37772 13580 37828 13636
rect 39004 13692 39060 13748
rect 38108 13186 38164 13188
rect 38108 13134 38110 13186
rect 38110 13134 38162 13186
rect 38162 13134 38164 13186
rect 38108 13132 38164 13134
rect 39228 13858 39284 13860
rect 39228 13806 39230 13858
rect 39230 13806 39282 13858
rect 39282 13806 39284 13858
rect 39228 13804 39284 13806
rect 39452 14252 39508 14308
rect 40012 24722 40068 24724
rect 40012 24670 40014 24722
rect 40014 24670 40066 24722
rect 40066 24670 40068 24722
rect 40012 24668 40068 24670
rect 39900 22482 39956 22484
rect 39900 22430 39902 22482
rect 39902 22430 39954 22482
rect 39954 22430 39956 22482
rect 39900 22428 39956 22430
rect 40236 23660 40292 23716
rect 40460 22428 40516 22484
rect 40012 20018 40068 20020
rect 40012 19966 40014 20018
rect 40014 19966 40066 20018
rect 40066 19966 40068 20018
rect 40012 19964 40068 19966
rect 40236 19906 40292 19908
rect 40236 19854 40238 19906
rect 40238 19854 40290 19906
rect 40290 19854 40292 19906
rect 40236 19852 40292 19854
rect 40348 19628 40404 19684
rect 40012 19068 40068 19124
rect 40796 26460 40852 26516
rect 40908 26402 40964 26404
rect 40908 26350 40910 26402
rect 40910 26350 40962 26402
rect 40962 26350 40964 26402
rect 40908 26348 40964 26350
rect 42140 27244 42196 27300
rect 42028 26572 42084 26628
rect 41580 26348 41636 26404
rect 41804 26460 41860 26516
rect 42028 26402 42084 26404
rect 42028 26350 42030 26402
rect 42030 26350 42082 26402
rect 42082 26350 42084 26402
rect 42028 26348 42084 26350
rect 41132 26012 41188 26068
rect 40684 25340 40740 25396
rect 42140 26290 42196 26292
rect 42140 26238 42142 26290
rect 42142 26238 42194 26290
rect 42194 26238 42196 26290
rect 42140 26236 42196 26238
rect 42252 25900 42308 25956
rect 42700 29538 42756 29540
rect 42700 29486 42702 29538
rect 42702 29486 42754 29538
rect 42754 29486 42756 29538
rect 42700 29484 42756 29486
rect 42476 28364 42532 28420
rect 43484 31724 43540 31780
rect 43708 31666 43764 31668
rect 43708 31614 43710 31666
rect 43710 31614 43762 31666
rect 43762 31614 43764 31666
rect 43708 31612 43764 31614
rect 43484 30268 43540 30324
rect 44268 34690 44324 34692
rect 44268 34638 44270 34690
rect 44270 34638 44322 34690
rect 44322 34638 44324 34690
rect 44268 34636 44324 34638
rect 44268 33516 44324 33572
rect 44156 32620 44212 32676
rect 45388 35644 45444 35700
rect 46172 38668 46228 38724
rect 46396 42028 46452 42084
rect 47404 45778 47460 45780
rect 47404 45726 47406 45778
rect 47406 45726 47458 45778
rect 47458 45726 47460 45778
rect 47404 45724 47460 45726
rect 47068 44044 47124 44100
rect 47628 45388 47684 45444
rect 48188 45388 48244 45444
rect 47628 44994 47684 44996
rect 47628 44942 47630 44994
rect 47630 44942 47682 44994
rect 47682 44942 47684 44994
rect 47628 44940 47684 44942
rect 46844 42924 46900 42980
rect 46956 43036 47012 43092
rect 46732 42700 46788 42756
rect 47516 42978 47572 42980
rect 47516 42926 47518 42978
rect 47518 42926 47570 42978
rect 47570 42926 47572 42978
rect 47516 42924 47572 42926
rect 47292 42140 47348 42196
rect 46956 42028 47012 42084
rect 48188 44098 48244 44100
rect 48188 44046 48190 44098
rect 48190 44046 48242 44098
rect 48242 44046 48244 44098
rect 48188 44044 48244 44046
rect 47740 43036 47796 43092
rect 47740 42754 47796 42756
rect 47740 42702 47742 42754
rect 47742 42702 47794 42754
rect 47794 42702 47796 42754
rect 47740 42700 47796 42702
rect 47852 42476 47908 42532
rect 47964 41132 48020 41188
rect 46508 40460 46564 40516
rect 47964 40514 48020 40516
rect 47964 40462 47966 40514
rect 47966 40462 48018 40514
rect 48018 40462 48020 40514
rect 47964 40460 48020 40462
rect 46396 39340 46452 39396
rect 46620 40124 46676 40180
rect 47068 39452 47124 39508
rect 46732 39228 46788 39284
rect 46844 39058 46900 39060
rect 46844 39006 46846 39058
rect 46846 39006 46898 39058
rect 46898 39006 46900 39058
rect 46844 39004 46900 39006
rect 46620 38946 46676 38948
rect 46620 38894 46622 38946
rect 46622 38894 46674 38946
rect 46674 38894 46676 38946
rect 46620 38892 46676 38894
rect 47068 38892 47124 38948
rect 46956 38834 47012 38836
rect 46956 38782 46958 38834
rect 46958 38782 47010 38834
rect 47010 38782 47012 38834
rect 46956 38780 47012 38782
rect 47740 39788 47796 39844
rect 48188 39116 48244 39172
rect 47740 38892 47796 38948
rect 47404 38834 47460 38836
rect 47404 38782 47406 38834
rect 47406 38782 47458 38834
rect 47458 38782 47460 38834
rect 47404 38780 47460 38782
rect 47292 38668 47348 38724
rect 47740 38444 47796 38500
rect 47404 38220 47460 38276
rect 46396 37884 46452 37940
rect 46284 37490 46340 37492
rect 46284 37438 46286 37490
rect 46286 37438 46338 37490
rect 46338 37438 46340 37490
rect 46284 37436 46340 37438
rect 46844 36204 46900 36260
rect 47068 37266 47124 37268
rect 47068 37214 47070 37266
rect 47070 37214 47122 37266
rect 47122 37214 47124 37266
rect 47068 37212 47124 37214
rect 47404 35810 47460 35812
rect 47404 35758 47406 35810
rect 47406 35758 47458 35810
rect 47458 35758 47460 35810
rect 47404 35756 47460 35758
rect 47628 37436 47684 37492
rect 47852 37266 47908 37268
rect 47852 37214 47854 37266
rect 47854 37214 47906 37266
rect 47906 37214 47908 37266
rect 47852 37212 47908 37214
rect 46172 35532 46228 35588
rect 45836 35474 45892 35476
rect 45836 35422 45838 35474
rect 45838 35422 45890 35474
rect 45890 35422 45892 35474
rect 45836 35420 45892 35422
rect 44380 33404 44436 33460
rect 44940 33516 44996 33572
rect 45500 33346 45556 33348
rect 45500 33294 45502 33346
rect 45502 33294 45554 33346
rect 45554 33294 45556 33346
rect 45500 33292 45556 33294
rect 45948 33292 46004 33348
rect 45388 33068 45444 33124
rect 44492 32786 44548 32788
rect 44492 32734 44494 32786
rect 44494 32734 44546 32786
rect 44546 32734 44548 32786
rect 44492 32732 44548 32734
rect 44940 32674 44996 32676
rect 44940 32622 44942 32674
rect 44942 32622 44994 32674
rect 44994 32622 44996 32674
rect 44940 32620 44996 32622
rect 45052 31948 45108 32004
rect 44044 31724 44100 31780
rect 44268 31724 44324 31780
rect 44156 31218 44212 31220
rect 44156 31166 44158 31218
rect 44158 31166 44210 31218
rect 44210 31166 44212 31218
rect 44156 31164 44212 31166
rect 44268 31106 44324 31108
rect 44268 31054 44270 31106
rect 44270 31054 44322 31106
rect 44322 31054 44324 31106
rect 44268 31052 44324 31054
rect 43932 30994 43988 30996
rect 43932 30942 43934 30994
rect 43934 30942 43986 30994
rect 43986 30942 43988 30994
rect 43932 30940 43988 30942
rect 45052 31778 45108 31780
rect 45052 31726 45054 31778
rect 45054 31726 45106 31778
rect 45106 31726 45108 31778
rect 45052 31724 45108 31726
rect 45164 31666 45220 31668
rect 45164 31614 45166 31666
rect 45166 31614 45218 31666
rect 45218 31614 45220 31666
rect 45164 31612 45220 31614
rect 45276 31052 45332 31108
rect 44828 30940 44884 30996
rect 43820 30156 43876 30212
rect 43372 29372 43428 29428
rect 43372 28642 43428 28644
rect 43372 28590 43374 28642
rect 43374 28590 43426 28642
rect 43426 28590 43428 28642
rect 43372 28588 43428 28590
rect 42700 28252 42756 28308
rect 43260 28418 43316 28420
rect 43260 28366 43262 28418
rect 43262 28366 43314 28418
rect 43314 28366 43316 28418
rect 43260 28364 43316 28366
rect 44156 29314 44212 29316
rect 44156 29262 44158 29314
rect 44158 29262 44210 29314
rect 44210 29262 44212 29314
rect 44156 29260 44212 29262
rect 43820 28364 43876 28420
rect 43036 27580 43092 27636
rect 43596 27580 43652 27636
rect 42476 27244 42532 27300
rect 42700 27244 42756 27300
rect 43148 27074 43204 27076
rect 43148 27022 43150 27074
rect 43150 27022 43202 27074
rect 43202 27022 43204 27074
rect 43148 27020 43204 27022
rect 42924 26962 42980 26964
rect 42924 26910 42926 26962
rect 42926 26910 42978 26962
rect 42978 26910 42980 26962
rect 42924 26908 42980 26910
rect 43932 26908 43988 26964
rect 42476 26684 42532 26740
rect 43932 26572 43988 26628
rect 42812 26402 42868 26404
rect 42812 26350 42814 26402
rect 42814 26350 42866 26402
rect 42866 26350 42868 26402
rect 42812 26348 42868 26350
rect 42588 26012 42644 26068
rect 42700 25900 42756 25956
rect 43484 26402 43540 26404
rect 43484 26350 43486 26402
rect 43486 26350 43538 26402
rect 43538 26350 43540 26402
rect 43484 26348 43540 26350
rect 46508 35420 46564 35476
rect 46396 35196 46452 35252
rect 47516 35196 47572 35252
rect 46620 34188 46676 34244
rect 46956 33068 47012 33124
rect 46060 32956 46116 33012
rect 48188 37212 48244 37268
rect 48412 37212 48468 37268
rect 48188 35922 48244 35924
rect 48188 35870 48190 35922
rect 48190 35870 48242 35922
rect 48242 35870 48244 35922
rect 48188 35868 48244 35870
rect 48076 35756 48132 35812
rect 48076 34188 48132 34244
rect 47516 33292 47572 33348
rect 47852 33068 47908 33124
rect 47068 31836 47124 31892
rect 47628 31948 47684 32004
rect 46172 31724 46228 31780
rect 45052 28642 45108 28644
rect 45052 28590 45054 28642
rect 45054 28590 45106 28642
rect 45106 28590 45108 28642
rect 45052 28588 45108 28590
rect 44940 27244 44996 27300
rect 45052 28364 45108 28420
rect 44380 26684 44436 26740
rect 44492 26908 44548 26964
rect 44828 26796 44884 26852
rect 43596 26290 43652 26292
rect 43596 26238 43598 26290
rect 43598 26238 43650 26290
rect 43650 26238 43652 26290
rect 43596 26236 43652 26238
rect 44940 26514 44996 26516
rect 44940 26462 44942 26514
rect 44942 26462 44994 26514
rect 44994 26462 44996 26514
rect 44940 26460 44996 26462
rect 43148 25788 43204 25844
rect 41692 24780 41748 24836
rect 41916 24108 41972 24164
rect 41804 23938 41860 23940
rect 41804 23886 41806 23938
rect 41806 23886 41858 23938
rect 41858 23886 41860 23938
rect 41804 23884 41860 23886
rect 41580 23436 41636 23492
rect 41468 23154 41524 23156
rect 41468 23102 41470 23154
rect 41470 23102 41522 23154
rect 41522 23102 41524 23154
rect 41468 23100 41524 23102
rect 42028 23324 42084 23380
rect 41804 22204 41860 22260
rect 41468 22146 41524 22148
rect 41468 22094 41470 22146
rect 41470 22094 41522 22146
rect 41522 22094 41524 22146
rect 41468 22092 41524 22094
rect 41916 21868 41972 21924
rect 41244 20690 41300 20692
rect 41244 20638 41246 20690
rect 41246 20638 41298 20690
rect 41298 20638 41300 20690
rect 41244 20636 41300 20638
rect 41804 21420 41860 21476
rect 42364 25228 42420 25284
rect 45388 28418 45444 28420
rect 45388 28366 45390 28418
rect 45390 28366 45442 28418
rect 45442 28366 45444 28418
rect 45388 28364 45444 28366
rect 45724 29260 45780 29316
rect 45836 28700 45892 28756
rect 45164 26236 45220 26292
rect 43596 25506 43652 25508
rect 43596 25454 43598 25506
rect 43598 25454 43650 25506
rect 43650 25454 43652 25506
rect 43596 25452 43652 25454
rect 43372 25340 43428 25396
rect 42476 24834 42532 24836
rect 42476 24782 42478 24834
rect 42478 24782 42530 24834
rect 42530 24782 42532 24834
rect 42476 24780 42532 24782
rect 43036 25282 43092 25284
rect 43036 25230 43038 25282
rect 43038 25230 43090 25282
rect 43090 25230 43092 25282
rect 43036 25228 43092 25230
rect 43148 24834 43204 24836
rect 43148 24782 43150 24834
rect 43150 24782 43202 24834
rect 43202 24782 43204 24834
rect 43148 24780 43204 24782
rect 42812 24108 42868 24164
rect 43148 23938 43204 23940
rect 43148 23886 43150 23938
rect 43150 23886 43202 23938
rect 43202 23886 43204 23938
rect 43148 23884 43204 23886
rect 42364 23548 42420 23604
rect 42476 23154 42532 23156
rect 42476 23102 42478 23154
rect 42478 23102 42530 23154
rect 42530 23102 42532 23154
rect 42476 23100 42532 23102
rect 42812 23436 42868 23492
rect 42700 23378 42756 23380
rect 42700 23326 42702 23378
rect 42702 23326 42754 23378
rect 42754 23326 42756 23378
rect 42700 23324 42756 23326
rect 43036 22428 43092 22484
rect 42924 22258 42980 22260
rect 42924 22206 42926 22258
rect 42926 22206 42978 22258
rect 42978 22206 42980 22258
rect 42924 22204 42980 22206
rect 42476 21474 42532 21476
rect 42476 21422 42478 21474
rect 42478 21422 42530 21474
rect 42530 21422 42532 21474
rect 42476 21420 42532 21422
rect 44044 25506 44100 25508
rect 44044 25454 44046 25506
rect 44046 25454 44098 25506
rect 44098 25454 44100 25506
rect 44044 25452 44100 25454
rect 43932 25282 43988 25284
rect 43932 25230 43934 25282
rect 43934 25230 43986 25282
rect 43986 25230 43988 25282
rect 43932 25228 43988 25230
rect 43596 24780 43652 24836
rect 44940 25394 44996 25396
rect 44940 25342 44942 25394
rect 44942 25342 44994 25394
rect 44994 25342 44996 25394
rect 44940 25340 44996 25342
rect 43596 23938 43652 23940
rect 43596 23886 43598 23938
rect 43598 23886 43650 23938
rect 43650 23886 43652 23938
rect 43596 23884 43652 23886
rect 44156 23884 44212 23940
rect 44044 23772 44100 23828
rect 43708 23660 43764 23716
rect 43596 23548 43652 23604
rect 43372 22540 43428 22596
rect 43484 22652 43540 22708
rect 43372 21868 43428 21924
rect 41580 20636 41636 20692
rect 41356 20300 41412 20356
rect 41468 20524 41524 20580
rect 41020 20076 41076 20132
rect 41580 20076 41636 20132
rect 41132 20018 41188 20020
rect 41132 19966 41134 20018
rect 41134 19966 41186 20018
rect 41186 19966 41188 20018
rect 41132 19964 41188 19966
rect 41468 19740 41524 19796
rect 40908 19628 40964 19684
rect 41020 19180 41076 19236
rect 40572 18956 40628 19012
rect 41132 18956 41188 19012
rect 40908 18450 40964 18452
rect 40908 18398 40910 18450
rect 40910 18398 40962 18450
rect 40962 18398 40964 18450
rect 40908 18396 40964 18398
rect 40348 18226 40404 18228
rect 40348 18174 40350 18226
rect 40350 18174 40402 18226
rect 40402 18174 40404 18226
rect 40348 18172 40404 18174
rect 40236 16716 40292 16772
rect 40348 17106 40404 17108
rect 40348 17054 40350 17106
rect 40350 17054 40402 17106
rect 40402 17054 40404 17106
rect 40348 17052 40404 17054
rect 39900 16604 39956 16660
rect 39788 16156 39844 16212
rect 40012 15538 40068 15540
rect 40012 15486 40014 15538
rect 40014 15486 40066 15538
rect 40066 15486 40068 15538
rect 40012 15484 40068 15486
rect 39900 14530 39956 14532
rect 39900 14478 39902 14530
rect 39902 14478 39954 14530
rect 39954 14478 39956 14530
rect 39900 14476 39956 14478
rect 40236 14028 40292 14084
rect 39676 13746 39732 13748
rect 39676 13694 39678 13746
rect 39678 13694 39730 13746
rect 39730 13694 39732 13746
rect 39676 13692 39732 13694
rect 40124 13634 40180 13636
rect 40124 13582 40126 13634
rect 40126 13582 40178 13634
rect 40178 13582 40180 13634
rect 40124 13580 40180 13582
rect 37548 12066 37604 12068
rect 37548 12014 37550 12066
rect 37550 12014 37602 12066
rect 37602 12014 37604 12066
rect 37548 12012 37604 12014
rect 37660 11340 37716 11396
rect 37660 10834 37716 10836
rect 37660 10782 37662 10834
rect 37662 10782 37714 10834
rect 37714 10782 37716 10834
rect 37660 10780 37716 10782
rect 38668 12124 38724 12180
rect 37996 11340 38052 11396
rect 38444 12012 38500 12068
rect 38220 11004 38276 11060
rect 38332 11116 38388 11172
rect 37884 10668 37940 10724
rect 38220 10668 38276 10724
rect 36652 8316 36708 8372
rect 37100 9602 37156 9604
rect 37100 9550 37102 9602
rect 37102 9550 37154 9602
rect 37154 9550 37156 9602
rect 37100 9548 37156 9550
rect 37100 8540 37156 8596
rect 37212 8370 37268 8372
rect 37212 8318 37214 8370
rect 37214 8318 37266 8370
rect 37266 8318 37268 8370
rect 37212 8316 37268 8318
rect 38332 9884 38388 9940
rect 40124 12738 40180 12740
rect 40124 12686 40126 12738
rect 40126 12686 40178 12738
rect 40178 12686 40180 12738
rect 40124 12684 40180 12686
rect 40236 12572 40292 12628
rect 39452 12178 39508 12180
rect 39452 12126 39454 12178
rect 39454 12126 39506 12178
rect 39506 12126 39508 12178
rect 39452 12124 39508 12126
rect 41804 20300 41860 20356
rect 42140 20188 42196 20244
rect 42028 19964 42084 20020
rect 42364 20578 42420 20580
rect 42364 20526 42366 20578
rect 42366 20526 42418 20578
rect 42418 20526 42420 20578
rect 42364 20524 42420 20526
rect 41692 18956 41748 19012
rect 41468 18172 41524 18228
rect 41020 16770 41076 16772
rect 41020 16718 41022 16770
rect 41022 16718 41074 16770
rect 41074 16718 41076 16770
rect 41020 16716 41076 16718
rect 41580 17612 41636 17668
rect 42924 20914 42980 20916
rect 42924 20862 42926 20914
rect 42926 20862 42978 20914
rect 42978 20862 42980 20914
rect 42924 20860 42980 20862
rect 42812 20690 42868 20692
rect 42812 20638 42814 20690
rect 42814 20638 42866 20690
rect 42866 20638 42868 20690
rect 42812 20636 42868 20638
rect 43372 20018 43428 20020
rect 43372 19966 43374 20018
rect 43374 19966 43426 20018
rect 43426 19966 43428 20018
rect 43372 19964 43428 19966
rect 42588 19852 42644 19908
rect 42700 19010 42756 19012
rect 42700 18958 42702 19010
rect 42702 18958 42754 19010
rect 42754 18958 42756 19010
rect 42700 18956 42756 18958
rect 43260 18620 43316 18676
rect 43708 23436 43764 23492
rect 44940 23548 44996 23604
rect 45164 25452 45220 25508
rect 46844 31666 46900 31668
rect 46844 31614 46846 31666
rect 46846 31614 46898 31666
rect 46898 31614 46900 31666
rect 46844 31612 46900 31614
rect 46508 31554 46564 31556
rect 46508 31502 46510 31554
rect 46510 31502 46562 31554
rect 46562 31502 46564 31554
rect 46508 31500 46564 31502
rect 46396 31164 46452 31220
rect 47180 31500 47236 31556
rect 47404 31388 47460 31444
rect 47964 32956 48020 33012
rect 48300 32620 48356 32676
rect 48524 31836 48580 31892
rect 47404 28642 47460 28644
rect 47404 28590 47406 28642
rect 47406 28590 47458 28642
rect 47458 28590 47460 28642
rect 47404 28588 47460 28590
rect 48076 28028 48132 28084
rect 48188 28642 48244 28644
rect 48188 28590 48190 28642
rect 48190 28590 48242 28642
rect 48242 28590 48244 28642
rect 48188 28588 48244 28590
rect 48188 27356 48244 27412
rect 47628 26908 47684 26964
rect 45836 26460 45892 26516
rect 45052 23772 45108 23828
rect 45388 23884 45444 23940
rect 44492 23436 44548 23492
rect 45164 23548 45220 23604
rect 45052 23042 45108 23044
rect 45052 22990 45054 23042
rect 45054 22990 45106 23042
rect 45106 22990 45108 23042
rect 45052 22988 45108 22990
rect 44268 22930 44324 22932
rect 44268 22878 44270 22930
rect 44270 22878 44322 22930
rect 44322 22878 44324 22930
rect 44268 22876 44324 22878
rect 43708 22482 43764 22484
rect 43708 22430 43710 22482
rect 43710 22430 43762 22482
rect 43762 22430 43764 22482
rect 43708 22428 43764 22430
rect 44268 21420 44324 21476
rect 44492 21698 44548 21700
rect 44492 21646 44494 21698
rect 44494 21646 44546 21698
rect 44546 21646 44548 21698
rect 44492 21644 44548 21646
rect 43708 20914 43764 20916
rect 43708 20862 43710 20914
rect 43710 20862 43762 20914
rect 43762 20862 43764 20914
rect 43708 20860 43764 20862
rect 44828 21586 44884 21588
rect 44828 21534 44830 21586
rect 44830 21534 44882 21586
rect 44882 21534 44884 21586
rect 44828 21532 44884 21534
rect 48188 27132 48244 27188
rect 46508 26290 46564 26292
rect 46508 26238 46510 26290
rect 46510 26238 46562 26290
rect 46562 26238 46564 26290
rect 46508 26236 46564 26238
rect 47068 25788 47124 25844
rect 47180 25340 47236 25396
rect 48188 25340 48244 25396
rect 46060 23212 46116 23268
rect 46396 23772 46452 23828
rect 45836 22988 45892 23044
rect 46060 22930 46116 22932
rect 46060 22878 46062 22930
rect 46062 22878 46114 22930
rect 46114 22878 46116 22930
rect 46060 22876 46116 22878
rect 45276 22652 45332 22708
rect 45276 22482 45332 22484
rect 45276 22430 45278 22482
rect 45278 22430 45330 22482
rect 45330 22430 45332 22482
rect 45276 22428 45332 22430
rect 45612 22204 45668 22260
rect 45388 21868 45444 21924
rect 45276 21474 45332 21476
rect 45276 21422 45278 21474
rect 45278 21422 45330 21474
rect 45330 21422 45332 21474
rect 45276 21420 45332 21422
rect 45500 21756 45556 21812
rect 46060 21756 46116 21812
rect 46396 21644 46452 21700
rect 46284 21362 46340 21364
rect 46284 21310 46286 21362
rect 46286 21310 46338 21362
rect 46338 21310 46340 21362
rect 46284 21308 46340 21310
rect 43932 19234 43988 19236
rect 43932 19182 43934 19234
rect 43934 19182 43986 19234
rect 43986 19182 43988 19234
rect 43932 19180 43988 19182
rect 44828 19234 44884 19236
rect 44828 19182 44830 19234
rect 44830 19182 44882 19234
rect 44882 19182 44884 19234
rect 44828 19180 44884 19182
rect 43708 18396 43764 18452
rect 43596 17836 43652 17892
rect 43820 17612 43876 17668
rect 41916 17052 41972 17108
rect 41356 16604 41412 16660
rect 40908 15202 40964 15204
rect 40908 15150 40910 15202
rect 40910 15150 40962 15202
rect 40962 15150 40964 15202
rect 40908 15148 40964 15150
rect 40572 14700 40628 14756
rect 41356 14588 41412 14644
rect 41468 15148 41524 15204
rect 40460 14530 40516 14532
rect 40460 14478 40462 14530
rect 40462 14478 40514 14530
rect 40514 14478 40516 14530
rect 40460 14476 40516 14478
rect 41580 14476 41636 14532
rect 41692 14252 41748 14308
rect 41020 14028 41076 14084
rect 40460 13074 40516 13076
rect 40460 13022 40462 13074
rect 40462 13022 40514 13074
rect 40514 13022 40516 13074
rect 40460 13020 40516 13022
rect 40908 12684 40964 12740
rect 41132 12572 41188 12628
rect 39340 11394 39396 11396
rect 39340 11342 39342 11394
rect 39342 11342 39394 11394
rect 39394 11342 39396 11394
rect 39340 11340 39396 11342
rect 39788 11340 39844 11396
rect 40236 11282 40292 11284
rect 40236 11230 40238 11282
rect 40238 11230 40290 11282
rect 40290 11230 40292 11282
rect 40236 11228 40292 11230
rect 40124 11170 40180 11172
rect 40124 11118 40126 11170
rect 40126 11118 40178 11170
rect 40178 11118 40180 11170
rect 40124 11116 40180 11118
rect 41580 12012 41636 12068
rect 40796 11394 40852 11396
rect 40796 11342 40798 11394
rect 40798 11342 40850 11394
rect 40850 11342 40852 11394
rect 40796 11340 40852 11342
rect 40684 10668 40740 10724
rect 40908 11228 40964 11284
rect 41020 11004 41076 11060
rect 39004 10498 39060 10500
rect 39004 10446 39006 10498
rect 39006 10446 39058 10498
rect 39058 10446 39060 10498
rect 39004 10444 39060 10446
rect 38892 9938 38948 9940
rect 38892 9886 38894 9938
rect 38894 9886 38946 9938
rect 38946 9886 38948 9938
rect 38892 9884 38948 9886
rect 38444 9772 38500 9828
rect 39676 9042 39732 9044
rect 39676 8990 39678 9042
rect 39678 8990 39730 9042
rect 39730 8990 39732 9042
rect 39676 8988 39732 8990
rect 38668 8540 38724 8596
rect 37436 8370 37492 8372
rect 37436 8318 37438 8370
rect 37438 8318 37490 8370
rect 37490 8318 37492 8370
rect 37436 8316 37492 8318
rect 38332 8370 38388 8372
rect 38332 8318 38334 8370
rect 38334 8318 38386 8370
rect 38386 8318 38388 8370
rect 38332 8316 38388 8318
rect 37660 8146 37716 8148
rect 37660 8094 37662 8146
rect 37662 8094 37714 8146
rect 37714 8094 37716 8146
rect 37660 8092 37716 8094
rect 37884 8146 37940 8148
rect 37884 8094 37886 8146
rect 37886 8094 37938 8146
rect 37938 8094 37940 8146
rect 37884 8092 37940 8094
rect 37660 7308 37716 7364
rect 37660 6748 37716 6804
rect 38332 7084 38388 7140
rect 36988 6690 37044 6692
rect 36988 6638 36990 6690
rect 36990 6638 37042 6690
rect 37042 6638 37044 6690
rect 36988 6636 37044 6638
rect 36092 6524 36148 6580
rect 41468 10780 41524 10836
rect 42588 16604 42644 16660
rect 43036 15202 43092 15204
rect 43036 15150 43038 15202
rect 43038 15150 43090 15202
rect 43090 15150 43092 15202
rect 43036 15148 43092 15150
rect 42028 14306 42084 14308
rect 42028 14254 42030 14306
rect 42030 14254 42082 14306
rect 42082 14254 42084 14306
rect 42028 14252 42084 14254
rect 42924 14588 42980 14644
rect 43148 14530 43204 14532
rect 43148 14478 43150 14530
rect 43150 14478 43202 14530
rect 43202 14478 43204 14530
rect 43148 14476 43204 14478
rect 41804 13020 41860 13076
rect 41804 12684 41860 12740
rect 41916 13132 41972 13188
rect 41916 12572 41972 12628
rect 41916 12348 41972 12404
rect 41804 10556 41860 10612
rect 43372 16268 43428 16324
rect 44156 16268 44212 16324
rect 46172 20412 46228 20468
rect 47404 23826 47460 23828
rect 47404 23774 47406 23826
rect 47406 23774 47458 23826
rect 47458 23774 47460 23826
rect 47404 23772 47460 23774
rect 47292 23212 47348 23268
rect 46732 21586 46788 21588
rect 46732 21534 46734 21586
rect 46734 21534 46786 21586
rect 46786 21534 46788 21586
rect 46732 21532 46788 21534
rect 46956 20412 47012 20468
rect 47628 23042 47684 23044
rect 47628 22990 47630 23042
rect 47630 22990 47682 23042
rect 47682 22990 47684 23042
rect 47628 22988 47684 22990
rect 48188 22988 48244 23044
rect 48188 22428 48244 22484
rect 47404 22258 47460 22260
rect 47404 22206 47406 22258
rect 47406 22206 47458 22258
rect 47458 22206 47460 22258
rect 47404 22204 47460 22206
rect 48076 21868 48132 21924
rect 47964 21810 48020 21812
rect 47964 21758 47966 21810
rect 47966 21758 48018 21810
rect 48018 21758 48020 21810
rect 47964 21756 48020 21758
rect 48188 21756 48244 21812
rect 47740 21474 47796 21476
rect 47740 21422 47742 21474
rect 47742 21422 47794 21474
rect 47794 21422 47796 21474
rect 47740 21420 47796 21422
rect 47852 21308 47908 21364
rect 48188 20914 48244 20916
rect 48188 20862 48190 20914
rect 48190 20862 48242 20914
rect 48242 20862 48244 20914
rect 48188 20860 48244 20862
rect 47180 20524 47236 20580
rect 45388 18396 45444 18452
rect 46844 18396 46900 18452
rect 45052 18284 45108 18340
rect 44940 17836 44996 17892
rect 45612 17724 45668 17780
rect 44828 15874 44884 15876
rect 44828 15822 44830 15874
rect 44830 15822 44882 15874
rect 44882 15822 44884 15874
rect 44828 15820 44884 15822
rect 43484 14700 43540 14756
rect 43596 14588 43652 14644
rect 42812 13746 42868 13748
rect 42812 13694 42814 13746
rect 42814 13694 42866 13746
rect 42866 13694 42868 13746
rect 42812 13692 42868 13694
rect 42476 13580 42532 13636
rect 42588 13468 42644 13524
rect 42140 12572 42196 12628
rect 42252 12684 42308 12740
rect 42476 12402 42532 12404
rect 42476 12350 42478 12402
rect 42478 12350 42530 12402
rect 42530 12350 42532 12402
rect 42476 12348 42532 12350
rect 42252 12124 42308 12180
rect 42140 12012 42196 12068
rect 43372 13692 43428 13748
rect 43036 13634 43092 13636
rect 43036 13582 43038 13634
rect 43038 13582 43090 13634
rect 43090 13582 43092 13634
rect 43036 13580 43092 13582
rect 42700 12572 42756 12628
rect 42812 12908 42868 12964
rect 42700 12178 42756 12180
rect 42700 12126 42702 12178
rect 42702 12126 42754 12178
rect 42754 12126 42756 12178
rect 42700 12124 42756 12126
rect 43036 12738 43092 12740
rect 43036 12686 43038 12738
rect 43038 12686 43090 12738
rect 43090 12686 43092 12738
rect 43036 12684 43092 12686
rect 42924 12012 42980 12068
rect 43036 12460 43092 12516
rect 42700 11228 42756 11284
rect 44044 13916 44100 13972
rect 43708 13580 43764 13636
rect 43932 13746 43988 13748
rect 43932 13694 43934 13746
rect 43934 13694 43986 13746
rect 43986 13694 43988 13746
rect 43932 13692 43988 13694
rect 43820 13468 43876 13524
rect 43596 12962 43652 12964
rect 43596 12910 43598 12962
rect 43598 12910 43650 12962
rect 43650 12910 43652 12962
rect 43596 12908 43652 12910
rect 44268 12962 44324 12964
rect 44268 12910 44270 12962
rect 44270 12910 44322 12962
rect 44322 12910 44324 12962
rect 44268 12908 44324 12910
rect 44268 12684 44324 12740
rect 42140 11004 42196 11060
rect 42028 10834 42084 10836
rect 42028 10782 42030 10834
rect 42030 10782 42082 10834
rect 42082 10782 42084 10834
rect 42028 10780 42084 10782
rect 41692 10108 41748 10164
rect 41468 9548 41524 9604
rect 40348 9154 40404 9156
rect 40348 9102 40350 9154
rect 40350 9102 40402 9154
rect 40402 9102 40404 9154
rect 40348 9100 40404 9102
rect 41132 9154 41188 9156
rect 41132 9102 41134 9154
rect 41134 9102 41186 9154
rect 41186 9102 41188 9154
rect 41132 9100 41188 9102
rect 39788 8316 39844 8372
rect 38780 8258 38836 8260
rect 38780 8206 38782 8258
rect 38782 8206 38834 8258
rect 38834 8206 38836 8258
rect 38780 8204 38836 8206
rect 39452 8092 39508 8148
rect 41356 8988 41412 9044
rect 40348 8482 40404 8484
rect 40348 8430 40350 8482
rect 40350 8430 40402 8482
rect 40402 8430 40404 8482
rect 40348 8428 40404 8430
rect 40124 8092 40180 8148
rect 40012 7644 40068 7700
rect 40012 7362 40068 7364
rect 40012 7310 40014 7362
rect 40014 7310 40066 7362
rect 40066 7310 40068 7362
rect 40012 7308 40068 7310
rect 40908 8316 40964 8372
rect 42140 9548 42196 9604
rect 41020 8204 41076 8260
rect 41244 7980 41300 8036
rect 41468 7698 41524 7700
rect 41468 7646 41470 7698
rect 41470 7646 41522 7698
rect 41522 7646 41524 7698
rect 41468 7644 41524 7646
rect 39228 5906 39284 5908
rect 39228 5854 39230 5906
rect 39230 5854 39282 5906
rect 39282 5854 39284 5906
rect 39228 5852 39284 5854
rect 36988 5628 37044 5684
rect 36316 5404 36372 5460
rect 36876 5292 36932 5348
rect 34972 4844 35028 4900
rect 34076 4338 34132 4340
rect 34076 4286 34078 4338
rect 34078 4286 34130 4338
rect 34130 4286 34132 4338
rect 34076 4284 34132 4286
rect 36092 4732 36148 4788
rect 38220 5404 38276 5460
rect 39228 5292 39284 5348
rect 39452 6130 39508 6132
rect 39452 6078 39454 6130
rect 39454 6078 39506 6130
rect 39506 6078 39508 6130
rect 39452 6076 39508 6078
rect 40236 6076 40292 6132
rect 39564 5628 39620 5684
rect 39788 5404 39844 5460
rect 39900 5852 39956 5908
rect 40236 5794 40292 5796
rect 40236 5742 40238 5794
rect 40238 5742 40290 5794
rect 40290 5742 40292 5794
rect 40236 5740 40292 5742
rect 40124 5628 40180 5684
rect 40236 5346 40292 5348
rect 40236 5294 40238 5346
rect 40238 5294 40290 5346
rect 40290 5294 40292 5346
rect 40236 5292 40292 5294
rect 41020 6076 41076 6132
rect 41132 6018 41188 6020
rect 41132 5966 41134 6018
rect 41134 5966 41186 6018
rect 41186 5966 41188 6018
rect 41132 5964 41188 5966
rect 40572 5292 40628 5348
rect 41692 7474 41748 7476
rect 41692 7422 41694 7474
rect 41694 7422 41746 7474
rect 41746 7422 41748 7474
rect 41692 7420 41748 7422
rect 42140 9042 42196 9044
rect 42140 8990 42142 9042
rect 42142 8990 42194 9042
rect 42194 8990 42196 9042
rect 42140 8988 42196 8990
rect 42252 8876 42308 8932
rect 43932 11282 43988 11284
rect 43932 11230 43934 11282
rect 43934 11230 43986 11282
rect 43986 11230 43988 11282
rect 43932 11228 43988 11230
rect 43596 11170 43652 11172
rect 43596 11118 43598 11170
rect 43598 11118 43650 11170
rect 43650 11118 43652 11170
rect 43596 11116 43652 11118
rect 43484 10610 43540 10612
rect 43484 10558 43486 10610
rect 43486 10558 43538 10610
rect 43538 10558 43540 10610
rect 43484 10556 43540 10558
rect 43372 9884 43428 9940
rect 43148 9602 43204 9604
rect 43148 9550 43150 9602
rect 43150 9550 43202 9602
rect 43202 9550 43204 9602
rect 43148 9548 43204 9550
rect 43372 9548 43428 9604
rect 42476 9212 42532 9268
rect 42924 9266 42980 9268
rect 42924 9214 42926 9266
rect 42926 9214 42978 9266
rect 42978 9214 42980 9266
rect 42924 9212 42980 9214
rect 43036 9154 43092 9156
rect 43036 9102 43038 9154
rect 43038 9102 43090 9154
rect 43090 9102 43092 9154
rect 43036 9100 43092 9102
rect 43148 9042 43204 9044
rect 43148 8990 43150 9042
rect 43150 8990 43202 9042
rect 43202 8990 43204 9042
rect 43148 8988 43204 8990
rect 42140 8258 42196 8260
rect 42140 8206 42142 8258
rect 42142 8206 42194 8258
rect 42194 8206 42196 8258
rect 42140 8204 42196 8206
rect 42364 8146 42420 8148
rect 42364 8094 42366 8146
rect 42366 8094 42418 8146
rect 42418 8094 42420 8146
rect 42364 8092 42420 8094
rect 42028 7532 42084 7588
rect 42252 7868 42308 7924
rect 42028 7250 42084 7252
rect 42028 7198 42030 7250
rect 42030 7198 42082 7250
rect 42082 7198 42084 7250
rect 42028 7196 42084 7198
rect 42588 8146 42644 8148
rect 42588 8094 42590 8146
rect 42590 8094 42642 8146
rect 42642 8094 42644 8146
rect 42588 8092 42644 8094
rect 42700 7980 42756 8036
rect 42924 7532 42980 7588
rect 41692 6300 41748 6356
rect 37436 5068 37492 5124
rect 41580 5794 41636 5796
rect 41580 5742 41582 5794
rect 41582 5742 41634 5794
rect 41634 5742 41636 5794
rect 41580 5740 41636 5742
rect 41244 5628 41300 5684
rect 40684 5122 40740 5124
rect 40684 5070 40686 5122
rect 40686 5070 40738 5122
rect 40738 5070 40740 5122
rect 40684 5068 40740 5070
rect 41020 5068 41076 5124
rect 37996 4898 38052 4900
rect 37996 4846 37998 4898
rect 37998 4846 38050 4898
rect 38050 4846 38052 4898
rect 37996 4844 38052 4846
rect 39564 4450 39620 4452
rect 39564 4398 39566 4450
rect 39566 4398 39618 4450
rect 39618 4398 39620 4450
rect 39564 4396 39620 4398
rect 40908 4450 40964 4452
rect 40908 4398 40910 4450
rect 40910 4398 40962 4450
rect 40962 4398 40964 4450
rect 40908 4396 40964 4398
rect 41356 5292 41412 5348
rect 41580 5516 41636 5572
rect 42364 6578 42420 6580
rect 42364 6526 42366 6578
rect 42366 6526 42418 6578
rect 42418 6526 42420 6578
rect 42364 6524 42420 6526
rect 42140 6466 42196 6468
rect 42140 6414 42142 6466
rect 42142 6414 42194 6466
rect 42194 6414 42196 6466
rect 42140 6412 42196 6414
rect 41804 5292 41860 5348
rect 41916 5852 41972 5908
rect 41692 5180 41748 5236
rect 41356 5122 41412 5124
rect 41356 5070 41358 5122
rect 41358 5070 41410 5122
rect 41410 5070 41412 5122
rect 41356 5068 41412 5070
rect 42252 5682 42308 5684
rect 42252 5630 42254 5682
rect 42254 5630 42306 5682
rect 42306 5630 42308 5682
rect 42252 5628 42308 5630
rect 42924 6578 42980 6580
rect 42924 6526 42926 6578
rect 42926 6526 42978 6578
rect 42978 6526 42980 6578
rect 42924 6524 42980 6526
rect 42812 6466 42868 6468
rect 42812 6414 42814 6466
rect 42814 6414 42866 6466
rect 42866 6414 42868 6466
rect 42812 6412 42868 6414
rect 42364 5516 42420 5572
rect 42252 5404 42308 5460
rect 42028 5068 42084 5124
rect 42140 5292 42196 5348
rect 40348 4338 40404 4340
rect 40348 4286 40350 4338
rect 40350 4286 40402 4338
rect 40402 4286 40404 4338
rect 40348 4284 40404 4286
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 39676 3836 39732 3892
rect 36540 3724 36596 3780
rect 35980 3554 36036 3556
rect 35980 3502 35982 3554
rect 35982 3502 36034 3554
rect 36034 3502 36036 3554
rect 35980 3500 36036 3502
rect 36988 3666 37044 3668
rect 36988 3614 36990 3666
rect 36990 3614 37042 3666
rect 37042 3614 37044 3666
rect 36988 3612 37044 3614
rect 38108 3276 38164 3332
rect 38892 3330 38948 3332
rect 38892 3278 38894 3330
rect 38894 3278 38946 3330
rect 38946 3278 38948 3330
rect 38892 3276 38948 3278
rect 42364 5180 42420 5236
rect 41580 3836 41636 3892
rect 40012 3778 40068 3780
rect 40012 3726 40014 3778
rect 40014 3726 40066 3778
rect 40066 3726 40068 3778
rect 40012 3724 40068 3726
rect 42812 5906 42868 5908
rect 42812 5854 42814 5906
rect 42814 5854 42866 5906
rect 42866 5854 42868 5906
rect 42812 5852 42868 5854
rect 43148 8146 43204 8148
rect 43148 8094 43150 8146
rect 43150 8094 43202 8146
rect 43202 8094 43204 8146
rect 43148 8092 43204 8094
rect 43260 7868 43316 7924
rect 43372 7586 43428 7588
rect 43372 7534 43374 7586
rect 43374 7534 43426 7586
rect 43426 7534 43428 7586
rect 43372 7532 43428 7534
rect 43260 7196 43316 7252
rect 43932 9884 43988 9940
rect 46284 16156 46340 16212
rect 46732 15372 46788 15428
rect 45388 14530 45444 14532
rect 45388 14478 45390 14530
rect 45390 14478 45442 14530
rect 45442 14478 45444 14530
rect 45388 14476 45444 14478
rect 45500 14700 45556 14756
rect 44492 14364 44548 14420
rect 45612 14530 45668 14532
rect 45612 14478 45614 14530
rect 45614 14478 45666 14530
rect 45666 14478 45668 14530
rect 45612 14476 45668 14478
rect 48076 18396 48132 18452
rect 47068 18338 47124 18340
rect 47068 18286 47070 18338
rect 47070 18286 47122 18338
rect 47122 18286 47124 18338
rect 47068 18284 47124 18286
rect 47852 18060 47908 18116
rect 47180 17778 47236 17780
rect 47180 17726 47182 17778
rect 47182 17726 47234 17778
rect 47234 17726 47236 17778
rect 47180 17724 47236 17726
rect 47404 16210 47460 16212
rect 47404 16158 47406 16210
rect 47406 16158 47458 16210
rect 47458 16158 47460 16210
rect 47404 16156 47460 16158
rect 48524 17724 48580 17780
rect 48188 17554 48244 17556
rect 48188 17502 48190 17554
rect 48190 17502 48242 17554
rect 48242 17502 48244 17554
rect 48188 17500 48244 17502
rect 47404 15426 47460 15428
rect 47404 15374 47406 15426
rect 47406 15374 47458 15426
rect 47458 15374 47460 15426
rect 47404 15372 47460 15374
rect 46732 14476 46788 14532
rect 46172 14418 46228 14420
rect 46172 14366 46174 14418
rect 46174 14366 46226 14418
rect 46226 14366 46228 14418
rect 46172 14364 46228 14366
rect 46508 14306 46564 14308
rect 46508 14254 46510 14306
rect 46510 14254 46562 14306
rect 46562 14254 46564 14306
rect 46508 14252 46564 14254
rect 47404 14252 47460 14308
rect 45164 14028 45220 14084
rect 45276 13132 45332 13188
rect 45388 12962 45444 12964
rect 45388 12910 45390 12962
rect 45390 12910 45442 12962
rect 45442 12910 45444 12962
rect 45388 12908 45444 12910
rect 47852 12850 47908 12852
rect 47852 12798 47854 12850
rect 47854 12798 47906 12850
rect 47906 12798 47908 12850
rect 47852 12796 47908 12798
rect 46396 12738 46452 12740
rect 46396 12686 46398 12738
rect 46398 12686 46450 12738
rect 46450 12686 46452 12738
rect 46396 12684 46452 12686
rect 47404 12684 47460 12740
rect 47628 12572 47684 12628
rect 48188 12572 48244 12628
rect 44604 11732 44660 11788
rect 44492 11340 44548 11396
rect 44268 9548 44324 9604
rect 44268 9042 44324 9044
rect 44268 8990 44270 9042
rect 44270 8990 44322 9042
rect 44322 8990 44324 9042
rect 44268 8988 44324 8990
rect 43820 8370 43876 8372
rect 43820 8318 43822 8370
rect 43822 8318 43874 8370
rect 43874 8318 43876 8370
rect 43820 8316 43876 8318
rect 43596 7980 43652 8036
rect 43596 7474 43652 7476
rect 43596 7422 43598 7474
rect 43598 7422 43650 7474
rect 43650 7422 43652 7474
rect 43596 7420 43652 7422
rect 43484 7308 43540 7364
rect 43372 6636 43428 6692
rect 43260 6578 43316 6580
rect 43260 6526 43262 6578
rect 43262 6526 43314 6578
rect 43314 6526 43316 6578
rect 43260 6524 43316 6526
rect 42812 5404 42868 5460
rect 43484 5234 43540 5236
rect 43484 5182 43486 5234
rect 43486 5182 43538 5234
rect 43538 5182 43540 5234
rect 43484 5180 43540 5182
rect 45276 12066 45332 12068
rect 45276 12014 45278 12066
rect 45278 12014 45330 12066
rect 45330 12014 45332 12066
rect 45276 12012 45332 12014
rect 45164 11564 45220 11620
rect 44604 9212 44660 9268
rect 45276 11394 45332 11396
rect 45276 11342 45278 11394
rect 45278 11342 45330 11394
rect 45330 11342 45332 11394
rect 45276 11340 45332 11342
rect 46732 11394 46788 11396
rect 46732 11342 46734 11394
rect 46734 11342 46786 11394
rect 46786 11342 46788 11394
rect 46732 11340 46788 11342
rect 44716 11116 44772 11172
rect 45164 11004 45220 11060
rect 45276 9938 45332 9940
rect 45276 9886 45278 9938
rect 45278 9886 45330 9938
rect 45330 9886 45332 9938
rect 45276 9884 45332 9886
rect 46284 9884 46340 9940
rect 47404 9938 47460 9940
rect 47404 9886 47406 9938
rect 47406 9886 47458 9938
rect 47458 9886 47460 9938
rect 47404 9884 47460 9886
rect 45276 8930 45332 8932
rect 45276 8878 45278 8930
rect 45278 8878 45330 8930
rect 45330 8878 45332 8930
rect 45276 8876 45332 8878
rect 46508 8876 46564 8932
rect 44716 8316 44772 8372
rect 44828 8428 44884 8484
rect 44716 8092 44772 8148
rect 43932 7308 43988 7364
rect 44044 7196 44100 7252
rect 43820 6690 43876 6692
rect 43820 6638 43822 6690
rect 43822 6638 43874 6690
rect 43874 6638 43876 6690
rect 43820 6636 43876 6638
rect 44156 7084 44212 7140
rect 43708 5180 43764 5236
rect 43596 3612 43652 3668
rect 45164 8204 45220 8260
rect 44604 7362 44660 7364
rect 44604 7310 44606 7362
rect 44606 7310 44658 7362
rect 44658 7310 44660 7362
rect 44604 7308 44660 7310
rect 44940 7084 44996 7140
rect 45052 7420 45108 7476
rect 44492 6860 44548 6916
rect 44828 6524 44884 6580
rect 47404 8930 47460 8932
rect 47404 8878 47406 8930
rect 47406 8878 47458 8930
rect 47458 8878 47460 8930
rect 47404 8876 47460 8878
rect 47180 8482 47236 8484
rect 47180 8430 47182 8482
rect 47182 8430 47234 8482
rect 47234 8430 47236 8482
rect 47180 8428 47236 8430
rect 46844 8370 46900 8372
rect 46844 8318 46846 8370
rect 46846 8318 46898 8370
rect 46898 8318 46900 8370
rect 46844 8316 46900 8318
rect 47852 8146 47908 8148
rect 47852 8094 47854 8146
rect 47854 8094 47906 8146
rect 47906 8094 47908 8146
rect 47852 8092 47908 8094
rect 45276 7980 45332 8036
rect 47068 8034 47124 8036
rect 47068 7982 47070 8034
rect 47070 7982 47122 8034
rect 47122 7982 47124 8034
rect 47068 7980 47124 7982
rect 45500 7084 45556 7140
rect 45276 6914 45332 6916
rect 45276 6862 45278 6914
rect 45278 6862 45330 6914
rect 45330 6862 45332 6914
rect 45276 6860 45332 6862
rect 46732 6860 46788 6916
rect 47852 6748 47908 6804
rect 47628 6690 47684 6692
rect 47628 6638 47630 6690
rect 47630 6638 47682 6690
rect 47682 6638 47684 6690
rect 47628 6636 47684 6638
rect 46284 6466 46340 6468
rect 46284 6414 46286 6466
rect 46286 6414 46338 6466
rect 46338 6414 46340 6466
rect 46284 6412 46340 6414
rect 47404 6412 47460 6468
rect 48188 7644 48244 7700
rect 48188 6690 48244 6692
rect 48188 6638 48190 6690
rect 48190 6638 48242 6690
rect 48242 6638 48244 6690
rect 48188 6636 48244 6638
rect 44828 5292 44884 5348
rect 44156 5068 44212 5124
rect 46956 5122 47012 5124
rect 46956 5070 46958 5122
rect 46958 5070 47010 5122
rect 47010 5070 47012 5122
rect 46956 5068 47012 5070
rect 45388 4284 45444 4340
rect 47628 4284 47684 4340
rect 45500 3666 45556 3668
rect 45500 3614 45502 3666
rect 45502 3614 45554 3666
rect 45554 3614 45556 3666
rect 45500 3612 45556 3614
rect 41244 1708 41300 1764
rect 42700 1708 42756 1764
rect 42812 3276 42868 3332
rect 44492 3330 44548 3332
rect 44492 3278 44494 3330
rect 44494 3278 44546 3330
rect 44546 3278 44548 3330
rect 44492 3276 44548 3278
rect 47852 3442 47908 3444
rect 47852 3390 47854 3442
rect 47854 3390 47906 3442
rect 47906 3390 47908 3442
rect 47852 3388 47908 3390
rect 47628 3276 47684 3332
rect 48188 3276 48244 3332
rect 48188 2716 48244 2772
<< metal3 >>
rect 49200 47124 50000 47152
rect 45266 47068 45276 47124
rect 45332 47068 50000 47124
rect 49200 47040 50000 47068
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 43250 45948 43260 46004
rect 43316 45948 43708 46004
rect 43652 45892 43708 45948
rect 17490 45836 17500 45892
rect 17556 45836 18060 45892
rect 18116 45836 19628 45892
rect 19684 45836 19694 45892
rect 43652 45836 43820 45892
rect 43876 45836 43886 45892
rect 24658 45724 24668 45780
rect 24724 45724 29148 45780
rect 29204 45724 29214 45780
rect 30594 45724 30604 45780
rect 30660 45724 33068 45780
rect 33124 45724 33134 45780
rect 38546 45724 38556 45780
rect 38612 45724 41692 45780
rect 41748 45724 41758 45780
rect 46610 45724 46620 45780
rect 46676 45724 47404 45780
rect 47460 45724 47470 45780
rect 31602 45612 31612 45668
rect 31668 45612 33852 45668
rect 33908 45612 33918 45668
rect 37986 45612 37996 45668
rect 38052 45612 39116 45668
rect 39172 45612 39182 45668
rect 39330 45612 39340 45668
rect 39396 45612 43596 45668
rect 43652 45612 43662 45668
rect 38434 45500 38444 45556
rect 38500 45500 46508 45556
rect 46564 45500 46574 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 32498 45388 32508 45444
rect 32564 45388 33404 45444
rect 33460 45388 33964 45444
rect 34020 45388 34030 45444
rect 40674 45388 40684 45444
rect 40740 45388 47628 45444
rect 47684 45388 48188 45444
rect 48244 45388 48254 45444
rect 25228 45276 31388 45332
rect 31444 45276 31454 45332
rect 31938 45276 31948 45332
rect 32004 45276 34412 45332
rect 34468 45276 34478 45332
rect 25228 45108 25284 45276
rect 18386 45052 18396 45108
rect 18452 45052 21420 45108
rect 21476 45052 21486 45108
rect 23202 45052 23212 45108
rect 23268 45052 25228 45108
rect 25284 45052 25294 45108
rect 25666 45052 25676 45108
rect 25732 45052 26348 45108
rect 26404 45052 27020 45108
rect 27076 45052 27086 45108
rect 31714 45052 31724 45108
rect 31780 45052 32284 45108
rect 32340 45052 32620 45108
rect 32676 45052 33740 45108
rect 33796 45052 33806 45108
rect 38612 45052 41020 45108
rect 41076 45052 41086 45108
rect 38612 44996 38668 45052
rect 16706 44940 16716 44996
rect 16772 44940 18172 44996
rect 18228 44940 19068 44996
rect 19124 44940 19134 44996
rect 24546 44940 24556 44996
rect 24612 44940 25564 44996
rect 25620 44940 25630 44996
rect 28466 44940 28476 44996
rect 28532 44940 31052 44996
rect 31108 44940 31118 44996
rect 33394 44940 33404 44996
rect 33460 44940 34636 44996
rect 34692 44940 34702 44996
rect 37202 44940 37212 44996
rect 37268 44940 38668 44996
rect 41682 44940 41692 44996
rect 41748 44940 42924 44996
rect 42980 44940 42990 44996
rect 43698 44940 43708 44996
rect 43764 44940 47628 44996
rect 47684 44940 47694 44996
rect 39666 44828 39676 44884
rect 39732 44828 40908 44884
rect 40964 44828 40974 44884
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 10434 44492 10444 44548
rect 10500 44492 10510 44548
rect 14578 44492 14588 44548
rect 14644 44492 16156 44548
rect 16212 44492 16222 44548
rect 31154 44492 31164 44548
rect 31220 44492 32284 44548
rect 32340 44492 33964 44548
rect 34020 44492 34030 44548
rect 34178 44492 34188 44548
rect 34244 44492 35532 44548
rect 35588 44492 35598 44548
rect 41570 44492 41580 44548
rect 41636 44492 43820 44548
rect 43876 44492 43886 44548
rect 10444 44436 10500 44492
rect 7634 44380 7644 44436
rect 7700 44380 11564 44436
rect 11620 44380 12012 44436
rect 12068 44380 12078 44436
rect 17378 44380 17388 44436
rect 17444 44380 17836 44436
rect 17892 44380 22540 44436
rect 22596 44380 22606 44436
rect 30930 44380 30940 44436
rect 30996 44380 33292 44436
rect 33348 44380 33358 44436
rect 15810 44268 15820 44324
rect 15876 44268 17276 44324
rect 17332 44268 17342 44324
rect 31938 44268 31948 44324
rect 32004 44268 33628 44324
rect 33684 44268 33694 44324
rect 36978 44268 36988 44324
rect 37044 44268 38556 44324
rect 38612 44268 38622 44324
rect 39890 44268 39900 44324
rect 39956 44268 41020 44324
rect 41076 44268 41468 44324
rect 41524 44268 44828 44324
rect 44884 44268 44894 44324
rect 10770 44156 10780 44212
rect 10836 44156 11452 44212
rect 11508 44156 11518 44212
rect 15026 44156 15036 44212
rect 15092 44156 16604 44212
rect 16660 44156 16670 44212
rect 17042 44156 17052 44212
rect 17108 44156 19516 44212
rect 19572 44156 19582 44212
rect 20290 44156 20300 44212
rect 20356 44156 20860 44212
rect 20916 44156 24556 44212
rect 24612 44156 24622 44212
rect 11330 44044 11340 44100
rect 11396 44044 14364 44100
rect 14420 44044 15820 44100
rect 15876 44044 15886 44100
rect 16034 44044 16044 44100
rect 16100 44044 16940 44100
rect 16996 44044 17006 44100
rect 47058 44044 47068 44100
rect 47124 44044 48188 44100
rect 48244 44044 48254 44100
rect 37426 43932 37436 43988
rect 37492 43932 39676 43988
rect 39732 43932 39742 43988
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 38612 43820 39060 43876
rect 39778 43820 39788 43876
rect 39844 43820 40348 43876
rect 40404 43820 42028 43876
rect 42084 43820 42094 43876
rect 38612 43764 38668 43820
rect 11666 43708 11676 43764
rect 11732 43652 11788 43764
rect 15250 43708 15260 43764
rect 15316 43708 16044 43764
rect 16100 43708 16110 43764
rect 19394 43708 19404 43764
rect 19460 43708 21420 43764
rect 21476 43708 21486 43764
rect 33618 43708 33628 43764
rect 33684 43708 35644 43764
rect 35700 43708 36652 43764
rect 36708 43708 36718 43764
rect 37202 43708 37212 43764
rect 37268 43708 38220 43764
rect 38276 43708 38668 43764
rect 39004 43652 39060 43820
rect 39218 43708 39228 43764
rect 39284 43708 40460 43764
rect 40516 43708 40526 43764
rect 9874 43596 9884 43652
rect 9940 43596 10892 43652
rect 10948 43596 10958 43652
rect 11732 43596 13580 43652
rect 13636 43596 13646 43652
rect 16594 43596 16604 43652
rect 16660 43596 16940 43652
rect 16996 43596 17836 43652
rect 17892 43596 17902 43652
rect 24322 43596 24332 43652
rect 24388 43596 27132 43652
rect 27188 43596 28476 43652
rect 28532 43596 28542 43652
rect 30258 43596 30268 43652
rect 30324 43596 31276 43652
rect 31332 43596 31342 43652
rect 38108 43596 38556 43652
rect 38612 43596 38622 43652
rect 38994 43596 39004 43652
rect 39060 43596 39070 43652
rect 40114 43596 40124 43652
rect 40180 43596 42476 43652
rect 42532 43596 42542 43652
rect 44818 43596 44828 43652
rect 44884 43596 46508 43652
rect 46564 43596 46574 43652
rect 38108 43540 38164 43596
rect 9762 43484 9772 43540
rect 9828 43484 11900 43540
rect 11956 43484 11966 43540
rect 16706 43484 16716 43540
rect 16772 43484 17500 43540
rect 17556 43484 17566 43540
rect 25666 43484 25676 43540
rect 25732 43484 26348 43540
rect 26404 43484 26414 43540
rect 30594 43484 30604 43540
rect 30660 43484 31164 43540
rect 31220 43484 33404 43540
rect 33460 43484 33470 43540
rect 34738 43484 34748 43540
rect 34804 43484 37100 43540
rect 37156 43484 38108 43540
rect 38164 43484 38174 43540
rect 38434 43484 38444 43540
rect 38500 43484 38668 43540
rect 26348 43428 26404 43484
rect 38612 43428 38668 43484
rect 40124 43428 40180 43596
rect 43652 43484 45724 43540
rect 45780 43484 45790 43540
rect 43652 43428 43708 43484
rect 6626 43372 6636 43428
rect 6692 43372 10444 43428
rect 10500 43372 10510 43428
rect 10994 43372 11004 43428
rect 11060 43372 11564 43428
rect 11620 43372 12236 43428
rect 12292 43372 12302 43428
rect 12562 43372 12572 43428
rect 12628 43372 20076 43428
rect 20132 43372 20142 43428
rect 20626 43372 20636 43428
rect 20692 43372 24220 43428
rect 24276 43372 24286 43428
rect 26348 43372 29596 43428
rect 29652 43372 29662 43428
rect 38612 43372 40180 43428
rect 42578 43372 42588 43428
rect 42644 43372 43372 43428
rect 43428 43372 43708 43428
rect 10770 43260 10780 43316
rect 10836 43260 12348 43316
rect 12404 43260 12414 43316
rect 12572 43204 12628 43372
rect 14130 43260 14140 43316
rect 14196 43260 22316 43316
rect 22372 43260 22382 43316
rect 24322 43260 24332 43316
rect 24388 43260 24780 43316
rect 24836 43260 25788 43316
rect 25844 43260 25854 43316
rect 29698 43260 29708 43316
rect 29764 43260 30604 43316
rect 30660 43260 31388 43316
rect 31444 43260 33068 43316
rect 33124 43260 33134 43316
rect 34514 43260 34524 43316
rect 34580 43260 35420 43316
rect 35476 43260 35486 43316
rect 40002 43260 40012 43316
rect 40068 43260 40908 43316
rect 40964 43260 40974 43316
rect 8866 43148 8876 43204
rect 8932 43148 9548 43204
rect 9604 43148 12628 43204
rect 24098 43148 24108 43204
rect 24164 43148 25452 43204
rect 25508 43148 25518 43204
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 10546 43036 10556 43092
rect 10612 43036 11788 43092
rect 11844 43036 11854 43092
rect 12114 43036 12124 43092
rect 12180 43036 23548 43092
rect 23604 43036 23614 43092
rect 40226 43036 40236 43092
rect 40292 43036 40572 43092
rect 40628 43036 40638 43092
rect 45602 43036 45612 43092
rect 45668 43036 46956 43092
rect 47012 43036 47740 43092
rect 47796 43036 47806 43092
rect 21634 42924 21644 42980
rect 21700 42924 24556 42980
rect 24612 42924 24622 42980
rect 37874 42924 37884 42980
rect 37940 42924 39788 42980
rect 39844 42924 42252 42980
rect 42308 42924 46844 42980
rect 46900 42924 47516 42980
rect 47572 42924 47582 42980
rect 20290 42812 20300 42868
rect 20356 42812 21308 42868
rect 21364 42812 22204 42868
rect 22260 42812 22270 42868
rect 23874 42812 23884 42868
rect 23940 42812 24892 42868
rect 24948 42812 24958 42868
rect 28466 42812 28476 42868
rect 28532 42812 39004 42868
rect 39060 42812 39070 42868
rect 18162 42700 18172 42756
rect 18228 42700 20188 42756
rect 20244 42700 20254 42756
rect 23986 42700 23996 42756
rect 24052 42700 24668 42756
rect 24724 42700 24734 42756
rect 29474 42700 29484 42756
rect 29540 42700 30380 42756
rect 30436 42700 30446 42756
rect 33618 42700 33628 42756
rect 33684 42700 36540 42756
rect 36596 42700 36606 42756
rect 40562 42700 40572 42756
rect 40628 42700 41356 42756
rect 41412 42700 41422 42756
rect 45714 42700 45724 42756
rect 45780 42700 46396 42756
rect 46452 42700 46462 42756
rect 46722 42700 46732 42756
rect 46788 42700 47740 42756
rect 47796 42700 47806 42756
rect 16706 42588 16716 42644
rect 16772 42588 17612 42644
rect 17668 42588 17678 42644
rect 20066 42588 20076 42644
rect 20132 42588 22092 42644
rect 22148 42588 22158 42644
rect 23538 42588 23548 42644
rect 23604 42588 24556 42644
rect 24612 42588 24622 42644
rect 26450 42588 26460 42644
rect 26516 42588 30044 42644
rect 30100 42588 30110 42644
rect 39890 42588 39900 42644
rect 39956 42588 42140 42644
rect 42196 42588 42206 42644
rect 44930 42588 44940 42644
rect 44996 42588 45612 42644
rect 45668 42588 45678 42644
rect 18498 42476 18508 42532
rect 18564 42476 25004 42532
rect 25060 42476 25070 42532
rect 40226 42476 40236 42532
rect 40292 42476 40684 42532
rect 40740 42476 40750 42532
rect 46274 42476 46284 42532
rect 46340 42476 47852 42532
rect 47908 42476 47918 42532
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 12674 42252 12684 42308
rect 12740 42252 13804 42308
rect 13860 42252 13870 42308
rect 33394 42252 33404 42308
rect 33460 42252 33964 42308
rect 34020 42252 36652 42308
rect 36708 42252 37548 42308
rect 37604 42252 37614 42308
rect 49200 42196 50000 42224
rect 17154 42140 17164 42196
rect 17220 42140 18396 42196
rect 18452 42140 19404 42196
rect 19460 42140 19470 42196
rect 24658 42140 24668 42196
rect 24724 42140 26684 42196
rect 26740 42140 26750 42196
rect 47282 42140 47292 42196
rect 47348 42140 50000 42196
rect 49200 42112 50000 42140
rect 6850 42028 6860 42084
rect 6916 42028 10780 42084
rect 10836 42028 10846 42084
rect 16034 42028 16044 42084
rect 16100 42028 16716 42084
rect 16772 42028 18732 42084
rect 18788 42028 18798 42084
rect 24546 42028 24556 42084
rect 24612 42028 25564 42084
rect 25620 42028 25630 42084
rect 31938 42028 31948 42084
rect 32004 42028 32396 42084
rect 32452 42028 33964 42084
rect 34020 42028 38668 42084
rect 45490 42028 45500 42084
rect 45556 42028 46396 42084
rect 46452 42028 46956 42084
rect 47012 42028 47022 42084
rect 38612 41972 38668 42028
rect 10322 41916 10332 41972
rect 10388 41916 10892 41972
rect 10948 41916 11676 41972
rect 11732 41916 11742 41972
rect 14130 41916 14140 41972
rect 14196 41916 15372 41972
rect 15428 41916 15438 41972
rect 18946 41916 18956 41972
rect 19012 41916 21084 41972
rect 21140 41916 21150 41972
rect 25778 41916 25788 41972
rect 25844 41916 27244 41972
rect 27300 41916 27310 41972
rect 29138 41916 29148 41972
rect 29204 41916 30492 41972
rect 30548 41916 30558 41972
rect 38612 41916 38892 41972
rect 38948 41916 38958 41972
rect 10434 41804 10444 41860
rect 10500 41804 11228 41860
rect 11284 41804 12012 41860
rect 12068 41804 12460 41860
rect 12516 41804 12526 41860
rect 13122 41804 13132 41860
rect 13188 41804 17836 41860
rect 17892 41804 17902 41860
rect 28018 41804 28028 41860
rect 28084 41804 32732 41860
rect 32788 41804 32798 41860
rect 38612 41804 39900 41860
rect 39956 41804 40124 41860
rect 40180 41804 40190 41860
rect 40562 41804 40572 41860
rect 40628 41804 43484 41860
rect 43540 41804 43550 41860
rect 38612 41748 38668 41804
rect 11106 41692 11116 41748
rect 11172 41692 11788 41748
rect 11844 41692 11854 41748
rect 26674 41692 26684 41748
rect 26740 41692 27692 41748
rect 27748 41692 27758 41748
rect 31276 41692 36988 41748
rect 37044 41692 38668 41748
rect 40338 41692 40348 41748
rect 40404 41692 41020 41748
rect 41076 41692 41086 41748
rect 41682 41692 41692 41748
rect 41748 41692 42364 41748
rect 42420 41692 42430 41748
rect 31276 41636 31332 41692
rect 8978 41580 8988 41636
rect 9044 41580 9884 41636
rect 9940 41580 11900 41636
rect 11956 41580 20524 41636
rect 20580 41580 20590 41636
rect 26450 41580 26460 41636
rect 26516 41580 29932 41636
rect 29988 41580 31276 41636
rect 31332 41580 31342 41636
rect 39442 41580 39452 41636
rect 39508 41580 40012 41636
rect 40068 41580 40908 41636
rect 40964 41580 40974 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 18050 41356 18060 41412
rect 18116 41356 19852 41412
rect 19908 41356 19918 41412
rect 4610 41244 4620 41300
rect 4676 41244 6076 41300
rect 6132 41244 6142 41300
rect 13682 41244 13692 41300
rect 13748 41244 14476 41300
rect 14532 41244 14542 41300
rect 20626 41244 20636 41300
rect 20692 41244 22764 41300
rect 22820 41244 22830 41300
rect 40226 41244 40236 41300
rect 40292 41244 40908 41300
rect 40964 41244 40974 41300
rect 10322 41132 10332 41188
rect 10388 41132 13580 41188
rect 13636 41132 13646 41188
rect 12898 41020 12908 41076
rect 12964 41020 13468 41076
rect 13524 41020 13534 41076
rect 13804 40964 13860 41244
rect 17826 41132 17836 41188
rect 17892 41132 19516 41188
rect 19572 41132 21420 41188
rect 21476 41132 21486 41188
rect 33730 41132 33740 41188
rect 33796 41132 34300 41188
rect 34356 41132 34366 41188
rect 36530 41132 36540 41188
rect 36596 41132 37324 41188
rect 37380 41132 37390 41188
rect 44258 41132 44268 41188
rect 44324 41132 47964 41188
rect 48020 41132 48030 41188
rect 21746 41020 21756 41076
rect 21812 41020 23996 41076
rect 24052 41020 24062 41076
rect 26786 41020 26796 41076
rect 26852 41020 29372 41076
rect 29428 41020 29438 41076
rect 32732 41020 33404 41076
rect 33460 41020 33470 41076
rect 33842 41020 33852 41076
rect 33908 41020 34636 41076
rect 34692 41020 35532 41076
rect 35588 41020 35598 41076
rect 32732 40964 32788 41020
rect 11330 40908 11340 40964
rect 11396 40908 13132 40964
rect 13188 40908 13198 40964
rect 13570 40908 13580 40964
rect 13636 40908 13860 40964
rect 17938 40908 17948 40964
rect 18004 40908 19068 40964
rect 19124 40908 19134 40964
rect 29698 40908 29708 40964
rect 29764 40908 30604 40964
rect 30660 40908 30670 40964
rect 31378 40908 31388 40964
rect 31444 40908 32060 40964
rect 32116 40908 32508 40964
rect 32564 40908 32574 40964
rect 32722 40908 32732 40964
rect 32788 40908 32798 40964
rect 39666 40908 39676 40964
rect 39732 40908 40572 40964
rect 40628 40908 40638 40964
rect 38658 40796 38668 40852
rect 38724 40796 45948 40852
rect 46004 40796 46014 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 20514 40684 20524 40740
rect 20580 40684 21420 40740
rect 21476 40684 21486 40740
rect 22754 40684 22764 40740
rect 22820 40684 25900 40740
rect 25956 40684 25966 40740
rect 30482 40684 30492 40740
rect 30548 40684 31444 40740
rect 12338 40572 12348 40628
rect 12404 40572 13132 40628
rect 13188 40572 20188 40628
rect 20244 40572 20254 40628
rect 24434 40572 24444 40628
rect 24500 40572 25452 40628
rect 25508 40572 31220 40628
rect 14130 40460 14140 40516
rect 14196 40460 14476 40516
rect 14532 40460 15148 40516
rect 15922 40460 15932 40516
rect 15988 40460 16044 40516
rect 16100 40460 16604 40516
rect 16660 40460 16670 40516
rect 24770 40460 24780 40516
rect 24836 40460 25564 40516
rect 25620 40460 25630 40516
rect 28018 40460 28028 40516
rect 28084 40460 28364 40516
rect 28420 40460 28924 40516
rect 28980 40460 28990 40516
rect 15092 40404 15148 40460
rect 31164 40404 31220 40572
rect 31388 40516 31444 40684
rect 32386 40572 32396 40628
rect 32452 40572 33740 40628
rect 33796 40572 33806 40628
rect 40338 40572 40348 40628
rect 40404 40572 43708 40628
rect 31378 40460 31388 40516
rect 31444 40460 31454 40516
rect 34402 40460 34412 40516
rect 34468 40460 34972 40516
rect 35028 40460 35038 40516
rect 39890 40460 39900 40516
rect 39956 40460 40684 40516
rect 40740 40460 41468 40516
rect 41524 40460 41534 40516
rect 43652 40404 43708 40572
rect 46498 40460 46508 40516
rect 46564 40460 47964 40516
rect 48020 40460 48030 40516
rect 15092 40348 15708 40404
rect 15764 40348 21532 40404
rect 21588 40348 21598 40404
rect 21756 40348 24220 40404
rect 24276 40348 24286 40404
rect 26114 40348 26124 40404
rect 26180 40348 26684 40404
rect 26740 40348 27804 40404
rect 27860 40348 28476 40404
rect 28532 40348 28542 40404
rect 30482 40348 30492 40404
rect 30548 40348 30716 40404
rect 30772 40348 30782 40404
rect 31154 40348 31164 40404
rect 31220 40348 31230 40404
rect 31490 40348 31500 40404
rect 31556 40348 33628 40404
rect 33684 40348 33694 40404
rect 38882 40348 38892 40404
rect 38948 40348 41916 40404
rect 41972 40348 42588 40404
rect 42644 40348 43036 40404
rect 43092 40348 43102 40404
rect 43652 40348 44604 40404
rect 44660 40348 44670 40404
rect 21756 40292 21812 40348
rect 10882 40236 10892 40292
rect 10948 40236 14140 40292
rect 14196 40236 14206 40292
rect 20738 40236 20748 40292
rect 20804 40236 21812 40292
rect 28914 40236 28924 40292
rect 28980 40236 31948 40292
rect 32004 40236 32014 40292
rect 21186 40124 21196 40180
rect 21252 40124 21644 40180
rect 21700 40124 21710 40180
rect 29138 40124 29148 40180
rect 29204 40124 31276 40180
rect 31332 40124 31342 40180
rect 31490 40124 31500 40180
rect 31556 40124 31836 40180
rect 31892 40124 31902 40180
rect 45714 40124 45724 40180
rect 45780 40124 46620 40180
rect 46676 40124 46686 40180
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 18722 39788 18732 39844
rect 18788 39788 19516 39844
rect 19572 39788 26908 39844
rect 26964 39788 28252 39844
rect 28308 39788 28318 39844
rect 30258 39788 30268 39844
rect 30324 39788 34076 39844
rect 34132 39788 34142 39844
rect 34402 39788 34412 39844
rect 34468 39788 34478 39844
rect 34626 39788 34636 39844
rect 34692 39788 36316 39844
rect 36372 39788 36382 39844
rect 44930 39788 44940 39844
rect 44996 39788 47740 39844
rect 47796 39788 47806 39844
rect 34412 39732 34468 39788
rect 34412 39676 35420 39732
rect 35476 39676 35486 39732
rect 36082 39676 36092 39732
rect 36148 39676 37324 39732
rect 37380 39676 37390 39732
rect 18834 39564 18844 39620
rect 18900 39564 19740 39620
rect 19796 39564 20076 39620
rect 20132 39564 20142 39620
rect 29250 39564 29260 39620
rect 29316 39564 30044 39620
rect 30100 39564 30110 39620
rect 30454 39564 30492 39620
rect 30548 39564 30558 39620
rect 31042 39564 31052 39620
rect 31108 39564 35308 39620
rect 35364 39564 35374 39620
rect 35634 39564 35644 39620
rect 35700 39564 37100 39620
rect 37156 39564 37166 39620
rect 1698 39452 1708 39508
rect 1764 39452 3388 39508
rect 3444 39452 4060 39508
rect 4116 39452 4126 39508
rect 7522 39452 7532 39508
rect 7588 39452 10108 39508
rect 10164 39452 10174 39508
rect 18274 39452 18284 39508
rect 18340 39452 18620 39508
rect 18676 39452 19628 39508
rect 19684 39452 19694 39508
rect 21074 39452 21084 39508
rect 21140 39452 27356 39508
rect 27412 39452 27422 39508
rect 29138 39452 29148 39508
rect 29204 39452 29708 39508
rect 29764 39452 29774 39508
rect 34850 39452 34860 39508
rect 34916 39452 35756 39508
rect 35812 39452 35822 39508
rect 39778 39452 39788 39508
rect 39844 39452 42476 39508
rect 42532 39452 42542 39508
rect 47058 39452 47068 39508
rect 47124 39452 47162 39508
rect 3042 39340 3052 39396
rect 3108 39340 4508 39396
rect 4564 39340 4574 39396
rect 8530 39340 8540 39396
rect 8596 39340 9996 39396
rect 10052 39340 10062 39396
rect 12898 39340 12908 39396
rect 12964 39340 15372 39396
rect 15428 39340 15438 39396
rect 18162 39340 18172 39396
rect 18228 39340 19852 39396
rect 19908 39340 19918 39396
rect 26226 39340 26236 39396
rect 26292 39340 26684 39396
rect 26740 39340 26750 39396
rect 32386 39340 32396 39396
rect 32452 39340 34972 39396
rect 35028 39340 35038 39396
rect 35410 39340 35420 39396
rect 35476 39340 36092 39396
rect 36148 39340 36158 39396
rect 42354 39340 42364 39396
rect 42420 39340 43484 39396
rect 43540 39340 43550 39396
rect 44370 39340 44380 39396
rect 44436 39340 46396 39396
rect 46452 39340 46462 39396
rect 3938 39228 3948 39284
rect 4004 39228 4620 39284
rect 4676 39228 4686 39284
rect 18386 39228 18396 39284
rect 18452 39228 18844 39284
rect 18900 39228 18910 39284
rect 38434 39228 38444 39284
rect 38500 39228 46732 39284
rect 46788 39228 46798 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 18946 39116 18956 39172
rect 19012 39116 19516 39172
rect 19572 39116 19582 39172
rect 21746 39116 21756 39172
rect 21812 39116 22540 39172
rect 22596 39116 22606 39172
rect 34178 39116 34188 39172
rect 34244 39116 35084 39172
rect 35140 39116 37212 39172
rect 37268 39116 37278 39172
rect 43810 39116 43820 39172
rect 43876 39116 48188 39172
rect 48244 39116 48254 39172
rect 8372 39004 8540 39060
rect 8596 39004 8606 39060
rect 10434 39004 10444 39060
rect 10500 39004 11004 39060
rect 11060 39004 11564 39060
rect 11620 39004 14084 39060
rect 15362 39004 15372 39060
rect 15428 39004 19852 39060
rect 19908 39004 22316 39060
rect 22372 39004 22382 39060
rect 24434 39004 24444 39060
rect 24500 39004 25340 39060
rect 25396 39004 32620 39060
rect 32676 39004 34076 39060
rect 34132 39004 34142 39060
rect 42130 39004 42140 39060
rect 42196 39004 43148 39060
rect 43204 39004 43214 39060
rect 45266 39004 45276 39060
rect 45332 39004 45836 39060
rect 45892 39004 46844 39060
rect 46900 39004 46910 39060
rect 8372 38948 8428 39004
rect 14028 38948 14084 39004
rect 6066 38892 6076 38948
rect 6132 38892 8428 38948
rect 9762 38892 9772 38948
rect 9828 38892 10332 38948
rect 10388 38892 10398 38948
rect 13122 38892 13132 38948
rect 13188 38892 13804 38948
rect 13860 38892 13870 38948
rect 14028 38892 32004 38948
rect 32162 38892 32172 38948
rect 32228 38892 36988 38948
rect 37044 38892 42700 38948
rect 42756 38892 42766 38948
rect 44930 38892 44940 38948
rect 44996 38892 46620 38948
rect 46676 38892 47068 38948
rect 47124 38892 47134 38948
rect 47730 38892 47740 38948
rect 47796 38892 47806 38948
rect 31948 38836 32004 38892
rect 2818 38780 2828 38836
rect 2884 38780 3388 38836
rect 3444 38780 3454 38836
rect 13570 38780 13580 38836
rect 13636 38780 14364 38836
rect 14420 38780 15932 38836
rect 15988 38780 15998 38836
rect 20066 38780 20076 38836
rect 20132 38780 21308 38836
rect 21364 38780 21374 38836
rect 22194 38780 22204 38836
rect 22260 38780 23212 38836
rect 23268 38780 23278 38836
rect 25778 38780 25788 38836
rect 25844 38780 26236 38836
rect 26292 38780 26302 38836
rect 26460 38780 29148 38836
rect 29204 38780 29214 38836
rect 30370 38780 30380 38836
rect 30436 38780 31612 38836
rect 31668 38780 31678 38836
rect 31938 38780 31948 38836
rect 32004 38780 33292 38836
rect 33348 38780 33358 38836
rect 33730 38780 33740 38836
rect 33796 38780 37996 38836
rect 38052 38780 38062 38836
rect 39778 38780 39788 38836
rect 39844 38780 40460 38836
rect 40516 38780 40526 38836
rect 43698 38780 43708 38836
rect 43764 38780 45724 38836
rect 45780 38780 45790 38836
rect 45938 38780 45948 38836
rect 46004 38780 46956 38836
rect 47012 38780 47404 38836
rect 47460 38780 47470 38836
rect 26460 38724 26516 38780
rect 2706 38668 2716 38724
rect 2772 38668 3836 38724
rect 3892 38668 3902 38724
rect 10770 38668 10780 38724
rect 10836 38668 11676 38724
rect 11732 38668 11742 38724
rect 12674 38668 12684 38724
rect 12740 38668 14252 38724
rect 14308 38668 14318 38724
rect 17826 38668 17836 38724
rect 17892 38668 21196 38724
rect 21252 38668 21262 38724
rect 23986 38668 23996 38724
rect 24052 38668 25340 38724
rect 25396 38668 25406 38724
rect 26114 38668 26124 38724
rect 26180 38668 26516 38724
rect 36418 38668 36428 38724
rect 36484 38668 38108 38724
rect 38164 38668 38174 38724
rect 46162 38668 46172 38724
rect 46228 38668 47292 38724
rect 47348 38668 47358 38724
rect 10546 38556 10556 38612
rect 10612 38556 11340 38612
rect 11396 38556 11406 38612
rect 18834 38556 18844 38612
rect 18900 38556 19628 38612
rect 19684 38556 20076 38612
rect 20132 38556 20142 38612
rect 28578 38556 28588 38612
rect 28644 38556 29596 38612
rect 29652 38556 29662 38612
rect 34290 38556 34300 38612
rect 34356 38556 35084 38612
rect 35140 38556 35150 38612
rect 41906 38556 41916 38612
rect 41972 38556 43036 38612
rect 43092 38556 43102 38612
rect 47740 38500 47796 38892
rect 16818 38444 16828 38500
rect 16884 38444 19404 38500
rect 19460 38444 21084 38500
rect 21140 38444 21150 38500
rect 21410 38444 21420 38500
rect 21476 38444 25676 38500
rect 25732 38444 25742 38500
rect 39778 38444 39788 38500
rect 39844 38444 40124 38500
rect 40180 38444 40190 38500
rect 47730 38444 47740 38500
rect 47796 38444 47806 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 16482 38332 16492 38388
rect 16548 38332 20300 38388
rect 20356 38332 20366 38388
rect 40226 38332 40236 38388
rect 40292 38332 41580 38388
rect 41636 38332 43148 38388
rect 43204 38332 45612 38388
rect 45668 38332 45678 38388
rect 16706 38220 16716 38276
rect 16772 38220 19404 38276
rect 19460 38220 19470 38276
rect 44146 38220 44156 38276
rect 44212 38220 47404 38276
rect 47460 38220 47470 38276
rect 7298 38108 7308 38164
rect 7364 38108 9884 38164
rect 9940 38108 11900 38164
rect 11956 38108 11966 38164
rect 12450 38108 12460 38164
rect 12516 38108 32172 38164
rect 32228 38108 32732 38164
rect 32788 38108 32798 38164
rect 36418 38108 36428 38164
rect 36484 38108 37436 38164
rect 37492 38108 37502 38164
rect 43138 38108 43148 38164
rect 43204 38108 43932 38164
rect 43988 38108 43998 38164
rect 1698 37996 1708 38052
rect 1764 37996 3836 38052
rect 3892 37996 3902 38052
rect 8082 37996 8092 38052
rect 8148 37996 8764 38052
rect 8820 37996 8830 38052
rect 12226 37996 12236 38052
rect 12292 37996 13692 38052
rect 13748 37996 13758 38052
rect 18834 37996 18844 38052
rect 18900 37996 19740 38052
rect 19796 37996 19806 38052
rect 24770 37996 24780 38052
rect 24836 37996 26572 38052
rect 26628 37996 26638 38052
rect 29586 37996 29596 38052
rect 29652 37996 30380 38052
rect 30436 37996 30446 38052
rect 33618 37996 33628 38052
rect 33684 37996 36204 38052
rect 36260 37996 36540 38052
rect 36596 37996 37100 38052
rect 37156 37996 37166 38052
rect 38098 37996 38108 38052
rect 38164 37996 40124 38052
rect 40180 37996 40190 38052
rect 40338 37996 40348 38052
rect 40404 37996 41916 38052
rect 41972 37996 41982 38052
rect 44930 37996 44940 38052
rect 44996 37996 45724 38052
rect 45780 37996 45790 38052
rect 7858 37884 7868 37940
rect 7924 37884 8428 37940
rect 8484 37884 9772 37940
rect 9828 37884 10332 37940
rect 10388 37884 10398 37940
rect 15138 37884 15148 37940
rect 15204 37884 19292 37940
rect 19348 37884 19358 37940
rect 30258 37884 30268 37940
rect 30324 37884 31388 37940
rect 31444 37884 31454 37940
rect 44146 37884 44156 37940
rect 44212 37884 45164 37940
rect 45220 37884 45230 37940
rect 45826 37884 45836 37940
rect 45892 37884 46396 37940
rect 46452 37884 46462 37940
rect 2594 37772 2604 37828
rect 2660 37772 3276 37828
rect 3332 37772 6076 37828
rect 6132 37772 6972 37828
rect 7028 37772 7038 37828
rect 18050 37772 18060 37828
rect 18116 37772 18396 37828
rect 18452 37772 19628 37828
rect 19684 37772 19694 37828
rect 43810 37772 43820 37828
rect 43876 37772 45052 37828
rect 45108 37772 45118 37828
rect 27234 37660 27244 37716
rect 27300 37660 27804 37716
rect 27860 37660 28588 37716
rect 28644 37660 38780 37716
rect 38836 37660 38846 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 27010 37548 27020 37604
rect 27076 37548 33740 37604
rect 33796 37548 35644 37604
rect 35700 37548 35710 37604
rect 17826 37436 17836 37492
rect 17892 37436 18620 37492
rect 18676 37436 18686 37492
rect 29474 37436 29484 37492
rect 29540 37436 34748 37492
rect 34804 37436 36092 37492
rect 36148 37436 38668 37492
rect 40114 37436 40124 37492
rect 40180 37436 41020 37492
rect 41076 37436 41086 37492
rect 45490 37436 45500 37492
rect 45556 37436 46284 37492
rect 46340 37436 47628 37492
rect 47684 37436 47694 37492
rect 8530 37324 8540 37380
rect 8596 37324 9884 37380
rect 9940 37324 9950 37380
rect 11330 37324 11340 37380
rect 11396 37324 23884 37380
rect 23940 37324 23950 37380
rect 35186 37324 35196 37380
rect 35252 37324 36428 37380
rect 36484 37324 36494 37380
rect 38612 37268 38668 37436
rect 43026 37324 43036 37380
rect 43092 37324 43708 37380
rect 43764 37324 43774 37380
rect 49200 37268 50000 37296
rect 5058 37212 5068 37268
rect 5124 37212 6748 37268
rect 6804 37212 9772 37268
rect 9828 37212 9838 37268
rect 16818 37212 16828 37268
rect 16884 37212 18396 37268
rect 18452 37212 19068 37268
rect 19124 37212 31164 37268
rect 31220 37212 31230 37268
rect 33618 37212 33628 37268
rect 33684 37212 34636 37268
rect 34692 37212 34702 37268
rect 38612 37212 41580 37268
rect 41636 37212 41646 37268
rect 47058 37212 47068 37268
rect 47124 37212 47162 37268
rect 47842 37212 47852 37268
rect 47908 37212 48188 37268
rect 48244 37212 48254 37268
rect 48402 37212 48412 37268
rect 48468 37212 50000 37268
rect 49200 37184 50000 37212
rect 13906 37100 13916 37156
rect 13972 37100 18172 37156
rect 18228 37100 18238 37156
rect 20066 37100 20076 37156
rect 20132 37100 21868 37156
rect 21924 37100 21934 37156
rect 30930 37100 30940 37156
rect 30996 37100 32060 37156
rect 32116 37100 32126 37156
rect 33170 37100 33180 37156
rect 33236 37100 33852 37156
rect 33908 37100 33918 37156
rect 35634 37100 35644 37156
rect 35700 37100 38780 37156
rect 38836 37100 38846 37156
rect 40002 37100 40012 37156
rect 40068 37100 40908 37156
rect 40964 37100 40974 37156
rect 21634 36988 21644 37044
rect 21700 36988 22764 37044
rect 22820 36988 22830 37044
rect 22978 36988 22988 37044
rect 23044 36988 23054 37044
rect 26534 36988 26572 37044
rect 26628 36988 26638 37044
rect 33180 36988 33628 37044
rect 33684 36988 33694 37044
rect 40338 36988 40348 37044
rect 40404 36988 41804 37044
rect 41860 36988 41870 37044
rect 22988 36932 23044 36988
rect 33180 36932 33236 36988
rect 17826 36876 17836 36932
rect 17892 36876 18844 36932
rect 18900 36876 18910 36932
rect 22530 36876 22540 36932
rect 22596 36876 23044 36932
rect 33170 36876 33180 36932
rect 33236 36876 33246 36932
rect 33954 36876 33964 36932
rect 34020 36876 34972 36932
rect 35028 36876 35038 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 44258 36652 44268 36708
rect 44324 36652 44334 36708
rect 2930 36540 2940 36596
rect 2996 36540 3836 36596
rect 3892 36540 3902 36596
rect 25666 36540 25676 36596
rect 25732 36540 29260 36596
rect 29316 36540 29820 36596
rect 29876 36540 29886 36596
rect 7298 36428 7308 36484
rect 7364 36428 8204 36484
rect 8260 36428 8270 36484
rect 19170 36428 19180 36484
rect 19236 36428 20524 36484
rect 20580 36428 20590 36484
rect 20850 36428 20860 36484
rect 20916 36428 21532 36484
rect 21588 36428 21598 36484
rect 24546 36428 24556 36484
rect 24612 36428 26908 36484
rect 39890 36428 39900 36484
rect 39956 36428 41132 36484
rect 41188 36428 41198 36484
rect 5730 36316 5740 36372
rect 5796 36316 6860 36372
rect 6916 36316 6926 36372
rect 8204 36260 8260 36428
rect 26852 36372 26908 36428
rect 23202 36316 23212 36372
rect 23268 36316 25564 36372
rect 25620 36316 25630 36372
rect 26852 36316 29708 36372
rect 29764 36316 31556 36372
rect 33058 36316 33068 36372
rect 33124 36316 33516 36372
rect 33572 36316 33582 36372
rect 38546 36316 38556 36372
rect 38612 36316 39788 36372
rect 39844 36316 39854 36372
rect 31500 36260 31556 36316
rect 8204 36204 8876 36260
rect 8932 36204 8942 36260
rect 12002 36204 12012 36260
rect 12068 36204 12572 36260
rect 12628 36204 16604 36260
rect 16660 36204 16670 36260
rect 17826 36204 17836 36260
rect 17892 36204 19964 36260
rect 20020 36204 20030 36260
rect 28242 36204 28252 36260
rect 28308 36204 29596 36260
rect 29652 36204 29662 36260
rect 31490 36204 31500 36260
rect 31556 36204 36428 36260
rect 36484 36204 37100 36260
rect 37156 36204 37166 36260
rect 30678 36092 30716 36148
rect 30772 36092 36092 36148
rect 36148 36092 36158 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 44268 36036 44324 36652
rect 44818 36204 44828 36260
rect 44884 36204 46844 36260
rect 46900 36204 46910 36260
rect 29138 35980 29148 36036
rect 29204 35980 29596 36036
rect 29652 35980 44324 36036
rect 6402 35868 6412 35924
rect 6468 35868 7196 35924
rect 7252 35868 7262 35924
rect 23986 35868 23996 35924
rect 24052 35868 26348 35924
rect 26404 35868 26414 35924
rect 26852 35868 37100 35924
rect 37156 35868 37660 35924
rect 37716 35868 40012 35924
rect 40068 35868 40078 35924
rect 41682 35868 41692 35924
rect 41748 35868 48188 35924
rect 48244 35868 48254 35924
rect 1698 35756 1708 35812
rect 1764 35756 3724 35812
rect 3780 35756 4396 35812
rect 4452 35756 4462 35812
rect 6850 35756 6860 35812
rect 6916 35756 8652 35812
rect 8708 35756 8718 35812
rect 26852 35700 26908 35868
rect 29474 35756 29484 35812
rect 29540 35756 30940 35812
rect 30996 35756 31388 35812
rect 31444 35756 31454 35812
rect 47394 35756 47404 35812
rect 47460 35756 48076 35812
rect 48132 35756 48142 35812
rect 23202 35644 23212 35700
rect 23268 35644 23772 35700
rect 23828 35644 23838 35700
rect 25330 35644 25340 35700
rect 25396 35644 26908 35700
rect 27682 35644 27692 35700
rect 27748 35644 27916 35700
rect 27972 35644 29148 35700
rect 29204 35644 29214 35700
rect 29362 35644 29372 35700
rect 29428 35644 30716 35700
rect 30772 35644 30782 35700
rect 31042 35644 31052 35700
rect 31108 35644 31836 35700
rect 31892 35644 32172 35700
rect 32228 35644 32238 35700
rect 35970 35644 35980 35700
rect 36036 35644 36988 35700
rect 37044 35644 37054 35700
rect 41234 35644 41244 35700
rect 41300 35644 42476 35700
rect 42532 35644 45388 35700
rect 45444 35644 45454 35700
rect 9650 35532 9660 35588
rect 9716 35532 10892 35588
rect 10948 35532 10958 35588
rect 15092 35532 17724 35588
rect 17780 35532 20300 35588
rect 20356 35532 20366 35588
rect 21746 35532 21756 35588
rect 21812 35532 22316 35588
rect 22372 35532 22764 35588
rect 22820 35532 26012 35588
rect 26068 35532 26078 35588
rect 31490 35532 31500 35588
rect 31556 35532 34524 35588
rect 34580 35532 34590 35588
rect 42690 35532 42700 35588
rect 42756 35532 43596 35588
rect 43652 35532 44940 35588
rect 44996 35532 46172 35588
rect 46228 35532 46238 35588
rect 7858 35308 7868 35364
rect 7924 35308 8204 35364
rect 8260 35308 8270 35364
rect 10546 35308 10556 35364
rect 10612 35308 13580 35364
rect 13636 35308 14028 35364
rect 14084 35308 14094 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 7074 35196 7084 35252
rect 7140 35196 9660 35252
rect 9716 35196 9726 35252
rect 10882 35196 10892 35252
rect 10948 35196 13468 35252
rect 13524 35196 13534 35252
rect 15092 35140 15148 35532
rect 26338 35420 26348 35476
rect 26404 35420 26908 35476
rect 30482 35420 30492 35476
rect 30548 35420 32172 35476
rect 32228 35420 32238 35476
rect 37538 35420 37548 35476
rect 37604 35420 39900 35476
rect 39956 35420 39966 35476
rect 40562 35420 40572 35476
rect 40628 35420 41244 35476
rect 41300 35420 42812 35476
rect 42868 35420 45836 35476
rect 45892 35420 46508 35476
rect 46564 35420 46574 35476
rect 26852 35364 26908 35420
rect 17266 35308 17276 35364
rect 17332 35308 26684 35364
rect 26740 35308 26750 35364
rect 26852 35308 30604 35364
rect 30660 35308 31500 35364
rect 31556 35308 31566 35364
rect 31714 35308 31724 35364
rect 31780 35308 32060 35364
rect 32116 35308 33068 35364
rect 33124 35308 33134 35364
rect 43250 35308 43260 35364
rect 43316 35308 44828 35364
rect 44884 35308 44894 35364
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 20738 35196 20748 35252
rect 20804 35196 21532 35252
rect 21588 35196 23548 35252
rect 23604 35196 23614 35252
rect 23762 35196 23772 35252
rect 23828 35196 25452 35252
rect 25508 35196 25518 35252
rect 46386 35196 46396 35252
rect 46452 35196 47516 35252
rect 47572 35196 47582 35252
rect 3490 35084 3500 35140
rect 3556 35084 4732 35140
rect 4788 35084 5404 35140
rect 5460 35084 5470 35140
rect 7746 35084 7756 35140
rect 7812 35084 10780 35140
rect 10836 35084 10846 35140
rect 11666 35084 11676 35140
rect 11732 35084 15148 35140
rect 21970 35084 21980 35140
rect 22036 35084 25004 35140
rect 25060 35084 25070 35140
rect 36306 35084 36316 35140
rect 36372 35084 36988 35140
rect 37044 35084 37054 35140
rect 4396 34972 5628 35028
rect 5684 34972 5694 35028
rect 18386 34972 18396 35028
rect 18452 34972 19964 35028
rect 20020 34972 20030 35028
rect 20290 34972 20300 35028
rect 20356 34972 22204 35028
rect 22260 34972 22270 35028
rect 23538 34972 23548 35028
rect 23604 34972 24668 35028
rect 24724 34972 24734 35028
rect 34178 34972 34188 35028
rect 34244 34972 35420 35028
rect 35476 34972 35486 35028
rect 4396 34916 4452 34972
rect 3266 34860 3276 34916
rect 3332 34860 4396 34916
rect 4452 34860 4462 34916
rect 5058 34860 5068 34916
rect 5124 34860 6636 34916
rect 6692 34860 8764 34916
rect 8820 34860 8830 34916
rect 9986 34860 9996 34916
rect 10052 34860 11452 34916
rect 11508 34860 11518 34916
rect 29446 34860 29484 34916
rect 29540 34860 29550 34916
rect 39778 34860 39788 34916
rect 39844 34860 41132 34916
rect 41188 34860 41198 34916
rect 3276 34804 3332 34860
rect 2930 34748 2940 34804
rect 2996 34748 3332 34804
rect 3602 34748 3612 34804
rect 3668 34748 7756 34804
rect 7812 34748 7822 34804
rect 8194 34748 8204 34804
rect 8260 34748 8876 34804
rect 8932 34748 8942 34804
rect 11218 34748 11228 34804
rect 11284 34748 12124 34804
rect 12180 34748 12460 34804
rect 12516 34748 12526 34804
rect 12786 34748 12796 34804
rect 12852 34748 13804 34804
rect 13860 34748 13870 34804
rect 25778 34748 25788 34804
rect 25844 34748 27972 34804
rect 28578 34748 28588 34804
rect 28644 34748 29932 34804
rect 29988 34748 31836 34804
rect 31892 34748 33068 34804
rect 33124 34748 33134 34804
rect 34514 34748 34524 34804
rect 34580 34748 38332 34804
rect 38388 34748 38668 34804
rect 43362 34748 43372 34804
rect 43428 34748 43596 34804
rect 43652 34748 43662 34804
rect 27916 34692 27972 34748
rect 38612 34692 38668 34748
rect 2370 34636 2380 34692
rect 2436 34636 3276 34692
rect 3332 34636 3500 34692
rect 3556 34636 3566 34692
rect 9090 34636 9100 34692
rect 9156 34636 9884 34692
rect 9940 34636 9950 34692
rect 13906 34636 13916 34692
rect 13972 34636 14700 34692
rect 14756 34636 14766 34692
rect 16482 34636 16492 34692
rect 16548 34636 18620 34692
rect 18676 34636 18686 34692
rect 20850 34636 20860 34692
rect 20916 34636 21980 34692
rect 22036 34636 23436 34692
rect 23492 34636 23502 34692
rect 24182 34636 24220 34692
rect 24276 34636 24286 34692
rect 25666 34636 25676 34692
rect 25732 34636 27468 34692
rect 27524 34636 27534 34692
rect 27906 34636 27916 34692
rect 27972 34636 27982 34692
rect 29362 34636 29372 34692
rect 29428 34636 29708 34692
rect 29764 34636 29774 34692
rect 38612 34636 38892 34692
rect 38948 34636 38958 34692
rect 43138 34636 43148 34692
rect 43204 34636 43708 34692
rect 43764 34636 44268 34692
rect 44324 34636 44334 34692
rect 31154 34524 31164 34580
rect 31220 34524 39228 34580
rect 39284 34524 39294 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4610 34412 4620 34468
rect 4676 34412 5964 34468
rect 6020 34412 7756 34468
rect 7812 34412 7822 34468
rect 36082 34412 36092 34468
rect 36148 34412 38220 34468
rect 38276 34412 44044 34468
rect 44100 34412 44110 34468
rect 13234 34300 13244 34356
rect 13300 34300 13692 34356
rect 13748 34300 14364 34356
rect 14420 34300 14430 34356
rect 23090 34300 23100 34356
rect 23156 34300 23996 34356
rect 24052 34300 24062 34356
rect 34066 34300 34076 34356
rect 34132 34300 36652 34356
rect 36708 34300 36718 34356
rect 38994 34300 39004 34356
rect 39060 34300 42476 34356
rect 42532 34300 42542 34356
rect 5954 34188 5964 34244
rect 6020 34188 6860 34244
rect 6916 34188 6926 34244
rect 13458 34188 13468 34244
rect 13524 34188 14140 34244
rect 14196 34188 18788 34244
rect 23762 34188 23772 34244
rect 23828 34188 25900 34244
rect 25956 34188 25966 34244
rect 38210 34188 38220 34244
rect 38276 34188 40012 34244
rect 40068 34188 40908 34244
rect 40964 34188 40974 34244
rect 46610 34188 46620 34244
rect 46676 34188 48076 34244
rect 48132 34188 48142 34244
rect 18732 34132 18788 34188
rect 18162 34076 18172 34132
rect 18228 34076 18508 34132
rect 18564 34076 18574 34132
rect 18722 34076 18732 34132
rect 18788 34076 19516 34132
rect 19572 34076 19582 34132
rect 29026 34076 29036 34132
rect 29092 34076 29932 34132
rect 29988 34076 29998 34132
rect 36754 34076 36764 34132
rect 36820 34076 42140 34132
rect 42196 34076 43932 34132
rect 43988 34076 43998 34132
rect 18508 34020 18564 34076
rect 11218 33964 11228 34020
rect 11284 33964 13356 34020
rect 13412 33964 13422 34020
rect 14690 33964 14700 34020
rect 14756 33964 15036 34020
rect 15092 33964 18060 34020
rect 18116 33964 18126 34020
rect 18508 33964 19180 34020
rect 19236 33964 19246 34020
rect 33842 33964 33852 34020
rect 33908 33964 36540 34020
rect 36596 33964 36606 34020
rect 39778 33964 39788 34020
rect 39844 33964 41020 34020
rect 41076 33964 41086 34020
rect 9874 33852 9884 33908
rect 9940 33852 12684 33908
rect 12740 33852 12750 33908
rect 14802 33852 14812 33908
rect 14868 33852 16436 33908
rect 17714 33852 17724 33908
rect 17780 33852 18284 33908
rect 18340 33852 18350 33908
rect 18946 33852 18956 33908
rect 19012 33852 20412 33908
rect 20468 33852 20478 33908
rect 24210 33852 24220 33908
rect 24276 33852 24332 33908
rect 24388 33852 24398 33908
rect 32162 33852 32172 33908
rect 32228 33852 36428 33908
rect 36484 33852 38220 33908
rect 38276 33852 38286 33908
rect 12450 33740 12460 33796
rect 12516 33740 16156 33796
rect 16212 33740 16222 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 16380 33684 16436 33852
rect 18498 33740 18508 33796
rect 18564 33740 19068 33796
rect 19124 33740 19134 33796
rect 23202 33740 23212 33796
rect 23268 33740 24892 33796
rect 24948 33740 24958 33796
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 16380 33628 19404 33684
rect 19460 33628 20076 33684
rect 20132 33628 20860 33684
rect 20916 33628 20926 33684
rect 24994 33628 25004 33684
rect 25060 33628 26796 33684
rect 26852 33628 26862 33684
rect 41570 33628 41580 33684
rect 41636 33628 42924 33684
rect 42980 33628 42990 33684
rect 14578 33516 14588 33572
rect 14644 33516 15708 33572
rect 15764 33516 15774 33572
rect 21858 33516 21868 33572
rect 21924 33516 22540 33572
rect 22596 33516 26236 33572
rect 26292 33516 26302 33572
rect 38770 33516 38780 33572
rect 38836 33516 44268 33572
rect 44324 33516 44940 33572
rect 44996 33516 45006 33572
rect 10322 33404 10332 33460
rect 10388 33404 13580 33460
rect 13636 33404 14140 33460
rect 14196 33404 14206 33460
rect 15138 33404 15148 33460
rect 15204 33404 16380 33460
rect 16436 33404 17500 33460
rect 17556 33404 20188 33460
rect 20244 33404 20254 33460
rect 21298 33404 21308 33460
rect 21364 33404 22428 33460
rect 22484 33404 22494 33460
rect 27010 33404 27020 33460
rect 27076 33404 29484 33460
rect 29540 33404 29550 33460
rect 31266 33404 31276 33460
rect 31332 33404 35868 33460
rect 35924 33404 35934 33460
rect 43698 33404 43708 33460
rect 43764 33404 44380 33460
rect 44436 33404 44446 33460
rect 22306 33292 22316 33348
rect 22372 33292 24556 33348
rect 24612 33292 24622 33348
rect 26002 33292 26012 33348
rect 26068 33292 27580 33348
rect 27636 33292 27646 33348
rect 29362 33292 29372 33348
rect 29428 33292 29484 33348
rect 29540 33292 29550 33348
rect 33058 33292 33068 33348
rect 33124 33292 33740 33348
rect 33796 33292 33806 33348
rect 37314 33292 37324 33348
rect 37380 33292 37996 33348
rect 38052 33292 38556 33348
rect 38612 33292 38780 33348
rect 38836 33292 38846 33348
rect 39106 33292 39116 33348
rect 39172 33292 41580 33348
rect 41636 33292 41646 33348
rect 45490 33292 45500 33348
rect 45556 33292 45948 33348
rect 46004 33292 47516 33348
rect 47572 33292 47582 33348
rect 19170 33180 19180 33236
rect 19236 33180 21308 33236
rect 21364 33180 21374 33236
rect 28242 33180 28252 33236
rect 28308 33180 30380 33236
rect 30436 33180 30446 33236
rect 37314 33180 37324 33236
rect 37380 33180 37548 33236
rect 37604 33180 37614 33236
rect 37874 33180 37884 33236
rect 37940 33180 39900 33236
rect 39956 33180 39966 33236
rect 5954 33068 5964 33124
rect 6020 33068 6748 33124
rect 6804 33068 6814 33124
rect 22866 33068 22876 33124
rect 22932 33068 23548 33124
rect 23604 33068 23614 33124
rect 27682 33068 27692 33124
rect 27748 33068 28588 33124
rect 28644 33068 31164 33124
rect 31220 33068 31230 33124
rect 35410 33068 35420 33124
rect 35476 33068 36428 33124
rect 36484 33068 38780 33124
rect 38836 33068 38846 33124
rect 39218 33068 39228 33124
rect 39284 33068 41692 33124
rect 41748 33068 41758 33124
rect 45378 33068 45388 33124
rect 45444 33068 46956 33124
rect 47012 33068 47852 33124
rect 47908 33068 47918 33124
rect 25778 32956 25788 33012
rect 25844 32956 28140 33012
rect 28196 32956 28206 33012
rect 28466 32956 28476 33012
rect 28532 32956 30268 33012
rect 30324 32956 30334 33012
rect 40338 32956 40348 33012
rect 40404 32956 46060 33012
rect 46116 32956 47964 33012
rect 48020 32956 48030 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 24546 32844 24556 32900
rect 24612 32844 26908 32900
rect 27346 32844 27356 32900
rect 27412 32844 29596 32900
rect 29652 32844 29662 32900
rect 26852 32788 26908 32844
rect 14018 32732 14028 32788
rect 14084 32732 14812 32788
rect 14868 32732 15148 32788
rect 15204 32732 15214 32788
rect 26852 32732 27468 32788
rect 27524 32732 27534 32788
rect 28018 32732 28028 32788
rect 28084 32732 28476 32788
rect 28532 32732 28542 32788
rect 30370 32732 30380 32788
rect 30436 32732 44492 32788
rect 44548 32732 44558 32788
rect 7746 32620 7756 32676
rect 7812 32620 8764 32676
rect 8820 32620 8830 32676
rect 16930 32620 16940 32676
rect 16996 32620 17836 32676
rect 17892 32620 17902 32676
rect 22642 32620 22652 32676
rect 22708 32620 27916 32676
rect 27972 32620 29820 32676
rect 29876 32620 29886 32676
rect 33170 32620 33180 32676
rect 33236 32620 33404 32676
rect 33460 32620 33470 32676
rect 44146 32620 44156 32676
rect 44212 32620 44940 32676
rect 44996 32620 45006 32676
rect 48290 32620 48300 32676
rect 48356 32620 48366 32676
rect 33404 32564 33460 32620
rect 13906 32508 13916 32564
rect 13972 32508 16828 32564
rect 16884 32508 18396 32564
rect 18452 32508 18462 32564
rect 23538 32508 23548 32564
rect 23604 32508 23642 32564
rect 24658 32508 24668 32564
rect 24724 32508 25228 32564
rect 25284 32508 25294 32564
rect 26002 32508 26012 32564
rect 26068 32508 28812 32564
rect 28868 32508 28878 32564
rect 32386 32508 32396 32564
rect 32452 32508 33068 32564
rect 33124 32508 33134 32564
rect 33404 32508 34300 32564
rect 34356 32508 36988 32564
rect 37044 32508 37054 32564
rect 39666 32508 39676 32564
rect 39732 32508 43708 32564
rect 43764 32508 43774 32564
rect 8306 32396 8316 32452
rect 8372 32396 9660 32452
rect 9716 32396 9726 32452
rect 11554 32396 11564 32452
rect 11620 32396 13244 32452
rect 13300 32396 13310 32452
rect 26226 32396 26236 32452
rect 26292 32396 26908 32452
rect 34178 32396 34188 32452
rect 34244 32396 35420 32452
rect 35476 32396 35486 32452
rect 15362 32284 15372 32340
rect 15428 32284 17388 32340
rect 17444 32284 17454 32340
rect 26852 32228 26908 32396
rect 48300 32340 48356 32620
rect 49200 32340 50000 32368
rect 48300 32284 50000 32340
rect 49200 32256 50000 32284
rect 26852 32172 27468 32228
rect 27524 32172 27916 32228
rect 27972 32172 29372 32228
rect 29428 32172 29438 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 32050 32060 32060 32116
rect 32116 32060 33404 32116
rect 33460 32060 33470 32116
rect 26870 31948 26908 32004
rect 26964 31948 26974 32004
rect 38658 31948 38668 32004
rect 38724 31948 38734 32004
rect 45042 31948 45052 32004
rect 45108 31948 47628 32004
rect 47684 31948 47694 32004
rect 38668 31892 38724 31948
rect 3714 31836 3724 31892
rect 3780 31836 4956 31892
rect 5012 31836 5022 31892
rect 6626 31836 6636 31892
rect 6692 31836 13356 31892
rect 13412 31836 13422 31892
rect 20962 31836 20972 31892
rect 21028 31836 21420 31892
rect 21476 31836 21486 31892
rect 24994 31836 25004 31892
rect 25060 31836 25676 31892
rect 25732 31836 26684 31892
rect 26740 31836 26750 31892
rect 37762 31836 37772 31892
rect 37828 31836 38724 31892
rect 41906 31836 41916 31892
rect 41972 31836 43036 31892
rect 43092 31836 43102 31892
rect 43698 31836 43708 31892
rect 43764 31836 47068 31892
rect 47124 31836 48524 31892
rect 48580 31836 48590 31892
rect 10546 31724 10556 31780
rect 10612 31724 13580 31780
rect 13636 31724 14588 31780
rect 14644 31724 14654 31780
rect 20626 31724 20636 31780
rect 20692 31724 22092 31780
rect 22148 31724 22158 31780
rect 27122 31724 27132 31780
rect 27188 31724 27356 31780
rect 27412 31724 27422 31780
rect 27794 31724 27804 31780
rect 27860 31724 28588 31780
rect 28644 31724 28654 31780
rect 36530 31724 36540 31780
rect 36596 31724 37548 31780
rect 37604 31724 39564 31780
rect 39620 31724 39630 31780
rect 42466 31724 42476 31780
rect 42532 31724 43484 31780
rect 43540 31724 44044 31780
rect 44100 31724 44110 31780
rect 44258 31724 44268 31780
rect 44324 31724 45052 31780
rect 45108 31724 46172 31780
rect 46228 31724 46238 31780
rect 2482 31612 2492 31668
rect 2548 31612 5740 31668
rect 5796 31612 5806 31668
rect 6178 31612 6188 31668
rect 6244 31612 7084 31668
rect 7140 31612 7150 31668
rect 8642 31612 8652 31668
rect 8708 31612 9884 31668
rect 9940 31612 9950 31668
rect 11106 31612 11116 31668
rect 11172 31612 11788 31668
rect 11844 31612 11854 31668
rect 12114 31612 12124 31668
rect 12180 31612 13804 31668
rect 13860 31612 13870 31668
rect 18610 31612 18620 31668
rect 18676 31612 19628 31668
rect 19684 31612 21308 31668
rect 21364 31612 21374 31668
rect 21634 31612 21644 31668
rect 21700 31612 23772 31668
rect 23828 31612 23838 31668
rect 27682 31612 27692 31668
rect 27748 31612 30268 31668
rect 30324 31612 30334 31668
rect 33954 31612 33964 31668
rect 34020 31612 39900 31668
rect 39956 31612 39966 31668
rect 40226 31612 40236 31668
rect 40292 31612 41916 31668
rect 41972 31612 41982 31668
rect 42914 31612 42924 31668
rect 42980 31612 43708 31668
rect 43764 31612 43774 31668
rect 45154 31612 45164 31668
rect 45220 31612 46844 31668
rect 46900 31612 46910 31668
rect 4386 31500 4396 31556
rect 4452 31500 6636 31556
rect 6692 31500 6702 31556
rect 25666 31500 25676 31556
rect 25732 31500 26572 31556
rect 26628 31500 26638 31556
rect 27794 31500 27804 31556
rect 27860 31500 29036 31556
rect 29092 31500 29102 31556
rect 33170 31500 33180 31556
rect 33236 31500 33516 31556
rect 33572 31500 33582 31556
rect 34738 31500 34748 31556
rect 34804 31500 37100 31556
rect 37156 31500 37166 31556
rect 37426 31500 37436 31556
rect 37492 31500 41356 31556
rect 41412 31500 43260 31556
rect 43316 31500 43326 31556
rect 46498 31500 46508 31556
rect 46564 31500 47180 31556
rect 47236 31500 47246 31556
rect 26786 31388 26796 31444
rect 26852 31388 30716 31444
rect 30772 31388 30782 31444
rect 31126 31388 31164 31444
rect 31220 31388 31230 31444
rect 35970 31388 35980 31444
rect 36036 31388 37772 31444
rect 37828 31388 37838 31444
rect 38658 31388 38668 31444
rect 38724 31388 47404 31444
rect 47460 31388 47470 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 30716 31332 30772 31388
rect 1810 31276 1820 31332
rect 1876 31276 3724 31332
rect 3780 31276 3790 31332
rect 7186 31276 7196 31332
rect 7252 31276 7756 31332
rect 7812 31276 7822 31332
rect 21410 31276 21420 31332
rect 21476 31276 22652 31332
rect 22708 31276 22718 31332
rect 26562 31276 26572 31332
rect 26628 31276 27916 31332
rect 27972 31276 28476 31332
rect 28532 31276 28542 31332
rect 30716 31276 36204 31332
rect 36260 31276 36270 31332
rect 16258 31164 16268 31220
rect 16324 31164 16828 31220
rect 16884 31164 16894 31220
rect 21186 31164 21196 31220
rect 21252 31164 21868 31220
rect 21924 31164 22540 31220
rect 22596 31164 23100 31220
rect 23156 31164 23166 31220
rect 23650 31164 23660 31220
rect 23716 31164 25564 31220
rect 25620 31164 26796 31220
rect 26852 31164 27020 31220
rect 27076 31164 27086 31220
rect 27356 31164 33964 31220
rect 34020 31164 34030 31220
rect 44146 31164 44156 31220
rect 44212 31164 46396 31220
rect 46452 31164 46462 31220
rect 27356 31108 27412 31164
rect 13682 31052 13692 31108
rect 13748 31052 14364 31108
rect 14420 31052 14924 31108
rect 14980 31052 14990 31108
rect 18274 31052 18284 31108
rect 18340 31052 20748 31108
rect 20804 31052 20814 31108
rect 23986 31052 23996 31108
rect 24052 31052 24780 31108
rect 24836 31052 27412 31108
rect 27570 31052 27580 31108
rect 27636 31052 27646 31108
rect 27906 31052 27916 31108
rect 27972 31052 32116 31108
rect 43250 31052 43260 31108
rect 43316 31052 44268 31108
rect 44324 31052 45276 31108
rect 45332 31052 45342 31108
rect 7074 30940 7084 30996
rect 7140 30940 8316 30996
rect 8372 30940 10780 30996
rect 10836 30940 10846 30996
rect 12114 30940 12124 30996
rect 12180 30940 22988 30996
rect 23044 30940 23054 30996
rect 23772 30940 25676 30996
rect 25732 30940 25742 30996
rect 11554 30828 11564 30884
rect 11620 30828 12572 30884
rect 12628 30828 12638 30884
rect 14130 30828 14140 30884
rect 14196 30828 14588 30884
rect 14644 30828 15148 30884
rect 15204 30828 15214 30884
rect 15586 30828 15596 30884
rect 15652 30828 16044 30884
rect 16100 30828 16604 30884
rect 16660 30828 16670 30884
rect 23772 30772 23828 30940
rect 27580 30884 27636 31052
rect 24658 30828 24668 30884
rect 24724 30828 26124 30884
rect 26180 30828 27636 30884
rect 32060 30884 32116 31052
rect 35074 30940 35084 30996
rect 35140 30940 36540 30996
rect 36596 30940 36606 30996
rect 41682 30940 41692 30996
rect 41748 30940 42364 30996
rect 42420 30940 42430 30996
rect 42802 30940 42812 30996
rect 42868 30940 43932 30996
rect 43988 30940 44828 30996
rect 44884 30940 44894 30996
rect 32060 30828 35980 30884
rect 36036 30828 36764 30884
rect 36820 30828 36830 30884
rect 41234 30828 41244 30884
rect 41300 30828 42028 30884
rect 42084 30828 42094 30884
rect 7186 30716 7196 30772
rect 7252 30716 7420 30772
rect 7476 30716 7486 30772
rect 22306 30716 22316 30772
rect 22372 30716 23772 30772
rect 23828 30716 23838 30772
rect 36082 30716 36092 30772
rect 36148 30716 41132 30772
rect 41188 30716 42476 30772
rect 42532 30716 42542 30772
rect 23090 30604 23100 30660
rect 23156 30604 33180 30660
rect 33236 30604 34860 30660
rect 34916 30604 34926 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 23874 30492 23884 30548
rect 23940 30492 25340 30548
rect 25396 30492 25406 30548
rect 34598 30492 34636 30548
rect 34692 30492 34702 30548
rect 26852 30380 31388 30436
rect 31444 30380 31454 30436
rect 34066 30380 34076 30436
rect 34132 30380 34748 30436
rect 34804 30380 34814 30436
rect 35410 30380 35420 30436
rect 35476 30380 40908 30436
rect 40964 30380 42812 30436
rect 42868 30380 42878 30436
rect 26852 30324 26908 30380
rect 12450 30268 12460 30324
rect 12516 30268 13804 30324
rect 13860 30268 13870 30324
rect 23958 30268 23996 30324
rect 24052 30268 24062 30324
rect 24210 30268 24220 30324
rect 24276 30268 26908 30324
rect 31042 30268 31052 30324
rect 31108 30268 31500 30324
rect 31556 30268 32060 30324
rect 32116 30268 32126 30324
rect 33506 30268 33516 30324
rect 33572 30268 34188 30324
rect 34244 30268 34636 30324
rect 34692 30268 34702 30324
rect 42354 30268 42364 30324
rect 42420 30268 43484 30324
rect 43540 30268 43550 30324
rect 5618 30156 5628 30212
rect 5684 30156 7588 30212
rect 9202 30156 9212 30212
rect 9268 30156 12124 30212
rect 12180 30156 12190 30212
rect 20738 30156 20748 30212
rect 20804 30156 21308 30212
rect 21364 30156 21374 30212
rect 26450 30156 26460 30212
rect 26516 30156 27244 30212
rect 27300 30156 27310 30212
rect 34262 30156 34300 30212
rect 34356 30156 34366 30212
rect 41794 30156 41804 30212
rect 41860 30156 43820 30212
rect 43876 30156 43886 30212
rect 7532 30100 7588 30156
rect 2482 30044 2492 30100
rect 2548 30044 5740 30100
rect 5796 30044 5806 30100
rect 5954 30044 5964 30100
rect 6020 30044 6972 30100
rect 7028 30044 7038 30100
rect 7522 30044 7532 30100
rect 7588 30044 7598 30100
rect 8418 30044 8428 30100
rect 8484 30044 9548 30100
rect 9604 30044 9614 30100
rect 16370 30044 16380 30100
rect 16436 30044 18732 30100
rect 18788 30044 19180 30100
rect 19236 30044 23660 30100
rect 23716 30044 25004 30100
rect 25060 30044 25070 30100
rect 25890 30044 25900 30100
rect 25956 30044 25966 30100
rect 26226 30044 26236 30100
rect 26292 30044 27692 30100
rect 27748 30044 27758 30100
rect 28914 30044 28924 30100
rect 28980 30044 32172 30100
rect 32228 30044 32238 30100
rect 33730 30044 33740 30100
rect 33796 30044 33852 30100
rect 33908 30044 35084 30100
rect 35140 30044 35150 30100
rect 25900 29988 25956 30044
rect 4834 29932 4844 29988
rect 4900 29932 6188 29988
rect 6244 29932 6254 29988
rect 6626 29932 6636 29988
rect 6692 29932 7308 29988
rect 7364 29932 7374 29988
rect 7858 29932 7868 29988
rect 7924 29932 7934 29988
rect 13010 29932 13020 29988
rect 13076 29932 13692 29988
rect 13748 29932 14588 29988
rect 14644 29932 14654 29988
rect 15092 29932 24556 29988
rect 24612 29932 24622 29988
rect 25900 29932 27468 29988
rect 27524 29932 27534 29988
rect 30370 29932 30380 29988
rect 30436 29932 31164 29988
rect 31220 29932 31724 29988
rect 31780 29932 31790 29988
rect 7868 29876 7924 29932
rect 15092 29876 15148 29932
rect 5730 29820 5740 29876
rect 5796 29820 7924 29876
rect 12898 29820 12908 29876
rect 12964 29820 14140 29876
rect 14196 29820 15148 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 6178 29708 6188 29764
rect 6244 29708 7196 29764
rect 7252 29708 7262 29764
rect 23986 29708 23996 29764
rect 24052 29708 28028 29764
rect 28084 29708 30492 29764
rect 30548 29708 31836 29764
rect 31892 29708 31902 29764
rect 4610 29596 4620 29652
rect 4676 29596 5068 29652
rect 5124 29596 7644 29652
rect 7700 29596 7710 29652
rect 18162 29596 18172 29652
rect 18228 29596 18956 29652
rect 19012 29596 19022 29652
rect 19180 29596 33628 29652
rect 33684 29596 35868 29652
rect 35924 29596 35934 29652
rect 38098 29596 38108 29652
rect 38164 29596 39900 29652
rect 39956 29596 39966 29652
rect 19180 29540 19236 29596
rect 6290 29484 6300 29540
rect 6356 29484 6860 29540
rect 6916 29484 7868 29540
rect 7924 29484 8540 29540
rect 8596 29484 8606 29540
rect 16818 29484 16828 29540
rect 16884 29484 18508 29540
rect 18564 29484 18574 29540
rect 18834 29484 18844 29540
rect 18900 29484 19236 29540
rect 26786 29484 26796 29540
rect 26852 29484 27356 29540
rect 27412 29484 28476 29540
rect 28532 29484 28542 29540
rect 33730 29484 33740 29540
rect 33796 29484 34972 29540
rect 35028 29484 35038 29540
rect 41234 29484 41244 29540
rect 41300 29484 42700 29540
rect 42756 29484 42766 29540
rect 3154 29372 3164 29428
rect 3220 29372 4620 29428
rect 4676 29372 5628 29428
rect 5684 29372 6076 29428
rect 6132 29372 6142 29428
rect 12450 29372 12460 29428
rect 12516 29372 13580 29428
rect 13636 29372 16044 29428
rect 16100 29372 17388 29428
rect 17444 29372 17454 29428
rect 34066 29372 34076 29428
rect 34132 29372 37324 29428
rect 37380 29372 40012 29428
rect 40068 29372 40078 29428
rect 43362 29372 43372 29428
rect 43428 29372 43596 29428
rect 43652 29372 43662 29428
rect 2482 29260 2492 29316
rect 2548 29260 3724 29316
rect 3780 29260 3790 29316
rect 8530 29260 8540 29316
rect 8596 29260 11676 29316
rect 11732 29260 11742 29316
rect 12786 29260 12796 29316
rect 12852 29260 14252 29316
rect 14308 29260 14318 29316
rect 14914 29260 14924 29316
rect 14980 29260 16380 29316
rect 16436 29260 17724 29316
rect 17780 29260 17790 29316
rect 21522 29260 21532 29316
rect 21588 29260 22428 29316
rect 22484 29260 22494 29316
rect 24434 29260 24444 29316
rect 24500 29260 29372 29316
rect 29428 29260 29438 29316
rect 36418 29260 36428 29316
rect 36484 29260 37884 29316
rect 37940 29260 37950 29316
rect 39106 29260 39116 29316
rect 39172 29260 40236 29316
rect 40292 29260 40302 29316
rect 44146 29260 44156 29316
rect 44212 29260 45724 29316
rect 45780 29260 45790 29316
rect 40012 29204 40068 29260
rect 3602 29148 3612 29204
rect 3668 29148 5628 29204
rect 5684 29148 5694 29204
rect 40002 29148 40012 29204
rect 40068 29148 40078 29204
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 3042 28812 3052 28868
rect 3108 28812 5180 28868
rect 5236 28812 5246 28868
rect 12002 28812 12012 28868
rect 12068 28812 12684 28868
rect 12740 28812 13580 28868
rect 13636 28812 13646 28868
rect 15708 28812 17948 28868
rect 18004 28812 18014 28868
rect 19730 28812 19740 28868
rect 19796 28812 20636 28868
rect 20692 28812 26908 28868
rect 26964 28812 26974 28868
rect 31602 28812 31612 28868
rect 31668 28812 33516 28868
rect 33572 28812 33582 28868
rect 33814 28812 33852 28868
rect 33908 28812 33918 28868
rect 15708 28756 15764 28812
rect 3826 28700 3836 28756
rect 3892 28700 5068 28756
rect 5124 28700 5134 28756
rect 10770 28700 10780 28756
rect 10836 28700 11676 28756
rect 11732 28700 11742 28756
rect 13122 28700 13132 28756
rect 13188 28700 13804 28756
rect 13860 28700 15764 28756
rect 18050 28700 18060 28756
rect 18116 28700 19180 28756
rect 19236 28700 19246 28756
rect 21410 28700 21420 28756
rect 21476 28700 22764 28756
rect 22820 28700 22830 28756
rect 23986 28700 23996 28756
rect 24052 28700 26012 28756
rect 26068 28700 26078 28756
rect 39778 28700 39788 28756
rect 39844 28700 45836 28756
rect 45892 28700 45902 28756
rect 18060 28644 18116 28700
rect 2482 28588 2492 28644
rect 2548 28588 3388 28644
rect 3490 28588 3500 28644
rect 3556 28588 4732 28644
rect 4788 28588 4798 28644
rect 9650 28588 9660 28644
rect 9716 28588 14924 28644
rect 14980 28588 18116 28644
rect 18834 28588 18844 28644
rect 18900 28588 19292 28644
rect 19348 28588 19358 28644
rect 21644 28588 22540 28644
rect 22596 28588 22606 28644
rect 26114 28588 26124 28644
rect 26180 28588 26684 28644
rect 26740 28588 27580 28644
rect 27636 28588 27646 28644
rect 34738 28588 34748 28644
rect 34804 28588 36428 28644
rect 36484 28588 36494 28644
rect 43362 28588 43372 28644
rect 43428 28588 45052 28644
rect 45108 28588 45118 28644
rect 47394 28588 47404 28644
rect 47460 28588 48188 28644
rect 48244 28588 48254 28644
rect 3332 28532 3388 28588
rect 21644 28532 21700 28588
rect 3332 28476 4620 28532
rect 4676 28476 4686 28532
rect 8082 28476 8092 28532
rect 8148 28476 9100 28532
rect 9156 28476 9166 28532
rect 10994 28476 11004 28532
rect 11060 28476 12460 28532
rect 12516 28476 12526 28532
rect 19058 28476 19068 28532
rect 19124 28476 19964 28532
rect 20020 28476 20030 28532
rect 20290 28476 20300 28532
rect 20356 28476 21644 28532
rect 21700 28476 21710 28532
rect 28242 28476 28252 28532
rect 28308 28476 29260 28532
rect 29316 28476 29484 28532
rect 29540 28476 29550 28532
rect 33852 28476 34300 28532
rect 34356 28476 34366 28532
rect 36978 28476 36988 28532
rect 37044 28476 38668 28532
rect 38724 28476 39676 28532
rect 39732 28476 39742 28532
rect 33852 28420 33908 28476
rect 5394 28364 5404 28420
rect 5460 28364 5964 28420
rect 6020 28364 6030 28420
rect 6626 28364 6636 28420
rect 6692 28364 8988 28420
rect 9044 28364 9054 28420
rect 18610 28364 18620 28420
rect 18676 28364 19516 28420
rect 19572 28364 19582 28420
rect 27794 28364 27804 28420
rect 27860 28364 28588 28420
rect 28644 28364 29148 28420
rect 29204 28364 29214 28420
rect 30258 28364 30268 28420
rect 30324 28364 30716 28420
rect 30772 28364 30782 28420
rect 31154 28364 31164 28420
rect 31220 28364 32172 28420
rect 32228 28364 32238 28420
rect 33842 28364 33852 28420
rect 33908 28364 33918 28420
rect 40338 28364 40348 28420
rect 40404 28364 41244 28420
rect 41300 28364 41310 28420
rect 42466 28364 42476 28420
rect 42532 28364 43260 28420
rect 43316 28364 43820 28420
rect 43876 28364 43886 28420
rect 45042 28364 45052 28420
rect 45108 28364 45388 28420
rect 45444 28364 45454 28420
rect 7074 28252 7084 28308
rect 7140 28252 8316 28308
rect 8372 28252 8382 28308
rect 37762 28252 37772 28308
rect 37828 28252 38332 28308
rect 38388 28252 42700 28308
rect 42756 28252 42766 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 10322 28140 10332 28196
rect 10388 28140 10780 28196
rect 10836 28140 11340 28196
rect 11396 28140 19684 28196
rect 27346 28140 27356 28196
rect 27412 28140 27916 28196
rect 27972 28140 32060 28196
rect 32116 28140 33292 28196
rect 33348 28140 33358 28196
rect 19628 28084 19684 28140
rect 8642 28028 8652 28084
rect 8708 28028 9660 28084
rect 9716 28028 9726 28084
rect 13682 28028 13692 28084
rect 13748 28028 15820 28084
rect 15876 28028 15886 28084
rect 19628 28028 24556 28084
rect 24612 28028 24892 28084
rect 24948 28028 24958 28084
rect 26198 28028 26236 28084
rect 26292 28028 26302 28084
rect 27122 28028 27132 28084
rect 27188 28028 28476 28084
rect 28532 28028 30044 28084
rect 30100 28028 30110 28084
rect 31266 28028 31276 28084
rect 31332 28028 31948 28084
rect 32004 28028 32014 28084
rect 14914 27916 14924 27972
rect 14980 27916 15932 27972
rect 15988 27916 17500 27972
rect 17556 27916 17566 27972
rect 26852 27916 38668 27972
rect 26852 27860 26908 27916
rect 9314 27804 9324 27860
rect 9380 27804 20412 27860
rect 20468 27804 20478 27860
rect 21410 27804 21420 27860
rect 21476 27804 21756 27860
rect 21812 27804 21822 27860
rect 26114 27804 26124 27860
rect 26180 27804 26908 27860
rect 30146 27804 30156 27860
rect 30212 27804 31836 27860
rect 31892 27804 31902 27860
rect 33730 27804 33740 27860
rect 33796 27804 34524 27860
rect 34580 27804 36988 27860
rect 37044 27804 37054 27860
rect 38612 27804 38668 27916
rect 41020 27860 41076 28252
rect 41458 28028 41468 28084
rect 41524 28028 42140 28084
rect 42196 28028 48076 28084
rect 48132 28028 48142 28084
rect 38724 27804 38734 27860
rect 41010 27804 41020 27860
rect 41076 27804 41086 27860
rect 1810 27692 1820 27748
rect 1876 27692 4172 27748
rect 4228 27692 4238 27748
rect 16146 27692 16156 27748
rect 16212 27692 16828 27748
rect 16884 27692 16894 27748
rect 17490 27692 17500 27748
rect 17556 27692 18956 27748
rect 19012 27692 19022 27748
rect 29138 27692 29148 27748
rect 29204 27692 29596 27748
rect 29652 27692 29662 27748
rect 33282 27692 33292 27748
rect 33348 27692 34412 27748
rect 34468 27692 34478 27748
rect 34822 27692 34860 27748
rect 34916 27692 34926 27748
rect 14354 27580 14364 27636
rect 14420 27580 15932 27636
rect 15988 27580 15998 27636
rect 16706 27580 16716 27636
rect 16772 27580 17388 27636
rect 17444 27580 17454 27636
rect 29698 27580 29708 27636
rect 29764 27580 34636 27636
rect 34692 27580 34702 27636
rect 43026 27580 43036 27636
rect 43092 27580 43596 27636
rect 43652 27580 43662 27636
rect 25442 27468 25452 27524
rect 25508 27468 26236 27524
rect 26292 27468 26302 27524
rect 26460 27468 30492 27524
rect 30548 27468 30558 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 26460 27412 26516 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 49200 27412 50000 27440
rect 15138 27356 15148 27412
rect 15204 27356 26516 27412
rect 26898 27356 26908 27412
rect 26964 27356 32284 27412
rect 32340 27356 32844 27412
rect 32900 27356 32910 27412
rect 48178 27356 48188 27412
rect 48244 27356 50000 27412
rect 49200 27328 50000 27356
rect 4610 27244 4620 27300
rect 4676 27244 5628 27300
rect 5684 27244 5694 27300
rect 20962 27244 20972 27300
rect 21028 27244 25788 27300
rect 25844 27244 27356 27300
rect 27412 27244 33012 27300
rect 33170 27244 33180 27300
rect 33236 27244 33964 27300
rect 34020 27244 34030 27300
rect 42130 27244 42140 27300
rect 42196 27244 42476 27300
rect 42532 27244 42542 27300
rect 42690 27244 42700 27300
rect 42756 27244 44940 27300
rect 44996 27244 48244 27300
rect 32956 27188 33012 27244
rect 48188 27188 48244 27244
rect 8194 27132 8204 27188
rect 8260 27132 8988 27188
rect 9044 27132 9054 27188
rect 20402 27132 20412 27188
rect 20468 27132 21084 27188
rect 21140 27132 21150 27188
rect 21308 27132 26012 27188
rect 26068 27132 27020 27188
rect 27076 27132 27086 27188
rect 31490 27132 31500 27188
rect 31556 27132 32508 27188
rect 32564 27132 32574 27188
rect 32956 27132 34076 27188
rect 34132 27132 35420 27188
rect 35476 27132 35486 27188
rect 48178 27132 48188 27188
rect 48244 27132 48254 27188
rect 21308 27076 21364 27132
rect 15138 27020 15148 27076
rect 15204 27020 15820 27076
rect 15876 27020 15886 27076
rect 18722 27020 18732 27076
rect 18788 27020 21364 27076
rect 23538 27020 23548 27076
rect 23604 27020 24220 27076
rect 24276 27020 26796 27076
rect 26852 27020 26862 27076
rect 32386 27020 32396 27076
rect 32452 27020 32462 27076
rect 32610 27020 32620 27076
rect 32676 27020 33404 27076
rect 33460 27020 33852 27076
rect 33908 27020 33918 27076
rect 34514 27020 34524 27076
rect 34580 27020 36540 27076
rect 36596 27020 39340 27076
rect 39396 27020 40348 27076
rect 40404 27020 40414 27076
rect 41346 27020 41356 27076
rect 41412 27020 43148 27076
rect 43204 27020 43214 27076
rect 32396 26964 32452 27020
rect 41356 26964 41412 27020
rect 4162 26908 4172 26964
rect 4228 26908 4620 26964
rect 4676 26908 6076 26964
rect 6132 26908 6142 26964
rect 13570 26908 13580 26964
rect 13636 26908 14588 26964
rect 14644 26908 14654 26964
rect 18610 26908 18620 26964
rect 18676 26908 25676 26964
rect 25732 26908 26572 26964
rect 26628 26908 26638 26964
rect 26908 26908 29820 26964
rect 29876 26908 29886 26964
rect 31490 26908 31500 26964
rect 31556 26908 32060 26964
rect 32116 26908 32126 26964
rect 32396 26908 32900 26964
rect 38546 26908 38556 26964
rect 38612 26908 39228 26964
rect 39284 26908 40124 26964
rect 40180 26908 40190 26964
rect 40348 26908 41412 26964
rect 42914 26908 42924 26964
rect 42980 26908 42990 26964
rect 43922 26908 43932 26964
rect 43988 26908 44492 26964
rect 44548 26908 47628 26964
rect 47684 26908 47694 26964
rect 26908 26852 26964 26908
rect 28028 26852 28084 26908
rect 32834 26852 32844 26908
rect 32900 26852 32910 26908
rect 19954 26796 19964 26852
rect 20020 26796 23996 26852
rect 24052 26796 24062 26852
rect 24322 26796 24332 26852
rect 24388 26796 24892 26852
rect 24948 26796 24958 26852
rect 26898 26796 26908 26852
rect 26964 26796 26974 26852
rect 28018 26796 28028 26852
rect 28084 26796 28094 26852
rect 33058 26796 33068 26852
rect 33124 26796 33852 26852
rect 33908 26796 33918 26852
rect 40348 26740 40404 26908
rect 42924 26852 42980 26908
rect 42924 26796 44828 26852
rect 44884 26796 44894 26852
rect 24658 26684 24668 26740
rect 24724 26684 25228 26740
rect 25284 26684 25294 26740
rect 28802 26684 28812 26740
rect 28868 26684 32732 26740
rect 32788 26684 37548 26740
rect 37604 26684 37614 26740
rect 40114 26684 40124 26740
rect 40180 26684 40404 26740
rect 42466 26684 42476 26740
rect 42532 26684 44380 26740
rect 44436 26684 44446 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 16258 26572 16268 26628
rect 16324 26572 18620 26628
rect 18676 26572 18686 26628
rect 20188 26572 33740 26628
rect 33796 26572 34636 26628
rect 34692 26572 34702 26628
rect 42018 26572 42028 26628
rect 42084 26572 43932 26628
rect 43988 26572 43998 26628
rect 6850 26460 6860 26516
rect 6916 26460 8428 26516
rect 8484 26460 8494 26516
rect 10546 26460 10556 26516
rect 10612 26460 11452 26516
rect 11508 26460 11518 26516
rect 16594 26460 16604 26516
rect 16660 26460 19068 26516
rect 19124 26460 19134 26516
rect 20188 26404 20244 26572
rect 23426 26460 23436 26516
rect 23492 26460 25788 26516
rect 25844 26460 25854 26516
rect 39442 26460 39452 26516
rect 39508 26460 40796 26516
rect 40852 26460 41804 26516
rect 41860 26460 41870 26516
rect 44930 26460 44940 26516
rect 44996 26460 45836 26516
rect 45892 26460 45902 26516
rect 16370 26348 16380 26404
rect 16436 26348 17836 26404
rect 17892 26348 20244 26404
rect 21858 26348 21868 26404
rect 21924 26348 25228 26404
rect 25284 26348 25294 26404
rect 40898 26348 40908 26404
rect 40964 26348 41580 26404
rect 41636 26348 42028 26404
rect 42084 26348 42094 26404
rect 42802 26348 42812 26404
rect 42868 26348 43484 26404
rect 43540 26348 43550 26404
rect 3714 26236 3724 26292
rect 3780 26236 4844 26292
rect 4900 26236 4910 26292
rect 12226 26236 12236 26292
rect 12292 26236 12908 26292
rect 12964 26236 13468 26292
rect 13524 26236 13534 26292
rect 16818 26236 16828 26292
rect 16884 26236 17388 26292
rect 17444 26236 18620 26292
rect 18676 26236 18686 26292
rect 20738 26236 20748 26292
rect 20804 26236 22204 26292
rect 22260 26236 22270 26292
rect 24546 26236 24556 26292
rect 24612 26236 26012 26292
rect 26068 26236 26078 26292
rect 37538 26236 37548 26292
rect 37604 26236 38892 26292
rect 38948 26236 39340 26292
rect 39396 26236 39406 26292
rect 42130 26236 42140 26292
rect 42196 26236 43596 26292
rect 43652 26236 43662 26292
rect 45154 26236 45164 26292
rect 45220 26236 46508 26292
rect 46564 26236 46574 26292
rect 3826 26124 3836 26180
rect 3892 26124 5068 26180
rect 5124 26124 5134 26180
rect 19058 26124 19068 26180
rect 19124 26124 28924 26180
rect 28980 26124 28990 26180
rect 41122 26012 41132 26068
rect 41188 26012 42588 26068
rect 42644 26012 42654 26068
rect 42242 25900 42252 25956
rect 42308 25900 42700 25956
rect 42756 25900 42766 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 16370 25788 16380 25844
rect 16436 25788 17948 25844
rect 18004 25788 24556 25844
rect 24612 25788 24622 25844
rect 43138 25788 43148 25844
rect 43204 25788 47068 25844
rect 47124 25788 47134 25844
rect 4162 25676 4172 25732
rect 4228 25676 5180 25732
rect 5236 25676 5246 25732
rect 7298 25676 7308 25732
rect 7364 25676 8540 25732
rect 8596 25676 8606 25732
rect 21522 25676 21532 25732
rect 21588 25676 22652 25732
rect 22708 25676 25452 25732
rect 25508 25676 25518 25732
rect 37986 25676 37996 25732
rect 38052 25676 38780 25732
rect 38836 25676 38846 25732
rect 24882 25564 24892 25620
rect 24948 25564 25172 25620
rect 32946 25564 32956 25620
rect 33012 25564 33180 25620
rect 33236 25564 33740 25620
rect 33796 25564 33806 25620
rect 3042 25452 3052 25508
rect 3108 25452 3948 25508
rect 4004 25452 4014 25508
rect 4722 25452 4732 25508
rect 4788 25452 5628 25508
rect 5684 25452 5694 25508
rect 6972 25452 7644 25508
rect 7700 25452 7710 25508
rect 8642 25452 8652 25508
rect 8708 25452 10444 25508
rect 10500 25452 10510 25508
rect 17490 25452 17500 25508
rect 17556 25452 20188 25508
rect 20244 25452 21980 25508
rect 22036 25452 23548 25508
rect 23604 25452 23614 25508
rect 4732 25396 4788 25452
rect 6972 25396 7028 25452
rect 25116 25396 25172 25564
rect 36418 25452 36428 25508
rect 36484 25452 37324 25508
rect 37380 25452 37660 25508
rect 37716 25452 37726 25508
rect 43558 25452 43596 25508
rect 43652 25452 43662 25508
rect 44034 25452 44044 25508
rect 44100 25452 45164 25508
rect 45220 25452 45230 25508
rect 3602 25340 3612 25396
rect 3668 25340 4788 25396
rect 6738 25340 6748 25396
rect 6804 25340 6972 25396
rect 7028 25340 7038 25396
rect 7410 25340 7420 25396
rect 7476 25340 8876 25396
rect 8932 25340 8942 25396
rect 11778 25340 11788 25396
rect 11844 25340 14252 25396
rect 14308 25340 14318 25396
rect 25116 25340 27804 25396
rect 27860 25340 28476 25396
rect 28532 25340 28542 25396
rect 36978 25340 36988 25396
rect 37044 25340 38108 25396
rect 38164 25340 39004 25396
rect 39060 25340 39070 25396
rect 39666 25340 39676 25396
rect 39732 25340 40684 25396
rect 40740 25340 40750 25396
rect 43334 25340 43372 25396
rect 43428 25340 43438 25396
rect 44930 25340 44940 25396
rect 44996 25340 47180 25396
rect 47236 25340 48188 25396
rect 48244 25340 48254 25396
rect 25116 25284 25172 25340
rect 1698 25228 1708 25284
rect 1764 25228 2940 25284
rect 2996 25228 3500 25284
rect 3556 25228 3566 25284
rect 6402 25228 6412 25284
rect 6468 25228 7084 25284
rect 7140 25228 7756 25284
rect 7812 25228 7822 25284
rect 8082 25228 8092 25284
rect 8148 25228 8372 25284
rect 8530 25228 8540 25284
rect 8596 25228 9324 25284
rect 9380 25228 9884 25284
rect 9940 25228 11228 25284
rect 11284 25228 11294 25284
rect 21746 25228 21756 25284
rect 21812 25228 23604 25284
rect 25106 25228 25116 25284
rect 25172 25228 25182 25284
rect 25442 25228 25452 25284
rect 25508 25228 32508 25284
rect 32564 25228 32574 25284
rect 33842 25228 33852 25284
rect 33908 25228 39452 25284
rect 39508 25228 39518 25284
rect 42354 25228 42364 25284
rect 42420 25228 43036 25284
rect 43092 25228 43932 25284
rect 43988 25228 43998 25284
rect 8316 25172 8372 25228
rect 23548 25172 23604 25228
rect 8316 25116 8876 25172
rect 8932 25116 9436 25172
rect 9492 25116 9502 25172
rect 9762 25116 9772 25172
rect 9828 25116 10332 25172
rect 10388 25116 11116 25172
rect 11172 25116 11182 25172
rect 23548 25116 26796 25172
rect 26852 25116 28588 25172
rect 28644 25116 36204 25172
rect 36260 25116 37212 25172
rect 37268 25116 37278 25172
rect 9436 25060 9492 25116
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 9436 25004 12236 25060
rect 12292 25004 12302 25060
rect 24322 25004 24332 25060
rect 24388 25004 31612 25060
rect 31668 25004 31678 25060
rect 37286 25004 37324 25060
rect 37380 25004 37390 25060
rect 16370 24892 16380 24948
rect 16436 24892 20580 24948
rect 24434 24892 24444 24948
rect 24500 24892 30492 24948
rect 30548 24892 30558 24948
rect 20524 24836 20580 24892
rect 2706 24780 2716 24836
rect 2772 24780 5180 24836
rect 5236 24780 5246 24836
rect 7858 24780 7868 24836
rect 7924 24780 9884 24836
rect 9940 24780 9950 24836
rect 19506 24780 19516 24836
rect 19572 24780 20300 24836
rect 20356 24780 20366 24836
rect 20524 24780 25452 24836
rect 25508 24780 25518 24836
rect 41682 24780 41692 24836
rect 41748 24780 42476 24836
rect 42532 24780 42542 24836
rect 43138 24780 43148 24836
rect 43204 24780 43596 24836
rect 43652 24780 43662 24836
rect 8306 24668 8316 24724
rect 8372 24668 9996 24724
rect 10052 24668 10062 24724
rect 13346 24668 13356 24724
rect 13412 24668 25340 24724
rect 25396 24668 25788 24724
rect 25844 24668 25854 24724
rect 38322 24668 38332 24724
rect 38388 24668 40012 24724
rect 40068 24668 40078 24724
rect 2482 24556 2492 24612
rect 2548 24556 5068 24612
rect 5124 24556 5134 24612
rect 16818 24556 16828 24612
rect 16884 24556 19516 24612
rect 19572 24556 19582 24612
rect 22194 24556 22204 24612
rect 22260 24556 22876 24612
rect 22932 24556 22942 24612
rect 34066 24556 34076 24612
rect 34132 24556 35980 24612
rect 36036 24556 37884 24612
rect 37940 24556 37950 24612
rect 19730 24444 19740 24500
rect 19796 24444 20636 24500
rect 20692 24444 20702 24500
rect 21970 24444 21980 24500
rect 22036 24444 22988 24500
rect 23044 24444 24444 24500
rect 24500 24444 25900 24500
rect 25956 24444 25966 24500
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 31126 24220 31164 24276
rect 31220 24220 31230 24276
rect 30454 24108 30492 24164
rect 30548 24108 30558 24164
rect 41906 24108 41916 24164
rect 41972 24108 42812 24164
rect 42868 24108 42878 24164
rect 6738 23996 6748 24052
rect 6804 23996 8316 24052
rect 8372 23996 8382 24052
rect 10546 23996 10556 24052
rect 10612 23996 12124 24052
rect 12180 23996 12190 24052
rect 18162 23996 18172 24052
rect 18228 23996 21756 24052
rect 21812 23996 21822 24052
rect 27234 23996 27244 24052
rect 27300 23996 27916 24052
rect 27972 23996 29372 24052
rect 29428 23996 29438 24052
rect 6178 23884 6188 23940
rect 6244 23884 7196 23940
rect 7252 23884 7262 23940
rect 8978 23884 8988 23940
rect 9044 23884 12460 23940
rect 12516 23884 12526 23940
rect 13570 23884 13580 23940
rect 13636 23884 16828 23940
rect 16884 23884 18060 23940
rect 18116 23884 18126 23940
rect 22978 23884 22988 23940
rect 23044 23884 26124 23940
rect 26180 23884 26190 23940
rect 27570 23884 27580 23940
rect 27636 23884 28140 23940
rect 28196 23884 29148 23940
rect 29204 23884 29214 23940
rect 37874 23884 37884 23940
rect 37940 23884 38444 23940
rect 38500 23884 39228 23940
rect 39284 23884 39294 23940
rect 39778 23884 39788 23940
rect 39844 23884 41804 23940
rect 41860 23884 41870 23940
rect 43138 23884 43148 23940
rect 43204 23884 43596 23940
rect 43652 23884 44156 23940
rect 44212 23884 45388 23940
rect 45444 23884 45454 23940
rect 5842 23772 5852 23828
rect 5908 23772 8428 23828
rect 8484 23772 8494 23828
rect 17602 23772 17612 23828
rect 17668 23772 23100 23828
rect 23156 23772 23166 23828
rect 25218 23772 25228 23828
rect 25284 23772 26684 23828
rect 26740 23772 27020 23828
rect 27076 23772 27086 23828
rect 28466 23772 28476 23828
rect 28532 23772 29484 23828
rect 29540 23772 29550 23828
rect 30146 23772 30156 23828
rect 30212 23772 31948 23828
rect 32004 23772 33068 23828
rect 33124 23772 33134 23828
rect 36418 23772 36428 23828
rect 36484 23772 38668 23828
rect 44034 23772 44044 23828
rect 44100 23772 45052 23828
rect 45108 23772 45118 23828
rect 46386 23772 46396 23828
rect 46452 23772 47404 23828
rect 47460 23772 47470 23828
rect 3266 23660 3276 23716
rect 3332 23660 4172 23716
rect 4228 23660 5684 23716
rect 21746 23660 21756 23716
rect 21812 23660 22988 23716
rect 23044 23660 23054 23716
rect 25778 23660 25788 23716
rect 25844 23660 27356 23716
rect 27412 23660 27422 23716
rect 28578 23660 28588 23716
rect 28644 23660 29372 23716
rect 29428 23660 29438 23716
rect 34626 23660 34636 23716
rect 34692 23660 34972 23716
rect 35028 23660 35038 23716
rect 38612 23660 38668 23772
rect 38724 23660 38734 23716
rect 39554 23660 39564 23716
rect 39620 23660 40236 23716
rect 40292 23660 40302 23716
rect 43698 23660 43708 23716
rect 43764 23660 44884 23716
rect 5628 23604 5684 23660
rect 44828 23604 44884 23660
rect 3602 23548 3612 23604
rect 3668 23548 4508 23604
rect 4564 23548 4574 23604
rect 5618 23548 5628 23604
rect 5684 23548 6748 23604
rect 6804 23548 6814 23604
rect 21634 23548 21644 23604
rect 21700 23548 22764 23604
rect 22820 23548 22830 23604
rect 27458 23548 27468 23604
rect 27524 23548 42364 23604
rect 42420 23548 43596 23604
rect 43652 23548 43662 23604
rect 44828 23548 44940 23604
rect 44996 23548 45164 23604
rect 45220 23548 45230 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 14354 23436 14364 23492
rect 14420 23436 15484 23492
rect 15540 23436 15550 23492
rect 23426 23436 23436 23492
rect 23492 23436 31108 23492
rect 31266 23436 31276 23492
rect 31332 23436 37324 23492
rect 37380 23436 37390 23492
rect 39442 23436 39452 23492
rect 39508 23436 41580 23492
rect 41636 23436 41646 23492
rect 42802 23436 42812 23492
rect 42868 23436 43708 23492
rect 43764 23436 44492 23492
rect 44548 23436 44558 23492
rect 31052 23380 31108 23436
rect 14578 23324 14588 23380
rect 14644 23324 15260 23380
rect 15316 23324 15326 23380
rect 18620 23324 20748 23380
rect 20804 23324 20814 23380
rect 22194 23324 22204 23380
rect 22260 23324 23212 23380
rect 23268 23324 23884 23380
rect 23940 23324 23950 23380
rect 24546 23324 24556 23380
rect 24612 23324 27132 23380
rect 27188 23324 27198 23380
rect 31052 23324 32004 23380
rect 33842 23324 33852 23380
rect 33908 23324 34748 23380
rect 34804 23324 34814 23380
rect 36866 23324 36876 23380
rect 36932 23324 36942 23380
rect 37426 23324 37436 23380
rect 37492 23324 38444 23380
rect 38500 23324 38510 23380
rect 42018 23324 42028 23380
rect 42084 23324 42700 23380
rect 42756 23324 42766 23380
rect 18620 23268 18676 23324
rect 31948 23268 32004 23324
rect 36876 23268 36932 23324
rect 8642 23212 8652 23268
rect 8708 23212 10892 23268
rect 10948 23212 10958 23268
rect 13458 23212 13468 23268
rect 13524 23212 14924 23268
rect 14980 23212 14990 23268
rect 16818 23212 16828 23268
rect 16884 23212 18620 23268
rect 18676 23212 18686 23268
rect 20402 23212 20412 23268
rect 20468 23212 23100 23268
rect 23156 23212 23166 23268
rect 23986 23212 23996 23268
rect 24052 23212 29260 23268
rect 29316 23212 31892 23268
rect 31948 23212 34804 23268
rect 36306 23212 36316 23268
rect 36372 23212 39564 23268
rect 39620 23212 39630 23268
rect 41244 23212 46060 23268
rect 46116 23212 47292 23268
rect 47348 23212 47358 23268
rect 31836 23156 31892 23212
rect 4050 23100 4060 23156
rect 4116 23100 5628 23156
rect 5684 23100 5694 23156
rect 12450 23100 12460 23156
rect 12516 23100 17500 23156
rect 17556 23100 21308 23156
rect 21364 23100 21374 23156
rect 22754 23100 22764 23156
rect 22820 23100 28028 23156
rect 28084 23100 28094 23156
rect 31826 23100 31836 23156
rect 31892 23100 31902 23156
rect 32498 23100 32508 23156
rect 32564 23100 33292 23156
rect 33348 23100 34300 23156
rect 34356 23100 34366 23156
rect 25106 22988 25116 23044
rect 25172 22988 26348 23044
rect 26404 22988 26414 23044
rect 13682 22876 13692 22932
rect 13748 22876 14476 22932
rect 14532 22876 14542 22932
rect 21858 22876 21868 22932
rect 21924 22876 25564 22932
rect 25620 22876 31276 22932
rect 31332 22876 31342 22932
rect 33740 22820 33796 23100
rect 34748 23044 34804 23212
rect 41244 23156 41300 23212
rect 35522 23100 35532 23156
rect 35588 23100 38780 23156
rect 38836 23100 38846 23156
rect 39442 23100 39452 23156
rect 39508 23100 41300 23156
rect 41458 23100 41468 23156
rect 41524 23100 42476 23156
rect 42532 23100 42542 23156
rect 34738 22988 34748 23044
rect 34804 22988 34814 23044
rect 35410 22988 35420 23044
rect 35476 22988 35644 23044
rect 35700 22988 35710 23044
rect 36082 22988 36092 23044
rect 36148 22988 36876 23044
rect 36932 22988 36942 23044
rect 37090 22988 37100 23044
rect 37156 22988 37772 23044
rect 37828 22988 37838 23044
rect 45042 22988 45052 23044
rect 45108 22988 45836 23044
rect 45892 22988 45902 23044
rect 47618 22988 47628 23044
rect 47684 22988 48188 23044
rect 48244 22988 48254 23044
rect 34962 22876 34972 22932
rect 35028 22876 35532 22932
rect 35588 22876 35598 22932
rect 35970 22876 35980 22932
rect 36036 22876 37884 22932
rect 37940 22876 37950 22932
rect 44258 22876 44268 22932
rect 44324 22876 46060 22932
rect 46116 22876 46126 22932
rect 15474 22764 15484 22820
rect 15540 22764 16380 22820
rect 16436 22764 18284 22820
rect 18340 22764 18350 22820
rect 33730 22764 33740 22820
rect 33796 22764 33806 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 38434 22652 38444 22708
rect 38500 22652 43484 22708
rect 43540 22652 45276 22708
rect 45332 22652 45342 22708
rect 3378 22540 3388 22596
rect 3444 22540 4620 22596
rect 4676 22540 5404 22596
rect 5460 22540 6300 22596
rect 6356 22540 6366 22596
rect 43334 22540 43372 22596
rect 43428 22540 43438 22596
rect 49200 22484 50000 22512
rect 15698 22428 15708 22484
rect 15764 22428 17276 22484
rect 17332 22428 17342 22484
rect 17826 22428 17836 22484
rect 17892 22428 20412 22484
rect 20468 22428 20478 22484
rect 24546 22428 24556 22484
rect 24612 22428 25676 22484
rect 25732 22428 25742 22484
rect 29138 22428 29148 22484
rect 29204 22428 30828 22484
rect 30884 22428 30894 22484
rect 39890 22428 39900 22484
rect 39956 22428 40460 22484
rect 40516 22428 40526 22484
rect 43026 22428 43036 22484
rect 43092 22428 43708 22484
rect 43764 22428 45276 22484
rect 45332 22428 45342 22484
rect 48178 22428 48188 22484
rect 48244 22428 50000 22484
rect 49200 22400 50000 22428
rect 5618 22316 5628 22372
rect 5684 22316 6412 22372
rect 6468 22316 7420 22372
rect 7476 22316 7486 22372
rect 29586 22316 29596 22372
rect 29652 22316 35980 22372
rect 36036 22316 36046 22372
rect 19954 22204 19964 22260
rect 20020 22204 22876 22260
rect 22932 22204 22942 22260
rect 31266 22204 31276 22260
rect 31332 22204 32284 22260
rect 32340 22204 32350 22260
rect 33926 22204 33964 22260
rect 34020 22204 34030 22260
rect 41794 22204 41804 22260
rect 41860 22204 42924 22260
rect 42980 22204 42990 22260
rect 45602 22204 45612 22260
rect 45668 22204 47404 22260
rect 47460 22204 47470 22260
rect 4946 22092 4956 22148
rect 5012 22092 6076 22148
rect 6132 22092 6142 22148
rect 16706 22092 16716 22148
rect 16772 22092 21868 22148
rect 21924 22092 21934 22148
rect 27794 22092 27804 22148
rect 27860 22092 28476 22148
rect 28532 22092 28542 22148
rect 31714 22092 31724 22148
rect 31780 22092 32620 22148
rect 32676 22092 32686 22148
rect 32844 22092 35644 22148
rect 35700 22092 41468 22148
rect 41524 22092 41534 22148
rect 28476 22036 28532 22092
rect 32844 22036 32900 22092
rect 22418 21980 22428 22036
rect 22484 21980 22876 22036
rect 22932 21980 22942 22036
rect 28476 21980 32060 22036
rect 32116 21980 32284 22036
rect 32340 21980 32350 22036
rect 32834 21980 32844 22036
rect 32900 21980 32910 22036
rect 34738 21980 34748 22036
rect 34804 21980 37548 22036
rect 37604 21980 37614 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 21970 21868 21980 21924
rect 22036 21868 22652 21924
rect 22708 21868 23324 21924
rect 23380 21868 23390 21924
rect 34374 21868 34412 21924
rect 34468 21868 34478 21924
rect 35252 21868 36092 21924
rect 36148 21868 41916 21924
rect 41972 21868 43372 21924
rect 43428 21868 43438 21924
rect 45378 21868 45388 21924
rect 45444 21868 48076 21924
rect 48132 21868 48142 21924
rect 2482 21756 2492 21812
rect 2548 21756 3836 21812
rect 3892 21756 3902 21812
rect 6850 21756 6860 21812
rect 6916 21756 7420 21812
rect 7476 21756 8540 21812
rect 8596 21756 8606 21812
rect 23090 21756 23100 21812
rect 23156 21756 23996 21812
rect 24052 21756 24062 21812
rect 27570 21756 27580 21812
rect 27636 21756 28812 21812
rect 28868 21756 28878 21812
rect 30818 21756 30828 21812
rect 30884 21756 31836 21812
rect 31892 21756 31902 21812
rect 35252 21700 35308 21868
rect 37426 21756 37436 21812
rect 37492 21756 38780 21812
rect 38836 21756 45500 21812
rect 45556 21756 46060 21812
rect 46116 21756 46126 21812
rect 47954 21756 47964 21812
rect 48020 21756 48188 21812
rect 48244 21756 48254 21812
rect 3490 21644 3500 21700
rect 3556 21644 4396 21700
rect 4452 21644 4462 21700
rect 7746 21644 7756 21700
rect 7812 21644 8428 21700
rect 8484 21644 8494 21700
rect 16594 21644 16604 21700
rect 16660 21644 19852 21700
rect 19908 21644 19918 21700
rect 22754 21644 22764 21700
rect 22820 21644 23436 21700
rect 23492 21644 24444 21700
rect 24500 21644 24510 21700
rect 30482 21644 30492 21700
rect 30548 21644 34188 21700
rect 34244 21644 34254 21700
rect 34626 21644 34636 21700
rect 34692 21644 35308 21700
rect 44482 21644 44492 21700
rect 44548 21644 46396 21700
rect 46452 21644 46462 21700
rect 4274 21532 4284 21588
rect 4340 21532 5180 21588
rect 5236 21532 5852 21588
rect 5908 21532 7532 21588
rect 7588 21532 8204 21588
rect 8260 21532 8270 21588
rect 10770 21532 10780 21588
rect 10836 21532 12796 21588
rect 12852 21532 12862 21588
rect 16370 21532 16380 21588
rect 16436 21532 19964 21588
rect 20020 21532 20030 21588
rect 31266 21532 31276 21588
rect 31332 21532 32508 21588
rect 32564 21532 32574 21588
rect 33618 21532 33628 21588
rect 33684 21532 34412 21588
rect 34468 21532 34478 21588
rect 44818 21532 44828 21588
rect 44884 21532 46732 21588
rect 46788 21532 46798 21588
rect 2482 21420 2492 21476
rect 2548 21420 4732 21476
rect 4788 21420 4798 21476
rect 11442 21420 11452 21476
rect 11508 21420 13916 21476
rect 13972 21420 13982 21476
rect 14140 21420 16156 21476
rect 16212 21420 16548 21476
rect 25218 21420 25228 21476
rect 25284 21420 26460 21476
rect 26516 21420 27804 21476
rect 27860 21420 28476 21476
rect 28532 21420 28542 21476
rect 31042 21420 31052 21476
rect 31108 21420 32284 21476
rect 32340 21420 35644 21476
rect 35700 21420 35710 21476
rect 36866 21420 36876 21476
rect 36932 21420 37212 21476
rect 37268 21420 37278 21476
rect 41794 21420 41804 21476
rect 41860 21420 42476 21476
rect 42532 21420 42542 21476
rect 44258 21420 44268 21476
rect 44324 21420 45276 21476
rect 45332 21420 47740 21476
rect 47796 21420 47806 21476
rect 14140 21364 14196 21420
rect 16492 21364 16548 21420
rect 7858 21308 7868 21364
rect 7924 21308 8204 21364
rect 8260 21308 9660 21364
rect 9716 21308 14196 21364
rect 14690 21308 14700 21364
rect 14756 21308 15484 21364
rect 15540 21308 15550 21364
rect 16482 21308 16492 21364
rect 16548 21308 16558 21364
rect 18386 21308 18396 21364
rect 18452 21308 26572 21364
rect 26628 21308 26638 21364
rect 31154 21308 31164 21364
rect 31220 21308 35980 21364
rect 36036 21308 36046 21364
rect 46274 21308 46284 21364
rect 46340 21308 47852 21364
rect 47908 21308 47918 21364
rect 17490 21196 17500 21252
rect 17556 21196 18060 21252
rect 18116 21196 18126 21252
rect 33954 21196 33964 21252
rect 34020 21196 34972 21252
rect 35028 21196 35038 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 14130 21084 14140 21140
rect 14196 21084 14812 21140
rect 14868 21084 14878 21140
rect 16930 21084 16940 21140
rect 16996 21084 19740 21140
rect 19796 21084 19806 21140
rect 3266 20972 3276 21028
rect 3332 20972 4620 21028
rect 4676 20972 5740 21028
rect 5796 20972 5806 21028
rect 10770 20972 10780 21028
rect 10836 20972 17164 21028
rect 17220 20972 19292 21028
rect 19348 20972 19358 21028
rect 24210 20972 24220 21028
rect 24276 20972 29484 21028
rect 29540 20972 30716 21028
rect 30772 20972 30782 21028
rect 13570 20860 13580 20916
rect 13636 20860 14588 20916
rect 14644 20860 15148 20916
rect 42914 20860 42924 20916
rect 42980 20860 43708 20916
rect 43764 20860 48188 20916
rect 48244 20860 48254 20916
rect 14018 20748 14028 20804
rect 14084 20748 14812 20804
rect 14868 20748 14878 20804
rect 15092 20748 15148 20860
rect 15204 20748 15214 20804
rect 20738 20748 20748 20804
rect 20804 20748 24892 20804
rect 24948 20748 24958 20804
rect 14812 20580 14868 20748
rect 18946 20636 18956 20692
rect 19012 20636 20636 20692
rect 20692 20636 20702 20692
rect 21410 20636 21420 20692
rect 21476 20636 23548 20692
rect 23604 20636 23772 20692
rect 23828 20636 23838 20692
rect 41234 20636 41244 20692
rect 41300 20636 41580 20692
rect 41636 20636 42812 20692
rect 42868 20636 42878 20692
rect 4946 20524 4956 20580
rect 5012 20524 9772 20580
rect 9828 20524 10444 20580
rect 10500 20524 10510 20580
rect 14812 20524 16604 20580
rect 16660 20524 16670 20580
rect 19730 20524 19740 20580
rect 19796 20524 22876 20580
rect 22932 20524 22942 20580
rect 29586 20524 29596 20580
rect 29652 20524 30268 20580
rect 30324 20524 30716 20580
rect 30772 20524 31164 20580
rect 31220 20524 31230 20580
rect 41458 20524 41468 20580
rect 41524 20524 42364 20580
rect 42420 20524 47180 20580
rect 47236 20524 47246 20580
rect 46162 20412 46172 20468
rect 46228 20412 46956 20468
rect 47012 20412 47022 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 20738 20300 20748 20356
rect 20804 20300 22540 20356
rect 22596 20300 22606 20356
rect 34514 20300 34524 20356
rect 34580 20300 35532 20356
rect 35588 20300 35598 20356
rect 41346 20300 41356 20356
rect 41412 20300 41804 20356
rect 41860 20300 41870 20356
rect 14578 20188 14588 20244
rect 14644 20188 16828 20244
rect 16884 20188 16894 20244
rect 27570 20188 27580 20244
rect 27636 20188 28364 20244
rect 28420 20188 29036 20244
rect 29092 20188 29484 20244
rect 29540 20188 29550 20244
rect 33282 20188 33292 20244
rect 33348 20188 34188 20244
rect 34244 20188 35084 20244
rect 35140 20188 35150 20244
rect 36530 20188 36540 20244
rect 36596 20188 37212 20244
rect 37268 20188 37278 20244
rect 42130 20188 42140 20244
rect 42196 20188 42206 20244
rect 42140 20132 42196 20188
rect 9762 20076 9772 20132
rect 9828 20076 10780 20132
rect 10836 20076 10846 20132
rect 12114 20076 12124 20132
rect 12180 20076 15596 20132
rect 15652 20076 15662 20132
rect 23874 20076 23884 20132
rect 23940 20076 25004 20132
rect 25060 20076 30380 20132
rect 30436 20076 30446 20132
rect 31826 20076 31836 20132
rect 31892 20076 33180 20132
rect 33236 20076 33246 20132
rect 33842 20076 33852 20132
rect 33908 20076 34748 20132
rect 34804 20076 41020 20132
rect 41076 20076 41086 20132
rect 41570 20076 41580 20132
rect 41636 20076 42196 20132
rect 9986 19964 9996 20020
rect 10052 19964 11004 20020
rect 11060 19964 11070 20020
rect 18834 19964 18844 20020
rect 18900 19964 26796 20020
rect 26852 19964 26862 20020
rect 27682 19964 27692 20020
rect 27748 19964 28364 20020
rect 28420 19964 28430 20020
rect 30930 19964 30940 20020
rect 30996 19964 33740 20020
rect 33796 19964 34300 20020
rect 34356 19964 34366 20020
rect 40002 19964 40012 20020
rect 40068 19964 41132 20020
rect 41188 19964 41198 20020
rect 42018 19964 42028 20020
rect 42084 19964 43372 20020
rect 43428 19964 43438 20020
rect 8194 19852 8204 19908
rect 8260 19852 8988 19908
rect 9044 19852 10892 19908
rect 10948 19852 15932 19908
rect 15988 19852 16380 19908
rect 16436 19852 22428 19908
rect 22484 19852 26348 19908
rect 26404 19852 26414 19908
rect 31490 19852 31500 19908
rect 31556 19852 31836 19908
rect 31892 19852 31902 19908
rect 32386 19852 32396 19908
rect 32452 19852 33516 19908
rect 33572 19852 33582 19908
rect 36082 19852 36092 19908
rect 36148 19852 37212 19908
rect 37268 19852 37278 19908
rect 40226 19852 40236 19908
rect 40292 19852 42588 19908
rect 42644 19852 42654 19908
rect 6514 19740 6524 19796
rect 6580 19740 7420 19796
rect 7476 19740 8764 19796
rect 8820 19740 8830 19796
rect 10434 19740 10444 19796
rect 10500 19740 11452 19796
rect 11508 19740 12012 19796
rect 12068 19740 12078 19796
rect 23090 19740 23100 19796
rect 23156 19740 24332 19796
rect 24388 19740 25004 19796
rect 25060 19740 25070 19796
rect 30482 19740 30492 19796
rect 30548 19740 31388 19796
rect 31444 19740 31454 19796
rect 31938 19740 31948 19796
rect 32004 19740 32284 19796
rect 32340 19740 32844 19796
rect 32900 19740 32910 19796
rect 39330 19740 39340 19796
rect 39396 19740 41468 19796
rect 41524 19740 41534 19796
rect 10546 19628 10556 19684
rect 10612 19628 13020 19684
rect 13076 19628 13086 19684
rect 30370 19628 30380 19684
rect 30436 19628 30446 19684
rect 40338 19628 40348 19684
rect 40404 19628 40908 19684
rect 40964 19628 40974 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 30380 19236 30436 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 1810 19180 1820 19236
rect 1876 19180 3388 19236
rect 3444 19180 5292 19236
rect 5348 19180 5740 19236
rect 5796 19180 5806 19236
rect 29250 19180 29260 19236
rect 29316 19180 30044 19236
rect 30100 19180 30110 19236
rect 30380 19180 30716 19236
rect 30772 19180 30782 19236
rect 33170 19180 33180 19236
rect 33236 19180 33516 19236
rect 33572 19180 33582 19236
rect 35410 19180 35420 19236
rect 35476 19180 36092 19236
rect 36148 19180 36158 19236
rect 41010 19180 41020 19236
rect 41076 19180 43932 19236
rect 43988 19180 44828 19236
rect 44884 19180 44894 19236
rect 2482 19068 2492 19124
rect 2548 19068 3388 19124
rect 4498 19068 4508 19124
rect 4564 19068 5628 19124
rect 5684 19068 5694 19124
rect 13794 19068 13804 19124
rect 13860 19068 14812 19124
rect 14868 19068 14878 19124
rect 30146 19068 30156 19124
rect 30212 19068 31556 19124
rect 33618 19068 33628 19124
rect 33684 19068 35532 19124
rect 35588 19068 35598 19124
rect 35746 19068 35756 19124
rect 35812 19068 40012 19124
rect 40068 19068 40078 19124
rect 3332 19012 3388 19068
rect 31500 19012 31556 19068
rect 3332 18956 5740 19012
rect 5796 18956 5806 19012
rect 6626 18956 6636 19012
rect 6692 18956 7644 19012
rect 7700 18956 7710 19012
rect 8194 18956 8204 19012
rect 8260 18956 8876 19012
rect 8932 18956 8942 19012
rect 13570 18956 13580 19012
rect 13636 18956 14364 19012
rect 14420 18956 15484 19012
rect 15540 18956 15550 19012
rect 29922 18956 29932 19012
rect 29988 18956 30940 19012
rect 30996 18956 31006 19012
rect 31490 18956 31500 19012
rect 31556 18956 40572 19012
rect 40628 18956 41132 19012
rect 41188 18956 41198 19012
rect 41682 18956 41692 19012
rect 41748 18956 42700 19012
rect 42756 18956 42766 19012
rect 28466 18844 28476 18900
rect 28532 18844 30044 18900
rect 30100 18844 30110 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 3602 18620 3612 18676
rect 3668 18620 4620 18676
rect 4676 18620 4686 18676
rect 18498 18620 18508 18676
rect 18564 18620 21868 18676
rect 21924 18620 21934 18676
rect 30706 18620 30716 18676
rect 30772 18620 35084 18676
rect 35140 18620 35150 18676
rect 43250 18620 43260 18676
rect 43316 18620 43326 18676
rect 22194 18508 22204 18564
rect 22260 18508 23212 18564
rect 23268 18508 23278 18564
rect 31462 18508 31500 18564
rect 31556 18508 31566 18564
rect 34290 18508 34300 18564
rect 34356 18508 34972 18564
rect 35028 18508 35420 18564
rect 35476 18508 35486 18564
rect 35858 18508 35868 18564
rect 35924 18508 39340 18564
rect 39396 18508 39406 18564
rect 43260 18452 43316 18620
rect 3154 18396 3164 18452
rect 3220 18396 4956 18452
rect 5012 18396 5628 18452
rect 5684 18396 5694 18452
rect 8306 18396 8316 18452
rect 8372 18396 9884 18452
rect 9940 18396 11452 18452
rect 11508 18396 12348 18452
rect 12404 18396 12796 18452
rect 12852 18396 12862 18452
rect 17826 18396 17836 18452
rect 17892 18396 19964 18452
rect 20020 18396 22316 18452
rect 22372 18396 22382 18452
rect 22642 18396 22652 18452
rect 22708 18396 22876 18452
rect 22932 18396 22942 18452
rect 25218 18396 25228 18452
rect 25284 18396 26348 18452
rect 26404 18396 26414 18452
rect 34626 18396 34636 18452
rect 34692 18396 34860 18452
rect 34916 18396 34926 18452
rect 37090 18396 37100 18452
rect 37156 18396 40908 18452
rect 40964 18396 40974 18452
rect 43260 18396 43708 18452
rect 43764 18396 43774 18452
rect 45378 18396 45388 18452
rect 45444 18396 46844 18452
rect 46900 18396 48076 18452
rect 48132 18396 48142 18452
rect 6962 18284 6972 18340
rect 7028 18284 8652 18340
rect 8708 18284 8718 18340
rect 16930 18284 16940 18340
rect 16996 18284 20860 18340
rect 20916 18284 20926 18340
rect 22876 18228 22932 18396
rect 24098 18284 24108 18340
rect 24164 18284 24556 18340
rect 24612 18284 27468 18340
rect 27524 18284 27534 18340
rect 34860 18228 34916 18396
rect 36306 18284 36316 18340
rect 36372 18284 37772 18340
rect 37828 18284 37838 18340
rect 45042 18284 45052 18340
rect 45108 18284 47068 18340
rect 47124 18284 47134 18340
rect 15922 18172 15932 18228
rect 15988 18172 17500 18228
rect 17556 18172 18620 18228
rect 18676 18172 18686 18228
rect 22876 18172 33180 18228
rect 33236 18172 33852 18228
rect 33908 18172 33918 18228
rect 34860 18172 38668 18228
rect 40338 18172 40348 18228
rect 40404 18172 41468 18228
rect 41524 18172 41534 18228
rect 38612 18116 38668 18172
rect 38612 18060 47852 18116
rect 47908 18060 47918 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 20850 17836 20860 17892
rect 20916 17836 23436 17892
rect 23492 17836 23502 17892
rect 28812 17836 34188 17892
rect 34244 17836 34254 17892
rect 43586 17836 43596 17892
rect 43652 17836 44940 17892
rect 44996 17836 45006 17892
rect 28812 17780 28868 17836
rect 14130 17724 14140 17780
rect 14196 17724 15708 17780
rect 15764 17724 15774 17780
rect 22754 17724 22764 17780
rect 22820 17724 23884 17780
rect 23940 17724 24332 17780
rect 24388 17724 24398 17780
rect 25750 17724 25788 17780
rect 25844 17724 26908 17780
rect 27682 17724 27692 17780
rect 27748 17724 28028 17780
rect 28084 17724 28812 17780
rect 28868 17724 28878 17780
rect 29138 17724 29148 17780
rect 29204 17724 30828 17780
rect 30884 17724 30894 17780
rect 34514 17724 34524 17780
rect 34580 17724 35644 17780
rect 35700 17724 35710 17780
rect 45602 17724 45612 17780
rect 45668 17724 47180 17780
rect 47236 17724 48524 17780
rect 48580 17724 48590 17780
rect 12002 17612 12012 17668
rect 12068 17612 13020 17668
rect 13076 17612 16156 17668
rect 16212 17612 17612 17668
rect 17668 17612 17678 17668
rect 19058 17612 19068 17668
rect 19124 17612 20524 17668
rect 20580 17612 20590 17668
rect 26852 17612 26908 17724
rect 26964 17612 28084 17668
rect 33954 17612 33964 17668
rect 34020 17612 35756 17668
rect 35812 17612 35822 17668
rect 41570 17612 41580 17668
rect 41636 17612 43820 17668
rect 43876 17612 43886 17668
rect 28028 17556 28084 17612
rect 49200 17556 50000 17584
rect 16258 17500 16268 17556
rect 16324 17500 17500 17556
rect 17556 17500 17566 17556
rect 19954 17500 19964 17556
rect 20020 17500 20300 17556
rect 20356 17500 21420 17556
rect 21476 17500 21486 17556
rect 26338 17500 26348 17556
rect 26404 17500 27244 17556
rect 27300 17500 27804 17556
rect 27860 17500 27870 17556
rect 28028 17500 34524 17556
rect 34580 17500 34590 17556
rect 35410 17500 35420 17556
rect 35476 17500 35644 17556
rect 35700 17500 35710 17556
rect 48178 17500 48188 17556
rect 48244 17500 50000 17556
rect 49200 17472 50000 17500
rect 4050 17388 4060 17444
rect 4116 17388 5628 17444
rect 5684 17388 5694 17444
rect 6850 17388 6860 17444
rect 6916 17388 9100 17444
rect 9156 17388 9166 17444
rect 22642 17388 22652 17444
rect 22708 17388 23660 17444
rect 23716 17388 23726 17444
rect 25442 17388 25452 17444
rect 25508 17388 27356 17444
rect 27412 17388 27422 17444
rect 32722 17388 32732 17444
rect 32788 17388 33180 17444
rect 33236 17388 33964 17444
rect 34020 17388 34030 17444
rect 31266 17276 31276 17332
rect 31332 17276 31836 17332
rect 31892 17276 31902 17332
rect 34850 17276 34860 17332
rect 34916 17276 36428 17332
rect 36484 17276 36494 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 16146 17052 16156 17108
rect 16212 17052 17388 17108
rect 17444 17052 17454 17108
rect 21858 17052 21868 17108
rect 21924 17052 22428 17108
rect 22484 17052 23100 17108
rect 23156 17052 25340 17108
rect 25396 17052 25406 17108
rect 31462 17052 31500 17108
rect 31556 17052 31566 17108
rect 31714 17052 31724 17108
rect 31780 17052 32284 17108
rect 32340 17052 32350 17108
rect 37426 17052 37436 17108
rect 37492 17052 38668 17108
rect 38724 17052 38734 17108
rect 40338 17052 40348 17108
rect 40404 17052 41916 17108
rect 41972 17052 41982 17108
rect 3378 16940 3388 16996
rect 3444 16940 4844 16996
rect 4900 16940 4910 16996
rect 11890 16940 11900 16996
rect 11956 16940 12908 16996
rect 12964 16940 12974 16996
rect 27346 16940 27356 16996
rect 27412 16940 28028 16996
rect 28084 16940 29708 16996
rect 29764 16940 29774 16996
rect 31154 16940 31164 16996
rect 31220 16940 31948 16996
rect 32004 16940 32014 16996
rect 40348 16884 40404 17052
rect 4274 16828 4284 16884
rect 4340 16828 4620 16884
rect 4676 16828 5404 16884
rect 5460 16828 5470 16884
rect 9202 16828 9212 16884
rect 9268 16828 9772 16884
rect 9828 16828 9838 16884
rect 10210 16828 10220 16884
rect 10276 16828 11340 16884
rect 11396 16828 11406 16884
rect 13906 16828 13916 16884
rect 13972 16828 15596 16884
rect 15652 16828 15662 16884
rect 18050 16828 18060 16884
rect 18116 16828 18396 16884
rect 18452 16828 21084 16884
rect 21140 16828 21150 16884
rect 24434 16828 24444 16884
rect 24500 16828 25228 16884
rect 25284 16828 27916 16884
rect 27972 16828 27982 16884
rect 30258 16828 30268 16884
rect 30324 16828 32060 16884
rect 32116 16828 33628 16884
rect 33684 16828 35084 16884
rect 35140 16828 35150 16884
rect 35634 16828 35644 16884
rect 35700 16828 36540 16884
rect 36596 16828 36606 16884
rect 37874 16828 37884 16884
rect 37940 16828 38556 16884
rect 38612 16828 40404 16884
rect 3714 16716 3724 16772
rect 3780 16716 4396 16772
rect 4452 16716 4462 16772
rect 11218 16716 11228 16772
rect 11284 16716 11900 16772
rect 11956 16716 11966 16772
rect 20962 16716 20972 16772
rect 21028 16716 21532 16772
rect 21588 16716 22764 16772
rect 22820 16716 23324 16772
rect 23380 16716 23390 16772
rect 31266 16716 31276 16772
rect 31332 16716 33292 16772
rect 33348 16716 33358 16772
rect 40226 16716 40236 16772
rect 40292 16716 41020 16772
rect 41076 16716 41086 16772
rect 19058 16604 19068 16660
rect 19124 16604 19740 16660
rect 19796 16604 20300 16660
rect 20356 16604 20366 16660
rect 28578 16604 28588 16660
rect 28644 16604 29708 16660
rect 29764 16604 29774 16660
rect 39890 16604 39900 16660
rect 39956 16604 41356 16660
rect 41412 16604 41422 16660
rect 42578 16604 42588 16660
rect 42644 16604 43372 16660
rect 43428 16604 43438 16660
rect 18274 16492 18284 16548
rect 18340 16492 19516 16548
rect 19572 16492 21308 16548
rect 21364 16492 21374 16548
rect 26898 16492 26908 16548
rect 26964 16492 33516 16548
rect 33572 16492 33582 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 4834 16380 4844 16436
rect 4900 16380 5180 16436
rect 5236 16380 5852 16436
rect 5908 16380 18060 16436
rect 18116 16380 18126 16436
rect 8866 16268 8876 16324
rect 8932 16268 9548 16324
rect 9604 16268 10108 16324
rect 10164 16268 10174 16324
rect 11778 16268 11788 16324
rect 11844 16268 12572 16324
rect 12628 16268 20020 16324
rect 20178 16268 20188 16324
rect 20244 16268 21196 16324
rect 21252 16268 21262 16324
rect 43362 16268 43372 16324
rect 43428 16268 44156 16324
rect 44212 16268 44222 16324
rect 19964 16212 20020 16268
rect 9202 16156 9212 16212
rect 9268 16156 9660 16212
rect 9716 16156 10780 16212
rect 10836 16156 12348 16212
rect 12404 16156 12414 16212
rect 18386 16156 18396 16212
rect 18452 16156 19628 16212
rect 19684 16156 19694 16212
rect 19964 16156 20860 16212
rect 20916 16156 21868 16212
rect 21924 16156 21934 16212
rect 27122 16156 27132 16212
rect 27188 16156 28140 16212
rect 28196 16156 29148 16212
rect 29204 16156 29214 16212
rect 36754 16156 36764 16212
rect 36820 16156 37772 16212
rect 37828 16156 37838 16212
rect 38882 16156 38892 16212
rect 38948 16156 39788 16212
rect 39844 16156 39854 16212
rect 46274 16156 46284 16212
rect 46340 16156 47404 16212
rect 47460 16156 47470 16212
rect 3378 16044 3388 16100
rect 3444 16044 3836 16100
rect 3892 16044 3902 16100
rect 5954 16044 5964 16100
rect 6020 16044 6412 16100
rect 6468 16044 12012 16100
rect 12068 16044 13580 16100
rect 13636 16044 15148 16100
rect 15204 16044 15214 16100
rect 18162 16044 18172 16100
rect 18228 16044 19068 16100
rect 19124 16044 19134 16100
rect 19282 16044 19292 16100
rect 19348 16044 21532 16100
rect 21588 16044 21598 16100
rect 22306 16044 22316 16100
rect 22372 16044 24668 16100
rect 24724 16044 24734 16100
rect 28578 16044 28588 16100
rect 28644 16044 29260 16100
rect 29316 16044 29326 16100
rect 36418 16044 36428 16100
rect 36484 16044 36876 16100
rect 36932 16044 36942 16100
rect 28466 15932 28476 15988
rect 28532 15932 30716 15988
rect 30772 15932 31276 15988
rect 31332 15932 31342 15988
rect 14466 15820 14476 15876
rect 14532 15820 15708 15876
rect 15764 15820 15774 15876
rect 17714 15820 17724 15876
rect 17780 15820 18396 15876
rect 18452 15820 18462 15876
rect 20402 15820 20412 15876
rect 20468 15820 23996 15876
rect 24052 15820 24062 15876
rect 27010 15820 27020 15876
rect 27076 15820 27356 15876
rect 27412 15820 29596 15876
rect 29652 15820 29662 15876
rect 29810 15820 29820 15876
rect 29876 15820 30268 15876
rect 30324 15820 30334 15876
rect 34514 15820 34524 15876
rect 34580 15820 37772 15876
rect 37828 15820 39116 15876
rect 39172 15820 39182 15876
rect 44790 15820 44828 15876
rect 44884 15820 44894 15876
rect 35410 15708 35420 15764
rect 35476 15708 35756 15764
rect 35812 15708 39564 15764
rect 39620 15708 39630 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 34178 15596 34188 15652
rect 34244 15596 37100 15652
rect 37156 15596 37166 15652
rect 9202 15484 9212 15540
rect 9268 15484 9772 15540
rect 9828 15484 9838 15540
rect 10658 15484 10668 15540
rect 10724 15484 11788 15540
rect 11844 15484 11854 15540
rect 17938 15484 17948 15540
rect 18004 15484 18844 15540
rect 18900 15484 19404 15540
rect 19460 15484 19470 15540
rect 19618 15484 19628 15540
rect 19684 15484 19964 15540
rect 20020 15484 20030 15540
rect 20178 15484 20188 15540
rect 20244 15484 20972 15540
rect 21028 15484 21038 15540
rect 23426 15484 23436 15540
rect 23492 15484 24444 15540
rect 24500 15484 24510 15540
rect 26002 15484 26012 15540
rect 26068 15484 27692 15540
rect 27748 15484 27758 15540
rect 31490 15484 31500 15540
rect 31556 15484 31836 15540
rect 31892 15484 31902 15540
rect 35746 15484 35756 15540
rect 35812 15484 40012 15540
rect 40068 15484 40078 15540
rect 18274 15372 18284 15428
rect 18340 15372 19740 15428
rect 19796 15372 20748 15428
rect 20804 15372 20814 15428
rect 31714 15372 31724 15428
rect 31780 15372 33404 15428
rect 33460 15372 33470 15428
rect 36082 15372 36092 15428
rect 36148 15372 37212 15428
rect 37268 15372 37278 15428
rect 46722 15372 46732 15428
rect 46788 15372 47404 15428
rect 47460 15372 47470 15428
rect 5506 15260 5516 15316
rect 5572 15260 6412 15316
rect 6468 15260 6478 15316
rect 6850 15260 6860 15316
rect 6916 15260 10556 15316
rect 10612 15260 10622 15316
rect 19506 15260 19516 15316
rect 19572 15260 20636 15316
rect 20692 15260 20702 15316
rect 22530 15260 22540 15316
rect 22596 15260 24780 15316
rect 24836 15260 24846 15316
rect 25890 15260 25900 15316
rect 25956 15260 27916 15316
rect 27972 15260 27982 15316
rect 28130 15260 28140 15316
rect 28196 15260 28588 15316
rect 28644 15260 28654 15316
rect 30594 15260 30604 15316
rect 30660 15260 33516 15316
rect 33572 15260 34804 15316
rect 36418 15260 36428 15316
rect 36484 15260 38332 15316
rect 38388 15260 38398 15316
rect 34748 15204 34804 15260
rect 1810 15148 1820 15204
rect 1876 15148 6076 15204
rect 6132 15148 7308 15204
rect 7364 15148 7374 15204
rect 9650 15148 9660 15204
rect 9716 15148 10444 15204
rect 10500 15148 10510 15204
rect 19618 15148 19628 15204
rect 19684 15148 20860 15204
rect 20916 15148 20926 15204
rect 25778 15148 25788 15204
rect 25844 15148 26236 15204
rect 26292 15148 28476 15204
rect 28532 15148 28542 15204
rect 34738 15148 34748 15204
rect 34804 15148 37660 15204
rect 37716 15148 37726 15204
rect 39554 15148 39564 15204
rect 39620 15148 40908 15204
rect 40964 15148 40974 15204
rect 41458 15148 41468 15204
rect 41524 15148 43036 15204
rect 43092 15148 43102 15204
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 40562 14700 40572 14756
rect 40628 14700 43484 14756
rect 43540 14700 45500 14756
rect 45556 14700 45566 14756
rect 15474 14588 15484 14644
rect 15540 14588 15708 14644
rect 15764 14588 24220 14644
rect 24276 14588 24286 14644
rect 24994 14588 25004 14644
rect 25060 14588 26460 14644
rect 26516 14588 26526 14644
rect 33730 14588 33740 14644
rect 33796 14588 34748 14644
rect 34804 14588 35308 14644
rect 35364 14588 35756 14644
rect 35812 14588 35822 14644
rect 41346 14588 41356 14644
rect 41412 14588 42924 14644
rect 42980 14588 43596 14644
rect 43652 14588 43662 14644
rect 4386 14476 4396 14532
rect 4452 14476 4956 14532
rect 5012 14476 5022 14532
rect 21746 14476 21756 14532
rect 21812 14476 24108 14532
rect 24164 14476 24174 14532
rect 32946 14476 32956 14532
rect 33012 14476 35868 14532
rect 35924 14476 35934 14532
rect 37202 14476 37212 14532
rect 37268 14476 38220 14532
rect 38276 14476 39004 14532
rect 39060 14476 39070 14532
rect 39890 14476 39900 14532
rect 39956 14476 40460 14532
rect 40516 14476 40526 14532
rect 41570 14476 41580 14532
rect 41636 14476 43148 14532
rect 43204 14476 45388 14532
rect 45444 14476 45454 14532
rect 45602 14476 45612 14532
rect 45668 14476 46732 14532
rect 46788 14476 46798 14532
rect 12562 14364 12572 14420
rect 12628 14364 13468 14420
rect 13524 14364 13534 14420
rect 14018 14364 14028 14420
rect 14084 14364 14924 14420
rect 14980 14364 14990 14420
rect 18386 14364 18396 14420
rect 18452 14364 20300 14420
rect 20356 14364 20366 14420
rect 28018 14364 28028 14420
rect 28084 14364 30156 14420
rect 30212 14364 30222 14420
rect 35970 14364 35980 14420
rect 36036 14364 37324 14420
rect 37380 14364 37390 14420
rect 44482 14364 44492 14420
rect 44548 14364 46172 14420
rect 46228 14364 46238 14420
rect 12236 14252 12908 14308
rect 12964 14252 14700 14308
rect 14756 14252 14766 14308
rect 16594 14252 16604 14308
rect 16660 14252 19516 14308
rect 19572 14252 19582 14308
rect 28354 14252 28364 14308
rect 28420 14252 29932 14308
rect 29988 14252 29998 14308
rect 36082 14252 36092 14308
rect 36148 14252 37436 14308
rect 37492 14252 37502 14308
rect 38770 14252 38780 14308
rect 38836 14252 39452 14308
rect 39508 14252 39518 14308
rect 41682 14252 41692 14308
rect 41748 14252 42028 14308
rect 42084 14252 42094 14308
rect 46498 14252 46508 14308
rect 46564 14252 47404 14308
rect 47460 14252 47470 14308
rect 12236 14196 12292 14252
rect 12226 14140 12236 14196
rect 12292 14140 12302 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 36642 14028 36652 14084
rect 36708 14028 40236 14084
rect 40292 14028 41020 14084
rect 41076 14028 45164 14084
rect 45220 14028 45230 14084
rect 26450 13916 26460 13972
rect 26516 13916 28364 13972
rect 28420 13916 28430 13972
rect 42812 13916 44044 13972
rect 44100 13916 44110 13972
rect 8372 13804 21308 13860
rect 21364 13804 22428 13860
rect 22484 13804 22494 13860
rect 38546 13804 38556 13860
rect 38612 13804 39228 13860
rect 39284 13804 39294 13860
rect 8372 13748 8428 13804
rect 42812 13748 42868 13916
rect 7074 13692 7084 13748
rect 7140 13692 7532 13748
rect 7588 13692 8428 13748
rect 15092 13692 15260 13748
rect 15316 13692 17948 13748
rect 18004 13692 23212 13748
rect 23268 13692 23278 13748
rect 24434 13692 24444 13748
rect 24500 13692 27356 13748
rect 27412 13692 27422 13748
rect 30146 13692 30156 13748
rect 30212 13692 31052 13748
rect 31108 13692 31388 13748
rect 31444 13692 31454 13748
rect 31826 13692 31836 13748
rect 31892 13692 33180 13748
rect 33236 13692 35644 13748
rect 35700 13692 35710 13748
rect 38994 13692 39004 13748
rect 39060 13692 39676 13748
rect 39732 13692 39742 13748
rect 42802 13692 42812 13748
rect 42868 13692 42878 13748
rect 43362 13692 43372 13748
rect 43428 13692 43932 13748
rect 43988 13692 43998 13748
rect 15092 13636 15148 13692
rect 9090 13580 9100 13636
rect 9156 13580 12012 13636
rect 12068 13580 12078 13636
rect 13794 13580 13804 13636
rect 13860 13580 15148 13636
rect 23874 13580 23884 13636
rect 23940 13580 24892 13636
rect 24948 13580 25340 13636
rect 25396 13580 25406 13636
rect 31714 13580 31724 13636
rect 31780 13580 32396 13636
rect 32452 13580 32462 13636
rect 17938 13468 17948 13524
rect 18004 13468 21084 13524
rect 21140 13468 21150 13524
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 34972 13300 35028 13692
rect 37426 13580 37436 13636
rect 37492 13580 37772 13636
rect 37828 13580 37838 13636
rect 40114 13580 40124 13636
rect 40180 13580 42476 13636
rect 42532 13580 43036 13636
rect 43092 13580 43708 13636
rect 43764 13580 43774 13636
rect 37090 13468 37100 13524
rect 37156 13468 42588 13524
rect 42644 13468 43820 13524
rect 43876 13468 43886 13524
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 11218 13244 11228 13300
rect 11284 13244 11676 13300
rect 11732 13244 11742 13300
rect 32050 13244 32060 13300
rect 32116 13244 34412 13300
rect 34468 13244 34478 13300
rect 34962 13244 34972 13300
rect 35028 13244 35038 13300
rect 2482 13132 2492 13188
rect 2548 13132 3724 13188
rect 3780 13132 3790 13188
rect 8372 13132 18508 13188
rect 18564 13132 19516 13188
rect 19572 13132 21308 13188
rect 21364 13132 21374 13188
rect 26572 13132 29484 13188
rect 29540 13132 29550 13188
rect 36530 13132 36540 13188
rect 36596 13132 37324 13188
rect 37380 13132 38108 13188
rect 38164 13132 38174 13188
rect 41906 13132 41916 13188
rect 41972 13132 45276 13188
rect 45332 13132 45342 13188
rect 8372 13076 8428 13132
rect 7074 13020 7084 13076
rect 7140 13020 7756 13076
rect 7812 13020 8428 13076
rect 12114 13020 12124 13076
rect 12180 13020 16268 13076
rect 16324 13020 16716 13076
rect 16772 13020 16782 13076
rect 26572 12964 26628 13132
rect 27682 13020 27692 13076
rect 27748 13020 29372 13076
rect 29428 13020 29438 13076
rect 40450 13020 40460 13076
rect 40516 13020 41804 13076
rect 41860 13020 41870 13076
rect 5282 12908 5292 12964
rect 5348 12908 6860 12964
rect 6916 12908 6926 12964
rect 7298 12908 7308 12964
rect 7364 12908 8316 12964
rect 8372 12908 8764 12964
rect 8820 12908 8830 12964
rect 17714 12908 17724 12964
rect 17780 12908 18844 12964
rect 18900 12908 19852 12964
rect 19908 12908 19918 12964
rect 20290 12908 20300 12964
rect 20356 12908 20524 12964
rect 20580 12908 20590 12964
rect 23314 12908 23324 12964
rect 23380 12908 26572 12964
rect 26628 12908 26638 12964
rect 42802 12908 42812 12964
rect 42868 12908 43596 12964
rect 43652 12908 43662 12964
rect 44258 12908 44268 12964
rect 44324 12908 45388 12964
rect 45444 12908 45454 12964
rect 20300 12852 20356 12908
rect 3826 12796 3836 12852
rect 3892 12796 4284 12852
rect 4340 12796 4732 12852
rect 4788 12796 5628 12852
rect 5684 12796 5694 12852
rect 15250 12796 15260 12852
rect 15316 12796 15596 12852
rect 15652 12796 15662 12852
rect 18162 12796 18172 12852
rect 18228 12796 18508 12852
rect 18564 12796 20356 12852
rect 25900 12796 26908 12852
rect 26964 12796 26974 12852
rect 27234 12796 27244 12852
rect 27300 12796 29708 12852
rect 29764 12796 30716 12852
rect 30772 12796 30782 12852
rect 34150 12796 34188 12852
rect 34244 12796 34254 12852
rect 34962 12796 34972 12852
rect 35028 12796 36204 12852
rect 36260 12796 36270 12852
rect 36866 12796 36876 12852
rect 36932 12796 47852 12852
rect 47908 12796 47918 12852
rect 25900 12740 25956 12796
rect 4834 12684 4844 12740
rect 4900 12684 5740 12740
rect 5796 12684 5806 12740
rect 7186 12684 7196 12740
rect 7252 12684 8092 12740
rect 8148 12684 8158 12740
rect 20850 12684 20860 12740
rect 20916 12684 21868 12740
rect 21924 12684 21934 12740
rect 22530 12684 22540 12740
rect 22596 12684 24108 12740
rect 24164 12684 24174 12740
rect 25890 12684 25900 12740
rect 25956 12684 25966 12740
rect 26236 12684 26460 12740
rect 26516 12684 26526 12740
rect 29138 12684 29148 12740
rect 29204 12684 29820 12740
rect 29876 12684 30604 12740
rect 30660 12684 30670 12740
rect 33618 12684 33628 12740
rect 33684 12684 33964 12740
rect 34020 12684 34524 12740
rect 34580 12684 34590 12740
rect 40114 12684 40124 12740
rect 40180 12684 40908 12740
rect 40964 12684 40974 12740
rect 41794 12684 41804 12740
rect 41860 12684 42252 12740
rect 42308 12684 42318 12740
rect 43026 12684 43036 12740
rect 43092 12684 44268 12740
rect 44324 12684 44334 12740
rect 46386 12684 46396 12740
rect 46452 12684 47404 12740
rect 47460 12684 47470 12740
rect 26236 12628 26292 12684
rect 49200 12628 50000 12656
rect 25442 12572 25452 12628
rect 25508 12572 26292 12628
rect 34402 12572 34412 12628
rect 34468 12572 35084 12628
rect 35140 12572 35150 12628
rect 40226 12572 40236 12628
rect 40292 12572 41132 12628
rect 41188 12572 41916 12628
rect 41972 12572 41982 12628
rect 42130 12572 42140 12628
rect 42196 12572 42700 12628
rect 42756 12572 43092 12628
rect 47618 12572 47628 12628
rect 47684 12572 48188 12628
rect 48244 12572 50000 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 43036 12516 43092 12572
rect 49200 12544 50000 12572
rect 25218 12460 25228 12516
rect 25284 12460 26124 12516
rect 26180 12460 26190 12516
rect 34290 12460 34300 12516
rect 34356 12460 34412 12516
rect 34468 12460 34478 12516
rect 43026 12460 43036 12516
rect 43092 12460 43102 12516
rect 6290 12348 6300 12404
rect 6356 12348 9604 12404
rect 9874 12348 9884 12404
rect 9940 12348 10332 12404
rect 10388 12348 11340 12404
rect 11396 12348 11406 12404
rect 31378 12348 31388 12404
rect 31444 12348 32060 12404
rect 32116 12348 32126 12404
rect 41906 12348 41916 12404
rect 41972 12348 42476 12404
rect 42532 12348 42542 12404
rect 9548 12292 9604 12348
rect 6962 12236 6972 12292
rect 7028 12236 8428 12292
rect 9538 12236 9548 12292
rect 9604 12236 9614 12292
rect 11666 12236 11676 12292
rect 11732 12236 12684 12292
rect 12740 12236 12750 12292
rect 24658 12236 24668 12292
rect 24724 12236 25788 12292
rect 25844 12236 25854 12292
rect 26674 12236 26684 12292
rect 26740 12236 27804 12292
rect 27860 12236 29036 12292
rect 29092 12236 29102 12292
rect 30482 12236 30492 12292
rect 30548 12236 31276 12292
rect 31332 12236 31342 12292
rect 34150 12236 34188 12292
rect 34244 12236 34254 12292
rect 8372 12180 8428 12236
rect 8372 12124 12012 12180
rect 12068 12124 12078 12180
rect 29810 12124 29820 12180
rect 29876 12124 30940 12180
rect 30996 12124 31006 12180
rect 37090 12124 37100 12180
rect 37156 12124 37324 12180
rect 37380 12124 37390 12180
rect 38658 12124 38668 12180
rect 38724 12124 39452 12180
rect 39508 12124 39518 12180
rect 42242 12124 42252 12180
rect 42308 12124 42700 12180
rect 42756 12124 42766 12180
rect 4610 12012 4620 12068
rect 4676 12012 5516 12068
rect 5572 12012 5582 12068
rect 13346 12012 13356 12068
rect 13412 12012 14028 12068
rect 14084 12012 14094 12068
rect 16706 12012 16716 12068
rect 16772 12012 17836 12068
rect 17892 12012 17902 12068
rect 23426 12012 23436 12068
rect 23492 12012 25676 12068
rect 25732 12012 26236 12068
rect 26292 12012 26302 12068
rect 36194 12012 36204 12068
rect 36260 12012 36988 12068
rect 37044 12012 37548 12068
rect 37604 12012 38444 12068
rect 38500 12012 38510 12068
rect 41570 12012 41580 12068
rect 41636 12012 42140 12068
rect 42196 12012 42924 12068
rect 42980 12012 45276 12068
rect 45332 12012 45342 12068
rect 15586 11900 15596 11956
rect 15652 11900 22204 11956
rect 22260 11900 22270 11956
rect 23762 11900 23772 11956
rect 23828 11900 25228 11956
rect 25284 11900 25294 11956
rect 44604 11900 44828 11956
rect 44884 11900 44894 11956
rect 5058 11788 5068 11844
rect 5124 11788 5964 11844
rect 6020 11788 6030 11844
rect 20188 11788 21420 11844
rect 21476 11788 21486 11844
rect 31938 11788 31948 11844
rect 32004 11788 33292 11844
rect 33348 11788 33358 11844
rect 44604 11788 44660 11900
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 20188 11732 20244 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 44594 11732 44604 11788
rect 44660 11732 44670 11788
rect 11666 11676 11676 11732
rect 11732 11676 13804 11732
rect 13860 11676 13870 11732
rect 16258 11676 16268 11732
rect 16324 11676 18172 11732
rect 18228 11676 20244 11732
rect 9874 11564 9884 11620
rect 9940 11564 10444 11620
rect 10500 11564 10892 11620
rect 10948 11564 10958 11620
rect 45126 11564 45164 11620
rect 45220 11564 45230 11620
rect 2482 11452 2492 11508
rect 2548 11452 4396 11508
rect 4452 11452 4462 11508
rect 33842 11452 33852 11508
rect 33908 11452 34748 11508
rect 34804 11452 34972 11508
rect 35028 11452 35038 11508
rect 37090 11452 37100 11508
rect 37156 11452 38668 11508
rect 38612 11396 38668 11452
rect 4610 11340 4620 11396
rect 4676 11340 5516 11396
rect 5572 11340 5582 11396
rect 11106 11340 11116 11396
rect 11172 11340 12124 11396
rect 12180 11340 15148 11396
rect 15362 11340 15372 11396
rect 15428 11340 19068 11396
rect 19124 11340 19134 11396
rect 33954 11340 33964 11396
rect 34020 11340 37660 11396
rect 37716 11340 37996 11396
rect 38052 11340 38062 11396
rect 38612 11340 39340 11396
rect 39396 11340 39406 11396
rect 39778 11340 39788 11396
rect 39844 11340 40796 11396
rect 40852 11340 40862 11396
rect 41916 11340 44492 11396
rect 44548 11340 45276 11396
rect 45332 11340 46732 11396
rect 46788 11340 46798 11396
rect 15092 11284 15148 11340
rect 8082 11228 8092 11284
rect 8148 11228 9660 11284
rect 9716 11228 9726 11284
rect 11554 11228 11564 11284
rect 11620 11228 12236 11284
rect 12292 11228 12302 11284
rect 15092 11228 15596 11284
rect 15652 11228 16604 11284
rect 16660 11228 16670 11284
rect 40226 11228 40236 11284
rect 40292 11228 40908 11284
rect 40964 11228 40974 11284
rect 9538 11116 9548 11172
rect 9604 11116 9996 11172
rect 10052 11116 10668 11172
rect 10724 11116 10734 11172
rect 30818 11116 30828 11172
rect 30884 11116 30894 11172
rect 35186 11116 35196 11172
rect 35252 11116 36652 11172
rect 36708 11116 36718 11172
rect 38322 11116 38332 11172
rect 38388 11116 40124 11172
rect 40180 11116 40190 11172
rect 21858 11004 21868 11060
rect 21924 11004 22764 11060
rect 22820 11004 26908 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 26852 10836 26908 11004
rect 30828 10948 30884 11116
rect 33394 11004 33404 11060
rect 33460 11004 34412 11060
rect 34468 11004 35532 11060
rect 35588 11004 35598 11060
rect 38210 11004 38220 11060
rect 38276 11004 41020 11060
rect 41076 11004 41086 11060
rect 41916 10948 41972 11340
rect 42690 11228 42700 11284
rect 42756 11228 43932 11284
rect 43988 11228 43998 11284
rect 43586 11116 43596 11172
rect 43652 11116 44716 11172
rect 44772 11116 44782 11172
rect 42130 11004 42140 11060
rect 42196 11004 45164 11060
rect 45220 11004 45230 11060
rect 30828 10892 41972 10948
rect 10098 10780 10108 10836
rect 10164 10780 11004 10836
rect 11060 10780 11070 10836
rect 20402 10780 20412 10836
rect 20468 10780 21532 10836
rect 21588 10780 21598 10836
rect 26852 10780 32284 10836
rect 32340 10780 32350 10836
rect 32610 10780 32620 10836
rect 32676 10780 33628 10836
rect 33684 10780 33694 10836
rect 36418 10780 36428 10836
rect 36484 10780 37660 10836
rect 37716 10780 38668 10836
rect 41458 10780 41468 10836
rect 41524 10780 42028 10836
rect 42084 10780 42094 10836
rect 38612 10724 38668 10780
rect 9538 10668 9548 10724
rect 9604 10668 11116 10724
rect 11172 10668 11182 10724
rect 30482 10668 30492 10724
rect 30548 10668 36652 10724
rect 36708 10668 36718 10724
rect 37874 10668 37884 10724
rect 37940 10668 38220 10724
rect 38276 10668 38286 10724
rect 38612 10668 40684 10724
rect 40740 10668 41860 10724
rect 41804 10612 41860 10668
rect 3938 10556 3948 10612
rect 4004 10556 5180 10612
rect 5236 10556 5246 10612
rect 7186 10556 7196 10612
rect 7252 10556 9996 10612
rect 10052 10556 10332 10612
rect 10388 10556 10398 10612
rect 10882 10556 10892 10612
rect 10948 10556 12236 10612
rect 12292 10556 12302 10612
rect 12674 10556 12684 10612
rect 12740 10556 15372 10612
rect 15428 10556 15438 10612
rect 35746 10556 35756 10612
rect 35812 10556 37100 10612
rect 37156 10556 37166 10612
rect 41794 10556 41804 10612
rect 41860 10556 43484 10612
rect 43540 10556 43550 10612
rect 1698 10444 1708 10500
rect 1764 10444 3612 10500
rect 3668 10444 3678 10500
rect 3826 10444 3836 10500
rect 3892 10444 5068 10500
rect 5124 10444 5134 10500
rect 24994 10444 25004 10500
rect 25060 10444 25676 10500
rect 25732 10444 25742 10500
rect 34290 10444 34300 10500
rect 34356 10444 34860 10500
rect 34916 10444 39004 10500
rect 39060 10444 39070 10500
rect 3490 10332 3500 10388
rect 3556 10332 4956 10388
rect 5012 10332 5022 10388
rect 31490 10332 31500 10388
rect 31556 10332 32396 10388
rect 32452 10332 32462 10388
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 13122 10108 13132 10164
rect 13188 10108 18452 10164
rect 32274 10108 32284 10164
rect 32340 10108 32350 10164
rect 38612 10108 41692 10164
rect 41748 10108 41758 10164
rect 18396 10052 18452 10108
rect 32284 10052 32340 10108
rect 38612 10052 38668 10108
rect 4386 9996 4396 10052
rect 4452 9996 5068 10052
rect 5124 9996 5964 10052
rect 6020 9996 6030 10052
rect 12450 9996 12460 10052
rect 12516 9996 13580 10052
rect 13636 9996 13646 10052
rect 18396 9996 23436 10052
rect 23492 9996 25116 10052
rect 25172 9996 25182 10052
rect 32284 9996 38668 10052
rect 4834 9884 4844 9940
rect 4900 9884 5628 9940
rect 5684 9884 5694 9940
rect 6738 9884 6748 9940
rect 6804 9884 7196 9940
rect 7252 9884 8540 9940
rect 8596 9884 8606 9940
rect 34412 9884 34636 9940
rect 34692 9884 35980 9940
rect 36036 9884 36046 9940
rect 38322 9884 38332 9940
rect 38388 9884 38892 9940
rect 38948 9884 38958 9940
rect 43362 9884 43372 9940
rect 43428 9884 43932 9940
rect 43988 9884 45276 9940
rect 45332 9884 45342 9940
rect 46274 9884 46284 9940
rect 46340 9884 47404 9940
rect 47460 9884 47470 9940
rect 3378 9772 3388 9828
rect 3444 9772 3724 9828
rect 3780 9772 3790 9828
rect 20962 9772 20972 9828
rect 21028 9772 21532 9828
rect 21588 9772 21868 9828
rect 21924 9772 21934 9828
rect 26226 9772 26236 9828
rect 26292 9772 27580 9828
rect 27636 9772 27646 9828
rect 10994 9660 11004 9716
rect 11060 9660 12572 9716
rect 12628 9660 12638 9716
rect 17266 9660 17276 9716
rect 17332 9660 18844 9716
rect 18900 9660 18910 9716
rect 27458 9660 27468 9716
rect 27524 9660 28700 9716
rect 28756 9660 28766 9716
rect 34412 9604 34468 9884
rect 34962 9772 34972 9828
rect 35028 9772 36204 9828
rect 36260 9772 36270 9828
rect 36418 9772 36428 9828
rect 36484 9772 38444 9828
rect 38500 9772 38510 9828
rect 35410 9660 35420 9716
rect 35476 9660 35756 9716
rect 35812 9660 35822 9716
rect 10434 9548 10444 9604
rect 10500 9548 10780 9604
rect 10836 9548 10846 9604
rect 18722 9548 18732 9604
rect 18788 9548 21644 9604
rect 21700 9548 21710 9604
rect 26114 9548 26124 9604
rect 26180 9548 27916 9604
rect 27972 9548 30716 9604
rect 30772 9548 31948 9604
rect 32004 9548 32014 9604
rect 34374 9548 34412 9604
rect 34468 9548 34478 9604
rect 35186 9548 35196 9604
rect 35252 9548 35868 9604
rect 35924 9548 37100 9604
rect 37156 9548 37166 9604
rect 41458 9548 41468 9604
rect 41524 9548 42140 9604
rect 42196 9548 43148 9604
rect 43204 9548 43214 9604
rect 43362 9548 43372 9604
rect 43428 9548 44268 9604
rect 44324 9548 44334 9604
rect 20514 9436 20524 9492
rect 20580 9436 21532 9492
rect 21588 9436 21598 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 6066 9212 6076 9268
rect 6132 9212 7308 9268
rect 7364 9212 7374 9268
rect 16818 9212 16828 9268
rect 16884 9212 17500 9268
rect 17556 9212 17566 9268
rect 32498 9212 32508 9268
rect 32564 9212 33516 9268
rect 33572 9212 33582 9268
rect 35186 9212 35196 9268
rect 35252 9212 36092 9268
rect 36148 9212 36158 9268
rect 42466 9212 42476 9268
rect 42532 9212 42924 9268
rect 42980 9212 44604 9268
rect 44660 9212 44670 9268
rect 6402 9100 6412 9156
rect 6468 9100 7196 9156
rect 7252 9100 7262 9156
rect 16034 9100 16044 9156
rect 16100 9100 17388 9156
rect 17444 9100 17454 9156
rect 25442 9100 25452 9156
rect 25508 9100 25900 9156
rect 25956 9100 25966 9156
rect 35298 9100 35308 9156
rect 35364 9100 36204 9156
rect 36260 9100 36270 9156
rect 40338 9100 40348 9156
rect 40404 9100 41132 9156
rect 41188 9100 43036 9156
rect 43092 9100 43102 9156
rect 27122 8988 27132 9044
rect 27188 8988 29596 9044
rect 29652 8988 30828 9044
rect 30884 8988 30894 9044
rect 32162 8988 32172 9044
rect 32228 8988 33292 9044
rect 33348 8988 33358 9044
rect 39666 8988 39676 9044
rect 39732 8988 41356 9044
rect 41412 8988 42140 9044
rect 42196 8988 42206 9044
rect 43138 8988 43148 9044
rect 43204 8988 44268 9044
rect 44324 8988 44334 9044
rect 21186 8876 21196 8932
rect 21252 8876 21980 8932
rect 22036 8876 22652 8932
rect 22708 8876 22718 8932
rect 26002 8876 26012 8932
rect 26068 8876 27020 8932
rect 27076 8876 29148 8932
rect 29204 8876 29214 8932
rect 34066 8876 34076 8932
rect 34132 8876 34972 8932
rect 35028 8876 35038 8932
rect 42242 8876 42252 8932
rect 42308 8876 45276 8932
rect 45332 8876 45342 8932
rect 46498 8876 46508 8932
rect 46564 8876 47404 8932
rect 47460 8876 47470 8932
rect 7746 8764 7756 8820
rect 7812 8764 8540 8820
rect 8596 8764 8606 8820
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 37090 8540 37100 8596
rect 37156 8540 38668 8596
rect 38724 8540 38734 8596
rect 12114 8428 12124 8484
rect 12180 8428 13580 8484
rect 13636 8428 13646 8484
rect 13794 8428 13804 8484
rect 13860 8428 14140 8484
rect 14196 8428 16044 8484
rect 16100 8428 16604 8484
rect 16660 8428 16670 8484
rect 20850 8428 20860 8484
rect 20916 8428 22428 8484
rect 22484 8428 22494 8484
rect 36530 8428 36540 8484
rect 36596 8428 40348 8484
rect 40404 8428 40414 8484
rect 44818 8428 44828 8484
rect 44884 8428 47180 8484
rect 47236 8428 47246 8484
rect 19170 8316 19180 8372
rect 19236 8316 21420 8372
rect 21476 8316 21486 8372
rect 23874 8316 23884 8372
rect 23940 8316 24556 8372
rect 24612 8316 24622 8372
rect 27794 8316 27804 8372
rect 27860 8316 29260 8372
rect 29316 8316 29326 8372
rect 34290 8316 34300 8372
rect 34356 8316 35196 8372
rect 35252 8316 35644 8372
rect 35700 8316 35710 8372
rect 36642 8316 36652 8372
rect 36708 8316 37212 8372
rect 37268 8316 37278 8372
rect 37426 8316 37436 8372
rect 37492 8316 38332 8372
rect 38388 8316 38398 8372
rect 39778 8316 39788 8372
rect 39844 8316 40908 8372
rect 40964 8316 40974 8372
rect 43810 8316 43820 8372
rect 43876 8316 44716 8372
rect 44772 8316 46844 8372
rect 46900 8316 46910 8372
rect 37212 8260 37268 8316
rect 1810 8204 1820 8260
rect 1876 8204 5516 8260
rect 5572 8204 5582 8260
rect 11890 8204 11900 8260
rect 11956 8204 12460 8260
rect 12516 8204 12526 8260
rect 12898 8204 12908 8260
rect 12964 8204 13692 8260
rect 13748 8204 13758 8260
rect 16258 8204 16268 8260
rect 16324 8204 16716 8260
rect 16772 8204 16782 8260
rect 18050 8204 18060 8260
rect 18116 8204 20188 8260
rect 20244 8204 20254 8260
rect 22978 8204 22988 8260
rect 23044 8204 23772 8260
rect 23828 8204 23838 8260
rect 25228 8204 25676 8260
rect 25732 8204 25742 8260
rect 37212 8204 38780 8260
rect 38836 8204 38846 8260
rect 41010 8204 41020 8260
rect 41076 8204 42140 8260
rect 42196 8204 42206 8260
rect 45126 8204 45164 8260
rect 45220 8204 45230 8260
rect 25228 8148 25284 8204
rect 8978 8092 8988 8148
rect 9044 8092 11228 8148
rect 11284 8092 11294 8148
rect 17266 8092 17276 8148
rect 17332 8092 17724 8148
rect 17780 8092 20300 8148
rect 20356 8092 20366 8148
rect 21410 8092 21420 8148
rect 21476 8092 22540 8148
rect 22596 8092 22606 8148
rect 23650 8092 23660 8148
rect 23716 8092 25228 8148
rect 25284 8092 25294 8148
rect 25442 8092 25452 8148
rect 25508 8092 25788 8148
rect 25844 8092 29484 8148
rect 29540 8092 29550 8148
rect 37650 8092 37660 8148
rect 37716 8092 37726 8148
rect 37874 8092 37884 8148
rect 37940 8092 39452 8148
rect 39508 8092 39518 8148
rect 40114 8092 40124 8148
rect 40180 8092 42364 8148
rect 42420 8092 42430 8148
rect 42578 8092 42588 8148
rect 42644 8092 43148 8148
rect 43204 8092 43214 8148
rect 44706 8092 44716 8148
rect 44772 8092 47852 8148
rect 47908 8092 47918 8148
rect 21420 8036 21476 8092
rect 14578 7980 14588 8036
rect 14644 7980 16156 8036
rect 16212 7980 16222 8036
rect 16706 7980 16716 8036
rect 16772 7980 17388 8036
rect 17444 7980 19404 8036
rect 19460 7980 19470 8036
rect 20178 7980 20188 8036
rect 20244 7980 21476 8036
rect 24098 7980 24108 8036
rect 24164 7980 25564 8036
rect 25620 7980 28252 8036
rect 28308 7980 28318 8036
rect 32498 7980 32508 8036
rect 32564 7980 34972 8036
rect 35028 7980 35038 8036
rect 37660 7924 37716 8092
rect 41234 7980 41244 8036
rect 41300 7980 42700 8036
rect 42756 7980 42766 8036
rect 43586 7980 43596 8036
rect 43652 7980 45276 8036
rect 45332 7980 47068 8036
rect 47124 7980 47134 8036
rect 16034 7868 16044 7924
rect 16100 7868 17276 7924
rect 17332 7868 17836 7924
rect 17892 7868 18396 7924
rect 18452 7868 18462 7924
rect 24546 7868 24556 7924
rect 24612 7868 32732 7924
rect 32788 7868 32798 7924
rect 33618 7868 33628 7924
rect 33684 7868 34860 7924
rect 34916 7868 34926 7924
rect 37660 7868 42252 7924
rect 42308 7868 42318 7924
rect 43250 7868 43260 7924
rect 43316 7868 43326 7924
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 43260 7700 43316 7868
rect 49200 7700 50000 7728
rect 19730 7644 19740 7700
rect 19796 7644 20300 7700
rect 20356 7644 20366 7700
rect 35746 7644 35756 7700
rect 35812 7644 38668 7700
rect 40002 7644 40012 7700
rect 40068 7644 41468 7700
rect 41524 7644 43316 7700
rect 48178 7644 48188 7700
rect 48244 7644 50000 7700
rect 4162 7532 4172 7588
rect 4228 7532 5068 7588
rect 5124 7532 5134 7588
rect 10770 7532 10780 7588
rect 10836 7532 12796 7588
rect 12852 7532 12862 7588
rect 23202 7532 23212 7588
rect 23268 7532 24108 7588
rect 24164 7532 24174 7588
rect 33618 7532 33628 7588
rect 33684 7532 34748 7588
rect 34804 7532 34814 7588
rect 38612 7476 38668 7644
rect 49200 7616 50000 7644
rect 41692 7532 42028 7588
rect 42084 7532 42094 7588
rect 42914 7532 42924 7588
rect 42980 7532 43372 7588
rect 43428 7532 43438 7588
rect 41692 7476 41748 7532
rect 2930 7420 2940 7476
rect 2996 7420 3388 7476
rect 3444 7420 4060 7476
rect 4116 7420 4396 7476
rect 4452 7420 4462 7476
rect 8194 7420 8204 7476
rect 8260 7420 9660 7476
rect 9716 7420 11564 7476
rect 11620 7420 11630 7476
rect 22642 7420 22652 7476
rect 22708 7420 26012 7476
rect 26068 7420 26078 7476
rect 31938 7420 31948 7476
rect 32004 7420 35532 7476
rect 35588 7420 35598 7476
rect 38612 7420 41692 7476
rect 41748 7420 41758 7476
rect 43586 7420 43596 7476
rect 43652 7420 45052 7476
rect 45108 7420 45118 7476
rect 8866 7308 8876 7364
rect 8932 7308 10332 7364
rect 10388 7308 10398 7364
rect 26226 7308 26236 7364
rect 26292 7308 26572 7364
rect 26628 7308 26638 7364
rect 37650 7308 37660 7364
rect 37716 7308 40012 7364
rect 40068 7308 43484 7364
rect 43540 7308 43550 7364
rect 43922 7308 43932 7364
rect 43988 7308 44604 7364
rect 44660 7308 44670 7364
rect 42018 7196 42028 7252
rect 42084 7196 43260 7252
rect 43316 7196 44044 7252
rect 44100 7196 44110 7252
rect 29026 7084 29036 7140
rect 29092 7084 29596 7140
rect 29652 7084 30268 7140
rect 30324 7084 30334 7140
rect 38322 7084 38332 7140
rect 38388 7084 44156 7140
rect 44212 7084 44940 7140
rect 44996 7084 45500 7140
rect 45556 7084 45566 7140
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 21868 6860 22428 6916
rect 22484 6860 22494 6916
rect 24546 6860 24556 6916
rect 24612 6860 28252 6916
rect 28308 6860 30940 6916
rect 30996 6860 31006 6916
rect 32946 6860 32956 6916
rect 33012 6860 33740 6916
rect 33796 6860 33806 6916
rect 34178 6860 34188 6916
rect 34244 6860 38668 6916
rect 44482 6860 44492 6916
rect 44548 6860 45276 6916
rect 45332 6860 46732 6916
rect 46788 6860 46798 6916
rect 6738 6748 6748 6804
rect 6804 6748 8204 6804
rect 8260 6748 8270 6804
rect 8978 6748 8988 6804
rect 9044 6748 10444 6804
rect 10500 6748 10510 6804
rect 11106 6748 11116 6804
rect 11172 6748 12124 6804
rect 12180 6748 13356 6804
rect 13412 6748 13422 6804
rect 16482 6748 16492 6804
rect 16548 6748 17052 6804
rect 17108 6748 17118 6804
rect 21868 6692 21924 6860
rect 38612 6804 38668 6860
rect 26450 6748 26460 6804
rect 26516 6748 30380 6804
rect 30436 6748 30446 6804
rect 32498 6748 32508 6804
rect 32564 6748 37660 6804
rect 37716 6748 37726 6804
rect 38612 6748 47852 6804
rect 47908 6748 47918 6804
rect 11218 6636 11228 6692
rect 11284 6636 15596 6692
rect 15652 6636 21924 6692
rect 24322 6636 24332 6692
rect 24388 6636 24780 6692
rect 24836 6636 26124 6692
rect 26180 6636 26684 6692
rect 26740 6636 26750 6692
rect 28354 6636 28364 6692
rect 28420 6636 29372 6692
rect 29428 6636 30044 6692
rect 30100 6636 30110 6692
rect 32162 6636 32172 6692
rect 32228 6636 33292 6692
rect 33348 6636 34188 6692
rect 34244 6636 34254 6692
rect 35522 6636 35532 6692
rect 35588 6636 36988 6692
rect 37044 6636 37054 6692
rect 43362 6636 43372 6692
rect 43428 6636 43820 6692
rect 43876 6636 43886 6692
rect 47618 6636 47628 6692
rect 47684 6636 48188 6692
rect 48244 6636 48254 6692
rect 4722 6524 4732 6580
rect 4788 6524 5628 6580
rect 5684 6524 5694 6580
rect 14242 6524 14252 6580
rect 14308 6524 16268 6580
rect 16324 6524 16334 6580
rect 17938 6524 17948 6580
rect 18004 6524 19964 6580
rect 20020 6524 20030 6580
rect 20738 6524 20748 6580
rect 20804 6524 21756 6580
rect 21812 6524 24220 6580
rect 24276 6524 24286 6580
rect 27458 6524 27468 6580
rect 27524 6524 29148 6580
rect 29204 6524 29214 6580
rect 34626 6524 34636 6580
rect 34692 6524 36092 6580
rect 36148 6524 36158 6580
rect 42354 6524 42364 6580
rect 42420 6524 42924 6580
rect 42980 6524 43260 6580
rect 43316 6524 44828 6580
rect 44884 6524 44894 6580
rect 5394 6412 5404 6468
rect 5460 6412 6300 6468
rect 6356 6412 7196 6468
rect 7252 6412 7262 6468
rect 16034 6412 16044 6468
rect 16100 6412 17164 6468
rect 17220 6412 17230 6468
rect 19282 6412 19292 6468
rect 19348 6412 21420 6468
rect 21476 6412 21486 6468
rect 28578 6412 28588 6468
rect 28644 6412 29596 6468
rect 29652 6412 30604 6468
rect 30660 6412 30670 6468
rect 34514 6412 34524 6468
rect 34580 6412 35868 6468
rect 35924 6412 35934 6468
rect 42130 6412 42140 6468
rect 42196 6412 42812 6468
rect 42868 6412 42878 6468
rect 46274 6412 46284 6468
rect 46340 6412 47404 6468
rect 47460 6412 47470 6468
rect 27346 6300 27356 6356
rect 27412 6300 31052 6356
rect 31108 6300 31612 6356
rect 31668 6300 31678 6356
rect 32722 6300 32732 6356
rect 32788 6300 41692 6356
rect 41748 6300 41758 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 5954 6188 5964 6244
rect 6020 6188 6636 6244
rect 6692 6188 7420 6244
rect 7476 6188 7980 6244
rect 8036 6188 8316 6244
rect 8372 6188 8382 6244
rect 2482 6076 2492 6132
rect 2548 6076 5180 6132
rect 5236 6076 5246 6132
rect 7858 6076 7868 6132
rect 7924 6076 8764 6132
rect 8820 6076 10220 6132
rect 10276 6076 10286 6132
rect 16930 6076 16940 6132
rect 16996 6076 17612 6132
rect 17668 6076 20860 6132
rect 20916 6076 20926 6132
rect 39442 6076 39452 6132
rect 39508 6076 40236 6132
rect 40292 6076 41020 6132
rect 41076 6076 41086 6132
rect 15026 5964 15036 6020
rect 15092 5964 15932 6020
rect 15988 5964 16156 6020
rect 16212 5964 17052 6020
rect 17108 5964 21532 6020
rect 21588 5964 21598 6020
rect 21970 5964 21980 6020
rect 22036 5964 25228 6020
rect 25284 5964 25294 6020
rect 33394 5964 33404 6020
rect 33460 5964 33852 6020
rect 33908 5964 33918 6020
rect 34962 5964 34972 6020
rect 35028 5964 41132 6020
rect 41188 5964 41198 6020
rect 6514 5852 6524 5908
rect 6580 5852 7084 5908
rect 7140 5852 7868 5908
rect 7924 5852 7934 5908
rect 9650 5852 9660 5908
rect 9716 5852 17948 5908
rect 18004 5852 18014 5908
rect 20066 5852 20076 5908
rect 20132 5852 21196 5908
rect 21252 5852 25340 5908
rect 25396 5852 25406 5908
rect 34178 5852 34188 5908
rect 34244 5852 34860 5908
rect 34916 5852 34926 5908
rect 39218 5852 39228 5908
rect 39284 5852 39900 5908
rect 39956 5852 39966 5908
rect 41906 5852 41916 5908
rect 41972 5852 42812 5908
rect 42868 5852 42878 5908
rect 8754 5740 8764 5796
rect 8820 5740 17612 5796
rect 17668 5740 21308 5796
rect 21364 5740 21374 5796
rect 21522 5740 21532 5796
rect 21588 5740 22428 5796
rect 22484 5740 22494 5796
rect 33170 5740 33180 5796
rect 33236 5740 33852 5796
rect 33908 5740 33918 5796
rect 40226 5740 40236 5796
rect 40292 5740 41580 5796
rect 41636 5740 41646 5796
rect 18162 5628 18172 5684
rect 18228 5628 18956 5684
rect 19012 5628 19022 5684
rect 22306 5628 22316 5684
rect 22372 5628 25900 5684
rect 25956 5628 25966 5684
rect 31042 5628 31052 5684
rect 31108 5628 36988 5684
rect 37044 5628 37054 5684
rect 38612 5628 39564 5684
rect 39620 5628 40124 5684
rect 40180 5628 40190 5684
rect 41234 5628 41244 5684
rect 41300 5628 42252 5684
rect 42308 5628 42318 5684
rect 15138 5516 15148 5572
rect 15204 5516 22204 5572
rect 22260 5516 22764 5572
rect 22820 5516 26908 5572
rect 26964 5516 26974 5572
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 31052 5460 31108 5628
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 38612 5460 38668 5628
rect 41570 5516 41580 5572
rect 41636 5516 42364 5572
rect 42420 5516 42430 5572
rect 26338 5404 26348 5460
rect 26404 5404 31108 5460
rect 36306 5404 36316 5460
rect 36372 5404 38220 5460
rect 38276 5404 38668 5460
rect 39778 5404 39788 5460
rect 39844 5404 42252 5460
rect 42308 5404 42812 5460
rect 42868 5404 42878 5460
rect 15708 5292 17948 5348
rect 18004 5292 18014 5348
rect 20290 5292 20300 5348
rect 20356 5292 20524 5348
rect 20580 5292 23660 5348
rect 23716 5292 23726 5348
rect 30034 5292 30044 5348
rect 30100 5292 31276 5348
rect 31332 5292 31342 5348
rect 35410 5292 35420 5348
rect 35476 5292 36876 5348
rect 36932 5292 39228 5348
rect 39284 5292 39294 5348
rect 40226 5292 40236 5348
rect 40292 5292 40572 5348
rect 40628 5292 41356 5348
rect 41412 5292 41422 5348
rect 41794 5292 41804 5348
rect 41860 5292 42140 5348
rect 42196 5292 44828 5348
rect 44884 5292 44894 5348
rect 15708 5012 15764 5292
rect 17826 5180 17836 5236
rect 17892 5180 19516 5236
rect 19572 5180 19582 5236
rect 23426 5180 23436 5236
rect 23492 5180 24668 5236
rect 24724 5180 24734 5236
rect 24892 5180 29148 5236
rect 29204 5180 29214 5236
rect 33506 5180 33516 5236
rect 33572 5180 34748 5236
rect 34804 5180 34814 5236
rect 35298 5180 35308 5236
rect 35364 5180 35756 5236
rect 35812 5180 35822 5236
rect 41682 5180 41692 5236
rect 41748 5180 42364 5236
rect 42420 5180 42430 5236
rect 43474 5180 43484 5236
rect 43540 5180 43708 5236
rect 43764 5180 43774 5236
rect 24892 5124 24948 5180
rect 16594 5068 16604 5124
rect 16660 5068 18508 5124
rect 18564 5068 18574 5124
rect 21634 5068 21644 5124
rect 21700 5068 23548 5124
rect 23604 5068 23614 5124
rect 23762 5068 23772 5124
rect 23828 5068 24948 5124
rect 26114 5068 26124 5124
rect 26180 5068 27804 5124
rect 27860 5068 27870 5124
rect 29474 5068 29484 5124
rect 29540 5068 30492 5124
rect 30548 5068 30558 5124
rect 33618 5068 33628 5124
rect 33684 5068 34636 5124
rect 34692 5068 35644 5124
rect 35700 5068 35710 5124
rect 37426 5068 37436 5124
rect 37492 5068 40684 5124
rect 40740 5068 40750 5124
rect 41010 5068 41020 5124
rect 41076 5068 41356 5124
rect 41412 5068 42028 5124
rect 42084 5068 42094 5124
rect 44146 5068 44156 5124
rect 44212 5068 46956 5124
rect 47012 5068 47022 5124
rect 1810 4956 1820 5012
rect 1876 4956 4172 5012
rect 4228 4956 4238 5012
rect 15698 4956 15708 5012
rect 15764 4956 15774 5012
rect 25778 4956 25788 5012
rect 25844 4956 29260 5012
rect 29316 4956 29326 5012
rect 34066 4956 34076 5012
rect 34132 4956 35532 5012
rect 35588 4956 35598 5012
rect 16034 4844 16044 4900
rect 16100 4844 17500 4900
rect 17556 4844 17566 4900
rect 23538 4844 23548 4900
rect 23604 4844 26348 4900
rect 26404 4844 26414 4900
rect 30370 4844 30380 4900
rect 30436 4844 32956 4900
rect 33012 4844 33022 4900
rect 34962 4844 34972 4900
rect 35028 4844 37996 4900
rect 38052 4844 38062 4900
rect 33954 4732 33964 4788
rect 34020 4732 36092 4788
rect 36148 4732 36158 4788
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 33282 4508 33292 4564
rect 33348 4508 34412 4564
rect 34468 4508 34860 4564
rect 34916 4508 34926 4564
rect 8978 4396 8988 4452
rect 9044 4396 11004 4452
rect 11060 4396 11070 4452
rect 16370 4396 16380 4452
rect 16436 4396 17388 4452
rect 17444 4396 17454 4452
rect 22418 4396 22428 4452
rect 22484 4396 25228 4452
rect 25284 4396 25294 4452
rect 39554 4396 39564 4452
rect 39620 4396 40908 4452
rect 40964 4396 40974 4452
rect 12898 4284 12908 4340
rect 12964 4284 21084 4340
rect 21140 4284 21150 4340
rect 32274 4284 32284 4340
rect 32340 4284 34076 4340
rect 34132 4284 34142 4340
rect 40338 4284 40348 4340
rect 40404 4284 45388 4340
rect 45444 4284 47628 4340
rect 47684 4284 47694 4340
rect 4946 4172 4956 4228
rect 5012 4172 7532 4228
rect 7588 4172 7598 4228
rect 20290 4172 20300 4228
rect 20356 4172 21420 4228
rect 21476 4172 25900 4228
rect 25956 4172 25966 4228
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 39666 3836 39676 3892
rect 39732 3836 41580 3892
rect 41636 3836 41646 3892
rect 22642 3724 22652 3780
rect 22708 3724 24556 3780
rect 24612 3724 24622 3780
rect 28690 3724 28700 3780
rect 28756 3724 29260 3780
rect 29316 3724 29326 3780
rect 36530 3724 36540 3780
rect 36596 3724 40012 3780
rect 40068 3724 40078 3780
rect 20850 3612 20860 3668
rect 20916 3612 22092 3668
rect 22148 3612 22158 3668
rect 31826 3612 31836 3668
rect 31892 3612 36988 3668
rect 37044 3612 37054 3668
rect 43586 3612 43596 3668
rect 43652 3612 45500 3668
rect 45556 3612 45566 3668
rect 13122 3500 13132 3556
rect 13188 3500 17612 3556
rect 17668 3500 17678 3556
rect 24658 3500 24668 3556
rect 24724 3500 29036 3556
rect 29092 3500 29102 3556
rect 32162 3500 32172 3556
rect 32228 3500 35980 3556
rect 36036 3500 36046 3556
rect 7746 3388 7756 3444
rect 7812 3388 8204 3444
rect 8260 3388 15148 3444
rect 15204 3388 15214 3444
rect 31490 3388 31500 3444
rect 31556 3388 47852 3444
rect 47908 3388 47918 3444
rect 23986 3276 23996 3332
rect 24052 3276 25228 3332
rect 25284 3276 25294 3332
rect 38098 3276 38108 3332
rect 38164 3276 38892 3332
rect 38948 3276 38958 3332
rect 42802 3276 42812 3332
rect 42868 3276 44492 3332
rect 44548 3276 44558 3332
rect 47618 3276 47628 3332
rect 47684 3276 48188 3332
rect 48244 3276 48254 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 49200 2772 50000 2800
rect 48178 2716 48188 2772
rect 48244 2716 50000 2772
rect 49200 2688 50000 2716
rect 41234 1708 41244 1764
rect 41300 1708 42700 1764
rect 42756 1708 42766 1764
<< via3 >>
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 16044 44044 16100 44100
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 16044 40460 16100 40516
rect 30492 40348 30548 40404
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 30492 39564 30548 39620
rect 47068 39452 47124 39508
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 25788 38780 25844 38836
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 47068 37212 47124 37268
rect 26572 36988 26628 37044
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 30716 36092 30772 36148
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 23548 34972 23604 35028
rect 29484 34860 29540 34916
rect 43372 34748 43428 34804
rect 24220 34636 24276 34692
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 24220 33852 24276 33908
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 26236 33516 26292 33572
rect 29484 33292 29540 33348
rect 37324 33180 37380 33236
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 23548 32508 23604 32564
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 26908 31948 26964 32004
rect 30716 31388 30772 31444
rect 31164 31388 31220 31444
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 34860 30604 34916 30660
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 34636 30492 34692 30548
rect 23996 30268 24052 30324
rect 34300 30156 34356 30212
rect 33852 30044 33908 30100
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 23996 29708 24052 29764
rect 30492 29708 30548 29764
rect 43596 29372 43652 29428
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 26908 28812 26964 28868
rect 33852 28812 33908 28868
rect 34300 28476 34356 28532
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 26236 28028 26292 28084
rect 34860 27692 34916 27748
rect 34636 27580 34692 27636
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 26908 27356 26964 27412
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 43596 25452 43652 25508
rect 43372 25340 43428 25396
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 37324 25004 37380 25060
rect 30492 24892 30548 24948
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 31164 24220 31220 24276
rect 30492 24108 30548 24164
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 33852 23324 33908 23380
rect 35644 22988 35700 23044
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 43372 22540 43428 22596
rect 33964 22204 34020 22260
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 34412 21868 34468 21924
rect 35644 21420 35700 21476
rect 26572 21308 26628 21364
rect 33964 21196 34020 21252
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 31500 18508 31556 18564
rect 33852 18172 33908 18228
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 25788 17724 25844 17780
rect 35756 17612 35812 17668
rect 35644 17500 35700 17556
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 31500 17052 31556 17108
rect 43372 16604 43428 16660
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 44828 15820 44884 15876
rect 35756 15708 35812 15764
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 35644 13692 35700 13748
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 34188 12796 34244 12852
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 34412 12460 34468 12516
rect 34188 12236 34244 12292
rect 44828 11900 44884 11956
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 45164 11564 45220 11620
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 34412 9548 34468 9604
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 45164 8204 45220 8260
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 34412 4508 34468 4564
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 46284 4768 46316
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 19808 45500 20128 46316
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 16044 44100 16100 44110
rect 16044 40516 16100 44044
rect 16044 40450 16100 40460
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 39228 20128 40740
rect 35168 46284 35488 46316
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 30492 40404 30548 40414
rect 30492 39620 30548 40348
rect 30492 39554 30548 39564
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 25788 38836 25844 38846
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 23548 35028 23604 35038
rect 23548 32564 23604 34972
rect 24220 34692 24276 34702
rect 24220 33908 24276 34636
rect 24220 33842 24276 33852
rect 23548 32498 23604 32508
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 23996 30324 24052 30334
rect 23996 29764 24052 30268
rect 23996 29698 24052 29708
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 25788 17780 25844 38780
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 26572 37044 26628 37054
rect 26236 33572 26292 33582
rect 26236 28084 26292 33516
rect 26236 28018 26292 28028
rect 26572 21364 26628 36988
rect 35168 36876 35488 38388
rect 47068 39508 47124 39518
rect 47068 37268 47124 39452
rect 47068 37202 47124 37212
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 30716 36148 30772 36158
rect 29484 34916 29540 34926
rect 29484 33348 29540 34860
rect 29484 33282 29540 33292
rect 26908 32004 26964 32014
rect 26908 28868 26964 31948
rect 30716 31444 30772 36092
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 43372 34804 43428 34814
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 30716 31378 30772 31388
rect 31164 31444 31220 31454
rect 26908 27412 26964 28812
rect 26908 27346 26964 27356
rect 30492 29764 30548 29774
rect 30492 24948 30548 29708
rect 30492 24164 30548 24892
rect 31164 24276 31220 31388
rect 34860 30660 34916 30670
rect 34636 30548 34692 30558
rect 34300 30212 34356 30222
rect 33852 30100 33908 30110
rect 33852 28868 33908 30044
rect 33852 28802 33908 28812
rect 34300 28532 34356 30156
rect 34300 28466 34356 28476
rect 34636 27636 34692 30492
rect 34860 27748 34916 30604
rect 34860 27682 34916 27692
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 34636 27570 34692 27580
rect 31164 24210 31220 24220
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 37324 33236 37380 33246
rect 37324 25060 37380 33180
rect 43372 25396 43428 34748
rect 43596 29428 43652 29438
rect 43596 25508 43652 29372
rect 43596 25442 43652 25452
rect 43372 25330 43428 25340
rect 37324 24994 37380 25004
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 30492 24098 30548 24108
rect 26572 21298 26628 21308
rect 33852 23380 33908 23390
rect 25788 17714 25844 17724
rect 31500 18564 31556 18574
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 31500 17108 31556 18508
rect 33852 18228 33908 23324
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 33964 22260 34020 22270
rect 33964 21252 34020 22204
rect 33964 21186 34020 21196
rect 34412 21924 34468 21934
rect 33852 18162 33908 18172
rect 31500 17042 31556 17052
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 34188 12852 34244 12862
rect 34188 12292 34244 12796
rect 34412 12516 34468 21868
rect 34412 12450 34468 12460
rect 35168 21196 35488 22708
rect 35644 23044 35700 23054
rect 35644 21476 35700 22988
rect 35644 21410 35700 21420
rect 43372 22596 43428 22606
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35756 17668 35812 17678
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35644 17556 35700 17566
rect 35644 13748 35700 17500
rect 35756 15764 35812 17612
rect 43372 16660 43428 22540
rect 43372 16594 43428 16604
rect 35756 15698 35812 15708
rect 44828 15876 44884 15886
rect 35644 13682 35700 13692
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 34188 12226 34244 12236
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 35168 11788 35488 13300
rect 44828 11956 44884 15820
rect 44828 11890 44884 11900
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 34412 9604 34468 9614
rect 34412 4564 34468 9548
rect 34412 4498 34468 4508
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 45164 11620 45220 11630
rect 45164 8260 45220 11564
rect 45164 8194 45220 8204
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _1024_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7392 0 1 32928
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1025_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20944 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1026_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1027_
timestamp 1698431365
transform 1 0 22960 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1028_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1029_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26096 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1030_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26992 0 1 20384
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1031_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 21728 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1032_
timestamp 1698431365
transform 1 0 19712 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1033_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19488 0 -1 28224
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1034_
timestamp 1698431365
transform 1 0 20384 0 -1 26656
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1035_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18144 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1036_
timestamp 1698431365
transform -1 0 28336 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1037_
timestamp 1698431365
transform 1 0 18256 0 -1 26656
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1038_
timestamp 1698431365
transform 1 0 18480 0 -1 23520
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1039_
timestamp 1698431365
transform 1 0 20496 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1040_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20720 0 -1 18816
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1041_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1042_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18032 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1043_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18256 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1044_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18368 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1045_
timestamp 1698431365
transform 1 0 20160 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1046_
timestamp 1698431365
transform 1 0 23856 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1047_
timestamp 1698431365
transform -1 0 30464 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1048_
timestamp 1698431365
transform 1 0 30016 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1049_
timestamp 1698431365
transform -1 0 30576 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1050_
timestamp 1698431365
transform 1 0 30576 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1051_
timestamp 1698431365
transform -1 0 28784 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1052_
timestamp 1698431365
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1053_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28672 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1054_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28000 0 1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1055_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31136 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1056_
timestamp 1698431365
transform -1 0 32032 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1057_
timestamp 1698431365
transform -1 0 23632 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1058_
timestamp 1698431365
transform 1 0 23408 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1059_
timestamp 1698431365
transform -1 0 31248 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1060_
timestamp 1698431365
transform 1 0 30688 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1061_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30688 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1062_
timestamp 1698431365
transform -1 0 32144 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1063_
timestamp 1698431365
transform -1 0 33488 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1064_
timestamp 1698431365
transform 1 0 31136 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1065_
timestamp 1698431365
transform 1 0 32144 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1066_
timestamp 1698431365
transform 1 0 34720 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1067_
timestamp 1698431365
transform 1 0 31248 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1068_
timestamp 1698431365
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1069_
timestamp 1698431365
transform -1 0 35056 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1070_
timestamp 1698431365
transform 1 0 30800 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1071_
timestamp 1698431365
transform 1 0 30240 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1072_
timestamp 1698431365
transform -1 0 48160 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1073_
timestamp 1698431365
transform 1 0 35280 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1074_
timestamp 1698431365
transform 1 0 29568 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1075_
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1076_
timestamp 1698431365
transform -1 0 26880 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1077_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27552 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1078_
timestamp 1698431365
transform -1 0 29680 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1079_
timestamp 1698431365
transform 1 0 31472 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1080_
timestamp 1698431365
transform 1 0 33040 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1081_
timestamp 1698431365
transform -1 0 22400 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1082_
timestamp 1698431365
transform -1 0 22624 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1083_
timestamp 1698431365
transform 1 0 33152 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1084_
timestamp 1698431365
transform -1 0 35504 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1085_
timestamp 1698431365
transform -1 0 32704 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1086_
timestamp 1698431365
transform -1 0 34384 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1087_
timestamp 1698431365
transform -1 0 33376 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1088_
timestamp 1698431365
transform -1 0 36512 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1089_
timestamp 1698431365
transform 1 0 34608 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1090_
timestamp 1698431365
transform -1 0 35504 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1091_
timestamp 1698431365
transform 1 0 33376 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1092_
timestamp 1698431365
transform -1 0 29792 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1093_
timestamp 1698431365
transform 1 0 30576 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1094_
timestamp 1698431365
transform -1 0 31920 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1095_
timestamp 1698431365
transform -1 0 24640 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1096_
timestamp 1698431365
transform 1 0 24080 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1097_
timestamp 1698431365
transform 1 0 22512 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1098_
timestamp 1698431365
transform 1 0 33376 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1099_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 24080 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1100_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23632 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1101_
timestamp 1698431365
transform 1 0 22176 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1102_
timestamp 1698431365
transform -1 0 25088 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1103_
timestamp 1698431365
transform 1 0 24752 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1104_
timestamp 1698431365
transform 1 0 25424 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1105_
timestamp 1698431365
transform -1 0 36624 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1106_
timestamp 1698431365
transform 1 0 24304 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1107_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1108_
timestamp 1698431365
transform -1 0 21504 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1109_
timestamp 1698431365
transform -1 0 11872 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1110_
timestamp 1698431365
transform 1 0 11424 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1111_
timestamp 1698431365
transform 1 0 20384 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1112_
timestamp 1698431365
transform -1 0 36848 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1113_
timestamp 1698431365
transform 1 0 24752 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1114_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21392 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1115_
timestamp 1698431365
transform 1 0 21952 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1116_
timestamp 1698431365
transform 1 0 37632 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1117_
timestamp 1698431365
transform -1 0 24304 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1118_
timestamp 1698431365
transform 1 0 22400 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1119_
timestamp 1698431365
transform 1 0 22960 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1120_
timestamp 1698431365
transform 1 0 22288 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1121_
timestamp 1698431365
transform -1 0 22064 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1122_
timestamp 1698431365
transform 1 0 18592 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1123_
timestamp 1698431365
transform -1 0 18592 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1124_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19376 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1125_
timestamp 1698431365
transform 1 0 20384 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1126_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20384 0 -1 15680
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1127_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19264 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1128_
timestamp 1698431365
transform 1 0 18592 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1129_
timestamp 1698431365
transform -1 0 19152 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1130_
timestamp 1698431365
transform 1 0 20160 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1131_
timestamp 1698431365
transform 1 0 11536 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1132_
timestamp 1698431365
transform 1 0 15008 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1133_
timestamp 1698431365
transform -1 0 18480 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1134_
timestamp 1698431365
transform 1 0 17696 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1135_
timestamp 1698431365
transform 1 0 21168 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1136_
timestamp 1698431365
transform -1 0 17920 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1137_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18480 0 1 12544
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1138_
timestamp 1698431365
transform 1 0 15120 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1139_
timestamp 1698431365
transform 1 0 16464 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1140_
timestamp 1698431365
transform -1 0 18144 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1141_
timestamp 1698431365
transform 1 0 10080 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1142_
timestamp 1698431365
transform -1 0 10080 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1143_
timestamp 1698431365
transform -1 0 11312 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1144_
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1145_
timestamp 1698431365
transform -1 0 13888 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1146_
timestamp 1698431365
transform -1 0 12880 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1147_
timestamp 1698431365
transform -1 0 13104 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1148_
timestamp 1698431365
transform 1 0 11984 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1149_
timestamp 1698431365
transform 1 0 11424 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1150_
timestamp 1698431365
transform 1 0 12096 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1151_
timestamp 1698431365
transform -1 0 11088 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1152_
timestamp 1698431365
transform -1 0 11088 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1153_
timestamp 1698431365
transform 1 0 11424 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1154_
timestamp 1698431365
transform -1 0 13888 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1155_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 12432 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1156_
timestamp 1698431365
transform -1 0 9184 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1157_
timestamp 1698431365
transform -1 0 12992 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1158_
timestamp 1698431365
transform -1 0 12544 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1159_
timestamp 1698431365
transform 1 0 11872 0 1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1160_
timestamp 1698431365
transform -1 0 13328 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1161_
timestamp 1698431365
transform 1 0 29904 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1162_
timestamp 1698431365
transform -1 0 28784 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1163_
timestamp 1698431365
transform 1 0 28448 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1164_
timestamp 1698431365
transform -1 0 30128 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1165_
timestamp 1698431365
transform -1 0 24192 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1166_
timestamp 1698431365
transform -1 0 21840 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1167_
timestamp 1698431365
transform 1 0 22512 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1168_
timestamp 1698431365
transform -1 0 23520 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1169_
timestamp 1698431365
transform -1 0 28784 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1170_
timestamp 1698431365
transform -1 0 24304 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1171_
timestamp 1698431365
transform -1 0 28336 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1172_
timestamp 1698431365
transform 1 0 23632 0 -1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1173_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22400 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1174_
timestamp 1698431365
transform 1 0 16128 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1175_
timestamp 1698431365
transform 1 0 15680 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1176_
timestamp 1698431365
transform -1 0 17808 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1177_
timestamp 1698431365
transform 1 0 24192 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1178_
timestamp 1698431365
transform -1 0 25760 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1179_
timestamp 1698431365
transform -1 0 22176 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1180_
timestamp 1698431365
transform -1 0 19376 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1181_
timestamp 1698431365
transform -1 0 22176 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1182_
timestamp 1698431365
transform -1 0 18928 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1183_
timestamp 1698431365
transform -1 0 20944 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1184_
timestamp 1698431365
transform -1 0 18256 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1185_
timestamp 1698431365
transform -1 0 19936 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1186_
timestamp 1698431365
transform -1 0 21392 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1187_
timestamp 1698431365
transform -1 0 17472 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1188_
timestamp 1698431365
transform -1 0 16464 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1189_
timestamp 1698431365
transform -1 0 16464 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1190_
timestamp 1698431365
transform 1 0 16576 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1191_
timestamp 1698431365
transform -1 0 16576 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1192_
timestamp 1698431365
transform -1 0 16464 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1193_
timestamp 1698431365
transform -1 0 15456 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1194_
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1195_
timestamp 1698431365
transform -1 0 17472 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1196_
timestamp 1698431365
transform 1 0 19712 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1197_
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1198_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20272 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1199_
timestamp 1698431365
transform -1 0 17024 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1200_
timestamp 1698431365
transform 1 0 16800 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1201_
timestamp 1698431365
transform -1 0 11200 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1202_
timestamp 1698431365
transform 1 0 9632 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1203_
timestamp 1698431365
transform -1 0 10192 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1204_
timestamp 1698431365
transform -1 0 3920 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1205_
timestamp 1698431365
transform -1 0 6160 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1206_
timestamp 1698431365
transform -1 0 4816 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1207_
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1208_
timestamp 1698431365
transform 1 0 4816 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1209_
timestamp 1698431365
transform -1 0 5264 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1210_
timestamp 1698431365
transform 1 0 4256 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1211_
timestamp 1698431365
transform -1 0 4256 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1212_
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1213_
timestamp 1698431365
transform 1 0 4144 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1214_
timestamp 1698431365
transform 1 0 4928 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1215_
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1216_
timestamp 1698431365
transform 1 0 6496 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1217_
timestamp 1698431365
transform 1 0 6384 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1218_
timestamp 1698431365
transform 1 0 5936 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1219_
timestamp 1698431365
transform 1 0 6832 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1220_
timestamp 1698431365
transform 1 0 8512 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1221_
timestamp 1698431365
transform -1 0 28560 0 -1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1222_
timestamp 1698431365
transform 1 0 30128 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1223_
timestamp 1698431365
transform -1 0 35616 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1224_
timestamp 1698431365
transform -1 0 23408 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1225_
timestamp 1698431365
transform 1 0 33488 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1226_
timestamp 1698431365
transform -1 0 35616 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1227_
timestamp 1698431365
transform -1 0 34160 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1228_
timestamp 1698431365
transform -1 0 32704 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1229_
timestamp 1698431365
transform -1 0 35168 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1230_
timestamp 1698431365
transform -1 0 34496 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1231_
timestamp 1698431365
transform 1 0 34608 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1232_
timestamp 1698431365
transform -1 0 36848 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1233_
timestamp 1698431365
transform -1 0 36624 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1234_
timestamp 1698431365
transform 1 0 35056 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1235_
timestamp 1698431365
transform 1 0 40096 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1236_
timestamp 1698431365
transform 1 0 39424 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1237_
timestamp 1698431365
transform -1 0 41776 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1238_
timestamp 1698431365
transform 1 0 40096 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1239_
timestamp 1698431365
transform 1 0 41888 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1240_
timestamp 1698431365
transform 1 0 42784 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1241_
timestamp 1698431365
transform -1 0 44352 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1242_
timestamp 1698431365
transform -1 0 45696 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1243_
timestamp 1698431365
transform 1 0 45024 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1244_
timestamp 1698431365
transform 1 0 46480 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1245_
timestamp 1698431365
transform -1 0 47824 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1246_
timestamp 1698431365
transform 1 0 45024 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1247_
timestamp 1698431365
transform 1 0 46032 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1248_
timestamp 1698431365
transform 1 0 29680 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1249_
timestamp 1698431365
transform 1 0 31584 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1250_
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1251_
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1252_
timestamp 1698431365
transform -1 0 34832 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1253_
timestamp 1698431365
transform -1 0 35280 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1254_
timestamp 1698431365
transform -1 0 34048 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1255_
timestamp 1698431365
transform 1 0 32256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1256_
timestamp 1698431365
transform -1 0 35952 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1257_
timestamp 1698431365
transform 1 0 36064 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1258_
timestamp 1698431365
transform -1 0 36064 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1259_
timestamp 1698431365
transform 1 0 35840 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1260_
timestamp 1698431365
transform -1 0 27552 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1261_
timestamp 1698431365
transform 1 0 33152 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1262_
timestamp 1698431365
transform -1 0 33600 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1263_
timestamp 1698431365
transform 1 0 33600 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1264_
timestamp 1698431365
transform -1 0 34944 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1265_
timestamp 1698431365
transform -1 0 33488 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1266_
timestamp 1698431365
transform -1 0 31696 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1267_
timestamp 1698431365
transform -1 0 34944 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1268_
timestamp 1698431365
transform -1 0 34272 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1269_
timestamp 1698431365
transform 1 0 33152 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1270_
timestamp 1698431365
transform -1 0 35056 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1271_
timestamp 1698431365
transform -1 0 34720 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1272_
timestamp 1698431365
transform 1 0 33040 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1273_
timestamp 1698431365
transform 1 0 35056 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1274_
timestamp 1698431365
transform -1 0 34272 0 -1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1275_
timestamp 1698431365
transform 1 0 34944 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1276_
timestamp 1698431365
transform 1 0 34944 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1277_
timestamp 1698431365
transform 1 0 36960 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1278_
timestamp 1698431365
transform -1 0 41776 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1279_
timestamp 1698431365
transform -1 0 42224 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1280_
timestamp 1698431365
transform -1 0 44688 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1281_
timestamp 1698431365
transform 1 0 46256 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1282_
timestamp 1698431365
transform -1 0 45696 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1283_
timestamp 1698431365
transform 1 0 46704 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1284_
timestamp 1698431365
transform -1 0 43680 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1285_
timestamp 1698431365
transform -1 0 43344 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1286_
timestamp 1698431365
transform -1 0 26208 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1287_
timestamp 1698431365
transform 1 0 25424 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1288_
timestamp 1698431365
transform 1 0 25984 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1289_
timestamp 1698431365
transform -1 0 27104 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1290_
timestamp 1698431365
transform 1 0 21728 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1291_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26208 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1292_
timestamp 1698431365
transform -1 0 25984 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1293_
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1294_
timestamp 1698431365
transform 1 0 26656 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1295_
timestamp 1698431365
transform -1 0 28224 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1296_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28112 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1297_
timestamp 1698431365
transform -1 0 26880 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1298_
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1299_
timestamp 1698431365
transform 1 0 29904 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1300_
timestamp 1698431365
transform -1 0 5600 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1301_
timestamp 1698431365
transform -1 0 4704 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1302_
timestamp 1698431365
transform -1 0 3808 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1303_
timestamp 1698431365
transform -1 0 4256 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1304_
timestamp 1698431365
transform 1 0 3584 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1305_
timestamp 1698431365
transform -1 0 3584 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1306_
timestamp 1698431365
transform 1 0 3248 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1307_
timestamp 1698431365
transform -1 0 6720 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1308_
timestamp 1698431365
transform 1 0 3248 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1309_
timestamp 1698431365
transform 1 0 4816 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1310_
timestamp 1698431365
transform -1 0 4256 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1311_
timestamp 1698431365
transform 1 0 3360 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1312_
timestamp 1698431365
transform -1 0 3360 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1313_
timestamp 1698431365
transform 1 0 4032 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1314_
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1315_
timestamp 1698431365
transform 1 0 4256 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1316_
timestamp 1698431365
transform 1 0 4928 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1317_
timestamp 1698431365
transform 1 0 10080 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1318_
timestamp 1698431365
transform 1 0 7056 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1319_
timestamp 1698431365
transform 1 0 6160 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1320_
timestamp 1698431365
transform 1 0 21616 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1321_
timestamp 1698431365
transform 1 0 5712 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1322_
timestamp 1698431365
transform 1 0 5824 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1323_
timestamp 1698431365
transform 1 0 7280 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1324_
timestamp 1698431365
transform -1 0 8400 0 -1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1325_
timestamp 1698431365
transform 1 0 7280 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1326_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31920 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1327_
timestamp 1698431365
transform -1 0 31584 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1328_
timestamp 1698431365
transform 1 0 24192 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1329_
timestamp 1698431365
transform -1 0 23184 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1330_
timestamp 1698431365
transform 1 0 21616 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1331_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1332_
timestamp 1698431365
transform 1 0 38528 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1333_
timestamp 1698431365
transform 1 0 20496 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1334_
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1335_
timestamp 1698431365
transform -1 0 24416 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1336_
timestamp 1698431365
transform -1 0 21840 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1337_
timestamp 1698431365
transform -1 0 23968 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1338_
timestamp 1698431365
transform -1 0 21840 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1339_
timestamp 1698431365
transform 1 0 18144 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1340_
timestamp 1698431365
transform -1 0 16688 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1341_
timestamp 1698431365
transform 1 0 17808 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1342_
timestamp 1698431365
transform -1 0 17696 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1343_
timestamp 1698431365
transform 1 0 18816 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1344_
timestamp 1698431365
transform -1 0 19600 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1345_
timestamp 1698431365
transform 1 0 17808 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1346_
timestamp 1698431365
transform -1 0 20944 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1347_
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1348_
timestamp 1698431365
transform 1 0 20272 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1349_
timestamp 1698431365
transform 1 0 23856 0 -1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1350_
timestamp 1698431365
transform -1 0 24304 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1351_
timestamp 1698431365
transform 1 0 23744 0 -1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1352_
timestamp 1698431365
transform 1 0 20496 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1353_
timestamp 1698431365
transform 1 0 25088 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1354_
timestamp 1698431365
transform 1 0 24416 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1355_
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1356_
timestamp 1698431365
transform 1 0 24416 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1357_
timestamp 1698431365
transform 1 0 21616 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1358_
timestamp 1698431365
transform 1 0 23408 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1359_
timestamp 1698431365
transform 1 0 30800 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1360_
timestamp 1698431365
transform -1 0 26208 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1361_
timestamp 1698431365
transform -1 0 25088 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1362_
timestamp 1698431365
transform 1 0 21840 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1363_
timestamp 1698431365
transform 1 0 30128 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1364_
timestamp 1698431365
transform -1 0 7280 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1365_
timestamp 1698431365
transform 1 0 5264 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1366_
timestamp 1698431365
transform -1 0 30576 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1367_
timestamp 1698431365
transform -1 0 27104 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1368_
timestamp 1698431365
transform -1 0 28224 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1369_
timestamp 1698431365
transform -1 0 27552 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1370_
timestamp 1698431365
transform -1 0 20384 0 1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1371_
timestamp 1698431365
transform -1 0 19264 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1372_
timestamp 1698431365
transform -1 0 17024 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1373_
timestamp 1698431365
transform 1 0 16576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1374_
timestamp 1698431365
transform -1 0 26432 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1375_
timestamp 1698431365
transform -1 0 25536 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1376_
timestamp 1698431365
transform -1 0 19488 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1377_
timestamp 1698431365
transform -1 0 17696 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1378_
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1379_
timestamp 1698431365
transform 1 0 28336 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1380_
timestamp 1698431365
transform 1 0 26880 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1381_
timestamp 1698431365
transform -1 0 25984 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1382_
timestamp 1698431365
transform 1 0 31360 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1383_
timestamp 1698431365
transform 1 0 38080 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1384_
timestamp 1698431365
transform 1 0 39872 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1385_
timestamp 1698431365
transform 1 0 39648 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1386_
timestamp 1698431365
transform 1 0 37184 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1387_
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1388_
timestamp 1698431365
transform -1 0 36624 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1389_
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1390_
timestamp 1698431365
transform 1 0 37408 0 1 36064
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1391_
timestamp 1698431365
transform 1 0 39648 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1392_
timestamp 1698431365
transform 1 0 35840 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1393_
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1394_
timestamp 1698431365
transform -1 0 42224 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1395_
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1396_
timestamp 1698431365
transform 1 0 38080 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1397_
timestamp 1698431365
transform 1 0 39648 0 1 36064
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1398_
timestamp 1698431365
transform 1 0 39536 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1399_
timestamp 1698431365
transform 1 0 38752 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1400_
timestamp 1698431365
transform 1 0 41888 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1401_
timestamp 1698431365
transform -1 0 45136 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1402_
timestamp 1698431365
transform 1 0 43904 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1403_
timestamp 1698431365
transform -1 0 44016 0 1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1404_
timestamp 1698431365
transform 1 0 47264 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1405_
timestamp 1698431365
transform -1 0 46256 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1406_
timestamp 1698431365
transform 1 0 45696 0 1 32928
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1407_
timestamp 1698431365
transform -1 0 47712 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1408_
timestamp 1698431365
transform 1 0 47824 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1409_
timestamp 1698431365
transform -1 0 46816 0 -1 36064
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1410_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1411_
timestamp 1698431365
transform -1 0 15680 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1412_
timestamp 1698431365
transform -1 0 6160 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1413_
timestamp 1698431365
transform -1 0 10640 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1414_
timestamp 1698431365
transform -1 0 8288 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1415_
timestamp 1698431365
transform -1 0 11760 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1416_
timestamp 1698431365
transform -1 0 8960 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1417_
timestamp 1698431365
transform -1 0 9184 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1418_
timestamp 1698431365
transform -1 0 5936 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1419_
timestamp 1698431365
transform -1 0 12768 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1420_
timestamp 1698431365
transform -1 0 12208 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1421_
timestamp 1698431365
transform 1 0 2800 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1422_
timestamp 1698431365
transform -1 0 2800 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1423_
timestamp 1698431365
transform -1 0 12656 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1424_
timestamp 1698431365
transform -1 0 7504 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1425_
timestamp 1698431365
transform 1 0 3024 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1426_
timestamp 1698431365
transform -1 0 4928 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1427_
timestamp 1698431365
transform -1 0 3696 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1428_
timestamp 1698431365
transform 1 0 3696 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1429_
timestamp 1698431365
transform -1 0 3696 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1430_
timestamp 1698431365
transform 1 0 2576 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1431_
timestamp 1698431365
transform 1 0 4368 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1432_
timestamp 1698431365
transform -1 0 4368 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1433_
timestamp 1698431365
transform -1 0 3024 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1434_
timestamp 1698431365
transform 1 0 3920 0 -1 36064
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1435_
timestamp 1698431365
transform 1 0 6496 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1436_
timestamp 1698431365
transform -1 0 6608 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1437_
timestamp 1698431365
transform -1 0 41216 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1438_
timestamp 1698431365
transform -1 0 36400 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1439_
timestamp 1698431365
transform 1 0 36176 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1440_
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1441_
timestamp 1698431365
transform -1 0 36288 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1442_
timestamp 1698431365
transform -1 0 35280 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1443_
timestamp 1698431365
transform 1 0 32928 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1444_
timestamp 1698431365
transform 1 0 32928 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1445_
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1446_
timestamp 1698431365
transform 1 0 33152 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1447_
timestamp 1698431365
transform 1 0 30128 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1448_
timestamp 1698431365
transform -1 0 32368 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1449_
timestamp 1698431365
transform -1 0 31136 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1450_
timestamp 1698431365
transform 1 0 30352 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1451_
timestamp 1698431365
transform 1 0 30576 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1452_
timestamp 1698431365
transform 1 0 28336 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1453_
timestamp 1698431365
transform 1 0 30128 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1454_
timestamp 1698431365
transform -1 0 26992 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1455_
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1456_
timestamp 1698431365
transform 1 0 30016 0 -1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1457_
timestamp 1698431365
transform -1 0 33152 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1458_
timestamp 1698431365
transform 1 0 31696 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1459_
timestamp 1698431365
transform 1 0 31248 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1460_
timestamp 1698431365
transform -1 0 34832 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1461_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33488 0 -1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1462_
timestamp 1698431365
transform 1 0 35728 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1463_
timestamp 1698431365
transform -1 0 45136 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1464_
timestamp 1698431365
transform 1 0 42896 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1465_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42784 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1466_
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1467_
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1468_
timestamp 1698431365
transform 1 0 40880 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1469_
timestamp 1698431365
transform -1 0 45360 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1470_
timestamp 1698431365
transform 1 0 40208 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1471_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 43344 0 1 37632
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1472_
timestamp 1698431365
transform 1 0 44688 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1473_
timestamp 1698431365
transform 1 0 45472 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1474_
timestamp 1698431365
transform 1 0 46592 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1475_
timestamp 1698431365
transform 1 0 46480 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1476_
timestamp 1698431365
transform -1 0 47264 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1477_
timestamp 1698431365
transform 1 0 44688 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1478_
timestamp 1698431365
transform 1 0 45248 0 -1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1479_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 45248 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1480_
timestamp 1698431365
transform -1 0 45808 0 -1 37632
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1481_
timestamp 1698431365
transform -1 0 38080 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1482_
timestamp 1698431365
transform 1 0 36848 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1483_
timestamp 1698431365
transform -1 0 40544 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1484_
timestamp 1698431365
transform 1 0 42000 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1485_
timestamp 1698431365
transform 1 0 43344 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1486_
timestamp 1698431365
transform 1 0 43904 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1487_
timestamp 1698431365
transform 1 0 46256 0 -1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1488_
timestamp 1698431365
transform 1 0 37744 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1489_
timestamp 1698431365
transform 1 0 32144 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1490_
timestamp 1698431365
transform -1 0 31584 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1491_
timestamp 1698431365
transform -1 0 29456 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1492_
timestamp 1698431365
transform 1 0 28336 0 -1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1493_
timestamp 1698431365
transform 1 0 34384 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1494_
timestamp 1698431365
transform 1 0 29680 0 1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1495_
timestamp 1698431365
transform -1 0 36176 0 1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1496_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32592 0 -1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1497_
timestamp 1698431365
transform 1 0 31696 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1498_
timestamp 1698431365
transform 1 0 32816 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1499_
timestamp 1698431365
transform 1 0 45696 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1500_
timestamp 1698431365
transform -1 0 18816 0 -1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1501_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26544 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1502_
timestamp 1698431365
transform 1 0 15008 0 1 20384
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1503_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25872 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1504_
timestamp 1698431365
transform -1 0 27888 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1505_
timestamp 1698431365
transform 1 0 32256 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1506_
timestamp 1698431365
transform 1 0 32928 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1507_
timestamp 1698431365
transform -1 0 34608 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1508_
timestamp 1698431365
transform 1 0 10640 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1509_
timestamp 1698431365
transform -1 0 10080 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1510_
timestamp 1698431365
transform -1 0 9072 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1511_
timestamp 1698431365
transform -1 0 10640 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1512_
timestamp 1698431365
transform 1 0 9856 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1513_
timestamp 1698431365
transform 1 0 33824 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1514_
timestamp 1698431365
transform -1 0 26544 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1515_
timestamp 1698431365
transform -1 0 24192 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1516_
timestamp 1698431365
transform 1 0 31920 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1517_
timestamp 1698431365
transform 1 0 36512 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1518_
timestamp 1698431365
transform -1 0 34048 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1519_
timestamp 1698431365
transform -1 0 30800 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1520_
timestamp 1698431365
transform 1 0 27440 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1521_
timestamp 1698431365
transform 1 0 26992 0 -1 39200
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1522_
timestamp 1698431365
transform -1 0 27104 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1523_
timestamp 1698431365
transform 1 0 29232 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1524_
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1525_
timestamp 1698431365
transform -1 0 30800 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1526_
timestamp 1698431365
transform -1 0 34272 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1527_
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1528_
timestamp 1698431365
transform 1 0 31024 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1529_
timestamp 1698431365
transform -1 0 32928 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1530_
timestamp 1698431365
transform 1 0 33600 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1531_
timestamp 1698431365
transform -1 0 32704 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1532_
timestamp 1698431365
transform -1 0 31808 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1533_
timestamp 1698431365
transform 1 0 34272 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1534_
timestamp 1698431365
transform 1 0 30800 0 1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1535_
timestamp 1698431365
transform 1 0 33488 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1536_
timestamp 1698431365
transform 1 0 36288 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1537_
timestamp 1698431365
transform -1 0 38864 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1538_
timestamp 1698431365
transform -1 0 35840 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1539_
timestamp 1698431365
transform -1 0 35168 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1540_
timestamp 1698431365
transform 1 0 37408 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1541_
timestamp 1698431365
transform -1 0 47040 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1542_
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1543_
timestamp 1698431365
transform 1 0 37744 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1544_
timestamp 1698431365
transform -1 0 40768 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1545_
timestamp 1698431365
transform 1 0 37968 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1546_
timestamp 1698431365
transform -1 0 40320 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1547_
timestamp 1698431365
transform 1 0 38528 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1548_
timestamp 1698431365
transform 1 0 39200 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1549_
timestamp 1698431365
transform -1 0 41216 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1550_
timestamp 1698431365
transform -1 0 39984 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1551_
timestamp 1698431365
transform -1 0 38976 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1552_
timestamp 1698431365
transform -1 0 40544 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1553_
timestamp 1698431365
transform 1 0 40432 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1554_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 42784 0 -1 43904
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1555_
timestamp 1698431365
transform -1 0 41216 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1556_
timestamp 1698431365
transform 1 0 41216 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1557_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 39424 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1558_
timestamp 1698431365
transform 1 0 41328 0 1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1559_
timestamp 1698431365
transform -1 0 42784 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1560_
timestamp 1698431365
transform 1 0 43120 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1561_
timestamp 1698431365
transform 1 0 44464 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1562_
timestamp 1698431365
transform 1 0 46368 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1563_
timestamp 1698431365
transform 1 0 45248 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1564_
timestamp 1698431365
transform -1 0 48160 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1565_
timestamp 1698431365
transform 1 0 45920 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1566_
timestamp 1698431365
transform 1 0 47264 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1567_
timestamp 1698431365
transform 1 0 46032 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1568_
timestamp 1698431365
transform 1 0 47264 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1569_
timestamp 1698431365
transform -1 0 10640 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1570_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10192 0 1 37632
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1571_
timestamp 1698431365
transform -1 0 10416 0 1 34496
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1572_
timestamp 1698431365
transform -1 0 8400 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1573_
timestamp 1698431365
transform -1 0 8624 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1574_
timestamp 1698431365
transform 1 0 6608 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1575_
timestamp 1698431365
transform -1 0 9072 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1576_
timestamp 1698431365
transform -1 0 7840 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1577_
timestamp 1698431365
transform 1 0 7280 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1578_
timestamp 1698431365
transform 1 0 10976 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1579_
timestamp 1698431365
transform 1 0 6384 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1580_
timestamp 1698431365
transform -1 0 6944 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1581_
timestamp 1698431365
transform 1 0 7616 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1582_
timestamp 1698431365
transform 1 0 12096 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1583_
timestamp 1698431365
transform 1 0 10080 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1584_
timestamp 1698431365
transform -1 0 12096 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1585_
timestamp 1698431365
transform 1 0 9744 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1586_
timestamp 1698431365
transform 1 0 9632 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1587_
timestamp 1698431365
transform 1 0 10304 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1588_
timestamp 1698431365
transform 1 0 10192 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1589_
timestamp 1698431365
transform 1 0 9632 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1590_
timestamp 1698431365
transform 1 0 10192 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1591_
timestamp 1698431365
transform -1 0 7280 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1592_
timestamp 1698431365
transform -1 0 7056 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1593_
timestamp 1698431365
transform 1 0 7280 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1594_
timestamp 1698431365
transform -1 0 8960 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1595_
timestamp 1698431365
transform -1 0 8064 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1596_
timestamp 1698431365
transform -1 0 8960 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1597_
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1598_
timestamp 1698431365
transform -1 0 6160 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1599_
timestamp 1698431365
transform 1 0 6608 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1600_
timestamp 1698431365
transform -1 0 6608 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1601_
timestamp 1698431365
transform -1 0 6608 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1602_
timestamp 1698431365
transform 1 0 3024 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1603_
timestamp 1698431365
transform 1 0 4480 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1604_
timestamp 1698431365
transform -1 0 4256 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1605_
timestamp 1698431365
transform 1 0 3136 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1606_
timestamp 1698431365
transform 1 0 3584 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1607_
timestamp 1698431365
transform -1 0 6496 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1608_
timestamp 1698431365
transform -1 0 3248 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1609_
timestamp 1698431365
transform 1 0 4032 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1610_
timestamp 1698431365
transform -1 0 6496 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1611_
timestamp 1698431365
transform 1 0 4816 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1612_
timestamp 1698431365
transform 1 0 3808 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1613_
timestamp 1698431365
transform -1 0 6160 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1614_
timestamp 1698431365
transform -1 0 3808 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1615_
timestamp 1698431365
transform 1 0 4816 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1616_
timestamp 1698431365
transform 1 0 2912 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1617_
timestamp 1698431365
transform -1 0 4928 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1618_
timestamp 1698431365
transform 1 0 4368 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1619_
timestamp 1698431365
transform -1 0 5376 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1620_
timestamp 1698431365
transform -1 0 5936 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1621_
timestamp 1698431365
transform 1 0 3472 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1622_
timestamp 1698431365
transform 1 0 6496 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1623_
timestamp 1698431365
transform -1 0 7504 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1624_
timestamp 1698431365
transform -1 0 8064 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1625_
timestamp 1698431365
transform -1 0 11312 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1626_
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1627_
timestamp 1698431365
transform -1 0 7280 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1628_
timestamp 1698431365
transform 1 0 7504 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1629_
timestamp 1698431365
transform -1 0 6496 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1630_
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1631_
timestamp 1698431365
transform -1 0 7504 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1632_
timestamp 1698431365
transform -1 0 6944 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1633_
timestamp 1698431365
transform 1 0 6384 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1634_
timestamp 1698431365
transform 1 0 7616 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1635_
timestamp 1698431365
transform -1 0 9072 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1636_
timestamp 1698431365
transform -1 0 9072 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1637_
timestamp 1698431365
transform 1 0 8176 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1638_
timestamp 1698431365
transform -1 0 8736 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1639_
timestamp 1698431365
transform 1 0 8288 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1640_
timestamp 1698431365
transform -1 0 6272 0 -1 23520
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1641_
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1642_
timestamp 1698431365
transform 1 0 7168 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1643_
timestamp 1698431365
transform -1 0 9296 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1644_
timestamp 1698431365
transform -1 0 8960 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1645_
timestamp 1698431365
transform 1 0 8064 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1646_
timestamp 1698431365
transform -1 0 9184 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1647_
timestamp 1698431365
transform -1 0 7616 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1648_
timestamp 1698431365
transform -1 0 8176 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1649_
timestamp 1698431365
transform 1 0 8176 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1650_
timestamp 1698431365
transform 1 0 26768 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1651_
timestamp 1698431365
transform 1 0 28336 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1652_
timestamp 1698431365
transform -1 0 29568 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1653_
timestamp 1698431365
transform -1 0 30576 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1654_
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1655_
timestamp 1698431365
transform -1 0 28784 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1656_
timestamp 1698431365
transform 1 0 28112 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1657_
timestamp 1698431365
transform 1 0 28112 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1658_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28672 0 -1 14112
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1659_
timestamp 1698431365
transform 1 0 28784 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1660_
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1661_
timestamp 1698431365
transform 1 0 27552 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1662_
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1663_
timestamp 1698431365
transform 1 0 22624 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1664_
timestamp 1698431365
transform -1 0 23744 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1665_
timestamp 1698431365
transform -1 0 26768 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1666_
timestamp 1698431365
transform -1 0 26880 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1667_
timestamp 1698431365
transform -1 0 26432 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1668_
timestamp 1698431365
transform 1 0 25424 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1669_
timestamp 1698431365
transform -1 0 27440 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1670_
timestamp 1698431365
transform -1 0 34944 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1671_
timestamp 1698431365
transform -1 0 27776 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1672_
timestamp 1698431365
transform 1 0 25424 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1673_
timestamp 1698431365
transform -1 0 26656 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1674_
timestamp 1698431365
transform 1 0 28336 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1675_
timestamp 1698431365
transform -1 0 28336 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1676_
timestamp 1698431365
transform -1 0 26208 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1677_
timestamp 1698431365
transform -1 0 25984 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1678_
timestamp 1698431365
transform 1 0 22960 0 1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1679_
timestamp 1698431365
transform -1 0 24640 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1680_
timestamp 1698431365
transform 1 0 26208 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1681_
timestamp 1698431365
transform -1 0 15904 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1682_
timestamp 1698431365
transform 1 0 12880 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1683_
timestamp 1698431365
transform -1 0 11424 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1684_
timestamp 1698431365
transform 1 0 14000 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1685_
timestamp 1698431365
transform 1 0 14336 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1686_
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1687_
timestamp 1698431365
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1688_
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1689_
timestamp 1698431365
transform -1 0 12096 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1690_
timestamp 1698431365
transform -1 0 39200 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1691_
timestamp 1698431365
transform -1 0 38192 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1692_
timestamp 1698431365
transform 1 0 33824 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1693_
timestamp 1698431365
transform -1 0 39760 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1694_
timestamp 1698431365
transform -1 0 42336 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1695_
timestamp 1698431365
transform -1 0 39984 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1696_
timestamp 1698431365
transform 1 0 39984 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1697_
timestamp 1698431365
transform 1 0 34720 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1698_
timestamp 1698431365
transform 1 0 39760 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1699_
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1700_
timestamp 1698431365
transform -1 0 41328 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1701_
timestamp 1698431365
transform -1 0 38416 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1702_
timestamp 1698431365
transform 1 0 37184 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1703_
timestamp 1698431365
transform -1 0 45136 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1704_
timestamp 1698431365
transform 1 0 35504 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1705_
timestamp 1698431365
transform 1 0 41664 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1706_
timestamp 1698431365
transform -1 0 39872 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1707_
timestamp 1698431365
transform 1 0 39872 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1708_
timestamp 1698431365
transform 1 0 40320 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1709_
timestamp 1698431365
transform -1 0 41776 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1710_
timestamp 1698431365
transform -1 0 39760 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1711_
timestamp 1698431365
transform -1 0 40320 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1712_
timestamp 1698431365
transform -1 0 39872 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1713_
timestamp 1698431365
transform -1 0 40096 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1714_
timestamp 1698431365
transform 1 0 38752 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1715_
timestamp 1698431365
transform -1 0 44128 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1716_
timestamp 1698431365
transform 1 0 42000 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1717_
timestamp 1698431365
transform 1 0 42000 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1718_
timestamp 1698431365
transform -1 0 44912 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1719_
timestamp 1698431365
transform 1 0 42336 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1720_
timestamp 1698431365
transform 1 0 42672 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1721_
timestamp 1698431365
transform 1 0 38864 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1722_
timestamp 1698431365
transform -1 0 39984 0 1 10976
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1723_
timestamp 1698431365
transform 1 0 40544 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1724_
timestamp 1698431365
transform -1 0 42224 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1725_
timestamp 1698431365
transform 1 0 42336 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1726_
timestamp 1698431365
transform -1 0 43792 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1727_
timestamp 1698431365
transform -1 0 40544 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1728_
timestamp 1698431365
transform -1 0 42448 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1729_
timestamp 1698431365
transform -1 0 43456 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1730_
timestamp 1698431365
transform 1 0 40096 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1731_
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1732_
timestamp 1698431365
transform 1 0 37968 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1733_
timestamp 1698431365
transform 1 0 39984 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1734_
timestamp 1698431365
transform -1 0 42336 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1735_
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1736_
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1737_
timestamp 1698431365
transform 1 0 42112 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1738_
timestamp 1698431365
transform -1 0 40768 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1739_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 42112 0 1 7840
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1740_
timestamp 1698431365
transform -1 0 36176 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1741_
timestamp 1698431365
transform 1 0 35952 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1742_
timestamp 1698431365
transform 1 0 36288 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1743_
timestamp 1698431365
transform 1 0 35616 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1744_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37968 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1745_
timestamp 1698431365
transform 1 0 31696 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1746_
timestamp 1698431365
transform 1 0 35728 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1747_
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1748_
timestamp 1698431365
transform -1 0 38864 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1749_
timestamp 1698431365
transform 1 0 38752 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1750_
timestamp 1698431365
transform 1 0 40096 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1751_
timestamp 1698431365
transform 1 0 40992 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1752_
timestamp 1698431365
transform 1 0 41664 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1753_
timestamp 1698431365
transform 1 0 38976 0 -1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1754_
timestamp 1698431365
transform 1 0 42672 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1755_
timestamp 1698431365
transform 1 0 43792 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1756_
timestamp 1698431365
transform 1 0 43568 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1757_
timestamp 1698431365
transform 1 0 46032 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1758_
timestamp 1698431365
transform 1 0 43120 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1759_
timestamp 1698431365
transform 1 0 45024 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1760_
timestamp 1698431365
transform 1 0 45920 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1761_
timestamp 1698431365
transform -1 0 36624 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1762_
timestamp 1698431365
transform 1 0 30128 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1763_
timestamp 1698431365
transform 1 0 42336 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1764_
timestamp 1698431365
transform 1 0 43792 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1765_
timestamp 1698431365
transform 1 0 42448 0 1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1766_
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1767_
timestamp 1698431365
transform 1 0 45808 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1768_
timestamp 1698431365
transform 1 0 34048 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1769_
timestamp 1698431365
transform 1 0 43456 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1770_
timestamp 1698431365
transform 1 0 46704 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1771_
timestamp 1698431365
transform -1 0 45024 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1772_
timestamp 1698431365
transform -1 0 48048 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1773_
timestamp 1698431365
transform 1 0 43792 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1774_
timestamp 1698431365
transform 1 0 45136 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1775_
timestamp 1698431365
transform 1 0 46032 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1776_
timestamp 1698431365
transform -1 0 43904 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1777_
timestamp 1698431365
transform -1 0 44240 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1778_
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1779_
timestamp 1698431365
transform 1 0 45808 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1780_
timestamp 1698431365
transform 1 0 41216 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1781_
timestamp 1698431365
transform -1 0 43120 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1782_
timestamp 1698431365
transform -1 0 43232 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1783_
timestamp 1698431365
transform -1 0 41440 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1784_
timestamp 1698431365
transform 1 0 42336 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1785_
timestamp 1698431365
transform 1 0 43344 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1786_
timestamp 1698431365
transform 1 0 43680 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1787_
timestamp 1698431365
transform -1 0 42560 0 1 6272
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1788_
timestamp 1698431365
transform -1 0 38080 0 1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1789_
timestamp 1698431365
transform -1 0 29232 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1790_
timestamp 1698431365
transform -1 0 28112 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1791_
timestamp 1698431365
transform 1 0 27216 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1792_
timestamp 1698431365
transform -1 0 40768 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1793_
timestamp 1698431365
transform 1 0 35728 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1794_
timestamp 1698431365
transform -1 0 43120 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1795_
timestamp 1698431365
transform -1 0 43232 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1796_
timestamp 1698431365
transform -1 0 42336 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1797_
timestamp 1698431365
transform -1 0 43120 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1798_
timestamp 1698431365
transform -1 0 44352 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1799_
timestamp 1698431365
transform -1 0 45136 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1800_
timestamp 1698431365
transform -1 0 44464 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1801_
timestamp 1698431365
transform -1 0 44688 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1802_
timestamp 1698431365
transform 1 0 42000 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1803_
timestamp 1698431365
transform -1 0 44240 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1804_
timestamp 1698431365
transform 1 0 41888 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1805_
timestamp 1698431365
transform -1 0 43792 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1806_
timestamp 1698431365
transform -1 0 40544 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1807_
timestamp 1698431365
transform 1 0 38192 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1808_
timestamp 1698431365
transform 1 0 38976 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1809_
timestamp 1698431365
transform -1 0 38640 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1810_
timestamp 1698431365
transform 1 0 37744 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1811_
timestamp 1698431365
transform 1 0 38640 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1812_
timestamp 1698431365
transform 1 0 33600 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1813_
timestamp 1698431365
transform 1 0 37184 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1814_
timestamp 1698431365
transform 1 0 39424 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1815_
timestamp 1698431365
transform 1 0 39984 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1816_
timestamp 1698431365
transform 1 0 39424 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1817_
timestamp 1698431365
transform -1 0 41888 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1818_
timestamp 1698431365
transform 1 0 40096 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1819_
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1820_
timestamp 1698431365
transform 1 0 40880 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1821_
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1822_
timestamp 1698431365
transform 1 0 40656 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1823_
timestamp 1698431365
transform 1 0 46368 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1824_
timestamp 1698431365
transform -1 0 48272 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1825_
timestamp 1698431365
transform -1 0 47824 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1826_
timestamp 1698431365
transform 1 0 42448 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1827_
timestamp 1698431365
transform -1 0 43568 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1828_
timestamp 1698431365
transform -1 0 43344 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1829_
timestamp 1698431365
transform -1 0 43344 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1830_
timestamp 1698431365
transform 1 0 42336 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1831_
timestamp 1698431365
transform 1 0 41888 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1832_
timestamp 1698431365
transform -1 0 47824 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1833_
timestamp 1698431365
transform -1 0 45136 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1834_
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1835_
timestamp 1698431365
transform 1 0 42000 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1836_
timestamp 1698431365
transform 1 0 39872 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1837_
timestamp 1698431365
transform 1 0 42448 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1838_
timestamp 1698431365
transform 1 0 40880 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1839_
timestamp 1698431365
transform 1 0 42336 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1840_
timestamp 1698431365
transform 1 0 42112 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1841_
timestamp 1698431365
transform 1 0 41776 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1842_
timestamp 1698431365
transform 1 0 39200 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1843_
timestamp 1698431365
transform -1 0 43344 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1844_
timestamp 1698431365
transform -1 0 42112 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1845_
timestamp 1698431365
transform -1 0 42448 0 -1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1846_
timestamp 1698431365
transform -1 0 42224 0 1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1847_
timestamp 1698431365
transform 1 0 41216 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1848_
timestamp 1698431365
transform -1 0 35840 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1849_
timestamp 1698431365
transform -1 0 39312 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1850_
timestamp 1698431365
transform 1 0 37072 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1851_
timestamp 1698431365
transform -1 0 38640 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1852_
timestamp 1698431365
transform -1 0 38976 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1853_
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1854_
timestamp 1698431365
transform 1 0 35840 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1855_
timestamp 1698431365
transform 1 0 36736 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1856_
timestamp 1698431365
transform 1 0 38640 0 -1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1857_
timestamp 1698431365
transform -1 0 41552 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1858_
timestamp 1698431365
transform 1 0 38192 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1859_
timestamp 1698431365
transform -1 0 38192 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1860_
timestamp 1698431365
transform 1 0 38976 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1861_
timestamp 1698431365
transform 1 0 38080 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1862_
timestamp 1698431365
transform 1 0 39424 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1863_
timestamp 1698431365
transform 1 0 42448 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1864_
timestamp 1698431365
transform 1 0 43008 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1865_
timestamp 1698431365
transform 1 0 45584 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1866_
timestamp 1698431365
transform 1 0 42672 0 1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1867_
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1868_
timestamp 1698431365
transform -1 0 44128 0 1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1869_
timestamp 1698431365
transform 1 0 44688 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1870_
timestamp 1698431365
transform 1 0 44352 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1871_
timestamp 1698431365
transform 1 0 45696 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1872_
timestamp 1698431365
transform 1 0 43344 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1873_
timestamp 1698431365
transform 1 0 44800 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1874_
timestamp 1698431365
transform 1 0 45696 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1875_
timestamp 1698431365
transform 1 0 43568 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1876_
timestamp 1698431365
transform 1 0 44128 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1877_
timestamp 1698431365
transform 1 0 44912 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1878_
timestamp 1698431365
transform 1 0 47600 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1879_
timestamp 1698431365
transform 1 0 43568 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1880_
timestamp 1698431365
transform -1 0 46704 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1881_
timestamp 1698431365
transform -1 0 44464 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1882_
timestamp 1698431365
transform -1 0 43904 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1883_
timestamp 1698431365
transform 1 0 44352 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1884_
timestamp 1698431365
transform 1 0 46704 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1885_
timestamp 1698431365
transform 1 0 30688 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1886_
timestamp 1698431365
transform -1 0 32704 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1887_
timestamp 1698431365
transform -1 0 33040 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1888_
timestamp 1698431365
transform 1 0 17360 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1889_
timestamp 1698431365
transform -1 0 19376 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1890_
timestamp 1698431365
transform 1 0 12656 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1891_
timestamp 1698431365
transform -1 0 26208 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1892_
timestamp 1698431365
transform -1 0 22960 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1893_
timestamp 1698431365
transform 1 0 13440 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1894_
timestamp 1698431365
transform -1 0 21840 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1895_
timestamp 1698431365
transform -1 0 20160 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1896_
timestamp 1698431365
transform 1 0 17584 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1897_
timestamp 1698431365
transform -1 0 20160 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1898_
timestamp 1698431365
transform -1 0 19936 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1899_
timestamp 1698431365
transform 1 0 17920 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1900_
timestamp 1698431365
transform -1 0 19712 0 1 36064
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1901_
timestamp 1698431365
transform -1 0 19264 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1902_
timestamp 1698431365
transform -1 0 17024 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1903_
timestamp 1698431365
transform -1 0 20832 0 1 42336
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1904_
timestamp 1698431365
transform 1 0 18480 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1905_
timestamp 1698431365
transform 1 0 19040 0 -1 42336
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1906_
timestamp 1698431365
transform -1 0 25312 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1907_
timestamp 1698431365
transform -1 0 18032 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1908_
timestamp 1698431365
transform -1 0 20384 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1909_
timestamp 1698431365
transform -1 0 18704 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1910_
timestamp 1698431365
transform 1 0 19600 0 -1 45472
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1911_
timestamp 1698431365
transform 1 0 11872 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1912_
timestamp 1698431365
transform 1 0 22176 0 1 42336
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1913_
timestamp 1698431365
transform -1 0 24864 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1914_
timestamp 1698431365
transform -1 0 23744 0 -1 43904
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1915_
timestamp 1698431365
transform -1 0 20944 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1916_
timestamp 1698431365
transform -1 0 23744 0 -1 40768
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1917_
timestamp 1698431365
transform -1 0 15680 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1918_
timestamp 1698431365
transform -1 0 21168 0 -1 39200
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1919_
timestamp 1698431365
transform 1 0 21952 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1920_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 -1 39200
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1921_
timestamp 1698431365
transform -1 0 21728 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1922_
timestamp 1698431365
transform -1 0 14672 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1923_
timestamp 1698431365
transform 1 0 13776 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1924_
timestamp 1698431365
transform 1 0 14672 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1925_
timestamp 1698431365
transform 1 0 15456 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1926_
timestamp 1698431365
transform 1 0 17920 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1927_
timestamp 1698431365
transform -1 0 19152 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1928_
timestamp 1698431365
transform -1 0 20048 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1929_
timestamp 1698431365
transform 1 0 20048 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1930_
timestamp 1698431365
transform -1 0 20272 0 1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1931_
timestamp 1698431365
transform -1 0 18144 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1932_
timestamp 1698431365
transform 1 0 16128 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1933_
timestamp 1698431365
transform -1 0 14336 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1934_
timestamp 1698431365
transform -1 0 16576 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1935_
timestamp 1698431365
transform -1 0 14336 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1936_
timestamp 1698431365
transform 1 0 16576 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1937_
timestamp 1698431365
transform -1 0 17024 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1938_
timestamp 1698431365
transform 1 0 16352 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1939_
timestamp 1698431365
transform -1 0 18480 0 -1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1940_
timestamp 1698431365
transform -1 0 15456 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1941_
timestamp 1698431365
transform 1 0 15456 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1942_
timestamp 1698431365
transform -1 0 14672 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1943_
timestamp 1698431365
transform -1 0 13104 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1944_
timestamp 1698431365
transform -1 0 11872 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1945_
timestamp 1698431365
transform -1 0 11424 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1946_
timestamp 1698431365
transform 1 0 11200 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1947_
timestamp 1698431365
transform 1 0 12096 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1948_
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1949_
timestamp 1698431365
transform -1 0 11200 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1950_
timestamp 1698431365
transform 1 0 11536 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1951_
timestamp 1698431365
transform 1 0 9744 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1952_
timestamp 1698431365
transform -1 0 11536 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1953_
timestamp 1698431365
transform 1 0 11760 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1954_
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1955_
timestamp 1698431365
transform 1 0 12320 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1956_
timestamp 1698431365
transform 1 0 12432 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1957_
timestamp 1698431365
transform 1 0 22176 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1958_
timestamp 1698431365
transform 1 0 21280 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1959_
timestamp 1698431365
transform -1 0 24304 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1960_
timestamp 1698431365
transform -1 0 22176 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1961_
timestamp 1698431365
transform 1 0 20496 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1962_
timestamp 1698431365
transform 1 0 21280 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1963_
timestamp 1698431365
transform 1 0 20496 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1964_
timestamp 1698431365
transform 1 0 22400 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1965_
timestamp 1698431365
transform -1 0 13328 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1966_
timestamp 1698431365
transform 1 0 11536 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1967_
timestamp 1698431365
transform -1 0 15120 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1968_
timestamp 1698431365
transform 1 0 13552 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1969_
timestamp 1698431365
transform -1 0 13104 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1970_
timestamp 1698431365
transform 1 0 14112 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1971_
timestamp 1698431365
transform 1 0 14448 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1972_
timestamp 1698431365
transform 1 0 15568 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1973_
timestamp 1698431365
transform -1 0 15680 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1974_
timestamp 1698431365
transform 1 0 13440 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1975_
timestamp 1698431365
transform -1 0 14784 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1976_
timestamp 1698431365
transform -1 0 13888 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1977_
timestamp 1698431365
transform 1 0 14448 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1978_
timestamp 1698431365
transform 1 0 14336 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1979_
timestamp 1698431365
transform -1 0 14448 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1980_
timestamp 1698431365
transform -1 0 17024 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1981_
timestamp 1698431365
transform -1 0 15008 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1982_
timestamp 1698431365
transform 1 0 15344 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1983_
timestamp 1698431365
transform -1 0 16128 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1984_
timestamp 1698431365
transform -1 0 14000 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1985_
timestamp 1698431365
transform 1 0 44240 0 -1 32928
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1986_
timestamp 1698431365
transform -1 0 28336 0 1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1987_
timestamp 1698431365
transform -1 0 26096 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1988_
timestamp 1698431365
transform -1 0 25984 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1989_
timestamp 1698431365
transform -1 0 25760 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1990_
timestamp 1698431365
transform -1 0 23968 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1991_
timestamp 1698431365
transform 1 0 25760 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1992_
timestamp 1698431365
transform 1 0 26992 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1993_
timestamp 1698431365
transform 1 0 25760 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1994_
timestamp 1698431365
transform -1 0 26992 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1995_
timestamp 1698431365
transform -1 0 27552 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1996_
timestamp 1698431365
transform -1 0 27216 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1997_
timestamp 1698431365
transform -1 0 28112 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1998_
timestamp 1698431365
transform -1 0 26320 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1999_
timestamp 1698431365
transform -1 0 29568 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2000_
timestamp 1698431365
transform 1 0 31584 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2001_
timestamp 1698431365
transform -1 0 32704 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2002_
timestamp 1698431365
transform -1 0 32480 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2003_
timestamp 1698431365
transform -1 0 31920 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2004_
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2005_
timestamp 1698431365
transform -1 0 27216 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2006_
timestamp 1698431365
transform 1 0 29120 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2007_
timestamp 1698431365
transform -1 0 28448 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2008_
timestamp 1698431365
transform -1 0 31360 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2009_
timestamp 1698431365
transform -1 0 30240 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2010_
timestamp 1698431365
transform -1 0 31248 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2011_
timestamp 1698431365
transform 1 0 29120 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2012_
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2013_
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2014_
timestamp 1698431365
transform 1 0 33600 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2015_
timestamp 1698431365
transform 1 0 34608 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2016_
timestamp 1698431365
transform 1 0 36176 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2017_
timestamp 1698431365
transform -1 0 34272 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2018_
timestamp 1698431365
transform -1 0 34384 0 -1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2019_
timestamp 1698431365
transform -1 0 33376 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2020_
timestamp 1698431365
transform -1 0 35392 0 -1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2021_
timestamp 1698431365
transform -1 0 35392 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2022_
timestamp 1698431365
transform 1 0 15568 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2023_
timestamp 1698431365
transform -1 0 16464 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2024_
timestamp 1698431365
transform 1 0 17248 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2025_
timestamp 1698431365
transform -1 0 13104 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2026_
timestamp 1698431365
transform -1 0 11424 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2027_
timestamp 1698431365
transform -1 0 12208 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2028_
timestamp 1698431365
transform -1 0 11200 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2029_
timestamp 1698431365
transform 1 0 8848 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2030_
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2031_
timestamp 1698431365
transform -1 0 9408 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2032_
timestamp 1698431365
transform 1 0 9744 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2033_
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2034_
timestamp 1698431365
transform 1 0 10304 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2035_
timestamp 1698431365
transform 1 0 11424 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2036_
timestamp 1698431365
transform 1 0 12432 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2037_
timestamp 1698431365
transform -1 0 11984 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2038_
timestamp 1698431365
transform 1 0 11760 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2039_
timestamp 1698431365
transform 1 0 14672 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2040_
timestamp 1698431365
transform 1 0 14112 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2041_
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2042_
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2043_
timestamp 1698431365
transform 1 0 14672 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2044_
timestamp 1698431365
transform 1 0 13664 0 -1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2045_
timestamp 1698431365
transform -1 0 15568 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2046_
timestamp 1698431365
transform -1 0 24864 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2047_
timestamp 1698431365
transform -1 0 23632 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2048_
timestamp 1698431365
transform 1 0 23632 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2049_
timestamp 1698431365
transform -1 0 23632 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2050_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32256 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2051_
timestamp 1698431365
transform -1 0 33824 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2052_
timestamp 1698431365
transform -1 0 34160 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2053_
timestamp 1698431365
transform -1 0 32256 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2054_
timestamp 1698431365
transform -1 0 30464 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2055_
timestamp 1698431365
transform 1 0 31248 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2056_
timestamp 1698431365
transform 1 0 31248 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2057_
timestamp 1698431365
transform 1 0 35168 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2058_
timestamp 1698431365
transform 1 0 33824 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2059_
timestamp 1698431365
transform 1 0 20384 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2060_
timestamp 1698431365
transform 1 0 22288 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2061_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22288 0 -1 36064
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2062_
timestamp 1698431365
transform -1 0 23184 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2063_
timestamp 1698431365
transform -1 0 24640 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2064_
timestamp 1698431365
transform 1 0 15680 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2065_
timestamp 1698431365
transform -1 0 21616 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2066_
timestamp 1698431365
transform 1 0 15792 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2067_
timestamp 1698431365
transform 1 0 7168 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2068_
timestamp 1698431365
transform 1 0 11424 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2069_
timestamp 1698431365
transform 1 0 8064 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2070_
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2071_
timestamp 1698431365
transform 1 0 9856 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2072_
timestamp 1698431365
transform 1 0 21504 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2073_
timestamp 1698431365
transform -1 0 24304 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2074_
timestamp 1698431365
transform 1 0 17920 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2075_
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2076_
timestamp 1698431365
transform -1 0 20944 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2077_
timestamp 1698431365
transform 1 0 13664 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2078_
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2079_
timestamp 1698431365
transform 1 0 13328 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2080_
timestamp 1698431365
transform 1 0 16464 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2081_
timestamp 1698431365
transform 1 0 18368 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2082_
timestamp 1698431365
transform 1 0 17248 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2083_
timestamp 1698431365
transform 1 0 8064 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2084_
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2085_
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2086_
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2087_
timestamp 1698431365
transform -1 0 9072 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2088_
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2089_
timestamp 1698431365
transform 1 0 10080 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2090_
timestamp 1698431365
transform 1 0 30576 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2091_
timestamp 1698431365
transform 1 0 33152 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2092_
timestamp 1698431365
transform -1 0 37408 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2093_
timestamp 1698431365
transform 1 0 35504 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2094_
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2095_
timestamp 1698431365
transform -1 0 44464 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2096_
timestamp 1698431365
transform -1 0 48384 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2097_
timestamp 1698431365
transform -1 0 48384 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2098_
timestamp 1698431365
transform 1 0 33040 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2099_
timestamp 1698431365
transform 1 0 31696 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2100_
timestamp 1698431365
transform 1 0 36848 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2101_
timestamp 1698431365
transform 1 0 36288 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2102_
timestamp 1698431365
transform 1 0 29904 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2103_
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2104_
timestamp 1698431365
transform 1 0 33488 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2105_
timestamp 1698431365
transform 1 0 34272 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2106_
timestamp 1698431365
transform 1 0 39312 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2107_
timestamp 1698431365
transform -1 0 48160 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2108_
timestamp 1698431365
transform -1 0 48384 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2109_
timestamp 1698431365
transform 1 0 40992 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2110_
timestamp 1698431365
transform 1 0 25648 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2111_
timestamp 1698431365
transform 1 0 24080 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2112_
timestamp 1698431365
transform 1 0 27776 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2113_
timestamp 1698431365
transform 1 0 25312 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2114_
timestamp 1698431365
transform -1 0 32144 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2115_
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2116_
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2117_
timestamp 1698431365
transform -1 0 4816 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2118_
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2119_
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2120_
timestamp 1698431365
transform 1 0 5264 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2121_
timestamp 1698431365
transform 1 0 4032 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2122_
timestamp 1698431365
transform 1 0 6608 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2123_
timestamp 1698431365
transform -1 0 24416 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2124_
timestamp 1698431365
transform 1 0 17248 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2125_
timestamp 1698431365
transform 1 0 14896 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2126_
timestamp 1698431365
transform 1 0 14448 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2127_
timestamp 1698431365
transform 1 0 17360 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2128_
timestamp 1698431365
transform -1 0 20944 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2129_
timestamp 1698431365
transform -1 0 24864 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2130_
timestamp 1698431365
transform 1 0 20608 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2131_
timestamp 1698431365
transform 1 0 28224 0 1 45472
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2132_
timestamp 1698431365
transform -1 0 27664 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2133_
timestamp 1698431365
transform 1 0 29120 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2134_
timestamp 1698431365
transform 1 0 21616 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2135_
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2136_
timestamp 1698431365
transform 1 0 5152 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2137_
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2138_
timestamp 1698431365
transform -1 0 20496 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2139_
timestamp 1698431365
transform 1 0 23632 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2140_
timestamp 1698431365
transform 1 0 15792 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2141_
timestamp 1698431365
transform -1 0 30576 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2142_
timestamp 1698431365
transform 1 0 23632 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2143_
timestamp 1698431365
transform 1 0 36288 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2144_
timestamp 1698431365
transform 1 0 36960 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2145_
timestamp 1698431365
transform 1 0 36400 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2146_
timestamp 1698431365
transform 1 0 39536 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2147_
timestamp 1698431365
transform 1 0 40656 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2148_
timestamp 1698431365
transform 1 0 42224 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2149_
timestamp 1698431365
transform 1 0 45136 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2150_
timestamp 1698431365
transform 1 0 45136 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2151_
timestamp 1698431365
transform 1 0 9632 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2152_
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2153_
timestamp 1698431365
transform -1 0 4816 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2154_
timestamp 1698431365
transform -1 0 4816 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2155_
timestamp 1698431365
transform -1 0 4816 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2156_
timestamp 1698431365
transform 1 0 4816 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2157_
timestamp 1698431365
transform 1 0 6608 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2158_
timestamp 1698431365
transform 1 0 22960 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2159_
timestamp 1698431365
transform 1 0 25536 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2160_
timestamp 1698431365
transform 1 0 25536 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2161_
timestamp 1698431365
transform 1 0 27104 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2162_
timestamp 1698431365
transform 1 0 27552 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2163_
timestamp 1698431365
transform -1 0 36512 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2164_
timestamp 1698431365
transform 1 0 33376 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2165_
timestamp 1698431365
transform -1 0 40096 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2166_
timestamp 1698431365
transform 1 0 41216 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2167_
timestamp 1698431365
transform 1 0 37184 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2168_
timestamp 1698431365
transform -1 0 44464 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2169_
timestamp 1698431365
transform 1 0 40768 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2170_
timestamp 1698431365
transform 1 0 44688 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2171_
timestamp 1698431365
transform -1 0 48384 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2172_
timestamp 1698431365
transform -1 0 48384 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2173_
timestamp 1698431365
transform -1 0 48384 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2174_
timestamp 1698431365
transform 1 0 5040 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2175_
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2176_
timestamp 1698431365
transform -1 0 13104 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2177_
timestamp 1698431365
transform -1 0 12432 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2178_
timestamp 1698431365
transform 1 0 7840 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2179_
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2180_
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2181_
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2182_
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2183_
timestamp 1698431365
transform -1 0 4816 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2184_
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2185_
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2186_
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2187_
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2188_
timestamp 1698431365
transform 1 0 3472 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2189_
timestamp 1698431365
transform -1 0 10864 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2190_
timestamp 1698431365
transform -1 0 12656 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2191_
timestamp 1698431365
transform 1 0 5936 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2192_
timestamp 1698431365
transform -1 0 24416 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2193_
timestamp 1698431365
transform 1 0 24752 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2194_
timestamp 1698431365
transform 1 0 25088 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2195_
timestamp 1698431365
transform -1 0 28112 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2196_
timestamp 1698431365
transform 1 0 21616 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2197_
timestamp 1698431365
transform 1 0 25536 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2198_
timestamp 1698431365
transform 1 0 5152 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2199_
timestamp 1698431365
transform 1 0 9632 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2200_
timestamp 1698431365
transform -1 0 16688 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2201_
timestamp 1698431365
transform -1 0 14000 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2202_
timestamp 1698431365
transform 1 0 10192 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2203_
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2204_
timestamp 1698431365
transform 1 0 35392 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2205_
timestamp 1698431365
transform -1 0 44016 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2206_
timestamp 1698431365
transform -1 0 48384 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2207_
timestamp 1698431365
transform -1 0 48384 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2208_
timestamp 1698431365
transform -1 0 48384 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2209_
timestamp 1698431365
transform -1 0 48384 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2210_
timestamp 1698431365
transform -1 0 48384 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2211_
timestamp 1698431365
transform -1 0 48384 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2212_
timestamp 1698431365
transform -1 0 40544 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2213_
timestamp 1698431365
transform -1 0 47936 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2214_
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2215_
timestamp 1698431365
transform -1 0 28336 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2216_
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2217_
timestamp 1698431365
transform 1 0 36176 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2218_
timestamp 1698431365
transform 1 0 36736 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2219_
timestamp 1698431365
transform 1 0 37184 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2220_
timestamp 1698431365
transform 1 0 45136 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2221_
timestamp 1698431365
transform 1 0 45024 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2222_
timestamp 1698431365
transform 1 0 45136 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2223_
timestamp 1698431365
transform -1 0 48384 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2224_
timestamp 1698431365
transform -1 0 48384 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2225_
timestamp 1698431365
transform 1 0 45136 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2226_
timestamp 1698431365
transform 1 0 44016 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2227_
timestamp 1698431365
transform 1 0 45136 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2228_
timestamp 1698431365
transform -1 0 32256 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2229_
timestamp 1698431365
transform 1 0 14000 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2230_
timestamp 1698431365
transform 1 0 14224 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2231_
timestamp 1698431365
transform 1 0 15792 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2232_
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2233_
timestamp 1698431365
transform -1 0 20496 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2234_
timestamp 1698431365
transform 1 0 13664 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2235_
timestamp 1698431365
transform -1 0 13664 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2236_
timestamp 1698431365
transform -1 0 10752 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2237_
timestamp 1698431365
transform 1 0 5712 0 -1 43904
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2238_
timestamp 1698431365
transform 1 0 5936 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2239_
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2240_
timestamp 1698431365
transform 1 0 13328 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2241_
timestamp 1698431365
transform -1 0 23408 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2242_
timestamp 1698431365
transform -1 0 23856 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2243_
timestamp 1698431365
transform 1 0 16688 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2244_
timestamp 1698431365
transform 1 0 10752 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2245_
timestamp 1698431365
transform 1 0 13328 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2246_
timestamp 1698431365
transform 1 0 12768 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2247_
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2248_
timestamp 1698431365
transform 1 0 10528 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2249_
timestamp 1698431365
transform 1 0 11200 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2250_
timestamp 1698431365
transform 1 0 12208 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2251_
timestamp 1698431365
transform 1 0 21952 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2252_
timestamp 1698431365
transform 1 0 23072 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2253_
timestamp 1698431365
transform 1 0 26432 0 -1 26656
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2254_
timestamp 1698431365
transform 1 0 28112 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2255_
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2256_
timestamp 1698431365
transform 1 0 25536 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2257_
timestamp 1698431365
transform -1 0 28784 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2258_
timestamp 1698431365
transform 1 0 29008 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2259_
timestamp 1698431365
transform 1 0 28784 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2260_
timestamp 1698431365
transform -1 0 36176 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2261_
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2262_
timestamp 1698431365
transform 1 0 31696 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2263_
timestamp 1698431365
transform 1 0 33376 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2264_
timestamp 1698431365
transform -1 0 17248 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2265_
timestamp 1698431365
transform 1 0 9632 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2266_
timestamp 1698431365
transform 1 0 5936 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2267_
timestamp 1698431365
transform 1 0 5936 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2268_
timestamp 1698431365
transform 1 0 8176 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2269_
timestamp 1698431365
transform -1 0 16688 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2270_
timestamp 1698431365
transform -1 0 16464 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2271_
timestamp 1698431365
transform 1 0 13888 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2272_
timestamp 1698431365
transform -1 0 24528 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2273_
timestamp 1698431365
transform -1 0 20944 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1025__A2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16800 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1034__B1
timestamp 1698431365
transform 1 0 20384 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1038__B1
timestamp 1698431365
transform -1 0 16352 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1040__A3
timestamp 1698431365
transform 1 0 18144 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1043__A2
timestamp 1698431365
transform 1 0 18032 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1047__I
timestamp 1698431365
transform 1 0 31136 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1052__I
timestamp 1698431365
transform 1 0 28560 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1053__A3
timestamp 1698431365
transform 1 0 30240 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1053__A4
timestamp 1698431365
transform 1 0 29792 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1057__I
timestamp 1698431365
transform -1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1059__A1
timestamp 1698431365
transform 1 0 30352 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1063__I
timestamp 1698431365
transform -1 0 32256 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1066__I
timestamp 1698431365
transform 1 0 36400 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1067__A1
timestamp 1698431365
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1069__I
timestamp 1698431365
transform 1 0 35280 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1070__A1
timestamp 1698431365
transform 1 0 32032 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1073__I
timestamp 1698431365
transform 1 0 36400 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1074__A1
timestamp 1698431365
transform 1 0 31472 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1082__I
timestamp 1698431365
transform 1 0 24640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1083__A1
timestamp 1698431365
transform 1 0 32480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1088__A1
timestamp 1698431365
transform 1 0 38640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1090__A1
timestamp 1698431365
transform -1 0 33376 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1092__I
timestamp 1698431365
transform 1 0 30688 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1097__I
timestamp 1698431365
transform 1 0 21392 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1098__I
timestamp 1698431365
transform 1 0 33152 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1100__A1
timestamp 1698431365
transform -1 0 23744 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1101__A1
timestamp 1698431365
transform -1 0 21952 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1102__I
timestamp 1698431365
transform -1 0 24416 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1103__I
timestamp 1698431365
transform -1 0 23296 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1105__I
timestamp 1698431365
transform -1 0 37968 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1106__A1
timestamp 1698431365
transform 1 0 24640 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1108__I
timestamp 1698431365
transform -1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1111__A1
timestamp 1698431365
transform 1 0 17696 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1112__I
timestamp 1698431365
transform -1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1115__A1
timestamp 1698431365
transform 1 0 20272 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1116__I
timestamp 1698431365
transform -1 0 38752 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1117__A1
timestamp 1698431365
transform -1 0 23632 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1119__A2
timestamp 1698431365
transform 1 0 25312 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1119__B
timestamp 1698431365
transform -1 0 24192 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1120__A2
timestamp 1698431365
transform 1 0 22848 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1121__I
timestamp 1698431365
transform -1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1127__A1
timestamp 1698431365
transform 1 0 18368 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1139__A1
timestamp 1698431365
transform 1 0 16240 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1153__I
timestamp 1698431365
transform 1 0 12544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1156__A1
timestamp 1698431365
transform 1 0 9632 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1158__I
timestamp 1698431365
transform 1 0 12768 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1165__A1
timestamp 1698431365
transform 1 0 26432 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1166__A1
timestamp 1698431365
transform 1 0 17584 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1170__A1
timestamp 1698431365
transform 1 0 24528 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1172__B
timestamp 1698431365
transform 1 0 23408 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1174__I
timestamp 1698431365
transform 1 0 16800 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1175__I
timestamp 1698431365
transform 1 0 16352 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1176__I
timestamp 1698431365
transform 1 0 18032 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1189__I
timestamp 1698431365
transform -1 0 16912 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1200__A1
timestamp 1698431365
transform 1 0 15680 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1202__B
timestamp 1698431365
transform 1 0 11424 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1216__A1
timestamp 1698431365
transform -1 0 7840 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1223__I
timestamp 1698431365
transform 1 0 34720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1225__A1
timestamp 1698431365
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1225__A2
timestamp 1698431365
transform 1 0 34272 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1231__A1
timestamp 1698431365
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1233__A1
timestamp 1698431365
transform 1 0 34384 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1235__I
timestamp 1698431365
transform 1 0 39984 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1237__A1
timestamp 1698431365
transform -1 0 41216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1240__A1
timestamp 1698431365
transform -1 0 42672 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1243__A1
timestamp 1698431365
transform 1 0 46928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1246__A1
timestamp 1698431365
transform 1 0 47152 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1251__A1
timestamp 1698431365
transform 1 0 32480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1256__A1
timestamp 1698431365
transform -1 0 36176 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1258__A1
timestamp 1698431365
transform -1 0 35056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1263__A1
timestamp 1698431365
transform 1 0 33376 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1265__A1
timestamp 1698431365
transform 1 0 32256 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1267__I
timestamp 1698431365
transform 1 0 34944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1268__A1
timestamp 1698431365
transform -1 0 34720 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1270__I
timestamp 1698431365
transform -1 0 35280 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1271__A1
timestamp 1698431365
transform 1 0 35392 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1273__I
timestamp 1698431365
transform 1 0 35952 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1274__A1
timestamp 1698431365
transform 1 0 35840 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1278__A1
timestamp 1698431365
transform 1 0 42448 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1280__A1
timestamp 1698431365
transform 1 0 43456 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1282__A1
timestamp 1698431365
transform 1 0 44240 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1284__A1
timestamp 1698431365
transform 1 0 43680 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1287__A1
timestamp 1698431365
transform 1 0 25200 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1291__C
timestamp 1698431365
transform -1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1300__A2
timestamp 1698431365
transform -1 0 5936 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1301__A2
timestamp 1698431365
transform -1 0 4928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1308__B
timestamp 1698431365
transform 1 0 4368 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1311__B
timestamp 1698431365
transform 1 0 5040 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1315__B
timestamp 1698431365
transform -1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1318__B
timestamp 1698431365
transform -1 0 8848 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1320__I
timestamp 1698431365
transform 1 0 22736 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1323__A1
timestamp 1698431365
transform 1 0 8176 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1329__A1
timestamp 1698431365
transform 1 0 22400 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1331__A1
timestamp 1698431365
transform 1 0 26208 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1332__I
timestamp 1698431365
transform -1 0 39424 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1334__A1
timestamp 1698431365
transform 1 0 23072 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1337__A1
timestamp 1698431365
transform -1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1339__A1
timestamp 1698431365
transform -1 0 18816 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1341__A1
timestamp 1698431365
transform -1 0 20048 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1343__A1
timestamp 1698431365
transform 1 0 20048 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1345__A1
timestamp 1698431365
transform 1 0 16800 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1349__A1
timestamp 1698431365
transform -1 0 25536 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1351__A1
timestamp 1698431365
transform -1 0 27216 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1353__A1
timestamp 1698431365
transform 1 0 26320 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1355__A1
timestamp 1698431365
transform 1 0 26320 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1357__I
timestamp 1698431365
transform 1 0 22512 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1358__I
timestamp 1698431365
transform 1 0 25312 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1359__A1
timestamp 1698431365
transform 1 0 31584 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1362__C
timestamp 1698431365
transform 1 0 26880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1364__A1
timestamp 1698431365
transform 1 0 7504 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1368__A1
timestamp 1698431365
transform 1 0 28448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1370__A1
timestamp 1698431365
transform 1 0 20608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1372__A1
timestamp 1698431365
transform -1 0 17696 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1374__A1
timestamp 1698431365
transform 1 0 27328 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1376__A1
timestamp 1698431365
transform -1 0 19712 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1378__A1
timestamp 1698431365
transform 1 0 29680 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1380__A1
timestamp 1698431365
transform 1 0 27104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1385__A1
timestamp 1698431365
transform 1 0 39312 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1386__A1
timestamp 1698431365
transform 1 0 37408 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1389__A1
timestamp 1698431365
transform 1 0 36400 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1396__A1
timestamp 1698431365
transform 1 0 38864 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1398__A1
timestamp 1698431365
transform 1 0 39648 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1399__A1
timestamp 1698431365
transform 1 0 41664 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1400__I
timestamp 1698431365
transform 1 0 41664 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1403__A1
timestamp 1698431365
transform -1 0 42784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1406__A1
timestamp 1698431365
transform 1 0 44912 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1409__A1
timestamp 1698431365
transform -1 0 42336 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1411__I
timestamp 1698431365
transform -1 0 15904 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1419__A1
timestamp 1698431365
transform -1 0 13776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1420__I
timestamp 1698431365
transform -1 0 12432 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1423__A1
timestamp 1698431365
transform -1 0 11312 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1501__A1
timestamp 1698431365
transform -1 0 28896 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1501__A2
timestamp 1698431365
transform 1 0 29120 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1503__A1
timestamp 1698431365
transform 1 0 28560 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1503__A2
timestamp 1698431365
transform 1 0 29568 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1503__A3
timestamp 1698431365
transform 1 0 26768 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1505__I
timestamp 1698431365
transform 1 0 32256 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1507__B
timestamp 1698431365
transform 1 0 34160 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1508__A2
timestamp 1698431365
transform 1 0 11536 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1511__A2
timestamp 1698431365
transform 1 0 10864 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1514__A2
timestamp 1698431365
transform -1 0 26768 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1516__A1
timestamp 1698431365
transform 1 0 32704 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1516__A2
timestamp 1698431365
transform 1 0 33152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1520__A2
timestamp 1698431365
transform 1 0 27216 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1522__A1
timestamp 1698431365
transform -1 0 26208 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1525__A1
timestamp 1698431365
transform 1 0 31248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1555__C
timestamp 1698431365
transform 1 0 39872 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1566__A1
timestamp 1698431365
transform 1 0 48160 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1576__A1
timestamp 1698431365
transform 1 0 8624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1579__A1
timestamp 1698431365
transform 1 0 6944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1583__I
timestamp 1698431365
transform 1 0 10752 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1595__I
timestamp 1698431365
transform 1 0 9632 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1610__I
timestamp 1698431365
transform 1 0 6720 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1625__I
timestamp 1698431365
transform 1 0 11312 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1639__B
timestamp 1698431365
transform 1 0 9184 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1648__B
timestamp 1698431365
transform 1 0 7056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1663__A1
timestamp 1698431365
transform 1 0 22400 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1664__A1
timestamp 1698431365
transform 1 0 24416 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1665__A1
timestamp 1698431365
transform 1 0 25424 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__A2
timestamp 1698431365
transform 1 0 26880 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1669__A3
timestamp 1698431365
transform -1 0 27552 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1671__A2
timestamp 1698431365
transform 1 0 28000 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1681__A1
timestamp 1698431365
transform -1 0 16128 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1681__A2
timestamp 1698431365
transform 1 0 14560 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1682__A1
timestamp 1698431365
transform 1 0 14112 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1684__A1
timestamp 1698431365
transform 1 0 15008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1686__A1
timestamp 1698431365
transform -1 0 14784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__A1
timestamp 1698431365
transform -1 0 14000 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__A2
timestamp 1698431365
transform 1 0 14112 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1691__A2
timestamp 1698431365
transform 1 0 39088 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1740__A1
timestamp 1698431365
transform 1 0 36512 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1740__B
timestamp 1698431365
transform 1 0 34944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1742__A2
timestamp 1698431365
transform -1 0 37296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1745__I
timestamp 1698431365
transform 1 0 31472 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1750__A1
timestamp 1698431365
transform 1 0 40992 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1753__A4
timestamp 1698431365
transform -1 0 38976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1759__A1
timestamp 1698431365
transform 1 0 44912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1762__A1
timestamp 1698431365
transform -1 0 29680 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1762__A2
timestamp 1698431365
transform 1 0 29904 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1766__A1
timestamp 1698431365
transform -1 0 45136 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1766__A2
timestamp 1698431365
transform 1 0 46704 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1768__I
timestamp 1698431365
transform -1 0 34048 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1771__A1
timestamp 1698431365
transform 1 0 44912 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1771__A2
timestamp 1698431365
transform -1 0 44688 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1774__A1
timestamp 1698431365
transform -1 0 45136 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1778__A1
timestamp 1698431365
transform -1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1778__A2
timestamp 1698431365
transform 1 0 46704 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1788__A1
timestamp 1698431365
transform 1 0 37520 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1788__A2
timestamp 1698431365
transform 1 0 38752 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1788__C
timestamp 1698431365
transform 1 0 38304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__A1
timestamp 1698431365
transform 1 0 29456 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__A2
timestamp 1698431365
transform 1 0 29456 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1790__A2
timestamp 1698431365
transform 1 0 28336 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1790__A3
timestamp 1698431365
transform 1 0 28336 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1791__B
timestamp 1698431365
transform -1 0 28560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1793__A2
timestamp 1698431365
transform 1 0 35504 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1848__B
timestamp 1698431365
transform 1 0 35504 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1853__A3
timestamp 1698431365
transform 1 0 36400 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1854__A2
timestamp 1698431365
transform 1 0 37856 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1856__A4
timestamp 1698431365
transform 1 0 37520 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1887__A1
timestamp 1698431365
transform 1 0 32032 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1889__A2
timestamp 1698431365
transform 1 0 16800 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1920__C
timestamp 1698431365
transform -1 0 25312 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1921__A1
timestamp 1698431365
transform -1 0 17920 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1926__A3
timestamp 1698431365
transform -1 0 16576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1927__A2
timestamp 1698431365
transform -1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1930__A4
timestamp 1698431365
transform -1 0 18480 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1957__B
timestamp 1698431365
transform 1 0 23408 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1960__A1
timestamp 1698431365
transform 1 0 24304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1962__A1
timestamp 1698431365
transform -1 0 16800 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1964__A1
timestamp 1698431365
transform 1 0 24304 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1968__B
timestamp 1698431365
transform 1 0 12880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1972__A1
timestamp 1698431365
transform -1 0 16912 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1984__A1
timestamp 1698431365
transform -1 0 14448 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1986__A1
timestamp 1698431365
transform 1 0 31136 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1986__A2
timestamp 1698431365
transform 1 0 30688 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1986__A3
timestamp 1698431365
transform -1 0 30464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1988__A1
timestamp 1698431365
transform 1 0 27440 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1988__A2
timestamp 1698431365
transform 1 0 27888 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1990__B
timestamp 1698431365
transform 1 0 22960 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1992__B
timestamp 1698431365
transform 1 0 24640 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1994__A1
timestamp 1698431365
transform 1 0 28336 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1994__B
timestamp 1698431365
transform 1 0 24528 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1996__B
timestamp 1698431365
transform -1 0 25536 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1998__A1
timestamp 1698431365
transform 1 0 26320 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1998__B
timestamp 1698431365
transform 1 0 24080 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2002__A1
timestamp 1698431365
transform 1 0 31584 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2006__A1
timestamp 1698431365
transform -1 0 31584 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2010__A1
timestamp 1698431365
transform 1 0 34496 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2014__A1
timestamp 1698431365
transform 1 0 34608 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2018__A1
timestamp 1698431365
transform 1 0 35616 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2020__A1
timestamp 1698431365
transform 1 0 36064 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2039__B
timestamp 1698431365
transform -1 0 15792 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2043__A1
timestamp 1698431365
transform 1 0 15568 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2047__A1
timestamp 1698431365
transform 1 0 23856 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2049__A1
timestamp 1698431365
transform -1 0 24752 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 25312 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_0__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 26768 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_1__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 21392 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_2__f_wb_clk_i_I
timestamp 1698431365
transform -1 0 37296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_3__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 36400 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 8960 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_1_wb_clk_i_I
timestamp 1698431365
transform 1 0 16352 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_2_wb_clk_i_I
timestamp 1698431365
transform 1 0 26320 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_3_wb_clk_i_I
timestamp 1698431365
transform 1 0 18032 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_4_wb_clk_i_I
timestamp 1698431365
transform 1 0 19152 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_5_wb_clk_i_I
timestamp 1698431365
transform 1 0 9632 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_6_wb_clk_i_I
timestamp 1698431365
transform 1 0 9632 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_7_wb_clk_i_I
timestamp 1698431365
transform 1 0 12544 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_8_wb_clk_i_I
timestamp 1698431365
transform 1 0 11312 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_9_wb_clk_i_I
timestamp 1698431365
transform 1 0 13104 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_10_wb_clk_i_I
timestamp 1698431365
transform 1 0 17808 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_11_wb_clk_i_I
timestamp 1698431365
transform 1 0 18704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_12_wb_clk_i_I
timestamp 1698431365
transform 1 0 21392 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_13_wb_clk_i_I
timestamp 1698431365
transform 1 0 16352 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_14_wb_clk_i_I
timestamp 1698431365
transform 1 0 24976 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_15_wb_clk_i_I
timestamp 1698431365
transform 1 0 35392 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_16_wb_clk_i_I
timestamp 1698431365
transform 1 0 32368 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_17_wb_clk_i_I
timestamp 1698431365
transform 1 0 41888 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_18_wb_clk_i_I
timestamp 1698431365
transform -1 0 41776 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_19_wb_clk_i_I
timestamp 1698431365
transform 1 0 42560 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_20_wb_clk_i_I
timestamp 1698431365
transform 1 0 44240 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_21_wb_clk_i_I
timestamp 1698431365
transform 1 0 44128 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_22_wb_clk_i_I
timestamp 1698431365
transform 1 0 43680 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_23_wb_clk_i_I
timestamp 1698431365
transform 1 0 38752 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_24_wb_clk_i_I
timestamp 1698431365
transform 1 0 42560 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_25_wb_clk_i_I
timestamp 1698431365
transform 1 0 43344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_26_wb_clk_i_I
timestamp 1698431365
transform 1 0 42112 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_27_wb_clk_i_I
timestamp 1698431365
transform 1 0 41776 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_28_wb_clk_i_I
timestamp 1698431365
transform 1 0 45472 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_29_wb_clk_i_I
timestamp 1698431365
transform 1 0 39984 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_30_wb_clk_i_I
timestamp 1698431365
transform 1 0 32480 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_31_wb_clk_i_I
timestamp 1698431365
transform 1 0 37632 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_32_wb_clk_i_I
timestamp 1698431365
transform 1 0 40320 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_33_wb_clk_i_I
timestamp 1698431365
transform 1 0 24864 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_34_wb_clk_i_I
timestamp 1698431365
transform 1 0 25312 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_35_wb_clk_i_I
timestamp 1698431365
transform 1 0 20832 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_36_wb_clk_i_I
timestamp 1698431365
transform 1 0 23856 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_37_wb_clk_i_I
timestamp 1698431365
transform 1 0 15568 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_38_wb_clk_i_I
timestamp 1698431365
transform 1 0 11312 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_39_wb_clk_i_I
timestamp 1698431365
transform 1 0 11088 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 48160 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 45024 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 47712 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 47712 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 47712 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 48272 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 47712 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 47488 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 41776 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform -1 0 43904 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform 1 0 33152 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform -1 0 43232 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform -1 0 18592 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output19_I
timestamp 1698431365
transform 1 0 31024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output20_I
timestamp 1698431365
transform 1 0 41552 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25536 0 -1 25088
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_wb_clk_i
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_wb_clk_i
timestamp 1698431365
transform -1 0 20944 0 1 29792
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_wb_clk_i
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_wb_clk_i
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_0_wb_clk_i
timestamp 1698431365
transform -1 0 8624 0 -1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_1_wb_clk_i
timestamp 1698431365
transform -1 0 16128 0 -1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_2_wb_clk_i
timestamp 1698431365
transform -1 0 22848 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_3_wb_clk_i
timestamp 1698431365
transform -1 0 26768 0 1 25088
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_4_wb_clk_i
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_5_wb_clk_i
timestamp 1698431365
transform -1 0 8848 0 -1 28224
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_6_wb_clk_i
timestamp 1698431365
transform -1 0 8512 0 -1 32928
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_7_wb_clk_i
timestamp 1698431365
transform -1 0 12320 0 1 36064
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_8_wb_clk_i
timestamp 1698431365
transform -1 0 11088 0 1 40768
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_9_wb_clk_i
timestamp 1698431365
transform -1 0 13104 0 1 42336
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_10_wb_clk_i
timestamp 1698431365
transform -1 0 19712 0 1 40768
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_11_wb_clk_i
timestamp 1698431365
transform -1 0 26768 0 1 43904
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_12_wb_clk_i
timestamp 1698431365
transform -1 0 28224 0 1 37632
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_13_wb_clk_i
timestamp 1698431365
transform -1 0 24416 0 -1 32928
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_14_wb_clk_i
timestamp 1698431365
transform 1 0 25200 0 -1 29792
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_15_wb_clk_i
timestamp 1698431365
transform -1 0 35168 0 1 34496
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_16_wb_clk_i
timestamp 1698431365
transform -1 0 32368 0 -1 43904
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_17_wb_clk_i
timestamp 1698431365
transform -1 0 40544 0 -1 40768
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_18_wb_clk_i
timestamp 1698431365
transform 1 0 41776 0 -1 45472
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_19_wb_clk_i
timestamp 1698431365
transform 1 0 42784 0 -1 42336
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_20_wb_clk_i
timestamp 1698431365
transform 1 0 42784 0 -1 34496
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_21_wb_clk_i
timestamp 1698431365
transform 1 0 42784 0 -1 28224
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_22_wb_clk_i
timestamp 1698431365
transform -1 0 42448 0 1 28224
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_23_wb_clk_i
timestamp 1698431365
transform -1 0 36624 0 1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_24_wb_clk_i
timestamp 1698431365
transform 1 0 37296 0 1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_25_wb_clk_i
timestamp 1698431365
transform 1 0 42784 0 -1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_26_wb_clk_i
timestamp 1698431365
transform 1 0 42784 0 -1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_27_wb_clk_i
timestamp 1698431365
transform 1 0 42784 0 -1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_28_wb_clk_i
timestamp 1698431365
transform 1 0 42448 0 -1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_29_wb_clk_i
timestamp 1698431365
transform -1 0 39312 0 -1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_30_wb_clk_i
timestamp 1698431365
transform -1 0 32480 0 -1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_31_wb_clk_i
timestamp 1698431365
transform -1 0 36624 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_32_wb_clk_i
timestamp 1698431365
transform -1 0 38528 0 -1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_33_wb_clk_i
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_34_wb_clk_i
timestamp 1698431365
transform -1 0 24752 0 -1 14112
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_35_wb_clk_i
timestamp 1698431365
transform -1 0 27664 0 1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_36_wb_clk_i
timestamp 1698431365
transform -1 0 22848 0 -1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_37_wb_clk_i
timestamp 1698431365
transform -1 0 15344 0 -1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_38_wb_clk_i
timestamp 1698431365
transform -1 0 11088 0 1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_39_wb_clk_i
timestamp 1698431365
transform -1 0 11088 0 1 14112
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_18 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3360 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_20 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3584 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_25 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4144 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_33
timestamp 1698431365
transform 1 0 5040 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_40
timestamp 1698431365
transform 1 0 5824 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_48
timestamp 1698431365
transform 1 0 6720 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_59
timestamp 1698431365
transform 1 0 7952 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_67
timestamp 1698431365
transform 1 0 8848 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_70 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_74
timestamp 1698431365
transform 1 0 9632 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_76
timestamp 1698431365
transform 1 0 9856 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_81
timestamp 1698431365
transform 1 0 10416 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_89
timestamp 1698431365
transform 1 0 11312 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_95
timestamp 1698431365
transform 1 0 11984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_97
timestamp 1698431365
transform 1 0 12208 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_174
timestamp 1698431365
transform 1 0 20832 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698431365
transform 1 0 23856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698431365
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_216
timestamp 1698431365
transform 1 0 25536 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_221
timestamp 1698431365
transform 1 0 26096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_223
timestamp 1698431365
transform 1 0 26320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_230
timestamp 1698431365
transform 1 0 27104 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_235
timestamp 1698431365
transform 1 0 27664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_237
timestamp 1698431365
transform 1 0 27888 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_303
timestamp 1698431365
transform 1 0 35280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_305
timestamp 1698431365
transform 1 0 35504 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_338
timestamp 1698431365
transform 1 0 39200 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_372
timestamp 1698431365
transform 1 0 43008 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_376
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_392
timestamp 1698431365
transform 1 0 45248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_396
timestamp 1698431365
transform 1 0 45696 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_398
timestamp 1698431365
transform 1 0 45920 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_403
timestamp 1698431365
transform 1 0 46480 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_407
timestamp 1698431365
transform 1 0 46928 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_410
timestamp 1698431365
transform 1 0 47264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_2
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_18
timestamp 1698431365
transform 1 0 3360 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_22
timestamp 1698431365
transform 1 0 3808 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_59
timestamp 1698431365
transform 1 0 7952 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_63
timestamp 1698431365
transform 1 0 8400 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_76
timestamp 1698431365
transform 1 0 9856 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_151
timestamp 1698431365
transform 1 0 18256 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_216
timestamp 1698431365
transform 1 0 25536 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_246
timestamp 1698431365
transform 1 0 28896 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_277
timestamp 1698431365
transform 1 0 32368 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698431365
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_319
timestamp 1698431365
transform 1 0 37072 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_366
timestamp 1698431365
transform 1 0 42336 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_417
timestamp 1698431365
transform 1 0 48048 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_419
timestamp 1698431365
transform 1 0 48272 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_44
timestamp 1698431365
transform 1 0 6272 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_46
timestamp 1698431365
transform 1 0 6496 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_115
timestamp 1698431365
transform 1 0 14224 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_119
timestamp 1698431365
transform 1 0 14672 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_173
timestamp 1698431365
transform 1 0 20720 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_193
timestamp 1698431365
transform 1 0 22960 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_214
timestamp 1698431365
transform 1 0 25312 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_222
timestamp 1698431365
transform 1 0 26208 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_226
timestamp 1698431365
transform 1 0 26656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_230
timestamp 1698431365
transform 1 0 27104 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_234
timestamp 1698431365
transform 1 0 27552 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_263
timestamp 1698431365
transform 1 0 30800 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_314
timestamp 1698431365
transform 1 0 36512 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_349
timestamp 1698431365
transform 1 0 40432 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_364
timestamp 1698431365
transform 1 0 42112 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_378
timestamp 1698431365
transform 1 0 43680 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_382
timestamp 1698431365
transform 1 0 44128 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_416
timestamp 1698431365
transform 1 0 47936 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_18
timestamp 1698431365
transform 1 0 3360 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_22
timestamp 1698431365
transform 1 0 3808 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_38
timestamp 1698431365
transform 1 0 5600 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_63
timestamp 1698431365
transform 1 0 8400 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_67
timestamp 1698431365
transform 1 0 8848 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_69
timestamp 1698431365
transform 1 0 9072 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_74
timestamp 1698431365
transform 1 0 9632 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_125
timestamp 1698431365
transform 1 0 15344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_129
timestamp 1698431365
transform 1 0 15792 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_144
timestamp 1698431365
transform 1 0 17472 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_179
timestamp 1698431365
transform 1 0 21392 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_209
timestamp 1698431365
transform 1 0 24752 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_278
timestamp 1698431365
transform 1 0 32480 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_295
timestamp 1698431365
transform 1 0 34384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_297
timestamp 1698431365
transform 1 0 34608 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_331
timestamp 1698431365
transform 1 0 38416 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_335
timestamp 1698431365
transform 1 0 38864 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_349
timestamp 1698431365
transform 1 0 40432 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_363
timestamp 1698431365
transform 1 0 42000 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_374
timestamp 1698431365
transform 1 0 43232 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_383
timestamp 1698431365
transform 1 0 44240 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_387
timestamp 1698431365
transform 1 0 44688 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_31
timestamp 1698431365
transform 1 0 4816 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_59
timestamp 1698431365
transform 1 0 7952 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_89
timestamp 1698431365
transform 1 0 11312 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_93
timestamp 1698431365
transform 1 0 11760 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_145
timestamp 1698431365
transform 1 0 17584 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_183
timestamp 1698431365
transform 1 0 21840 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_235
timestamp 1698431365
transform 1 0 27664 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_268
timestamp 1698431365
transform 1 0 31360 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_272
timestamp 1698431365
transform 1 0 31808 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_276
timestamp 1698431365
transform 1 0 32256 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_280
timestamp 1698431365
transform 1 0 32704 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_313
timestamp 1698431365
transform 1 0 36400 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_357
timestamp 1698431365
transform 1 0 41328 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_383
timestamp 1698431365
transform 1 0 44240 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_403
timestamp 1698431365
transform 1 0 46480 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_407
timestamp 1698431365
transform 1 0 46928 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_411
timestamp 1698431365
transform 1 0 47376 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_10
timestamp 1698431365
transform 1 0 2464 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_34
timestamp 1698431365
transform 1 0 5152 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_107
timestamp 1698431365
transform 1 0 13328 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_109
timestamp 1698431365
transform 1 0 13552 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_139
timestamp 1698431365
transform 1 0 16912 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_198
timestamp 1698431365
transform 1 0 23520 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_243
timestamp 1698431365
transform 1 0 28560 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_245
timestamp 1698431365
transform 1 0 28784 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_275
timestamp 1698431365
transform 1 0 32144 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_343
timestamp 1698431365
transform 1 0 39760 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_347
timestamp 1698431365
transform 1 0 40208 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_349
timestamp 1698431365
transform 1 0 40432 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_352
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_354
timestamp 1698431365
transform 1 0 40992 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_365
timestamp 1698431365
transform 1 0 42224 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_390
timestamp 1698431365
transform 1 0 45024 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_31
timestamp 1698431365
transform 1 0 4816 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_112
timestamp 1698431365
transform 1 0 13888 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_128
timestamp 1698431365
transform 1 0 15680 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_144
timestamp 1698431365
transform 1 0 17472 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_157
timestamp 1698431365
transform 1 0 18928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_159
timestamp 1698431365
transform 1 0 19152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_186
timestamp 1698431365
transform 1 0 22176 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_198
timestamp 1698431365
transform 1 0 23520 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_205
timestamp 1698431365
transform 1 0 24304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_209
timestamp 1698431365
transform 1 0 24752 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_239
timestamp 1698431365
transform 1 0 28112 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_261
timestamp 1698431365
transform 1 0 30576 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_265
timestamp 1698431365
transform 1 0 31024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_328
timestamp 1698431365
transform 1 0 38080 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_332
timestamp 1698431365
transform 1 0 38528 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_336
timestamp 1698431365
transform 1 0 38976 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_340
timestamp 1698431365
transform 1 0 39424 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_384
timestamp 1698431365
transform 1 0 44352 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_387
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_417
timestamp 1698431365
transform 1 0 48048 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_419
timestamp 1698431365
transform 1 0 48272 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_26
timestamp 1698431365
transform 1 0 4256 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_34
timestamp 1698431365
transform 1 0 5152 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_38
timestamp 1698431365
transform 1 0 5600 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_40
timestamp 1698431365
transform 1 0 5824 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_59
timestamp 1698431365
transform 1 0 7952 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_67
timestamp 1698431365
transform 1 0 8848 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_69
timestamp 1698431365
transform 1 0 9072 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_76
timestamp 1698431365
transform 1 0 9856 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_78
timestamp 1698431365
transform 1 0 10080 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_87
timestamp 1698431365
transform 1 0 11088 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_89
timestamp 1698431365
transform 1 0 11312 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_119
timestamp 1698431365
transform 1 0 14672 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_127
timestamp 1698431365
transform 1 0 15568 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_135
timestamp 1698431365
transform 1 0 16464 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_139
timestamp 1698431365
transform 1 0 16912 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_171
timestamp 1698431365
transform 1 0 20496 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_173
timestamp 1698431365
transform 1 0 20720 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_205
timestamp 1698431365
transform 1 0 24304 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_207
timestamp 1698431365
transform 1 0 24528 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_222
timestamp 1698431365
transform 1 0 26208 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_265
timestamp 1698431365
transform 1 0 31024 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_273
timestamp 1698431365
transform 1 0 31920 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_277
timestamp 1698431365
transform 1 0 32368 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_294
timestamp 1698431365
transform 1 0 34272 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_296
timestamp 1698431365
transform 1 0 34496 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_334
timestamp 1698431365
transform 1 0 38752 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_338
timestamp 1698431365
transform 1 0 39200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_10
timestamp 1698431365
transform 1 0 2464 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_14
timestamp 1698431365
transform 1 0 2912 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_16
timestamp 1698431365
transform 1 0 3136 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_25
timestamp 1698431365
transform 1 0 4144 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_29
timestamp 1698431365
transform 1 0 4592 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_33
timestamp 1698431365
transform 1 0 5040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_66
timestamp 1698431365
transform 1 0 8736 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_74
timestamp 1698431365
transform 1 0 9632 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_78
timestamp 1698431365
transform 1 0 10080 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_87
timestamp 1698431365
transform 1 0 11088 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_91
timestamp 1698431365
transform 1 0 11536 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_95
timestamp 1698431365
transform 1 0 11984 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_102
timestamp 1698431365
transform 1 0 12768 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_104
timestamp 1698431365
transform 1 0 12992 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_147
timestamp 1698431365
transform 1 0 17808 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_151
timestamp 1698431365
transform 1 0 18256 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_161
timestamp 1698431365
transform 1 0 19376 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_169
timestamp 1698431365
transform 1 0 20272 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_173
timestamp 1698431365
transform 1 0 20720 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_186
timestamp 1698431365
transform 1 0 22176 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_188
timestamp 1698431365
transform 1 0 22400 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_193
timestamp 1698431365
transform 1 0 22960 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_199
timestamp 1698431365
transform 1 0 23632 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_240
timestamp 1698431365
transform 1 0 28224 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_244
timestamp 1698431365
transform 1 0 28672 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_255
timestamp 1698431365
transform 1 0 29904 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_259
timestamp 1698431365
transform 1 0 30352 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_290
timestamp 1698431365
transform 1 0 33824 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_294
timestamp 1698431365
transform 1 0 34272 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_321
timestamp 1698431365
transform 1 0 37296 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_325
timestamp 1698431365
transform 1 0 37744 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_333
timestamp 1698431365
transform 1 0 38640 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_344
timestamp 1698431365
transform 1 0 39872 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_348
timestamp 1698431365
transform 1 0 40320 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_350
timestamp 1698431365
transform 1 0 40544 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_367
timestamp 1698431365
transform 1 0 42448 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_387
timestamp 1698431365
transform 1 0 44688 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_37
timestamp 1698431365
transform 1 0 5488 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_53
timestamp 1698431365
transform 1 0 7280 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_69
timestamp 1698431365
transform 1 0 9072 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_80
timestamp 1698431365
transform 1 0 10304 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_88
timestamp 1698431365
transform 1 0 11200 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_92
timestamp 1698431365
transform 1 0 11648 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_94
timestamp 1698431365
transform 1 0 11872 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_103
timestamp 1698431365
transform 1 0 12880 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_119
timestamp 1698431365
transform 1 0 14672 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_127
timestamp 1698431365
transform 1 0 15568 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_135
timestamp 1698431365
transform 1 0 16464 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_139
timestamp 1698431365
transform 1 0 16912 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_146
timestamp 1698431365
transform 1 0 17696 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_183
timestamp 1698431365
transform 1 0 21840 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_199
timestamp 1698431365
transform 1 0 23632 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_207
timestamp 1698431365
transform 1 0 24528 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_209
timestamp 1698431365
transform 1 0 24752 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_220
timestamp 1698431365
transform 1 0 25984 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_236
timestamp 1698431365
transform 1 0 27776 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_244
timestamp 1698431365
transform 1 0 28672 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_246
timestamp 1698431365
transform 1 0 28896 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_322
timestamp 1698431365
transform 1 0 37408 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_326
timestamp 1698431365
transform 1 0 37856 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_360
timestamp 1698431365
transform 1 0 41664 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_10
timestamp 1698431365
transform 1 0 2464 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_14
timestamp 1698431365
transform 1 0 2912 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_16
timestamp 1698431365
transform 1 0 3136 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_33
timestamp 1698431365
transform 1 0 5040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_47
timestamp 1698431365
transform 1 0 6608 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_51
timestamp 1698431365
transform 1 0 7056 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_89
timestamp 1698431365
transform 1 0 11312 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_103
timestamp 1698431365
transform 1 0 12880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_158
timestamp 1698431365
transform 1 0 19040 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_174
timestamp 1698431365
transform 1 0 20832 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_189
timestamp 1698431365
transform 1 0 22512 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_204
timestamp 1698431365
transform 1 0 24192 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_212
timestamp 1698431365
transform 1 0 25088 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_253
timestamp 1698431365
transform 1 0 29680 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_353
timestamp 1698431365
transform 1 0 40880 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_382
timestamp 1698431365
transform 1 0 44128 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_384
timestamp 1698431365
transform 1 0 44352 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_403
timestamp 1698431365
transform 1 0 46480 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_407
timestamp 1698431365
transform 1 0 46928 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_415
timestamp 1698431365
transform 1 0 47824 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_419
timestamp 1698431365
transform 1 0 48272 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_31
timestamp 1698431365
transform 1 0 4816 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_69
timestamp 1698431365
transform 1 0 9072 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_86
timestamp 1698431365
transform 1 0 10976 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_100
timestamp 1698431365
transform 1 0 12544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_104
timestamp 1698431365
transform 1 0 12992 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_150
timestamp 1698431365
transform 1 0 18144 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_220
timestamp 1698431365
transform 1 0 25984 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_230
timestamp 1698431365
transform 1 0 27104 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_238
timestamp 1698431365
transform 1 0 28000 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_242
timestamp 1698431365
transform 1 0 28448 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_244
timestamp 1698431365
transform 1 0 28672 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_249
timestamp 1698431365
transform 1 0 29232 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_257
timestamp 1698431365
transform 1 0 30128 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_262
timestamp 1698431365
transform 1 0 30688 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_272
timestamp 1698431365
transform 1 0 31808 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698431365
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_317
timestamp 1698431365
transform 1 0 36848 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_319
timestamp 1698431365
transform 1 0 37072 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_330
timestamp 1698431365
transform 1 0 38304 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_334
timestamp 1698431365
transform 1 0 38752 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_348
timestamp 1698431365
transform 1 0 40320 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_361
timestamp 1698431365
transform 1 0 41776 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_387
timestamp 1698431365
transform 1 0 44688 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_18
timestamp 1698431365
transform 1 0 3360 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_26
timestamp 1698431365
transform 1 0 4256 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_28
timestamp 1698431365
transform 1 0 4480 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_45
timestamp 1698431365
transform 1 0 6384 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_54
timestamp 1698431365
transform 1 0 7392 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_58
timestamp 1698431365
transform 1 0 7840 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_60
timestamp 1698431365
transform 1 0 8064 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_104
timestamp 1698431365
transform 1 0 12992 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_125
timestamp 1698431365
transform 1 0 15344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_129
timestamp 1698431365
transform 1 0 15792 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_135
timestamp 1698431365
transform 1 0 16464 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_143
timestamp 1698431365
transform 1 0 17360 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_171
timestamp 1698431365
transform 1 0 20496 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_185
timestamp 1698431365
transform 1 0 22064 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_187
timestamp 1698431365
transform 1 0 22288 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_208
timestamp 1698431365
transform 1 0 24640 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_212
timestamp 1698431365
transform 1 0 25088 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_214
timestamp 1698431365
transform 1 0 25312 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_231
timestamp 1698431365
transform 1 0 27216 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_239
timestamp 1698431365
transform 1 0 28112 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_243
timestamp 1698431365
transform 1 0 28560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_257
timestamp 1698431365
transform 1 0 30128 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_261
timestamp 1698431365
transform 1 0 30576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_263
timestamp 1698431365
transform 1 0 30800 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_302
timestamp 1698431365
transform 1 0 35168 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_310
timestamp 1698431365
transform 1 0 36064 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_314
timestamp 1698431365
transform 1 0 36512 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_325
timestamp 1698431365
transform 1 0 37744 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_331
timestamp 1698431365
transform 1 0 38416 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_333
timestamp 1698431365
transform 1 0 38640 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_336
timestamp 1698431365
transform 1 0 38976 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_352
timestamp 1698431365
transform 1 0 40768 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_387
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_389
timestamp 1698431365
transform 1 0 44912 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_404
timestamp 1698431365
transform 1 0 46592 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_39
timestamp 1698431365
transform 1 0 5712 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_43
timestamp 1698431365
transform 1 0 6160 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_53
timestamp 1698431365
transform 1 0 7280 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_57
timestamp 1698431365
transform 1 0 7728 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_65
timestamp 1698431365
transform 1 0 8624 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_69
timestamp 1698431365
transform 1 0 9072 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_76
timestamp 1698431365
transform 1 0 9856 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_82
timestamp 1698431365
transform 1 0 10528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_90
timestamp 1698431365
transform 1 0 11424 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_92
timestamp 1698431365
transform 1 0 11648 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_99
timestamp 1698431365
transform 1 0 12432 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_107
timestamp 1698431365
transform 1 0 13328 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_109
timestamp 1698431365
transform 1 0 13552 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_121
timestamp 1698431365
transform 1 0 14896 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_125
timestamp 1698431365
transform 1 0 15344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_129
timestamp 1698431365
transform 1 0 15792 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_137
timestamp 1698431365
transform 1 0 16688 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_139
timestamp 1698431365
transform 1 0 16912 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698431365
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_216
timestamp 1698431365
transform 1 0 25536 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_226
timestamp 1698431365
transform 1 0 26656 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_230
timestamp 1698431365
transform 1 0 27104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_286
timestamp 1698431365
transform 1 0 33376 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_290
timestamp 1698431365
transform 1 0 33824 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_296
timestamp 1698431365
transform 1 0 34496 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_333
timestamp 1698431365
transform 1 0 38640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_335
timestamp 1698431365
transform 1 0 38864 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_347
timestamp 1698431365
transform 1 0 40208 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_349
timestamp 1698431365
transform 1 0 40432 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_356
timestamp 1698431365
transform 1 0 41216 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_362
timestamp 1698431365
transform 1 0 41888 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_366
timestamp 1698431365
transform 1 0 42336 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_387
timestamp 1698431365
transform 1 0 44688 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_87
timestamp 1698431365
transform 1 0 11088 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_89
timestamp 1698431365
transform 1 0 11312 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_98
timestamp 1698431365
transform 1 0 12320 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_112
timestamp 1698431365
transform 1 0 13888 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_116
timestamp 1698431365
transform 1 0 14336 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_118
timestamp 1698431365
transform 1 0 14560 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_127
timestamp 1698431365
transform 1 0 15568 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_157
timestamp 1698431365
transform 1 0 18928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_159
timestamp 1698431365
transform 1 0 19152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698431365
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_206
timestamp 1698431365
transform 1 0 24416 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_265
timestamp 1698431365
transform 1 0 31024 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_297
timestamp 1698431365
transform 1 0 34608 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_306
timestamp 1698431365
transform 1 0 35616 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_360
timestamp 1698431365
transform 1 0 41664 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_384
timestamp 1698431365
transform 1 0 44352 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_387
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_389
timestamp 1698431365
transform 1 0 44912 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_405
timestamp 1698431365
transform 1 0 46704 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_409
timestamp 1698431365
transform 1 0 47152 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_417
timestamp 1698431365
transform 1 0 48048 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_419
timestamp 1698431365
transform 1 0 48272 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_31
timestamp 1698431365
transform 1 0 4816 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_86
timestamp 1698431365
transform 1 0 10976 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_95
timestamp 1698431365
transform 1 0 11984 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_103
timestamp 1698431365
transform 1 0 12880 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_107
timestamp 1698431365
transform 1 0 13328 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_137
timestamp 1698431365
transform 1 0 16688 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698431365
transform 1 0 16912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_150
timestamp 1698431365
transform 1 0 18144 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_158
timestamp 1698431365
transform 1 0 19040 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_179
timestamp 1698431365
transform 1 0 21392 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_181
timestamp 1698431365
transform 1 0 21616 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_190
timestamp 1698431365
transform 1 0 22624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_194
timestamp 1698431365
transform 1 0 23072 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_200
timestamp 1698431365
transform 1 0 23744 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_204
timestamp 1698431365
transform 1 0 24192 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_208
timestamp 1698431365
transform 1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_214
timestamp 1698431365
transform 1 0 25312 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_252
timestamp 1698431365
transform 1 0 29568 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_254
timestamp 1698431365
transform 1 0 29792 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_263
timestamp 1698431365
transform 1 0 30800 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_265
timestamp 1698431365
transform 1 0 31024 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_275
timestamp 1698431365
transform 1 0 32144 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698431365
transform 1 0 32592 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_312
timestamp 1698431365
transform 1 0 36288 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_316
timestamp 1698431365
transform 1 0 36736 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_335
timestamp 1698431365
transform 1 0 38864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_343
timestamp 1698431365
transform 1 0 39760 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_347
timestamp 1698431365
transform 1 0 40208 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_349
timestamp 1698431365
transform 1 0 40432 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_381
timestamp 1698431365
transform 1 0 44016 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_389
timestamp 1698431365
transform 1 0 44912 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_10
timestamp 1698431365
transform 1 0 2464 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_28
timestamp 1698431365
transform 1 0 4480 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_32
timestamp 1698431365
transform 1 0 4928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_41
timestamp 1698431365
transform 1 0 5936 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_48
timestamp 1698431365
transform 1 0 6720 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_64
timestamp 1698431365
transform 1 0 8512 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_66
timestamp 1698431365
transform 1 0 8736 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_83
timestamp 1698431365
transform 1 0 10640 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_89
timestamp 1698431365
transform 1 0 11312 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_128
timestamp 1698431365
transform 1 0 15680 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_144
timestamp 1698431365
transform 1 0 17472 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698431365
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_190
timestamp 1698431365
transform 1 0 22624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_192
timestamp 1698431365
transform 1 0 22848 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_209
timestamp 1698431365
transform 1 0 24752 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_211
timestamp 1698431365
transform 1 0 24976 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_298
timestamp 1698431365
transform 1 0 34720 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_302
timestamp 1698431365
transform 1 0 35168 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_311
timestamp 1698431365
transform 1 0 36176 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_352
timestamp 1698431365
transform 1 0 40768 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_10
timestamp 1698431365
transform 1 0 2464 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_14
timestamp 1698431365
transform 1 0 2912 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_38
timestamp 1698431365
transform 1 0 5600 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_40
timestamp 1698431365
transform 1 0 5824 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_80
timestamp 1698431365
transform 1 0 10304 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_88
timestamp 1698431365
transform 1 0 11200 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_126
timestamp 1698431365
transform 1 0 15456 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_135
timestamp 1698431365
transform 1 0 16464 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698431365
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_146
timestamp 1698431365
transform 1 0 17696 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_148
timestamp 1698431365
transform 1 0 17920 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_208
timestamp 1698431365
transform 1 0 24640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_224
timestamp 1698431365
transform 1 0 26432 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_230
timestamp 1698431365
transform 1 0 27104 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_260
timestamp 1698431365
transform 1 0 30464 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698431365
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_338
timestamp 1698431365
transform 1 0 39200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698431365
transform 1 0 40096 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_361
timestamp 1698431365
transform 1 0 41776 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_363
timestamp 1698431365
transform 1 0 42000 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_366
timestamp 1698431365
transform 1 0 42336 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_31
timestamp 1698431365
transform 1 0 4816 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_43
timestamp 1698431365
transform 1 0 6160 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_47
timestamp 1698431365
transform 1 0 6608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_49
timestamp 1698431365
transform 1 0 6832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_52
timestamp 1698431365
transform 1 0 7168 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_60
timestamp 1698431365
transform 1 0 8064 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_64
timestamp 1698431365
transform 1 0 8512 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_72
timestamp 1698431365
transform 1 0 9408 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_103
timestamp 1698431365
transform 1 0 12880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_111
timestamp 1698431365
transform 1 0 13776 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_148
timestamp 1698431365
transform 1 0 17920 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_168
timestamp 1698431365
transform 1 0 20160 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_172
timestamp 1698431365
transform 1 0 20608 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_185
timestamp 1698431365
transform 1 0 22064 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_199
timestamp 1698431365
transform 1 0 23632 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_203
timestamp 1698431365
transform 1 0 24080 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_207
timestamp 1698431365
transform 1 0 24528 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_209
timestamp 1698431365
transform 1 0 24752 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_212
timestamp 1698431365
transform 1 0 25088 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_236
timestamp 1698431365
transform 1 0 27776 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_306
timestamp 1698431365
transform 1 0 35616 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_308
timestamp 1698431365
transform 1 0 35840 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_371
timestamp 1698431365
transform 1 0 42896 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_373
timestamp 1698431365
transform 1 0 43120 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_384
timestamp 1698431365
transform 1 0 44352 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_387
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_389
timestamp 1698431365
transform 1 0 44912 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_407
timestamp 1698431365
transform 1 0 46928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_411
timestamp 1698431365
transform 1 0 47376 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_413
timestamp 1698431365
transform 1 0 47600 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_10
timestamp 1698431365
transform 1 0 2464 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_14
timestamp 1698431365
transform 1 0 2912 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_31
timestamp 1698431365
transform 1 0 4816 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_33
timestamp 1698431365
transform 1 0 5040 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_63
timestamp 1698431365
transform 1 0 8400 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_67
timestamp 1698431365
transform 1 0 8848 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_69
timestamp 1698431365
transform 1 0 9072 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_80
timestamp 1698431365
transform 1 0 10304 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_117
timestamp 1698431365
transform 1 0 14448 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_125
timestamp 1698431365
transform 1 0 15344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_135
timestamp 1698431365
transform 1 0 16464 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_137
timestamp 1698431365
transform 1 0 16688 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_173
timestamp 1698431365
transform 1 0 20720 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_180
timestamp 1698431365
transform 1 0 21504 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_188
timestamp 1698431365
transform 1 0 22400 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_205
timestamp 1698431365
transform 1 0 24304 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698431365
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_274
timestamp 1698431365
transform 1 0 32032 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_278
timestamp 1698431365
transform 1 0 32480 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_286
timestamp 1698431365
transform 1 0 33376 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_310
timestamp 1698431365
transform 1 0 36064 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_410
timestamp 1698431365
transform 1 0 47264 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_415
timestamp 1698431365
transform 1 0 47824 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_419
timestamp 1698431365
transform 1 0 48272 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_31
timestamp 1698431365
transform 1 0 4816 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_43
timestamp 1698431365
transform 1 0 6160 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_58
timestamp 1698431365
transform 1 0 7840 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_89
timestamp 1698431365
transform 1 0 11312 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_113
timestamp 1698431365
transform 1 0 14000 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_117
timestamp 1698431365
transform 1 0 14448 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_132
timestamp 1698431365
transform 1 0 16128 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_136
timestamp 1698431365
transform 1 0 16576 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_140
timestamp 1698431365
transform 1 0 17024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_207
timestamp 1698431365
transform 1 0 24528 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_238
timestamp 1698431365
transform 1 0 28000 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_242
timestamp 1698431365
transform 1 0 28448 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698431365
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_251
timestamp 1698431365
transform 1 0 29456 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_267
timestamp 1698431365
transform 1 0 31248 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_309
timestamp 1698431365
transform 1 0 35952 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698431365
transform 1 0 36512 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_10
timestamp 1698431365
transform 1 0 2464 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_14
timestamp 1698431365
transform 1 0 2912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_69
timestamp 1698431365
transform 1 0 9072 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_192
timestamp 1698431365
transform 1 0 22848 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_196
timestamp 1698431365
transform 1 0 23296 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_203
timestamp 1698431365
transform 1 0 24080 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_207
timestamp 1698431365
transform 1 0 24528 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698431365
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_214
timestamp 1698431365
transform 1 0 25312 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_221
timestamp 1698431365
transform 1 0 26096 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_225
timestamp 1698431365
transform 1 0 26544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_229
timestamp 1698431365
transform 1 0 26992 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_237
timestamp 1698431365
transform 1 0 27888 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_243
timestamp 1698431365
transform 1 0 28560 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_253
timestamp 1698431365
transform 1 0 29680 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_257
timestamp 1698431365
transform 1 0 30128 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_261
timestamp 1698431365
transform 1 0 30576 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_275
timestamp 1698431365
transform 1 0 32144 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_292
timestamp 1698431365
transform 1 0 34048 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_296
timestamp 1698431365
transform 1 0 34496 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_298
timestamp 1698431365
transform 1 0 34720 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_301
timestamp 1698431365
transform 1 0 35056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_305
timestamp 1698431365
transform 1 0 35504 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_307
timestamp 1698431365
transform 1 0 35728 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_341
timestamp 1698431365
transform 1 0 39536 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_343
timestamp 1698431365
transform 1 0 39760 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_369
timestamp 1698431365
transform 1 0 42672 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_31
timestamp 1698431365
transform 1 0 4816 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_66
timestamp 1698431365
transform 1 0 8736 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_70
timestamp 1698431365
transform 1 0 9184 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_72
timestamp 1698431365
transform 1 0 9408 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_79
timestamp 1698431365
transform 1 0 10192 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_88
timestamp 1698431365
transform 1 0 11200 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_92
timestamp 1698431365
transform 1 0 11648 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_100
timestamp 1698431365
transform 1 0 12544 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_104
timestamp 1698431365
transform 1 0 12992 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_111
timestamp 1698431365
transform 1 0 13776 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_113
timestamp 1698431365
transform 1 0 14000 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_169
timestamp 1698431365
transform 1 0 20272 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_186
timestamp 1698431365
transform 1 0 22176 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_188
timestamp 1698431365
transform 1 0 22400 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_239
timestamp 1698431365
transform 1 0 28112 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_243
timestamp 1698431365
transform 1 0 28560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_249
timestamp 1698431365
transform 1 0 29232 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_260
timestamp 1698431365
transform 1 0 30464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_264
timestamp 1698431365
transform 1 0 30912 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_268
timestamp 1698431365
transform 1 0 31360 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_272
timestamp 1698431365
transform 1 0 31808 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_276
timestamp 1698431365
transform 1 0 32256 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_284
timestamp 1698431365
transform 1 0 33152 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_288
timestamp 1698431365
transform 1 0 33600 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_292
timestamp 1698431365
transform 1 0 34048 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_300
timestamp 1698431365
transform 1 0 34944 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_304
timestamp 1698431365
transform 1 0 35392 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_307
timestamp 1698431365
transform 1 0 35728 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698431365
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_321
timestamp 1698431365
transform 1 0 37296 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_373
timestamp 1698431365
transform 1 0 43120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_387
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_10
timestamp 1698431365
transform 1 0 2464 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_14
timestamp 1698431365
transform 1 0 2912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_36
timestamp 1698431365
transform 1 0 5376 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_38
timestamp 1698431365
transform 1 0 5600 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_52
timestamp 1698431365
transform 1 0 7168 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698431365
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_76
timestamp 1698431365
transform 1 0 9856 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_80
timestamp 1698431365
transform 1 0 10304 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_131
timestamp 1698431365
transform 1 0 16016 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_192
timestamp 1698431365
transform 1 0 22848 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698431365
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_249
timestamp 1698431365
transform 1 0 29232 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_253
timestamp 1698431365
transform 1 0 29680 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_255
timestamp 1698431365
transform 1 0 29904 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_288
timestamp 1698431365
transform 1 0 33600 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_303
timestamp 1698431365
transform 1 0 35280 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_339
timestamp 1698431365
transform 1 0 39312 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_347
timestamp 1698431365
transform 1 0 40208 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_349
timestamp 1698431365
transform 1 0 40432 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_356
timestamp 1698431365
transform 1 0 41216 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_374
timestamp 1698431365
transform 1 0 43232 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_382
timestamp 1698431365
transform 1 0 44128 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_419
timestamp 1698431365
transform 1 0 48272 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_31
timestamp 1698431365
transform 1 0 4816 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_47
timestamp 1698431365
transform 1 0 6608 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_51
timestamp 1698431365
transform 1 0 7056 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_87
timestamp 1698431365
transform 1 0 11088 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_103
timestamp 1698431365
transform 1 0 12880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_115
timestamp 1698431365
transform 1 0 14224 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_124
timestamp 1698431365
transform 1 0 15232 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_130
timestamp 1698431365
transform 1 0 15904 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_134
timestamp 1698431365
transform 1 0 16352 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_188
timestamp 1698431365
transform 1 0 22400 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_228
timestamp 1698431365
transform 1 0 26880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_230
timestamp 1698431365
transform 1 0 27104 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_239
timestamp 1698431365
transform 1 0 28112 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_243
timestamp 1698431365
transform 1 0 28560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_312
timestamp 1698431365
transform 1 0 36288 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_314
timestamp 1698431365
transform 1 0 36512 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_352
timestamp 1698431365
transform 1 0 40768 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_387
timestamp 1698431365
transform 1 0 44688 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_10
timestamp 1698431365
transform 1 0 2464 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_14
timestamp 1698431365
transform 1 0 2912 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_44
timestamp 1698431365
transform 1 0 6272 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_51
timestamp 1698431365
transform 1 0 7056 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_59
timestamp 1698431365
transform 1 0 7952 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698431365
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_104
timestamp 1698431365
transform 1 0 12992 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_134
timestamp 1698431365
transform 1 0 16352 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_150
timestamp 1698431365
transform 1 0 18144 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_152
timestamp 1698431365
transform 1 0 18368 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_197
timestamp 1698431365
transform 1 0 23408 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_199
timestamp 1698431365
transform 1 0 23632 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_220
timestamp 1698431365
transform 1 0 25984 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_227
timestamp 1698431365
transform 1 0 26768 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_229
timestamp 1698431365
transform 1 0 26992 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698431365
transform 1 0 32368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698431365
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_324
timestamp 1698431365
transform 1 0 37632 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_328
timestamp 1698431365
transform 1 0 38080 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_342
timestamp 1698431365
transform 1 0 39648 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_352
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_372
timestamp 1698431365
transform 1 0 43008 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_380
timestamp 1698431365
transform 1 0 43904 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_404
timestamp 1698431365
transform 1 0 46592 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_18
timestamp 1698431365
transform 1 0 3360 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_22
timestamp 1698431365
transform 1 0 3808 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_29
timestamp 1698431365
transform 1 0 4592 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_33
timestamp 1698431365
transform 1 0 5040 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_43
timestamp 1698431365
transform 1 0 6160 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_59
timestamp 1698431365
transform 1 0 7952 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_70
timestamp 1698431365
transform 1 0 9184 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_74
timestamp 1698431365
transform 1 0 9632 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_136
timestamp 1698431365
transform 1 0 16576 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_187
timestamp 1698431365
transform 1 0 22288 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_198
timestamp 1698431365
transform 1 0 23520 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_256
timestamp 1698431365
transform 1 0 30016 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_319
timestamp 1698431365
transform 1 0 37072 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_332
timestamp 1698431365
transform 1 0 38528 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_336
timestamp 1698431365
transform 1 0 38976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_346
timestamp 1698431365
transform 1 0 40096 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_365
timestamp 1698431365
transform 1 0 42224 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_387
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_39
timestamp 1698431365
transform 1 0 5712 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_46
timestamp 1698431365
transform 1 0 6496 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_50
timestamp 1698431365
transform 1 0 6944 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698431365
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_74
timestamp 1698431365
transform 1 0 9632 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_101
timestamp 1698431365
transform 1 0 12656 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_133
timestamp 1698431365
transform 1 0 16240 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_171
timestamp 1698431365
transform 1 0 20496 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_201
timestamp 1698431365
transform 1 0 23856 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_203
timestamp 1698431365
transform 1 0 24080 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698431365
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_274
timestamp 1698431365
transform 1 0 32032 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_348
timestamp 1698431365
transform 1 0 40320 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_352
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_360
timestamp 1698431365
transform 1 0 41664 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_364
timestamp 1698431365
transform 1 0 42112 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_370
timestamp 1698431365
transform 1 0 42784 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_375
timestamp 1698431365
transform 1 0 43344 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_379
timestamp 1698431365
transform 1 0 43792 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_402
timestamp 1698431365
transform 1 0 46368 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_418
timestamp 1698431365
transform 1 0 48160 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_10
timestamp 1698431365
transform 1 0 2464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698431365
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_43
timestamp 1698431365
transform 1 0 6160 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_70
timestamp 1698431365
transform 1 0 9184 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_84
timestamp 1698431365
transform 1 0 10752 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_91
timestamp 1698431365
transform 1 0 11536 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_99
timestamp 1698431365
transform 1 0 12432 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_103
timestamp 1698431365
transform 1 0 12880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_138
timestamp 1698431365
transform 1 0 16800 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_227
timestamp 1698431365
transform 1 0 26768 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_240
timestamp 1698431365
transform 1 0 28224 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698431365
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_251
timestamp 1698431365
transform 1 0 29456 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_292
timestamp 1698431365
transform 1 0 34048 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_308
timestamp 1698431365
transform 1 0 35840 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_312
timestamp 1698431365
transform 1 0 36288 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_339
timestamp 1698431365
transform 1 0 39312 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_348
timestamp 1698431365
transform 1 0 40320 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_350
timestamp 1698431365
transform 1 0 40544 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_359
timestamp 1698431365
transform 1 0 41552 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_361
timestamp 1698431365
transform 1 0 41776 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_375
timestamp 1698431365
transform 1 0 43344 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_39
timestamp 1698431365
transform 1 0 5712 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_46
timestamp 1698431365
transform 1 0 6496 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_50
timestamp 1698431365
transform 1 0 6944 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_67
timestamp 1698431365
transform 1 0 8848 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_69
timestamp 1698431365
transform 1 0 9072 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_87
timestamp 1698431365
transform 1 0 11088 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_95
timestamp 1698431365
transform 1 0 11984 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_99
timestamp 1698431365
transform 1 0 12432 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_101
timestamp 1698431365
transform 1 0 12656 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_146
timestamp 1698431365
transform 1 0 17696 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_148
timestamp 1698431365
transform 1 0 17920 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_222
timestamp 1698431365
transform 1 0 26208 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_255
timestamp 1698431365
transform 1 0 29904 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_271
timestamp 1698431365
transform 1 0 31696 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698431365
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_284
timestamp 1698431365
transform 1 0 33152 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_294
timestamp 1698431365
transform 1 0 34272 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_298
timestamp 1698431365
transform 1 0 34720 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698431365
transform 1 0 36512 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698431365
transform 1 0 37408 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_344
timestamp 1698431365
transform 1 0 39872 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_348
timestamp 1698431365
transform 1 0 40320 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_395
timestamp 1698431365
transform 1 0 45584 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_399
timestamp 1698431365
transform 1 0 46032 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_401
timestamp 1698431365
transform 1 0 46256 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_419
timestamp 1698431365
transform 1 0 48272 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_31
timestamp 1698431365
transform 1 0 4816 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_99
timestamp 1698431365
transform 1 0 12432 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_103
timestamp 1698431365
transform 1 0 12880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_111
timestamp 1698431365
transform 1 0 13776 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_113
timestamp 1698431365
transform 1 0 14000 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_122
timestamp 1698431365
transform 1 0 15008 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_126
timestamp 1698431365
transform 1 0 15456 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_128
timestamp 1698431365
transform 1 0 15680 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_158
timestamp 1698431365
transform 1 0 19040 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_168
timestamp 1698431365
transform 1 0 20160 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_172
timestamp 1698431365
transform 1 0 20608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698431365
transform 1 0 20832 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_212
timestamp 1698431365
transform 1 0 25088 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_214
timestamp 1698431365
transform 1 0 25312 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_230
timestamp 1698431365
transform 1 0 27104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_234
timestamp 1698431365
transform 1 0 27552 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698431365
transform 1 0 28448 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698431365
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_251
timestamp 1698431365
transform 1 0 29456 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_261
timestamp 1698431365
transform 1 0 30576 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_265
timestamp 1698431365
transform 1 0 31024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_271
timestamp 1698431365
transform 1 0 31696 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_275
timestamp 1698431365
transform 1 0 32144 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_287
timestamp 1698431365
transform 1 0 33488 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_298
timestamp 1698431365
transform 1 0 34720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_302
timestamp 1698431365
transform 1 0 35168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_306
timestamp 1698431365
transform 1 0 35616 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_314
timestamp 1698431365
transform 1 0 36512 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_335
timestamp 1698431365
transform 1 0 38864 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_359
timestamp 1698431365
transform 1 0 41552 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_361
timestamp 1698431365
transform 1 0 41776 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_382
timestamp 1698431365
transform 1 0 44128 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_384
timestamp 1698431365
transform 1 0 44352 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_387
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_389
timestamp 1698431365
transform 1 0 44912 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_419
timestamp 1698431365
transform 1 0 48272 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_10
timestamp 1698431365
transform 1 0 2464 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_14
timestamp 1698431365
transform 1 0 2912 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_16
timestamp 1698431365
transform 1 0 3136 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_67
timestamp 1698431365
transform 1 0 8848 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_69
timestamp 1698431365
transform 1 0 9072 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_76
timestamp 1698431365
transform 1 0 9856 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_113
timestamp 1698431365
transform 1 0 14000 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_135
timestamp 1698431365
transform 1 0 16464 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_139
timestamp 1698431365
transform 1 0 16912 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_146
timestamp 1698431365
transform 1 0 17696 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_150
timestamp 1698431365
transform 1 0 18144 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_152
timestamp 1698431365
transform 1 0 18368 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_185
timestamp 1698431365
transform 1 0 22064 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_187
timestamp 1698431365
transform 1 0 22288 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_195
timestamp 1698431365
transform 1 0 23184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_199
timestamp 1698431365
transform 1 0 23632 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_203
timestamp 1698431365
transform 1 0 24080 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698431365
transform 1 0 24416 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_216
timestamp 1698431365
transform 1 0 25536 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_220
timestamp 1698431365
transform 1 0 25984 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_228
timestamp 1698431365
transform 1 0 26880 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_243
timestamp 1698431365
transform 1 0 28560 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_259
timestamp 1698431365
transform 1 0 30352 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_278
timestamp 1698431365
transform 1 0 32480 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_345
timestamp 1698431365
transform 1 0 39984 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_352
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_362
timestamp 1698431365
transform 1 0 41888 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_369
timestamp 1698431365
transform 1 0 42672 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_10
timestamp 1698431365
transform 1 0 2464 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_71
timestamp 1698431365
transform 1 0 9296 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_79
timestamp 1698431365
transform 1 0 10192 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_83
timestamp 1698431365
transform 1 0 10640 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_86
timestamp 1698431365
transform 1 0 10976 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_90
timestamp 1698431365
transform 1 0 11424 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_157
timestamp 1698431365
transform 1 0 18928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_170
timestamp 1698431365
transform 1 0 20384 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698431365
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_223
timestamp 1698431365
transform 1 0 26320 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_238
timestamp 1698431365
transform 1 0 28000 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_240
timestamp 1698431365
transform 1 0 28224 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_304
timestamp 1698431365
transform 1 0 35392 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_306
timestamp 1698431365
transform 1 0 35616 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_367
timestamp 1698431365
transform 1 0 42448 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_376
timestamp 1698431365
transform 1 0 43456 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_380
timestamp 1698431365
transform 1 0 43904 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_384
timestamp 1698431365
transform 1 0 44352 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_401
timestamp 1698431365
transform 1 0 46256 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_409
timestamp 1698431365
transform 1 0 47152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_136
timestamp 1698431365
transform 1 0 16576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_160
timestamp 1698431365
transform 1 0 19264 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_197
timestamp 1698431365
transform 1 0 23408 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_199
timestamp 1698431365
transform 1 0 23632 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_208
timestamp 1698431365
transform 1 0 24640 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_263
timestamp 1698431365
transform 1 0 30800 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_267
timestamp 1698431365
transform 1 0 31248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_269
timestamp 1698431365
transform 1 0 31472 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_278
timestamp 1698431365
transform 1 0 32480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_284
timestamp 1698431365
transform 1 0 33152 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_323
timestamp 1698431365
transform 1 0 37520 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_327
timestamp 1698431365
transform 1 0 37968 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_362
timestamp 1698431365
transform 1 0 41888 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_366
timestamp 1698431365
transform 1 0 42336 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_384
timestamp 1698431365
transform 1 0 44352 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_388
timestamp 1698431365
transform 1 0 44800 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_390
timestamp 1698431365
transform 1 0 45024 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_31
timestamp 1698431365
transform 1 0 4816 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_60
timestamp 1698431365
transform 1 0 8064 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_66
timestamp 1698431365
transform 1 0 8736 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_72
timestamp 1698431365
transform 1 0 9408 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_88
timestamp 1698431365
transform 1 0 11200 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_91
timestamp 1698431365
transform 1 0 11536 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_99
timestamp 1698431365
transform 1 0 12432 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_123
timestamp 1698431365
transform 1 0 15120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_181
timestamp 1698431365
transform 1 0 21616 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_191
timestamp 1698431365
transform 1 0 22736 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_195
timestamp 1698431365
transform 1 0 23184 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_205
timestamp 1698431365
transform 1 0 24304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_209
timestamp 1698431365
transform 1 0 24752 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_242
timestamp 1698431365
transform 1 0 28448 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_244
timestamp 1698431365
transform 1 0 28672 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_255
timestamp 1698431365
transform 1 0 29904 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_279
timestamp 1698431365
transform 1 0 32592 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_281
timestamp 1698431365
transform 1 0 32816 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_306
timestamp 1698431365
transform 1 0 35616 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_310
timestamp 1698431365
transform 1 0 36064 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_312
timestamp 1698431365
transform 1 0 36288 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_367
timestamp 1698431365
transform 1 0 42448 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_375
timestamp 1698431365
transform 1 0 43344 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_378
timestamp 1698431365
transform 1 0 43680 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_382
timestamp 1698431365
transform 1 0 44128 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_384
timestamp 1698431365
transform 1 0 44352 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_387
timestamp 1698431365
transform 1 0 44688 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_18
timestamp 1698431365
transform 1 0 3360 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_48
timestamp 1698431365
transform 1 0 6720 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_55
timestamp 1698431365
transform 1 0 7504 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_69
timestamp 1698431365
transform 1 0 9072 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_80
timestamp 1698431365
transform 1 0 10304 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_82
timestamp 1698431365
transform 1 0 10528 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_89
timestamp 1698431365
transform 1 0 11312 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_98
timestamp 1698431365
transform 1 0 12320 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_102
timestamp 1698431365
transform 1 0 12768 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_110
timestamp 1698431365
transform 1 0 13664 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_116
timestamp 1698431365
transform 1 0 14336 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_130
timestamp 1698431365
transform 1 0 15904 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_175
timestamp 1698431365
transform 1 0 20944 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_197
timestamp 1698431365
transform 1 0 23408 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_206
timestamp 1698431365
transform 1 0 24416 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_214
timestamp 1698431365
transform 1 0 25312 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_237
timestamp 1698431365
transform 1 0 27888 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_278
timestamp 1698431365
transform 1 0 32480 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_288
timestamp 1698431365
transform 1 0 33600 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_292
timestamp 1698431365
transform 1 0 34048 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_317
timestamp 1698431365
transform 1 0 36848 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_319
timestamp 1698431365
transform 1 0 37072 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_349
timestamp 1698431365
transform 1 0 40432 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_365
timestamp 1698431365
transform 1 0 42224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_387
timestamp 1698431365
transform 1 0 44688 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_418
timestamp 1698431365
transform 1 0 48160 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_31
timestamp 1698431365
transform 1 0 4816 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_53
timestamp 1698431365
transform 1 0 7280 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_55
timestamp 1698431365
transform 1 0 7504 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_85
timestamp 1698431365
transform 1 0 10864 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_89
timestamp 1698431365
transform 1 0 11312 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_91
timestamp 1698431365
transform 1 0 11536 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_96
timestamp 1698431365
transform 1 0 12096 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_104
timestamp 1698431365
transform 1 0 12992 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_116
timestamp 1698431365
transform 1 0 14336 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_183
timestamp 1698431365
transform 1 0 21840 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_213
timestamp 1698431365
transform 1 0 25200 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_239
timestamp 1698431365
transform 1 0 28112 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_243
timestamp 1698431365
transform 1 0 28560 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_276
timestamp 1698431365
transform 1 0 32256 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_294
timestamp 1698431365
transform 1 0 34272 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_296
timestamp 1698431365
transform 1 0 34496 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_299
timestamp 1698431365
transform 1 0 34832 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_303
timestamp 1698431365
transform 1 0 35280 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_307
timestamp 1698431365
transform 1 0 35728 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_311
timestamp 1698431365
transform 1 0 36176 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_338
timestamp 1698431365
transform 1 0 39200 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_368
timestamp 1698431365
transform 1 0 42560 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_370
timestamp 1698431365
transform 1 0 42784 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_375
timestamp 1698431365
transform 1 0 43344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_377
timestamp 1698431365
transform 1 0 43568 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_380
timestamp 1698431365
transform 1 0 43904 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_382
timestamp 1698431365
transform 1 0 44128 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_409
timestamp 1698431365
transform 1 0 47152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_418
timestamp 1698431365
transform 1 0 48160 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_10
timestamp 1698431365
transform 1 0 2464 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_69
timestamp 1698431365
transform 1 0 9072 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_76
timestamp 1698431365
transform 1 0 9856 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_78
timestamp 1698431365
transform 1 0 10080 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_108
timestamp 1698431365
transform 1 0 13440 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_110
timestamp 1698431365
transform 1 0 13664 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_128
timestamp 1698431365
transform 1 0 15680 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_132
timestamp 1698431365
transform 1 0 16128 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_136
timestamp 1698431365
transform 1 0 16576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_146
timestamp 1698431365
transform 1 0 17696 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_252
timestamp 1698431365
transform 1 0 29568 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_256
timestamp 1698431365
transform 1 0 30016 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_260
timestamp 1698431365
transform 1 0 30464 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698431365
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_301
timestamp 1698431365
transform 1 0 35056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_311
timestamp 1698431365
transform 1 0 36176 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_349
timestamp 1698431365
transform 1 0 40432 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_45
timestamp 1698431365
transform 1 0 6384 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_47
timestamp 1698431365
transform 1 0 6608 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_53
timestamp 1698431365
transform 1 0 7280 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_83
timestamp 1698431365
transform 1 0 10640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_85
timestamp 1698431365
transform 1 0 10864 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_90
timestamp 1698431365
transform 1 0 11424 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_98
timestamp 1698431365
transform 1 0 12320 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_102
timestamp 1698431365
transform 1 0 12768 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_104
timestamp 1698431365
transform 1 0 12992 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_137
timestamp 1698431365
transform 1 0 16688 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_141
timestamp 1698431365
transform 1 0 17136 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_172
timestamp 1698431365
transform 1 0 20608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_174
timestamp 1698431365
transform 1 0 20832 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_183
timestamp 1698431365
transform 1 0 21840 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_185
timestamp 1698431365
transform 1 0 22064 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_202
timestamp 1698431365
transform 1 0 23968 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_215
timestamp 1698431365
transform 1 0 25424 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_217
timestamp 1698431365
transform 1 0 25648 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_224
timestamp 1698431365
transform 1 0 26432 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_241
timestamp 1698431365
transform 1 0 28336 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_256
timestamp 1698431365
transform 1 0 30016 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_260
timestamp 1698431365
transform 1 0 30464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_264
timestamp 1698431365
transform 1 0 30912 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_268
timestamp 1698431365
transform 1 0 31360 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_278
timestamp 1698431365
transform 1 0 32480 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_311
timestamp 1698431365
transform 1 0 36176 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_319
timestamp 1698431365
transform 1 0 37072 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_350
timestamp 1698431365
transform 1 0 40544 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_387
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_31
timestamp 1698431365
transform 1 0 4816 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_62
timestamp 1698431365
transform 1 0 8288 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_112
timestamp 1698431365
transform 1 0 13888 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_120
timestamp 1698431365
transform 1 0 14784 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_124
timestamp 1698431365
transform 1 0 15232 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_130
timestamp 1698431365
transform 1 0 15904 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_132
timestamp 1698431365
transform 1 0 16128 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_137
timestamp 1698431365
transform 1 0 16688 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_139
timestamp 1698431365
transform 1 0 16912 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_146
timestamp 1698431365
transform 1 0 17696 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_165
timestamp 1698431365
transform 1 0 19824 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_169
timestamp 1698431365
transform 1 0 20272 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_207
timestamp 1698431365
transform 1 0 24528 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_209
timestamp 1698431365
transform 1 0 24752 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_320
timestamp 1698431365
transform 1 0 37184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_324
timestamp 1698431365
transform 1 0 37632 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_334
timestamp 1698431365
transform 1 0 38752 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_340
timestamp 1698431365
transform 1 0 39424 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_358
timestamp 1698431365
transform 1 0 41440 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_4
timestamp 1698431365
transform 1 0 1792 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_21
timestamp 1698431365
transform 1 0 3696 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_32
timestamp 1698431365
transform 1 0 4928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_43
timestamp 1698431365
transform 1 0 6160 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_81
timestamp 1698431365
transform 1 0 10416 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_85
timestamp 1698431365
transform 1 0 10864 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_116
timestamp 1698431365
transform 1 0 14336 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_120
timestamp 1698431365
transform 1 0 14784 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_163
timestamp 1698431365
transform 1 0 19600 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_167
timestamp 1698431365
transform 1 0 20048 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_171
timestamp 1698431365
transform 1 0 20496 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_181
timestamp 1698431365
transform 1 0 21616 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_189
timestamp 1698431365
transform 1 0 22512 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_193
timestamp 1698431365
transform 1 0 22960 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_202
timestamp 1698431365
transform 1 0 23968 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_214
timestamp 1698431365
transform 1 0 25312 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_220
timestamp 1698431365
transform 1 0 25984 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_222
timestamp 1698431365
transform 1 0 26208 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_225
timestamp 1698431365
transform 1 0 26544 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_231
timestamp 1698431365
transform 1 0 27216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_235
timestamp 1698431365
transform 1 0 27664 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_239
timestamp 1698431365
transform 1 0 28112 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_243
timestamp 1698431365
transform 1 0 28560 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_302
timestamp 1698431365
transform 1 0 35168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_306
timestamp 1698431365
transform 1 0 35616 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_308
timestamp 1698431365
transform 1 0 35840 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_333
timestamp 1698431365
transform 1 0 38640 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_337
timestamp 1698431365
transform 1 0 39088 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_381
timestamp 1698431365
transform 1 0 44016 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_387
timestamp 1698431365
transform 1 0 44688 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_10
timestamp 1698431365
transform 1 0 2464 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_14
timestamp 1698431365
transform 1 0 2912 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_34
timestamp 1698431365
transform 1 0 5152 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_42
timestamp 1698431365
transform 1 0 6048 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_56
timestamp 1698431365
transform 1 0 7616 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_80
timestamp 1698431365
transform 1 0 10304 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_113
timestamp 1698431365
transform 1 0 14000 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_129
timestamp 1698431365
transform 1 0 15792 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_137
timestamp 1698431365
transform 1 0 16688 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_139
timestamp 1698431365
transform 1 0 16912 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_152
timestamp 1698431365
transform 1 0 18368 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_187
timestamp 1698431365
transform 1 0 22288 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_196
timestamp 1698431365
transform 1 0 23296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_223
timestamp 1698431365
transform 1 0 26320 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_242
timestamp 1698431365
transform 1 0 28448 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_246
timestamp 1698431365
transform 1 0 28896 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_250
timestamp 1698431365
transform 1 0 29344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_277
timestamp 1698431365
transform 1 0 32368 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_279
timestamp 1698431365
transform 1 0 32592 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_288
timestamp 1698431365
transform 1 0 33600 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_294
timestamp 1698431365
transform 1 0 34272 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_298
timestamp 1698431365
transform 1 0 34720 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_306
timestamp 1698431365
transform 1 0 35616 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_346
timestamp 1698431365
transform 1 0 40096 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_356
timestamp 1698431365
transform 1 0 41216 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_358
timestamp 1698431365
transform 1 0 41440 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_394
timestamp 1698431365
transform 1 0 45472 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_31
timestamp 1698431365
transform 1 0 4816 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_41
timestamp 1698431365
transform 1 0 5936 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_45
timestamp 1698431365
transform 1 0 6384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_47
timestamp 1698431365
transform 1 0 6608 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_98
timestamp 1698431365
transform 1 0 12320 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_102
timestamp 1698431365
transform 1 0 12768 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_104
timestamp 1698431365
transform 1 0 12992 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_111
timestamp 1698431365
transform 1 0 13776 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_142
timestamp 1698431365
transform 1 0 17248 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_144
timestamp 1698431365
transform 1 0 17472 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_168
timestamp 1698431365
transform 1 0 20160 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_257
timestamp 1698431365
transform 1 0 30128 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_268
timestamp 1698431365
transform 1 0 31360 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_270
timestamp 1698431365
transform 1 0 31584 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_300
timestamp 1698431365
transform 1 0 34944 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_308
timestamp 1698431365
transform 1 0 35840 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_312
timestamp 1698431365
transform 1 0 36288 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_333
timestamp 1698431365
transform 1 0 38640 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_341
timestamp 1698431365
transform 1 0 39536 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_359
timestamp 1698431365
transform 1 0 41552 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_363
timestamp 1698431365
transform 1 0 42000 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_366
timestamp 1698431365
transform 1 0 42336 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_10
timestamp 1698431365
transform 1 0 2464 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_12
timestamp 1698431365
transform 1 0 2688 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_21
timestamp 1698431365
transform 1 0 3696 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_29
timestamp 1698431365
transform 1 0 4592 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_68
timestamp 1698431365
transform 1 0 8960 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_103
timestamp 1698431365
transform 1 0 12880 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_125
timestamp 1698431365
transform 1 0 15344 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_133
timestamp 1698431365
transform 1 0 16240 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_136
timestamp 1698431365
transform 1 0 16576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_195
timestamp 1698431365
transform 1 0 23184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_204
timestamp 1698431365
transform 1 0 24192 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_214
timestamp 1698431365
transform 1 0 25312 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_245
timestamp 1698431365
transform 1 0 28784 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698431365
transform 1 0 32256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_304
timestamp 1698431365
transform 1 0 35392 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_308
timestamp 1698431365
transform 1 0 35840 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_312
timestamp 1698431365
transform 1 0 36288 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_316
timestamp 1698431365
transform 1 0 36736 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_347
timestamp 1698431365
transform 1 0 40208 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_349
timestamp 1698431365
transform 1 0 40432 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_358
timestamp 1698431365
transform 1 0 41440 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_397
timestamp 1698431365
transform 1 0 45808 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_6
timestamp 1698431365
transform 1 0 2016 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_8
timestamp 1698431365
transform 1 0 2240 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_27
timestamp 1698431365
transform 1 0 4368 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_47
timestamp 1698431365
transform 1 0 6608 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_55
timestamp 1698431365
transform 1 0 7504 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_83
timestamp 1698431365
transform 1 0 10640 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_87
timestamp 1698431365
transform 1 0 11088 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_93
timestamp 1698431365
transform 1 0 11760 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_95
timestamp 1698431365
transform 1 0 11984 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_102
timestamp 1698431365
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_104
timestamp 1698431365
transform 1 0 12992 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_111
timestamp 1698431365
transform 1 0 13776 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_144
timestamp 1698431365
transform 1 0 17472 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_173
timestamp 1698431365
transform 1 0 20720 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_182
timestamp 1698431365
transform 1 0 21728 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_189
timestamp 1698431365
transform 1 0 22512 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_240
timestamp 1698431365
transform 1 0 28224 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_242
timestamp 1698431365
transform 1 0 28448 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_266
timestamp 1698431365
transform 1 0 31136 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_270
timestamp 1698431365
transform 1 0 31584 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_272
timestamp 1698431365
transform 1 0 31808 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_278
timestamp 1698431365
transform 1 0 32480 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_282
timestamp 1698431365
transform 1 0 32928 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_325
timestamp 1698431365
transform 1 0 37744 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_329
timestamp 1698431365
transform 1 0 38192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_331
timestamp 1698431365
transform 1 0 38416 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_383
timestamp 1698431365
transform 1 0 44240 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_419
timestamp 1698431365
transform 1 0 48272 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_31
timestamp 1698431365
transform 1 0 4816 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_33
timestamp 1698431365
transform 1 0 5040 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_69
timestamp 1698431365
transform 1 0 9072 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_97
timestamp 1698431365
transform 1 0 12208 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_136
timestamp 1698431365
transform 1 0 16576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_225
timestamp 1698431365
transform 1 0 26544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_279
timestamp 1698431365
transform 1 0 32592 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_297
timestamp 1698431365
transform 1 0 34608 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_299
timestamp 1698431365
transform 1 0 34832 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_304
timestamp 1698431365
transform 1 0 35392 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_306
timestamp 1698431365
transform 1 0 35616 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_315
timestamp 1698431365
transform 1 0 36624 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_333
timestamp 1698431365
transform 1 0 38640 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_337
timestamp 1698431365
transform 1 0 39088 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_339
timestamp 1698431365
transform 1 0 39312 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_2
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_10
timestamp 1698431365
transform 1 0 2464 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_33
timestamp 1698431365
transform 1 0 5040 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_45
timestamp 1698431365
transform 1 0 6384 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_84
timestamp 1698431365
transform 1 0 10752 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_92
timestamp 1698431365
transform 1 0 11648 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_96
timestamp 1698431365
transform 1 0 12096 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_99
timestamp 1698431365
transform 1 0 12432 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_103
timestamp 1698431365
transform 1 0 12880 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_111
timestamp 1698431365
transform 1 0 13776 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_119
timestamp 1698431365
transform 1 0 14672 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_123
timestamp 1698431365
transform 1 0 15120 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_128
timestamp 1698431365
transform 1 0 15680 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_222
timestamp 1698431365
transform 1 0 26208 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_224
timestamp 1698431365
transform 1 0 26432 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_237
timestamp 1698431365
transform 1 0 27888 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_251
timestamp 1698431365
transform 1 0 29456 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_264
timestamp 1698431365
transform 1 0 30912 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_268
timestamp 1698431365
transform 1 0 31360 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_270
timestamp 1698431365
transform 1 0 31584 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_285
timestamp 1698431365
transform 1 0 33264 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_326
timestamp 1698431365
transform 1 0 37856 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_330
timestamp 1698431365
transform 1 0 38304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_332
timestamp 1698431365
transform 1 0 38528 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_345
timestamp 1698431365
transform 1 0 39984 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_371
timestamp 1698431365
transform 1 0 42896 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_375
timestamp 1698431365
transform 1 0 43344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_377
timestamp 1698431365
transform 1 0 43568 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_31
timestamp 1698431365
transform 1 0 4816 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_63
timestamp 1698431365
transform 1 0 8400 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_67
timestamp 1698431365
transform 1 0 8848 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_69
timestamp 1698431365
transform 1 0 9072 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_107
timestamp 1698431365
transform 1 0 13328 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_109
timestamp 1698431365
transform 1 0 13552 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_116
timestamp 1698431365
transform 1 0 14336 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_124
timestamp 1698431365
transform 1 0 15232 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_200
timestamp 1698431365
transform 1 0 23744 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_222
timestamp 1698431365
transform 1 0 26208 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_229
timestamp 1698431365
transform 1 0 26992 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_250
timestamp 1698431365
transform 1 0 29344 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_254
timestamp 1698431365
transform 1 0 29792 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_265
timestamp 1698431365
transform 1 0 31024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_286
timestamp 1698431365
transform 1 0 33376 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_298
timestamp 1698431365
transform 1 0 34720 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_360
timestamp 1698431365
transform 1 0 41664 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_364
timestamp 1698431365
transform 1 0 42112 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_370
timestamp 1698431365
transform 1 0 42784 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_378
timestamp 1698431365
transform 1 0 43680 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_382
timestamp 1698431365
transform 1 0 44128 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_384
timestamp 1698431365
transform 1 0 44352 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_393
timestamp 1698431365
transform 1 0 45360 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_418
timestamp 1698431365
transform 1 0 48160 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_87
timestamp 1698431365
transform 1 0 11088 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_91
timestamp 1698431365
transform 1 0 11536 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_113
timestamp 1698431365
transform 1 0 14000 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_168
timestamp 1698431365
transform 1 0 20160 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_210
timestamp 1698431365
transform 1 0 24864 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_214
timestamp 1698431365
transform 1 0 25312 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_255
timestamp 1698431365
transform 1 0 29904 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_259
timestamp 1698431365
transform 1 0 30352 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_303
timestamp 1698431365
transform 1 0 35280 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_307
timestamp 1698431365
transform 1 0 35728 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_312
timestamp 1698431365
transform 1 0 36288 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_314
timestamp 1698431365
transform 1 0 36512 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_319
timestamp 1698431365
transform 1 0 37072 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_354
timestamp 1698431365
transform 1 0 40992 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_387
timestamp 1698431365
transform 1 0 44688 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_34
timestamp 1698431365
transform 1 0 5152 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_38
timestamp 1698431365
transform 1 0 5600 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_40
timestamp 1698431365
transform 1 0 5824 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_74
timestamp 1698431365
transform 1 0 9632 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_97
timestamp 1698431365
transform 1 0 12208 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_103
timestamp 1698431365
transform 1 0 12880 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_107
timestamp 1698431365
transform 1 0 13328 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_109
timestamp 1698431365
transform 1 0 13552 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_116
timestamp 1698431365
transform 1 0 14336 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_142
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_146
timestamp 1698431365
transform 1 0 17696 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_149
timestamp 1698431365
transform 1 0 18032 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_205
timestamp 1698431365
transform 1 0 24304 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_212
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_216
timestamp 1698431365
transform 1 0 25536 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_265
timestamp 1698431365
transform 1 0 31024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_269
timestamp 1698431365
transform 1 0 31472 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_277
timestamp 1698431365
transform 1 0 32368 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_279
timestamp 1698431365
transform 1 0 32592 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_286
timestamp 1698431365
transform 1 0 33376 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_302
timestamp 1698431365
transform 1 0 35168 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_310
timestamp 1698431365
transform 1 0 36064 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_328
timestamp 1698431365
transform 1 0 38080 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_336
timestamp 1698431365
transform 1 0 38976 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_2
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698431365
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_37
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_53
timestamp 1698431365
transform 1 0 7280 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_150
timestamp 1698431365
transform 1 0 18144 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_154
timestamp 1698431365
transform 1 0 18592 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_174
timestamp 1698431365
transform 1 0 20832 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_183
timestamp 1698431365
transform 1 0 21840 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_185
timestamp 1698431365
transform 1 0 22064 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_214
timestamp 1698431365
transform 1 0 25312 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_263
timestamp 1698431365
transform 1 0 30800 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_273
timestamp 1698431365
transform 1 0 31920 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_279
timestamp 1698431365
transform 1 0 32592 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_281
timestamp 1698431365
transform 1 0 32816 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_317
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_321
timestamp 1698431365
transform 1 0 37296 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_328
timestamp 1698431365
transform 1 0 38080 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_336
timestamp 1698431365
transform 1 0 38976 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_391
timestamp 1698431365
transform 1 0 45136 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_418
timestamp 1698431365
transform 1 0 48160 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_2
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_34
timestamp 1698431365
transform 1 0 5152 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_38
timestamp 1698431365
transform 1 0 5600 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_102
timestamp 1698431365
transform 1 0 12768 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_106
timestamp 1698431365
transform 1 0 13216 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_114
timestamp 1698431365
transform 1 0 14112 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_153
timestamp 1698431365
transform 1 0 18480 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_209
timestamp 1698431365
transform 1 0 24752 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_221
timestamp 1698431365
transform 1 0 26096 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_225
timestamp 1698431365
transform 1 0 26544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_277
timestamp 1698431365
transform 1 0 32368 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_279
timestamp 1698431365
transform 1 0 32592 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_308
timestamp 1698431365
transform 1 0 35840 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_320
timestamp 1698431365
transform 1 0 37184 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_324
timestamp 1698431365
transform 1 0 37632 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_326
timestamp 1698431365
transform 1 0 37856 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_370
timestamp 1698431365
transform 1 0 42784 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_372
timestamp 1698431365
transform 1 0 43008 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_2
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698431365
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_37
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_53
timestamp 1698431365
transform 1 0 7280 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_98
timestamp 1698431365
transform 1 0 12320 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_119
timestamp 1698431365
transform 1 0 14672 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_227
timestamp 1698431365
transform 1 0 26768 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_231
timestamp 1698431365
transform 1 0 27216 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_239
timestamp 1698431365
transform 1 0 28112 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_243
timestamp 1698431365
transform 1 0 28560 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_247
timestamp 1698431365
transform 1 0 29008 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_255
timestamp 1698431365
transform 1 0 29904 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_282
timestamp 1698431365
transform 1 0 32928 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_286
timestamp 1698431365
transform 1 0 33376 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_295
timestamp 1698431365
transform 1 0 34384 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_303
timestamp 1698431365
transform 1 0 35280 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_313
timestamp 1698431365
transform 1 0 36400 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_335
timestamp 1698431365
transform 1 0 38864 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_337
timestamp 1698431365
transform 1 0 39088 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_381
timestamp 1698431365
transform 1 0 44016 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_416
timestamp 1698431365
transform 1 0 47936 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_66
timestamp 1698431365
transform 1 0 8736 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_72
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_80
timestamp 1698431365
transform 1 0 10304 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_139
timestamp 1698431365
transform 1 0 16912 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_142
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_203
timestamp 1698431365
transform 1 0 24080 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_205
timestamp 1698431365
transform 1 0 24304 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_221
timestamp 1698431365
transform 1 0 26096 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_225
timestamp 1698431365
transform 1 0 26544 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_233
timestamp 1698431365
transform 1 0 27440 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_263
timestamp 1698431365
transform 1 0 30800 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_282
timestamp 1698431365
transform 1 0 32928 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_284
timestamp 1698431365
transform 1 0 33152 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_314
timestamp 1698431365
transform 1 0 36512 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_316
timestamp 1698431365
transform 1 0 36736 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_346
timestamp 1698431365
transform 1 0 40096 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_356
timestamp 1698431365
transform 1 0 41216 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_358
timestamp 1698431365
transform 1 0 41440 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_411
timestamp 1698431365
transform 1 0 47376 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_2
timestamp 1698431365
transform 1 0 1568 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_36
timestamp 1698431365
transform 1 0 5376 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_70
timestamp 1698431365
transform 1 0 9184 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_78
timestamp 1698431365
transform 1 0 10080 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_90
timestamp 1698431365
transform 1 0 11424 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_98
timestamp 1698431365
transform 1 0 12320 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_104
timestamp 1698431365
transform 1 0 12992 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_138
timestamp 1698431365
transform 1 0 16800 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_146
timestamp 1698431365
transform 1 0 17696 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_150
timestamp 1698431365
transform 1 0 18144 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_201
timestamp 1698431365
transform 1 0 23856 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_203
timestamp 1698431365
transform 1 0 24080 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_235
timestamp 1698431365
transform 1 0 27664 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_237
timestamp 1698431365
transform 1 0 27888 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_271
timestamp 1698431365
transform 1 0 31696 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_300
timestamp 1698431365
transform 1 0 34944 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_304
timestamp 1698431365
transform 1 0 35392 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_308
timestamp 1698431365
transform 1 0 35840 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_324
timestamp 1698431365
transform 1 0 37632 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_331
timestamp 1698431365
transform 1 0 38416 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_339
timestamp 1698431365
transform 1 0 39312 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_342
timestamp 1698431365
transform 1 0 39648 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_350
timestamp 1698431365
transform 1 0 40544 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_354
timestamp 1698431365
transform 1 0 40992 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_356
timestamp 1698431365
transform 1 0 41216 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_367
timestamp 1698431365
transform 1 0 42448 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_371
timestamp 1698431365
transform 1 0 42896 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_382
timestamp 1698431365
transform 1 0 44128 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_386
timestamp 1698431365
transform 1 0 44576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_416
timestamp 1698431365
transform 1 0 47936 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input1
timestamp 1698431365
transform -1 0 48384 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform 1 0 45024 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input3
timestamp 1698431365
transform -1 0 48384 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input4
timestamp 1698431365
transform -1 0 48384 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input5
timestamp 1698431365
transform -1 0 48384 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input6
timestamp 1698431365
transform -1 0 48384 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input7
timestamp 1698431365
transform -1 0 48384 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input8
timestamp 1698431365
transform -1 0 48384 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input9
timestamp 1698431365
transform -1 0 48384 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input10
timestamp 1698431365
transform -1 0 48384 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input11
timestamp 1698431365
transform -1 0 32928 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input12
timestamp 1698431365
transform -1 0 44128 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input13
timestamp 1698431365
transform 1 0 18704 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17472 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698431365
transform 1 0 20944 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698431365
transform 1 0 28896 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698431365
transform -1 0 36400 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698431365
transform -1 0 42560 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698431365
transform -1 0 16576 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698431365
transform 1 0 17808 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_55 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 48608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_56
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 48608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_57
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 48608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_58
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 48608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_59
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 48608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_60
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 48608 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_61
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 48608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_62
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 48608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_63
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 48608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_64
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 48608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_65
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 48608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_66
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 48608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_67
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 48608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_68
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 48608 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_69
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 48608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_70
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 48608 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_71
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 48608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_72
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 48608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_73
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 48608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_74
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 48608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_75
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 48608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_76
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 48608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_77
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 48608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_78
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 48608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_79
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 48608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_80
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 48608 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_81
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 48608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_82
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 48608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_83
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 48608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_84
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 48608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_85
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 48608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_86
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 48608 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_87
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 48608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_88
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 48608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_89
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 48608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_90
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 48608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_91
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 48608 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_92
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 48608 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_93
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 48608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_94
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 48608 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_95
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 48608 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_96
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 48608 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_97
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 48608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_98
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 48608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_99
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 48608 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_100
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 48608 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_101
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 48608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_102
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 48608 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_103
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 48608 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_104
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 48608 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_105
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 48608 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_106
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 48608 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_107
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 48608 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_108
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 48608 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_109
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 48608 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_110 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_111
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_112
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_113
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_114
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_115
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_116
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_117
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_118
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_119
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_120
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_121
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_122
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_123
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_124
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_125
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_126
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_127
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_128
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_129
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_130
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_131
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_132
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_133
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_134
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_135
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_136
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_137
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_138
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_139
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_140
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_141
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_142
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_143
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_144
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_145
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_146
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_147
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_148
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_149
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_150
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_151
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_152
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_153
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_154
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_155
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_156
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_157
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_158
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_159
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_160
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_161
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_162
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_163
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_164
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_165
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_166
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_167
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_168
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_169
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_170
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_171
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_172
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_173
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_174
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_175
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_176
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_177
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_178
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_179
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_180
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_181
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_182
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_183
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_184
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_185
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_186
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_187
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_188
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_189
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_190
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_191
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_192
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_193
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_194
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_195
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_196
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_197
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_198
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_199
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_200
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_201
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_202
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_203
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_204
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_205
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_206
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_207
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_208
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_209
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_210
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_211
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_212
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_213
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_214
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_215
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_216
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_217
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_218
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_219
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_220
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_221
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_222
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_223
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_224
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_225
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_226
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_227
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_228
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_229
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_230
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_231
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_232
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_233
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_234
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_235
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_236
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_237
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_238
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_239
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_240
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_241
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_242
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_243
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_244
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_245
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_246
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_247
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_248
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_249
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_250
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_251
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_252
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_253
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_254
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_255
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_256
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_257
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_258
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_259
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_260
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_261
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_262
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_263
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_264
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_265
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_266
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_267
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_268
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_269
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_270
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_271
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_272
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_273
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_274
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_275
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_276
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_277
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_278
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_279
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_280
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_281
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_282
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_283
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_284
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_285
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_286
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_287
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_288
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_289
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_290
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_291
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_292
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_293
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_294
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_295
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_296
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_297
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_298
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_299
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_300
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_301
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_302
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_303
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_304
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_305
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_306
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_307
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_308
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_309
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_310
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_311
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_312
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_313
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_314
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_315
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_316
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_317
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_318
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_319
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_320
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_321
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_322
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_323
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_324
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_325
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_326
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_327
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_328
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_329
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_330
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_331
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_332
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_333
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_334
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_335
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_336
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_337
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_338
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_339
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_340
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_341
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_342
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_343
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_344
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_345
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_346
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_347
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_348
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_349
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_350
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_351
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_352
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_353
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_354
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_355
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_356
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_357
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_358
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_359
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_360
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_361
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_362
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_363
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_364
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_365
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_366
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_367
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_368
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_369
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_370
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_371
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_372
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_373
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_374
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_375
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_376
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_377
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_378
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_379
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_380
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_381
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_382
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_383
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_384
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_385
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_386
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_387
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_388
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_389
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_390
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_391
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_392
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_393
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_394
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_395
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_396
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_397
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_398
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_399
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_400
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_401
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_402
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_403
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_404
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_405
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_406
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_407
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_408
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_409
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_410
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_411
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_412
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_413
timestamp 1698431365
transform 1 0 5152 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_414
timestamp 1698431365
transform 1 0 8960 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_415
timestamp 1698431365
transform 1 0 12768 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_416
timestamp 1698431365
transform 1 0 16576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_417
timestamp 1698431365
transform 1 0 20384 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_418
timestamp 1698431365
transform 1 0 24192 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_419
timestamp 1698431365
transform 1 0 28000 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_420
timestamp 1698431365
transform 1 0 31808 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_421
timestamp 1698431365
transform 1 0 35616 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_422
timestamp 1698431365
transform 1 0 39424 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_423
timestamp 1698431365
transform 1 0 43232 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_424
timestamp 1698431365
transform 1 0 47040 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_23 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 4144 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_24
timestamp 1698431365
transform -1 0 5824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_25
timestamp 1698431365
transform -1 0 7280 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_26
timestamp 1698431365
transform -1 0 8848 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_27
timestamp 1698431365
transform -1 0 10416 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_28
timestamp 1698431365
transform -1 0 11984 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_29
timestamp 1698431365
transform 1 0 12320 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_30
timestamp 1698431365
transform 1 0 13216 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_31
timestamp 1698431365
transform -1 0 25536 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_32
timestamp 1698431365
transform -1 0 25536 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_33
timestamp 1698431365
transform -1 0 26096 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_34
timestamp 1698431365
transform -1 0 27664 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_35
timestamp 1698431365
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_36
timestamp 1698431365
transform -1 0 41888 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_37
timestamp 1698431365
transform -1 0 43008 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_38
timestamp 1698431365
transform -1 0 44800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_39
timestamp 1698431365
transform -1 0 45248 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_40
timestamp 1698431365
transform -1 0 46480 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_41
timestamp 1698431365
transform -1 0 39200 0 1 3136
box -86 -86 534 870
<< labels >>
flabel metal3 s 49200 42112 50000 42224 0 FreeSans 448 0 0 0 custom_settings[0]
port 0 nsew signal input
flabel metal3 s 49200 47040 50000 47152 0 FreeSans 448 0 0 0 custom_settings[1]
port 1 nsew signal input
flabel metal3 s 49200 2688 50000 2800 0 FreeSans 448 0 0 0 io_in_1[0]
port 2 nsew signal input
flabel metal3 s 49200 7616 50000 7728 0 FreeSans 448 0 0 0 io_in_1[1]
port 3 nsew signal input
flabel metal3 s 49200 12544 50000 12656 0 FreeSans 448 0 0 0 io_in_1[2]
port 4 nsew signal input
flabel metal3 s 49200 17472 50000 17584 0 FreeSans 448 0 0 0 io_in_1[3]
port 5 nsew signal input
flabel metal3 s 49200 22400 50000 22512 0 FreeSans 448 0 0 0 io_in_1[4]
port 6 nsew signal input
flabel metal3 s 49200 27328 50000 27440 0 FreeSans 448 0 0 0 io_in_1[5]
port 7 nsew signal input
flabel metal3 s 49200 32256 50000 32368 0 FreeSans 448 0 0 0 io_in_1[6]
port 8 nsew signal input
flabel metal3 s 49200 37184 50000 37296 0 FreeSans 448 0 0 0 io_in_1[7]
port 9 nsew signal input
flabel metal2 s 30912 49200 31024 50000 0 FreeSans 448 90 0 0 io_in_2[0]
port 10 nsew signal input
flabel metal2 s 43232 49200 43344 50000 0 FreeSans 448 90 0 0 io_in_2[1]
port 11 nsew signal input
flabel metal2 s 3584 0 3696 800 0 FreeSans 448 90 0 0 io_out[0]
port 12 nsew signal tristate
flabel metal2 s 19264 0 19376 800 0 FreeSans 448 90 0 0 io_out[10]
port 13 nsew signal tristate
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 io_out[11]
port 14 nsew signal tristate
flabel metal2 s 22400 0 22512 800 0 FreeSans 448 90 0 0 io_out[12]
port 15 nsew signal tristate
flabel metal2 s 23968 0 24080 800 0 FreeSans 448 90 0 0 io_out[13]
port 16 nsew signal tristate
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 io_out[14]
port 17 nsew signal tristate
flabel metal2 s 27104 0 27216 800 0 FreeSans 448 90 0 0 io_out[15]
port 18 nsew signal tristate
flabel metal2 s 28672 0 28784 800 0 FreeSans 448 90 0 0 io_out[16]
port 19 nsew signal tristate
flabel metal2 s 30240 0 30352 800 0 FreeSans 448 90 0 0 io_out[17]
port 20 nsew signal tristate
flabel metal2 s 31808 0 31920 800 0 FreeSans 448 90 0 0 io_out[18]
port 21 nsew signal tristate
flabel metal2 s 33376 0 33488 800 0 FreeSans 448 90 0 0 io_out[19]
port 22 nsew signal tristate
flabel metal2 s 5152 0 5264 800 0 FreeSans 448 90 0 0 io_out[1]
port 23 nsew signal tristate
flabel metal2 s 34944 0 35056 800 0 FreeSans 448 90 0 0 io_out[20]
port 24 nsew signal tristate
flabel metal2 s 36512 0 36624 800 0 FreeSans 448 90 0 0 io_out[21]
port 25 nsew signal tristate
flabel metal2 s 38080 0 38192 800 0 FreeSans 448 90 0 0 io_out[22]
port 26 nsew signal tristate
flabel metal2 s 39648 0 39760 800 0 FreeSans 448 90 0 0 io_out[23]
port 27 nsew signal tristate
flabel metal2 s 41216 0 41328 800 0 FreeSans 448 90 0 0 io_out[24]
port 28 nsew signal tristate
flabel metal2 s 42784 0 42896 800 0 FreeSans 448 90 0 0 io_out[25]
port 29 nsew signal tristate
flabel metal2 s 44352 0 44464 800 0 FreeSans 448 90 0 0 io_out[26]
port 30 nsew signal tristate
flabel metal2 s 45920 0 46032 800 0 FreeSans 448 90 0 0 io_out[27]
port 31 nsew signal tristate
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 io_out[2]
port 32 nsew signal tristate
flabel metal2 s 8288 0 8400 800 0 FreeSans 448 90 0 0 io_out[3]
port 33 nsew signal tristate
flabel metal2 s 9856 0 9968 800 0 FreeSans 448 90 0 0 io_out[4]
port 34 nsew signal tristate
flabel metal2 s 11424 0 11536 800 0 FreeSans 448 90 0 0 io_out[5]
port 35 nsew signal tristate
flabel metal2 s 12992 0 13104 800 0 FreeSans 448 90 0 0 io_out[6]
port 36 nsew signal tristate
flabel metal2 s 14560 0 14672 800 0 FreeSans 448 90 0 0 io_out[7]
port 37 nsew signal tristate
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 io_out[8]
port 38 nsew signal tristate
flabel metal2 s 17696 0 17808 800 0 FreeSans 448 90 0 0 io_out[9]
port 39 nsew signal tristate
flabel metal2 s 18592 49200 18704 50000 0 FreeSans 448 90 0 0 rst_n
port 40 nsew signal input
flabel metal4 s 4448 3076 4768 46316 0 FreeSans 1280 90 0 0 vdd
port 41 nsew power bidirectional
flabel metal4 s 35168 3076 35488 46316 0 FreeSans 1280 90 0 0 vdd
port 41 nsew power bidirectional
flabel metal4 s 19808 3076 20128 46316 0 FreeSans 1280 90 0 0 vss
port 42 nsew ground bidirectional
flabel metal2 s 6272 49200 6384 50000 0 FreeSans 448 90 0 0 wb_clk_i
port 43 nsew signal input
rlabel metal1 24976 46256 24976 46256 0 vdd
rlabel metal1 24976 45472 24976 45472 0 vss
rlabel metal2 31864 17192 31864 17192 0 _0000_
rlabel metal2 32872 16408 32872 16408 0 _0001_
rlabel metal2 33152 13048 33152 13048 0 _0002_
rlabel metal2 31304 11312 31304 11312 0 _0003_
rlabel metal2 29512 17976 29512 17976 0 _0004_
rlabel metal2 32424 7896 32424 7896 0 _0005_
rlabel metal2 32200 5432 32200 5432 0 _0006_
rlabel metal2 36120 6272 36120 6272 0 _0007_
rlabel metal2 34776 4144 34776 4144 0 _0008_
rlabel metal3 21896 33432 21896 33432 0 _0009_
rlabel metal3 24416 36344 24416 36344 0 _0010_
rlabel metal2 21504 35784 21504 35784 0 _0011_
rlabel metal2 22680 36512 22680 36512 0 _0012_
rlabel metal2 23688 17192 23688 17192 0 _0013_
rlabel metal2 16632 14336 16632 14336 0 _0014_
rlabel metal2 21448 10416 21448 10416 0 _0015_
rlabel metal2 16744 11760 16744 11760 0 _0016_
rlabel metal2 9688 11032 9688 11032 0 _0017_
rlabel metal2 12376 9352 12376 9352 0 _0018_
rlabel metal2 9016 6720 9016 6720 0 _0019_
rlabel metal3 9632 7336 9632 7336 0 _0020_
rlabel metal2 10808 6384 10808 6384 0 _0021_
rlabel metal2 21560 5488 21560 5488 0 _0022_
rlabel metal2 23352 8456 23352 8456 0 _0023_
rlabel metal2 18872 10248 18872 10248 0 _0024_
rlabel metal2 18424 8680 18424 8680 0 _0025_
rlabel metal3 18984 6552 18984 6552 0 _0026_
rlabel metal2 14616 7784 14616 7784 0 _0027_
rlabel metal2 16296 6328 16296 6328 0 _0028_
rlabel metal2 14280 4816 14280 4816 0 _0029_
rlabel metal2 17192 4312 17192 4312 0 _0030_
rlabel metal2 19320 5432 19320 5432 0 _0031_
rlabel metal2 17696 22232 17696 22232 0 _0032_
rlabel metal2 9072 19320 9072 19320 0 _0033_
rlabel metal3 2940 19096 2940 19096 0 _0034_
rlabel metal3 3136 13160 3136 13160 0 _0035_
rlabel metal3 3472 11480 3472 11480 0 _0036_
rlabel metal2 7224 12768 7224 12768 0 _0037_
rlabel metal2 6328 9464 6328 9464 0 _0038_
rlabel metal3 10024 4424 10024 4424 0 _0039_
rlabel metal2 31528 10136 31528 10136 0 _0040_
rlabel metal2 34160 12152 34160 12152 0 _0041_
rlabel metal2 36512 10584 36512 10584 0 _0042_
rlabel metal2 36344 9128 36344 9128 0 _0043_
rlabel metal2 41720 18256 41720 18256 0 _0044_
rlabel metal2 43512 16520 43512 16520 0 _0045_
rlabel metal3 47096 15400 47096 15400 0 _0046_
rlabel metal3 46872 16184 46872 16184 0 _0047_
rlabel metal2 35000 21280 35000 21280 0 _0048_
rlabel metal2 32592 19320 32592 19320 0 _0049_
rlabel metal3 37072 18312 37072 18312 0 _0050_
rlabel metal3 36680 19880 36680 19880 0 _0051_
rlabel metal2 31416 26208 31416 26208 0 _0052_
rlabel metal2 33880 24864 33880 24864 0 _0053_
rlabel metal3 33880 27720 33880 27720 0 _0054_
rlabel metal2 35168 28840 35168 28840 0 _0055_
rlabel metal2 41944 31416 41944 31416 0 _0056_
rlabel metal2 47208 31304 47208 31304 0 _0057_
rlabel metal2 47208 30184 47208 30184 0 _0058_
rlabel metal3 42504 31864 42504 31864 0 _0059_
rlabel metal2 26600 3976 26600 3976 0 _0060_
rlabel metal2 25032 10192 25032 10192 0 _0061_
rlabel metal2 28728 9408 28728 9408 0 _0062_
rlabel metal2 26600 6720 26600 6720 0 _0063_
rlabel metal2 31192 7952 31192 7952 0 _0064_
rlabel metal2 3304 17136 3304 17136 0 _0065_
rlabel metal2 2520 15792 2520 15792 0 _0066_
rlabel metal3 4480 10472 4480 10472 0 _0067_
rlabel metal2 2856 7728 2856 7728 0 _0068_
rlabel metal3 3864 6104 3864 6104 0 _0069_
rlabel metal2 6440 7056 6440 7056 0 _0070_
rlabel metal2 7560 3920 7560 3920 0 _0071_
rlabel metal2 7784 4760 7784 4760 0 _0072_
rlabel metal3 24640 26488 24640 26488 0 _0073_
rlabel metal2 21840 23912 21840 23912 0 _0074_
rlabel metal2 16408 34552 16408 34552 0 _0075_
rlabel metal2 15400 32088 15400 32088 0 _0076_
rlabel metal2 18368 33208 18368 33208 0 _0077_
rlabel metal2 20608 31192 20608 31192 0 _0078_
rlabel metal2 23968 41272 23968 41272 0 _0079_
rlabel metal2 20776 45304 20776 45304 0 _0080_
rlabel metal2 24696 45528 24696 45528 0 _0081_
rlabel metal2 24696 42056 24696 42056 0 _0082_
rlabel metal2 30072 4872 30072 4872 0 _0083_
rlabel metal2 22568 4648 22568 4648 0 _0084_
rlabel metal2 32984 4256 32984 4256 0 _0085_
rlabel metal2 5768 16912 5768 16912 0 _0086_
rlabel metal3 18592 29624 18592 29624 0 _0087_
rlabel metal3 18200 24584 18200 24584 0 _0088_
rlabel metal2 24584 24752 24584 24752 0 _0089_
rlabel metal2 16744 27384 16744 27384 0 _0090_
rlabel metal2 29512 23240 29512 23240 0 _0091_
rlabel metal3 25144 22456 25144 22456 0 _0092_
rlabel metal2 37240 32704 37240 32704 0 _0093_
rlabel metal2 37912 36848 37912 36848 0 _0094_
rlabel metal2 37352 35280 37352 35280 0 _0095_
rlabel metal2 40376 35000 40376 35000 0 _0096_
rlabel metal2 39144 33208 39144 33208 0 _0097_
rlabel metal2 43512 35280 43512 35280 0 _0098_
rlabel metal2 46088 34104 46088 34104 0 _0099_
rlabel metal2 46312 36064 46312 36064 0 _0100_
rlabel metal2 14056 35112 14056 35112 0 _0101_
rlabel metal2 2520 34440 2520 34440 0 _0102_
rlabel metal2 2968 36792 2968 36792 0 _0103_
rlabel metal2 4648 39312 4648 39312 0 _0104_
rlabel metal2 2744 38416 2744 38416 0 _0105_
rlabel metal2 5768 37744 5768 37744 0 _0106_
rlabel metal3 8848 39480 8848 39480 0 _0107_
rlabel metal2 23912 39060 23912 39060 0 _0108_
rlabel metal2 26432 41272 26432 41272 0 _0109_
rlabel metal3 28280 42616 28280 42616 0 _0110_
rlabel metal3 30408 41832 30408 41832 0 _0111_
rlabel metal3 29792 44968 29792 44968 0 _0112_
rlabel metal3 34888 44520 34888 44520 0 _0113_
rlabel metal2 34328 43064 34328 43064 0 _0114_
rlabel metal2 39144 45416 39144 45416 0 _0115_
rlabel metal3 41048 42616 41048 42616 0 _0116_
rlabel metal2 38136 41496 38136 41496 0 _0117_
rlabel metal2 43512 41552 43512 41552 0 _0118_
rlabel metal2 41720 43932 41720 43932 0 _0119_
rlabel metal2 45640 43932 45640 43932 0 _0120_
rlabel metal2 47432 43176 47432 43176 0 _0121_
rlabel metal2 47544 44660 47544 44660 0 _0122_
rlabel metal2 47488 39704 47488 39704 0 _0123_
rlabel metal3 6440 34216 6440 34216 0 _0124_
rlabel metal2 11816 25144 11816 25144 0 _0125_
rlabel metal3 11368 24024 11368 24024 0 _0126_
rlabel metal3 11032 26488 11032 26488 0 _0127_
rlabel metal2 8736 21784 8736 21784 0 _0128_
rlabel metal2 6384 20888 6384 20888 0 _0129_
rlabel metal2 2520 21168 2520 21168 0 _0130_
rlabel metal2 2520 22008 2520 22008 0 _0131_
rlabel metal3 3808 24584 3808 24584 0 _0132_
rlabel metal3 4480 26152 4480 26152 0 _0133_
rlabel metal2 2520 27888 2520 27888 0 _0134_
rlabel metal2 3752 29008 3752 29008 0 _0135_
rlabel metal3 4144 30072 4144 30072 0 _0136_
rlabel metal3 4144 31640 4144 31640 0 _0137_
rlabel metal2 4424 31304 4424 31304 0 _0138_
rlabel metal2 8680 31416 8680 31416 0 _0139_
rlabel metal3 10136 29288 10136 29288 0 _0140_
rlabel metal3 7672 26488 7672 26488 0 _0141_
rlabel metal2 23464 14840 23464 14840 0 _0142_
rlabel metal2 25704 19712 25704 19712 0 _0143_
rlabel metal2 26152 15680 26152 15680 0 _0144_
rlabel metal2 27608 14840 27608 14840 0 _0145_
rlabel metal2 22568 12488 22568 12488 0 _0146_
rlabel metal2 26488 11760 26488 11760 0 _0147_
rlabel metal3 7252 38920 7252 38920 0 _0148_
rlabel metal2 11144 33768 11144 33768 0 _0149_
rlabel metal2 15736 33488 15736 33488 0 _0150_
rlabel metal2 12992 35112 12992 35112 0 _0151_
rlabel metal3 11480 31640 11480 31640 0 _0152_
rlabel metal3 37296 16184 37296 16184 0 _0153_
rlabel metal3 37408 15288 37408 15288 0 _0154_
rlabel metal3 42280 15176 42280 15176 0 _0155_
rlabel metal2 47432 14056 47432 14056 0 _0156_
rlabel metal2 47432 12488 47432 12488 0 _0157_
rlabel metal3 46872 9912 46872 9912 0 _0158_
rlabel metal2 47432 7784 47432 7784 0 _0159_
rlabel metal2 46536 8512 46536 8512 0 _0160_
rlabel metal2 47432 6216 47432 6216 0 _0161_
rlabel metal3 40264 4424 40264 4424 0 _0162_
rlabel metal2 44184 4256 44184 4256 0 _0163_
rlabel metal2 37800 7224 37800 7224 0 _0164_
rlabel metal2 27440 21672 27440 21672 0 _0165_
rlabel metal2 38136 22008 38136 22008 0 _0166_
rlabel metal2 37072 23352 37072 23352 0 _0167_
rlabel metal2 37464 27496 37464 27496 0 _0168_
rlabel metal2 39928 29456 39928 29456 0 _0169_
rlabel metal2 46088 29064 46088 29064 0 _0170_
rlabel metal3 45416 26488 45416 26488 0 _0171_
rlabel metal2 45976 25144 45976 25144 0 _0172_
rlabel metal2 46424 23520 46424 23520 0 _0173_
rlabel metal2 45640 21952 45640 21952 0 _0174_
rlabel metal2 46032 20888 46032 20888 0 _0175_
rlabel metal2 43624 17808 43624 17808 0 _0176_
rlabel metal2 46088 19880 46088 19880 0 _0177_
rlabel metal3 31808 22232 31808 22232 0 _0178_
rlabel metal2 14952 36960 14952 36960 0 _0179_
rlabel metal3 17248 37912 17248 37912 0 _0180_
rlabel metal2 16744 39816 16744 39816 0 _0181_
rlabel metal2 14056 42392 14056 42392 0 _0182_
rlabel metal3 18312 44184 18312 44184 0 _0183_
rlabel metal2 14616 44744 14616 44744 0 _0184_
rlabel metal2 12712 44688 12712 44688 0 _0185_
rlabel metal3 10864 43512 10864 43512 0 _0186_
rlabel metal3 8568 43400 8568 43400 0 _0187_
rlabel metal2 6888 42000 6888 42000 0 _0188_
rlabel metal2 10360 40824 10360 40824 0 _0189_
rlabel metal3 13496 38696 13496 38696 0 _0190_
rlabel metal2 21560 29008 21560 29008 0 _0191_
rlabel metal2 22064 22456 22064 22456 0 _0192_
rlabel metal3 20384 23800 20384 23800 0 _0193_
rlabel metal2 11704 28112 11704 28112 0 _0194_
rlabel metal2 12824 29008 12824 29008 0 _0195_
rlabel metal2 13720 27216 13720 27216 0 _0196_
rlabel metal2 13664 23352 13664 23352 0 _0197_
rlabel metal3 12712 21448 12712 21448 0 _0198_
rlabel metal2 15624 20776 15624 20776 0 _0199_
rlabel metal2 13160 18144 13160 18144 0 _0200_
rlabel metal2 22904 32480 22904 32480 0 _0201_
rlabel metal3 25032 28728 25032 28728 0 _0202_
rlabel metal2 27440 26376 27440 26376 0 _0203_
rlabel metal2 29064 31304 29064 31304 0 _0204_
rlabel metal2 29960 31920 29960 31920 0 _0205_
rlabel metal2 26488 34440 26488 34440 0 _0206_
rlabel metal2 28168 36120 28168 36120 0 _0207_
rlabel metal2 29960 36512 29960 36512 0 _0208_
rlabel metal2 29736 34440 29736 34440 0 _0209_
rlabel metal2 34888 32984 34888 32984 0 _0210_
rlabel metal2 33936 34216 33936 34216 0 _0211_
rlabel metal2 32648 36792 32648 36792 0 _0212_
rlabel metal2 34328 38360 34328 38360 0 _0213_
rlabel metal3 16912 17528 16912 17528 0 _0214_
rlabel metal2 10584 17976 10584 17976 0 _0215_
rlabel metal2 6888 17192 6888 17192 0 _0216_
rlabel metal3 8736 15288 8736 15288 0 _0217_
rlabel metal2 9128 13328 9128 13328 0 _0218_
rlabel metal2 15736 15624 15736 15624 0 _0219_
rlabel metal2 15512 12656 15512 12656 0 _0220_
rlabel metal2 14840 10304 14840 10304 0 _0221_
rlabel metal2 23576 19376 23576 19376 0 _0222_
rlabel metal3 21448 22232 21448 22232 0 _0223_
rlabel metal3 47040 45752 47040 45752 0 _0224_
rlabel metal2 46144 38696 46144 38696 0 _0225_
rlabel metal2 9464 34216 9464 34216 0 _0226_
rlabel metal2 9240 36400 9240 36400 0 _0227_
rlabel metal3 8568 34776 8568 34776 0 _0228_
rlabel metal2 8064 35448 8064 35448 0 _0229_
rlabel metal2 7392 34888 7392 34888 0 _0230_
rlabel metal2 7448 19600 7448 19600 0 _0231_
rlabel metal2 7112 21616 7112 21616 0 _0232_
rlabel metal2 7952 26264 7952 26264 0 _0233_
rlabel metal2 11592 25032 11592 25032 0 _0234_
rlabel metal3 6888 25368 6888 25368 0 _0235_
rlabel metal2 6048 25256 6048 25256 0 _0236_
rlabel metal3 8232 25256 8232 25256 0 _0237_
rlabel metal2 12040 24584 12040 24584 0 _0238_
rlabel metal2 10920 25480 10920 25480 0 _0239_
rlabel metal2 10472 24920 10472 24920 0 _0240_
rlabel metal2 10248 24696 10248 24696 0 _0241_
rlabel metal2 10696 25872 10696 25872 0 _0242_
rlabel metal2 10192 26376 10192 26376 0 _0243_
rlabel metal2 6832 23800 6832 23800 0 _0244_
rlabel metal2 5656 22736 5656 22736 0 _0245_
rlabel metal3 8120 21672 8120 21672 0 _0246_
rlabel metal2 8904 22232 8904 22232 0 _0247_
rlabel metal2 7560 21616 7560 21616 0 _0248_
rlabel metal2 6048 21672 6048 21672 0 _0249_
rlabel metal2 3304 23464 3304 23464 0 _0250_
rlabel metal2 6552 21448 6552 21448 0 _0251_
rlabel metal2 4984 21896 4984 21896 0 _0252_
rlabel metal2 4536 21616 4536 21616 0 _0253_
rlabel metal2 3976 22232 3976 22232 0 _0254_
rlabel metal2 3640 22344 3640 22344 0 _0255_
rlabel metal2 3080 28672 3080 28672 0 _0256_
rlabel metal2 2744 25032 2744 25032 0 _0257_
rlabel metal2 4536 24024 4536 24024 0 _0258_
rlabel metal2 5432 25480 5432 25480 0 _0259_
rlabel metal2 4312 25536 4312 25536 0 _0260_
rlabel metal3 5208 25480 5208 25480 0 _0261_
rlabel metal2 3528 25984 3528 25984 0 _0262_
rlabel metal2 3416 28560 3416 28560 0 _0263_
rlabel metal2 4424 25592 4424 25592 0 _0264_
rlabel metal2 3976 28448 3976 28448 0 _0265_
rlabel metal2 3640 28896 3640 28896 0 _0266_
rlabel metal2 7336 32144 7336 32144 0 _0267_
rlabel metal3 6496 30072 6496 30072 0 _0268_
rlabel metal3 6608 30184 6608 30184 0 _0269_
rlabel metal3 9576 30968 9576 30968 0 _0270_
rlabel metal2 5992 32424 5992 32424 0 _0271_
rlabel metal2 8568 30240 8568 30240 0 _0272_
rlabel metal2 5936 29624 5936 29624 0 _0273_
rlabel metal2 6944 31192 6944 31192 0 _0274_
rlabel metal2 6440 30968 6440 30968 0 _0275_
rlabel metal2 8288 31192 8288 31192 0 _0276_
rlabel metal2 8848 31080 8848 31080 0 _0277_
rlabel metal2 8680 29008 8680 29008 0 _0278_
rlabel metal2 8344 29680 8344 29680 0 _0279_
rlabel metal3 7168 23800 7168 23800 0 _0280_
rlabel metal3 7840 28392 7840 28392 0 _0281_
rlabel metal3 8624 28504 8624 28504 0 _0282_
rlabel metal2 8792 26544 8792 26544 0 _0283_
rlabel metal2 8232 24416 8232 24416 0 _0284_
rlabel metal2 8456 24808 8456 24808 0 _0285_
rlabel metal3 8176 25368 8176 25368 0 _0286_
rlabel metal2 7336 25648 7336 25648 0 _0287_
rlabel metal2 8344 26432 8344 26432 0 _0288_
rlabel metal2 29624 12768 29624 12768 0 _0289_
rlabel metal2 29400 16128 29400 16128 0 _0290_
rlabel metal2 29064 15904 29064 15904 0 _0291_
rlabel metal3 30072 15848 30072 15848 0 _0292_
rlabel metal2 29736 16408 29736 16408 0 _0293_
rlabel metal2 28280 14280 28280 14280 0 _0294_
rlabel metal2 28728 13720 28728 13720 0 _0295_
rlabel metal3 29176 14280 29176 14280 0 _0296_
rlabel metal2 29400 14224 29400 14224 0 _0297_
rlabel metal2 29120 12936 29120 12936 0 _0298_
rlabel metal2 29736 13832 29736 13832 0 _0299_
rlabel metal2 28056 14168 28056 14168 0 _0300_
rlabel metal2 23352 12208 23352 12208 0 _0301_
rlabel metal2 23576 15204 23576 15204 0 _0302_
rlabel metal2 25984 15624 25984 15624 0 _0303_
rlabel metal2 25872 16856 25872 16856 0 _0304_
rlabel metal2 25648 16632 25648 16632 0 _0305_
rlabel metal2 26376 15176 26376 15176 0 _0306_
rlabel metal2 36008 23016 36008 23016 0 _0307_
rlabel metal2 25536 15288 25536 15288 0 _0308_
rlabel metal2 26040 13440 26040 13440 0 _0309_
rlabel metal3 28392 15288 28392 15288 0 _0310_
rlabel metal2 25704 12376 25704 12376 0 _0311_
rlabel metal2 23800 11648 23800 11648 0 _0312_
rlabel metal2 24192 11592 24192 11592 0 _0313_
rlabel metal2 13720 31304 13720 31304 0 _0314_
rlabel metal2 11256 33712 11256 33712 0 _0315_
rlabel metal2 14504 33376 14504 33376 0 _0316_
rlabel metal3 13328 34776 13328 34776 0 _0317_
rlabel metal2 12040 31640 12040 31640 0 _0318_
rlabel metal2 38696 17024 38696 17024 0 _0319_
rlabel metal2 37016 16128 37016 16128 0 _0320_
rlabel metal2 18424 38724 18424 38724 0 _0321_
rlabel metal2 39480 7896 39480 7896 0 _0322_
rlabel metal2 42168 4200 42168 4200 0 _0323_
rlabel metal2 40264 6384 40264 6384 0 _0324_
rlabel metal3 40936 5768 40936 5768 0 _0325_
rlabel metal2 41384 6664 41384 6664 0 _0326_
rlabel metal2 41384 5488 41384 5488 0 _0327_
rlabel metal2 41272 6328 41272 6328 0 _0328_
rlabel metal2 41272 7560 41272 7560 0 _0329_
rlabel metal3 39004 11368 39004 11368 0 _0330_
rlabel metal2 38304 10584 38304 10584 0 _0331_
rlabel metal3 43792 9240 43792 9240 0 _0332_
rlabel metal2 42056 8288 42056 8288 0 _0333_
rlabel metal2 41384 9072 41384 9072 0 _0334_
rlabel metal2 39592 9520 39592 9520 0 _0335_
rlabel metal2 40936 12432 40936 12432 0 _0336_
rlabel metal2 41384 12656 41384 12656 0 _0337_
rlabel metal2 40824 11424 40824 11424 0 _0338_
rlabel metal2 39256 11480 39256 11480 0 _0339_
rlabel metal2 39872 12152 39872 12152 0 _0340_
rlabel metal2 39928 11144 39928 11144 0 _0341_
rlabel metal2 39424 10024 39424 10024 0 _0342_
rlabel metal2 39816 8960 39816 8960 0 _0343_
rlabel metal2 43960 12208 43960 12208 0 _0344_
rlabel metal2 42784 12152 42784 12152 0 _0345_
rlabel metal2 42000 9800 42000 9800 0 _0346_
rlabel metal2 44352 9800 44352 9800 0 _0347_
rlabel metal2 42952 9968 42952 9968 0 _0348_
rlabel metal2 42168 10024 42168 10024 0 _0349_
rlabel metal2 38696 10416 38696 10416 0 _0350_
rlabel metal2 41104 9688 41104 9688 0 _0351_
rlabel metal3 41216 5096 41216 5096 0 _0352_
rlabel metal3 40768 7672 40768 7672 0 _0353_
rlabel metal3 43736 9016 43736 9016 0 _0354_
rlabel metal3 42112 9128 42112 9128 0 _0355_
rlabel metal2 40264 9520 40264 9520 0 _0356_
rlabel metal2 41608 9184 41608 9184 0 _0357_
rlabel metal3 42896 8120 42896 8120 0 _0358_
rlabel metal2 40432 10472 40432 10472 0 _0359_
rlabel metal2 38024 10472 38024 10472 0 _0360_
rlabel metal2 38360 10976 38360 10976 0 _0361_
rlabel metal2 40936 10976 40936 10976 0 _0362_
rlabel metal2 41496 10752 41496 10752 0 _0363_
rlabel metal2 40936 9576 40936 9576 0 _0364_
rlabel metal3 41608 8232 41608 8232 0 _0365_
rlabel metal2 40152 8176 40152 8176 0 _0366_
rlabel metal2 40264 7616 40264 7616 0 _0367_
rlabel metal2 36008 15540 36008 15540 0 _0368_
rlabel metal2 35896 16800 35896 16800 0 _0369_
rlabel metal2 45080 12040 45080 12040 0 _0370_
rlabel metal2 43848 13608 43848 13608 0 _0371_
rlabel metal2 38248 14560 38248 14560 0 _0372_
rlabel metal2 32312 21504 32312 21504 0 _0373_
rlabel metal3 36680 14392 36680 14392 0 _0374_
rlabel metal2 38528 15288 38528 15288 0 _0375_
rlabel metal3 40208 14504 40208 14504 0 _0376_
rlabel metal2 40992 14392 40992 14392 0 _0377_
rlabel metal3 42840 13832 42840 13832 0 _0378_
rlabel metal2 42504 13272 42504 13272 0 _0379_
rlabel metal3 43680 13720 43680 13720 0 _0380_
rlabel metal2 44072 13328 44072 13328 0 _0381_
rlabel metal2 44520 14168 44520 14168 0 _0382_
rlabel metal3 44856 12936 44856 12936 0 _0383_
rlabel metal2 45920 12824 45920 12824 0 _0384_
rlabel metal2 29736 11256 29736 11256 0 _0385_
rlabel metal3 30856 11032 30856 11032 0 _0386_
rlabel metal2 44240 12152 44240 12152 0 _0387_
rlabel metal2 45080 11676 45080 11676 0 _0388_
rlabel metal3 45360 8344 45360 8344 0 _0389_
rlabel metal2 45808 11256 45808 11256 0 _0390_
rlabel metal2 23408 23464 23408 23464 0 _0391_
rlabel metal2 44184 8680 44184 8680 0 _0392_
rlabel metal2 44856 7952 44856 7952 0 _0393_
rlabel metal2 44744 7896 44744 7896 0 _0394_
rlabel metal2 45472 8344 45472 8344 0 _0395_
rlabel metal2 46032 8120 46032 8120 0 _0396_
rlabel metal2 45080 7168 45080 7168 0 _0397_
rlabel metal2 42392 6048 42392 6048 0 _0398_
rlabel metal2 45808 6552 45808 6552 0 _0399_
rlabel metal2 41944 5600 41944 5600 0 _0400_
rlabel metal2 42728 5544 42728 5544 0 _0401_
rlabel metal2 41272 5040 41272 5040 0 _0402_
rlabel metal3 43624 5208 43624 5208 0 _0403_
rlabel metal2 43960 4592 43960 4592 0 _0404_
rlabel metal2 42280 7392 42280 7392 0 _0405_
rlabel metal3 28224 21784 28224 21784 0 _0406_
rlabel metal2 27160 21560 27160 21560 0 _0407_
rlabel metal2 36344 22344 36344 22344 0 _0408_
rlabel metal3 37072 21448 37072 21448 0 _0409_
rlabel metal3 42056 20664 42056 20664 0 _0410_
rlabel metal2 42168 21392 42168 21392 0 _0411_
rlabel metal2 41832 22008 41832 22008 0 _0412_
rlabel metal3 42000 23128 42000 23128 0 _0413_
rlabel metal2 44072 24976 44072 24976 0 _0414_
rlabel metal2 44576 25368 44576 25368 0 _0415_
rlabel metal3 43512 25256 43512 25256 0 _0416_
rlabel metal2 44408 27552 44408 27552 0 _0417_
rlabel metal2 43848 27104 43848 27104 0 _0418_
rlabel metal2 43960 26544 43960 26544 0 _0419_
rlabel metal2 42168 26768 42168 26768 0 _0420_
rlabel metal3 43176 26376 43176 26376 0 _0421_
rlabel metal2 38808 29344 38808 29344 0 _0422_
rlabel metal2 39256 26992 39256 26992 0 _0423_
rlabel metal2 41832 26432 41832 26432 0 _0424_
rlabel metal2 39032 25816 39032 25816 0 _0425_
rlabel metal2 38024 25872 38024 25872 0 _0426_
rlabel metal2 39816 25536 39816 25536 0 _0427_
rlabel metal2 39480 24976 39480 24976 0 _0428_
rlabel metal2 38360 24360 38360 24360 0 _0429_
rlabel metal2 39816 24416 39816 24416 0 _0430_
rlabel metal2 40096 23912 40096 23912 0 _0431_
rlabel metal2 40712 25424 40712 25424 0 _0432_
rlabel metal2 41608 28616 41608 28616 0 _0433_
rlabel metal2 40376 28224 40376 28224 0 _0434_
rlabel metal2 43064 28000 43064 28000 0 _0435_
rlabel metal3 41496 26376 41496 26376 0 _0436_
rlabel metal2 41384 25872 41384 25872 0 _0437_
rlabel metal2 41104 25256 41104 25256 0 _0438_
rlabel metal2 46816 26264 46816 26264 0 _0439_
rlabel metal2 47768 26152 47768 26152 0 _0440_
rlabel metal2 47096 25984 47096 25984 0 _0441_
rlabel metal2 42056 25704 42056 25704 0 _0442_
rlabel metal2 43232 22344 43232 22344 0 _0443_
rlabel metal2 42952 24136 42952 24136 0 _0444_
rlabel metal3 42112 24808 42112 24808 0 _0445_
rlabel metal2 42616 25144 42616 25144 0 _0446_
rlabel metal2 42280 24304 42280 24304 0 _0447_
rlabel metal2 47208 20104 47208 20104 0 _0448_
rlabel metal3 44408 19208 44408 19208 0 _0449_
rlabel metal2 41328 20216 41328 20216 0 _0450_
rlabel metal2 42224 19992 42224 19992 0 _0451_
rlabel metal2 42616 19656 42616 19656 0 _0452_
rlabel metal3 42224 18984 42224 18984 0 _0453_
rlabel metal2 41832 21168 41832 21168 0 _0454_
rlabel metal3 42392 23352 42392 23352 0 _0455_
rlabel metal2 42392 22624 42392 22624 0 _0456_
rlabel metal2 42504 20440 42504 20440 0 _0457_
rlabel metal2 41664 23128 41664 23128 0 _0458_
rlabel metal2 41944 23632 41944 23632 0 _0459_
rlabel metal2 41776 23352 41776 23352 0 _0460_
rlabel metal2 41272 24976 41272 24976 0 _0461_
rlabel metal2 41328 22344 41328 22344 0 _0462_
rlabel metal2 35672 22624 35672 22624 0 _0463_
rlabel metal2 39144 22400 39144 22400 0 _0464_
rlabel metal2 45528 21672 45528 21672 0 _0465_
rlabel metal2 38360 21504 38360 21504 0 _0466_
rlabel metal2 43400 18088 43400 18088 0 _0467_
rlabel metal2 37800 24136 37800 24136 0 _0468_
rlabel metal2 36904 23072 36904 23072 0 _0469_
rlabel metal2 39816 26600 39816 26600 0 _0470_
rlabel metal2 41048 27384 41048 27384 0 _0471_
rlabel metal2 38360 27160 38360 27160 0 _0472_
rlabel metal2 46088 24024 46088 24024 0 _0473_
rlabel metal2 39424 29288 39424 29288 0 _0474_
rlabel metal2 43120 29400 43120 29400 0 _0475_
rlabel metal2 45752 29064 45752 29064 0 _0476_
rlabel metal3 44240 28616 44240 28616 0 _0477_
rlabel metal3 45248 28392 45248 28392 0 _0478_
rlabel metal2 44856 26544 44856 26544 0 _0479_
rlabel metal2 45696 24584 45696 24584 0 _0480_
rlabel metal3 45192 22904 45192 22904 0 _0481_
rlabel metal2 45864 23072 45864 23072 0 _0482_
rlabel metal3 46536 21448 46536 21448 0 _0483_
rlabel metal2 45024 21560 45024 21560 0 _0484_
rlabel metal2 47880 21392 47880 21392 0 _0485_
rlabel metal3 45472 21672 45472 21672 0 _0486_
rlabel metal2 43736 18144 43736 18144 0 _0487_
rlabel metal3 45808 21560 45808 21560 0 _0488_
rlabel metal2 31752 21952 31752 21952 0 _0489_
rlabel metal2 32592 21784 32592 21784 0 _0490_
rlabel metal2 18312 39200 18312 39200 0 _0491_
rlabel metal3 16072 37128 16072 37128 0 _0492_
rlabel metal2 13160 40544 13160 40544 0 _0493_
rlabel metal2 22736 39368 22736 39368 0 _0494_
rlabel metal2 22456 39928 22456 39928 0 _0495_
rlabel metal2 14056 43400 14056 43400 0 _0496_
rlabel metal3 20832 42840 20832 42840 0 _0497_
rlabel metal2 19880 41440 19880 41440 0 _0498_
rlabel metal2 18200 39144 18200 39144 0 _0499_
rlabel metal2 19824 36680 19824 36680 0 _0500_
rlabel metal2 19488 37464 19488 37464 0 _0501_
rlabel metal2 18200 36232 18200 36232 0 _0502_
rlabel metal2 18536 38528 18536 38528 0 _0503_
rlabel metal2 18760 40880 18760 40880 0 _0504_
rlabel metal2 18816 42056 18816 42056 0 _0505_
rlabel metal2 19656 42280 19656 42280 0 _0506_
rlabel metal3 20048 41944 20048 41944 0 _0507_
rlabel metal2 20552 44184 20552 44184 0 _0508_
rlabel metal2 18536 43680 18536 43680 0 _0509_
rlabel metal2 17528 45584 17528 45584 0 _0510_
rlabel metal2 19712 45080 19712 45080 0 _0511_
rlabel metal3 19936 45080 19936 45080 0 _0512_
rlabel metal2 22008 44352 22008 44352 0 _0513_
rlabel metal2 12152 43568 12152 43568 0 _0514_
rlabel metal2 22680 43232 22680 43232 0 _0515_
rlabel metal3 23128 42952 23128 42952 0 _0516_
rlabel metal2 23240 41888 23240 41888 0 _0517_
rlabel metal2 20664 40768 20664 40768 0 _0518_
rlabel metal2 22568 38976 22568 38976 0 _0519_
rlabel metal2 12936 39144 12936 39144 0 _0520_
rlabel metal3 20720 38808 20720 38808 0 _0521_
rlabel metal3 22736 38808 22736 38808 0 _0522_
rlabel metal2 21616 38024 21616 38024 0 _0523_
rlabel metal2 14504 40040 14504 40040 0 _0524_
rlabel metal2 10864 41720 10864 41720 0 _0525_
rlabel metal2 14840 37184 14840 37184 0 _0526_
rlabel metal2 16688 40152 16688 40152 0 _0527_
rlabel metal2 19656 38416 19656 38416 0 _0528_
rlabel metal3 19320 38024 19320 38024 0 _0529_
rlabel metal2 20328 38248 20328 38248 0 _0530_
rlabel metal2 17976 41720 17976 41720 0 _0531_
rlabel metal2 16296 41104 16296 41104 0 _0532_
rlabel metal2 13832 42112 13832 42112 0 _0533_
rlabel metal3 14784 41944 14784 41944 0 _0534_
rlabel metal2 16856 43288 16856 43288 0 _0535_
rlabel metal3 15680 43736 15680 43736 0 _0536_
rlabel metal2 14392 44184 14392 44184 0 _0537_
rlabel metal2 15288 44408 15288 44408 0 _0538_
rlabel metal2 13216 44184 13216 44184 0 _0539_
rlabel metal3 10416 43624 10416 43624 0 _0540_
rlabel metal2 11144 44660 11144 44660 0 _0541_
rlabel metal2 12376 43344 12376 43344 0 _0542_
rlabel metal2 10248 41944 10248 41944 0 _0543_
rlabel metal2 11816 41776 11816 41776 0 _0544_
rlabel metal3 10864 41832 10864 41832 0 _0545_
rlabel metal3 13216 41048 13216 41048 0 _0546_
rlabel metal2 12488 39424 12488 39424 0 _0547_
rlabel metal2 22120 28672 22120 28672 0 _0548_
rlabel metal2 22120 21448 22120 21448 0 _0549_
rlabel metal2 21672 23016 21672 23016 0 _0550_
rlabel metal2 20888 20552 20888 20552 0 _0551_
rlabel metal2 20776 19880 20776 19880 0 _0552_
rlabel metal2 12712 28728 12712 28728 0 _0553_
rlabel metal3 14168 29960 14168 29960 0 _0554_
rlabel metal2 12376 29456 12376 29456 0 _0555_
rlabel metal2 14392 27384 14392 27384 0 _0556_
rlabel metal2 15288 23240 15288 23240 0 _0557_
rlabel metal3 14224 23240 14224 23240 0 _0558_
rlabel metal2 13944 16408 13944 16408 0 _0559_
rlabel metal3 14112 22904 14112 22904 0 _0560_
rlabel metal2 16632 20272 16632 20272 0 _0561_
rlabel metal2 14280 21728 14280 21728 0 _0562_
rlabel metal2 16296 20272 16296 20272 0 _0563_
rlabel metal2 14728 21112 14728 21112 0 _0564_
rlabel metal3 14336 19096 14336 19096 0 _0565_
rlabel metal2 30408 32928 30408 32928 0 _0566_
rlabel metal2 26152 32536 26152 32536 0 _0567_
rlabel metal3 24640 31192 24640 31192 0 _0568_
rlabel metal2 25592 30520 25592 30520 0 _0569_
rlabel metal2 25480 30464 25480 30464 0 _0570_
rlabel metal2 26264 32760 26264 32760 0 _0571_
rlabel metal2 27272 30520 27272 30520 0 _0572_
rlabel metal2 26768 30184 26768 30184 0 _0573_
rlabel metal2 27048 31752 27048 31752 0 _0574_
rlabel metal2 26040 32200 26040 32200 0 _0575_
rlabel metal2 32368 33208 32368 33208 0 _0576_
rlabel metal2 29848 34776 29848 34776 0 _0577_
rlabel metal2 31752 35504 31752 35504 0 _0578_
rlabel metal2 30856 35840 30856 35840 0 _0579_
rlabel metal3 28280 33432 28280 33432 0 _0580_
rlabel metal2 28280 36008 28280 36008 0 _0581_
rlabel metal2 30072 36176 30072 36176 0 _0582_
rlabel metal2 29288 35336 29288 35336 0 _0583_
rlabel metal3 34160 37240 34160 37240 0 _0584_
rlabel metal2 33544 35896 33544 35896 0 _0585_
rlabel metal2 34776 32704 34776 32704 0 _0586_
rlabel metal3 35392 34328 35392 34328 0 _0587_
rlabel metal3 33544 37128 33544 37128 0 _0588_
rlabel metal2 34888 37688 34888 37688 0 _0589_
rlabel metal2 16240 18200 16240 18200 0 _0590_
rlabel metal2 16184 16912 16184 16912 0 _0591_
rlabel via2 10808 16184 10808 16184 0 _0592_
rlabel metal2 10920 14112 10920 14112 0 _0593_
rlabel metal3 11592 16744 11592 16744 0 _0594_
rlabel metal3 9240 16296 9240 16296 0 _0595_
rlabel metal2 9688 17192 9688 17192 0 _0596_
rlabel metal2 10696 15680 10696 15680 0 _0597_
rlabel metal3 10080 15176 10080 15176 0 _0598_
rlabel metal2 12376 14392 12376 14392 0 _0599_
rlabel metal2 14784 14392 14784 14392 0 _0600_
rlabel metal2 11816 13832 11816 13832 0 _0601_
rlabel metal2 14896 14616 14896 14616 0 _0602_
rlabel metal2 13720 13664 13720 13664 0 _0603_
rlabel metal2 14672 12824 14672 12824 0 _0604_
rlabel metal2 14952 12768 14952 12768 0 _0605_
rlabel metal2 24472 22344 24472 22344 0 _0606_
rlabel metal2 23128 22064 23128 22064 0 _0607_
rlabel metal2 16856 22736 16856 22736 0 _0608_
rlabel metal3 20720 17528 20720 17528 0 _0609_
rlabel metal3 23688 20664 23688 20664 0 _0610_
rlabel metal2 23352 22344 23352 22344 0 _0611_
rlabel metal2 25368 21784 25368 21784 0 _0612_
rlabel metal2 25144 21896 25144 21896 0 _0613_
rlabel metal2 19768 20608 19768 20608 0 _0614_
rlabel metal2 21224 16184 21224 16184 0 _0615_
rlabel metal3 22008 26824 22008 26824 0 _0616_
rlabel metal3 21504 26264 21504 26264 0 _0617_
rlabel metal2 19992 18368 19992 18368 0 _0618_
rlabel metal2 17528 23072 17528 23072 0 _0619_
rlabel metal2 28056 23408 28056 23408 0 _0620_
rlabel metal2 19544 25424 19544 25424 0 _0621_
rlabel metal3 19824 17640 19824 17640 0 _0622_
rlabel metal2 18088 16632 18088 16632 0 _0623_
rlabel metal2 21336 16968 21336 16968 0 _0624_
rlabel metal2 16296 17192 16296 17192 0 _0625_
rlabel metal2 19096 16352 19096 16352 0 _0626_
rlabel metal2 19824 16856 19824 16856 0 _0627_
rlabel metal3 22232 15848 22232 15848 0 _0628_
rlabel metal2 30128 21784 30128 21784 0 _0629_
rlabel metal2 33544 10920 33544 10920 0 _0630_
rlabel metal2 30856 30184 30856 30184 0 _0631_
rlabel metal2 30408 27216 30408 27216 0 _0632_
rlabel metal2 28504 28336 28504 28336 0 _0633_
rlabel metal3 24976 32536 24976 32536 0 _0634_
rlabel metal2 27944 30464 27944 30464 0 _0635_
rlabel metal3 25872 23352 25872 23352 0 _0636_
rlabel metal2 31080 20104 31080 20104 0 _0637_
rlabel metal2 31528 16968 31528 16968 0 _0638_
rlabel metal2 23240 19208 23240 19208 0 _0639_
rlabel metal3 25144 25312 25144 25312 0 _0640_
rlabel metal3 30464 18984 30464 18984 0 _0641_
rlabel metal2 31080 17136 31080 17136 0 _0642_
rlabel metal3 31584 16968 31584 16968 0 _0643_
rlabel metal3 32592 15400 32592 15400 0 _0644_
rlabel metal2 31640 16296 31640 16296 0 _0645_
rlabel metal2 38696 7336 38696 7336 0 _0646_
rlabel metal3 32088 13608 32088 13608 0 _0647_
rlabel metal3 34888 18536 34888 18536 0 _0648_
rlabel metal2 30408 12208 30408 12208 0 _0649_
rlabel metal2 38696 31528 38696 31528 0 _0650_
rlabel metal2 25480 41216 25480 41216 0 _0651_
rlabel metal2 29176 19152 29176 19152 0 _0652_
rlabel metal2 26264 29848 26264 29848 0 _0653_
rlabel metal3 28784 28504 28784 28504 0 _0654_
rlabel metal3 31864 23184 31864 23184 0 _0655_
rlabel metal3 32760 9016 32760 9016 0 _0656_
rlabel metal3 35168 5096 35168 5096 0 _0657_
rlabel metal3 20216 18648 20216 18648 0 _0658_
rlabel metal2 22008 15652 22008 15652 0 _0659_
rlabel metal2 35112 8568 35112 8568 0 _0660_
rlabel metal2 32536 7784 32536 7784 0 _0661_
rlabel metal3 33544 5768 33544 5768 0 _0662_
rlabel metal2 35896 5824 35896 5824 0 _0663_
rlabel metal2 33544 4816 33544 4816 0 _0664_
rlabel metal2 24248 21280 24248 21280 0 _0665_
rlabel metal3 19320 22120 19320 22120 0 _0666_
rlabel metal2 24248 30576 24248 30576 0 _0667_
rlabel metal2 24360 31248 24360 31248 0 _0668_
rlabel metal2 22792 35616 22792 35616 0 _0669_
rlabel metal3 19544 38696 19544 38696 0 _0670_
rlabel metal2 23800 17696 23800 17696 0 _0671_
rlabel metal2 24304 35672 24304 35672 0 _0672_
rlabel metal2 22960 33320 22960 33320 0 _0673_
rlabel metal2 24584 27496 24584 27496 0 _0674_
rlabel metal2 25368 35280 25368 35280 0 _0675_
rlabel metal2 21336 40320 21336 40320 0 _0676_
rlabel metal2 26600 31248 26600 31248 0 _0677_
rlabel metal2 25032 35672 25032 35672 0 _0678_
rlabel metal2 12712 13776 12712 13776 0 _0679_
rlabel metal2 11704 13104 11704 13104 0 _0680_
rlabel metal2 12152 13608 12152 13608 0 _0681_
rlabel metal3 21224 36456 21224 36456 0 _0682_
rlabel metal2 26824 32704 26824 32704 0 _0683_
rlabel metal3 23520 35112 23520 35112 0 _0684_
rlabel metal2 22456 35280 22456 35280 0 _0685_
rlabel metal2 24024 36512 24024 36512 0 _0686_
rlabel metal3 23520 35672 23520 35672 0 _0687_
rlabel metal2 23240 16856 23240 16856 0 _0688_
rlabel metal3 7448 13048 7448 13048 0 _0689_
rlabel metal2 19432 16408 19432 16408 0 _0690_
rlabel metal3 19040 15400 19040 15400 0 _0691_
rlabel metal2 20664 15960 20664 15960 0 _0692_
rlabel metal3 20272 15176 20272 15176 0 _0693_
rlabel metal2 18760 13272 18760 13272 0 _0694_
rlabel metal2 19040 13832 19040 13832 0 _0695_
rlabel metal2 18424 14168 18424 14168 0 _0696_
rlabel metal3 21000 10808 21000 10808 0 _0697_
rlabel metal3 6216 16072 6216 16072 0 _0698_
rlabel metal2 13832 12656 13832 12656 0 _0699_
rlabel metal2 17920 12936 17920 12936 0 _0700_
rlabel metal2 21280 10584 21280 10584 0 _0701_
rlabel metal2 17640 12488 17640 12488 0 _0702_
rlabel metal3 17248 11368 17248 11368 0 _0703_
rlabel metal3 11648 11368 11648 11368 0 _0704_
rlabel metal2 17192 12152 17192 12152 0 _0705_
rlabel metal2 10920 11480 10920 11480 0 _0706_
rlabel metal2 6328 12656 6328 12656 0 _0707_
rlabel metal2 10136 10752 10136 10752 0 _0708_
rlabel metal2 12488 10192 12488 10192 0 _0709_
rlabel metal3 13328 8232 13328 8232 0 _0710_
rlabel metal2 12600 7336 12600 7336 0 _0711_
rlabel metal3 11928 11256 11928 11256 0 _0712_
rlabel metal2 12152 10024 12152 10024 0 _0713_
rlabel metal2 10752 9240 10752 9240 0 _0714_
rlabel metal2 8680 6608 8680 6608 0 _0715_
rlabel metal3 12880 8456 12880 8456 0 _0716_
rlabel metal2 9016 7840 9016 7840 0 _0717_
rlabel metal2 12824 11872 12824 11872 0 _0718_
rlabel metal2 8120 7140 8120 7140 0 _0719_
rlabel metal2 13048 7168 13048 7168 0 _0720_
rlabel via2 29624 6440 29624 6440 0 _0721_
rlabel metal2 24584 7056 24584 7056 0 _0722_
rlabel metal2 29512 4424 29512 4424 0 _0723_
rlabel metal2 23800 5040 23800 5040 0 _0724_
rlabel metal2 23576 5152 23576 5152 0 _0725_
rlabel metal2 22792 8904 22792 8904 0 _0726_
rlabel metal2 22568 7896 22568 7896 0 _0727_
rlabel metal2 25592 8064 25592 8064 0 _0728_
rlabel metal2 23800 8288 23800 8288 0 _0729_
rlabel metal2 24360 6944 24360 6944 0 _0730_
rlabel metal2 23240 7896 23240 7896 0 _0731_
rlabel metal3 18480 24920 18480 24920 0 _0732_
rlabel metal3 16520 21392 16520 21392 0 _0733_
rlabel metal2 17864 7952 17864 7952 0 _0734_
rlabel metal2 25256 5208 25256 5208 0 _0735_
rlabel metal2 22008 5488 22008 5488 0 _0736_
rlabel metal3 20328 8344 20328 8344 0 _0737_
rlabel metal2 18760 8960 18760 8960 0 _0738_
rlabel metal2 20216 8288 20216 8288 0 _0739_
rlabel metal3 18088 8008 18088 8008 0 _0740_
rlabel metal2 16968 6272 16968 6272 0 _0741_
rlabel metal2 16744 8288 16744 8288 0 _0742_
rlabel metal2 15064 5488 15064 5488 0 _0743_
rlabel metal2 16464 5992 16464 5992 0 _0744_
rlabel metal2 15512 5208 15512 5208 0 _0745_
rlabel metal2 17304 3808 17304 3808 0 _0746_
rlabel metal2 20440 5432 20440 5432 0 _0747_
rlabel metal2 17192 21672 17192 21672 0 _0748_
rlabel metal2 16744 21840 16744 21840 0 _0749_
rlabel metal3 10136 20552 10136 20552 0 _0750_
rlabel metal2 9968 20216 9968 20216 0 _0751_
rlabel metal3 4704 14504 4704 14504 0 _0752_
rlabel metal2 4872 14756 4872 14756 0 _0753_
rlabel metal2 4536 18760 4536 18760 0 _0754_
rlabel metal2 5096 12320 5096 12320 0 _0755_
rlabel via2 4312 12824 4312 12824 0 _0756_
rlabel metal2 4088 13328 4088 13328 0 _0757_
rlabel metal2 4872 12040 4872 12040 0 _0758_
rlabel metal2 5320 12656 5320 12656 0 _0759_
rlabel metal2 6440 11648 6440 11648 0 _0760_
rlabel metal2 6664 9800 6664 9800 0 _0761_
rlabel metal2 8624 4424 8624 4424 0 _0762_
rlabel metal2 28056 28896 28056 28896 0 _0763_
rlabel metal2 40264 15680 40264 15680 0 _0764_
rlabel metal2 34440 12656 34440 12656 0 _0765_
rlabel metal3 22792 18424 22792 18424 0 _0766_
rlabel metal2 33992 17920 33992 17920 0 _0767_
rlabel metal2 35112 15260 35112 15260 0 _0768_
rlabel metal2 32536 10752 32536 10752 0 _0769_
rlabel metal2 34384 13048 34384 13048 0 _0770_
rlabel metal2 35112 10528 35112 10528 0 _0771_
rlabel metal2 35224 9184 35224 9184 0 _0772_
rlabel metal2 40600 16408 40600 16408 0 _0773_
rlabel via2 41384 16632 41384 16632 0 _0774_
rlabel metal3 40656 16744 40656 16744 0 _0775_
rlabel metal2 42448 25592 42448 25592 0 _0776_
rlabel metal3 43792 16296 43792 16296 0 _0777_
rlabel metal3 26040 45080 26040 45080 0 _0778_
rlabel metal2 46648 16324 46648 16324 0 _0779_
rlabel metal3 26040 43512 26040 43512 0 _0780_
rlabel metal2 45976 17752 45976 17752 0 _0781_
rlabel metal2 31920 27832 31920 27832 0 _0782_
rlabel metal2 32984 23128 32984 23128 0 _0783_
rlabel metal2 35224 18704 35224 18704 0 _0784_
rlabel metal2 35616 18648 35616 18648 0 _0785_
rlabel metal2 35000 21560 35000 21560 0 _0786_
rlabel metal3 32984 19880 32984 19880 0 _0787_
rlabel metal2 36232 19152 36232 19152 0 _0788_
rlabel metal2 35560 18368 35560 18368 0 _0789_
rlabel metal2 20664 28784 20664 28784 0 _0790_
rlabel metal3 34440 30072 34440 30072 0 _0791_
rlabel metal2 33376 29400 33376 29400 0 _0792_
rlabel metal2 34776 30856 34776 30856 0 _0793_
rlabel metal2 33880 29792 33880 29792 0 _0794_
rlabel metal2 32760 27216 32760 27216 0 _0795_
rlabel metal3 19040 26376 19040 26376 0 _0796_
rlabel metal2 33432 25592 33432 25592 0 _0797_
rlabel metal2 20104 33824 20104 33824 0 _0798_
rlabel metal2 33992 27216 33992 27216 0 _0799_
rlabel metal2 18872 28784 18872 28784 0 _0800_
rlabel metal2 35056 28616 35056 28616 0 _0801_
rlabel metal2 40936 30688 40936 30688 0 _0802_
rlabel metal2 41384 31360 41384 31360 0 _0803_
rlabel metal3 41664 30856 41664 30856 0 _0804_
rlabel metal3 45304 31192 45304 31192 0 _0805_
rlabel metal3 46032 31640 46032 31640 0 _0806_
rlabel metal2 43176 31416 43176 31416 0 _0807_
rlabel metal2 25704 4200 25704 4200 0 _0808_
rlabel metal2 26264 9016 26264 9016 0 _0809_
rlabel metal2 26488 5880 26488 5880 0 _0810_
rlabel metal2 23352 21840 23352 21840 0 _0811_
rlabel metal2 25368 9856 25368 9856 0 _0812_
rlabel metal3 28560 8344 28560 8344 0 _0813_
rlabel metal2 27496 7448 27496 7448 0 _0814_
rlabel metal2 26768 5992 26768 5992 0 _0815_
rlabel metal2 29288 7056 29288 7056 0 _0816_
rlabel metal2 3864 14924 3864 14924 0 _0817_
rlabel metal2 3640 16688 3640 16688 0 _0818_
rlabel metal2 3416 14728 3416 14728 0 _0819_
rlabel metal3 3640 16072 3640 16072 0 _0820_
rlabel metal2 3584 7672 3584 7672 0 _0821_
rlabel metal2 5096 7112 5096 7112 0 _0822_
rlabel metal2 3528 10136 3528 10136 0 _0823_
rlabel metal3 4256 7448 4256 7448 0 _0824_
rlabel metal2 3416 7224 3416 7224 0 _0825_
rlabel metal2 4760 6328 4760 6328 0 _0826_
rlabel metal2 7224 6160 7224 6160 0 _0827_
rlabel metal2 5040 5992 5040 5992 0 _0828_
rlabel metal2 7896 6384 7896 6384 0 _0829_
rlabel metal2 7112 6664 7112 6664 0 _0830_
rlabel metal2 7784 3472 7784 3472 0 _0831_
rlabel metal2 6216 5432 6216 5432 0 _0832_
rlabel metal2 7448 3864 7448 3864 0 _0833_
rlabel metal2 7448 5040 7448 5040 0 _0834_
rlabel metal2 32200 30016 32200 30016 0 _0835_
rlabel metal2 24360 24920 24360 24920 0 _0836_
rlabel metal3 23240 24472 23240 24472 0 _0837_
rlabel metal3 22120 25704 22120 25704 0 _0838_
rlabel metal2 25256 26320 25256 26320 0 _0839_
rlabel metal3 24584 23912 24584 23912 0 _0840_
rlabel metal2 21336 24696 21336 24696 0 _0841_
rlabel metal2 23800 35168 23800 35168 0 _0842_
rlabel metal2 18648 32088 18648 32088 0 _0843_
rlabel metal2 20552 39368 20552 39368 0 _0844_
rlabel metal2 19208 33656 19208 33656 0 _0845_
rlabel metal2 16520 34440 16520 34440 0 _0846_
rlabel metal2 17584 32424 17584 32424 0 _0847_
rlabel metal2 19376 34328 19376 34328 0 _0848_
rlabel metal3 19544 31080 19544 31080 0 _0849_
rlabel metal2 25816 44408 25816 44408 0 _0850_
rlabel metal3 23016 40376 23016 40376 0 _0851_
rlabel metal2 24360 40208 24360 40208 0 _0852_
rlabel metal3 22456 43400 22456 43400 0 _0853_
rlabel metal3 25088 44968 25088 44968 0 _0854_
rlabel metal2 24584 42000 24584 42000 0 _0855_
rlabel metal2 23576 18760 23576 18760 0 _0856_
rlabel metal2 24472 15960 24472 15960 0 _0857_
rlabel metal2 22344 5376 22344 5376 0 _0858_
rlabel metal3 23632 3752 23632 3752 0 _0859_
rlabel metal2 6552 14532 6552 14532 0 _0860_
rlabel metal2 28056 26264 28056 26264 0 _0861_
rlabel metal3 17472 26600 17472 26600 0 _0862_
rlabel metal2 27272 23968 27272 23968 0 _0863_
rlabel metal3 17864 26488 17864 26488 0 _0864_
rlabel metal2 19656 28784 19656 28784 0 _0865_
rlabel metal2 16744 25144 16744 25144 0 _0866_
rlabel metal2 25704 27440 25704 27440 0 _0867_
rlabel metal3 18256 27720 18256 27720 0 _0868_
rlabel metal3 29008 23800 29008 23800 0 _0869_
rlabel metal2 25816 23464 25816 23464 0 _0870_
rlabel metal3 40488 34216 40488 34216 0 _0871_
rlabel metal2 37800 35168 37800 35168 0 _0872_
rlabel metal2 46088 32368 46088 32368 0 _0873_
rlabel metal3 38920 33208 38920 33208 0 _0874_
rlabel metal2 39760 38808 39760 38808 0 _0875_
rlabel metal2 44072 33880 44072 33880 0 _0876_
rlabel metal2 37464 36344 37464 36344 0 _0877_
rlabel metal2 41272 39200 41272 39200 0 _0878_
rlabel metal3 36680 35112 36680 35112 0 _0879_
rlabel metal3 42504 38584 42504 38584 0 _0880_
rlabel metal3 46200 35448 46200 35448 0 _0881_
rlabel metal2 38584 35616 38584 35616 0 _0882_
rlabel metal2 39760 32760 39760 32760 0 _0883_
rlabel metal2 45528 11256 45528 11256 0 _0884_
rlabel metal3 45864 36232 45864 36232 0 _0885_
rlabel metal2 44184 34160 44184 34160 0 _0886_
rlabel metal2 47544 36960 47544 36960 0 _0887_
rlabel metal2 45752 32480 45752 32480 0 _0888_
rlabel metal3 46480 38808 46480 38808 0 _0889_
rlabel metal2 48104 33880 48104 33880 0 _0890_
rlabel metal2 15176 29120 15176 29120 0 _0891_
rlabel metal2 2352 34776 2352 34776 0 _0892_
rlabel metal2 9688 38780 9688 38780 0 _0893_
rlabel metal2 7336 36176 7336 36176 0 _0894_
rlabel metal3 10752 34888 10752 34888 0 _0895_
rlabel metal2 9016 36120 9016 36120 0 _0896_
rlabel metal2 6888 36008 6888 36008 0 _0897_
rlabel metal2 3248 35672 3248 35672 0 _0898_
rlabel metal2 12376 39088 12376 39088 0 _0899_
rlabel metal3 3136 38808 3136 38808 0 _0900_
rlabel metal2 2184 34944 2184 34944 0 _0901_
rlabel metal3 10920 38136 10920 38136 0 _0902_
rlabel metal2 3192 37240 3192 37240 0 _0903_
rlabel metal2 3304 36456 3304 36456 0 _0904_
rlabel metal2 3696 39480 3696 39480 0 _0905_
rlabel metal2 4480 39704 4480 39704 0 _0906_
rlabel metal2 3248 39368 3248 39368 0 _0907_
rlabel metal2 4536 39424 4536 39424 0 _0908_
rlabel metal2 3024 37912 3024 37912 0 _0909_
rlabel metal2 6664 35168 6664 35168 0 _0910_
rlabel metal3 6832 35896 6832 35896 0 _0911_
rlabel metal3 40320 44856 40320 44856 0 _0912_
rlabel metal2 35448 43904 35448 43904 0 _0913_
rlabel metal2 36736 39480 36736 39480 0 _0914_
rlabel metal2 36064 39704 36064 39704 0 _0915_
rlabel metal2 35896 39928 35896 39928 0 _0916_
rlabel metal2 34328 40432 34328 40432 0 _0917_
rlabel metal2 33768 41328 33768 41328 0 _0918_
rlabel metal2 33096 41664 33096 41664 0 _0919_
rlabel metal2 33320 41440 33320 41440 0 _0920_
rlabel metal2 33824 40488 33824 40488 0 _0921_
rlabel metal2 31192 43176 31192 43176 0 _0922_
rlabel metal3 32312 40936 32312 40936 0 _0923_
rlabel metal2 30520 38920 30520 38920 0 _0924_
rlabel metal2 30800 41384 30800 41384 0 _0925_
rlabel metal2 31640 40656 31640 40656 0 _0926_
rlabel metal2 29680 38920 29680 38920 0 _0927_
rlabel metal2 31752 38864 31752 38864 0 _0928_
rlabel metal2 26096 38808 26096 38808 0 _0929_
rlabel metal2 30184 39508 30184 39508 0 _0930_
rlabel metal2 30520 40656 30520 40656 0 _0931_
rlabel metal2 32704 41160 32704 41160 0 _0932_
rlabel metal2 32256 40488 32256 40488 0 _0933_
rlabel metal3 32592 40376 32592 40376 0 _0934_
rlabel metal2 34104 39984 34104 39984 0 _0935_
rlabel metal2 36120 39088 36120 39088 0 _0936_
rlabel metal2 38136 38752 38136 38752 0 _0937_
rlabel metal2 44800 42504 44800 42504 0 _0938_
rlabel metal2 43344 36456 43344 36456 0 _0939_
rlabel metal2 43064 37016 43064 37016 0 _0940_
rlabel metal2 42616 39116 42616 39116 0 _0941_
rlabel metal2 40712 40712 40712 40712 0 _0942_
rlabel metal2 40152 38668 40152 38668 0 _0943_
rlabel metal3 39872 43736 39872 43736 0 _0944_
rlabel metal2 41720 39648 41720 39648 0 _0945_
rlabel metal2 43960 37688 43960 37688 0 _0946_
rlabel metal2 47768 39648 47768 39648 0 _0947_
rlabel metal2 46648 39928 46648 39928 0 _0948_
rlabel metal2 44968 38864 44968 38864 0 _0949_
rlabel metal2 44184 39088 44184 39088 0 _0950_
rlabel metal2 46984 35616 46984 35616 0 _0951_
rlabel metal2 45136 38920 45136 38920 0 _0952_
rlabel metal3 44744 38808 44744 38808 0 _0953_
rlabel metal2 44464 38584 44464 38584 0 _0954_
rlabel metal2 42672 37464 42672 37464 0 _0955_
rlabel metal2 37184 38808 37184 38808 0 _0956_
rlabel metal2 37688 38808 37688 38808 0 _0957_
rlabel metal2 39816 39256 39816 39256 0 _0958_
rlabel metal3 42952 39368 42952 39368 0 _0959_
rlabel metal2 44016 39480 44016 39480 0 _0960_
rlabel metal2 46424 39144 46424 39144 0 _0961_
rlabel metal2 46760 39144 46760 39144 0 _0962_
rlabel metal3 35896 38808 35896 38808 0 _0963_
rlabel metal2 32088 39984 32088 39984 0 _0964_
rlabel metal2 31304 39592 31304 39592 0 _0965_
rlabel metal2 29176 39872 29176 39872 0 _0966_
rlabel metal2 31976 39648 31976 39648 0 _0967_
rlabel metal3 35336 39480 35336 39480 0 _0968_
rlabel metal2 30912 39368 30912 39368 0 _0969_
rlabel metal2 32424 39144 32424 39144 0 _0970_
rlabel metal2 32312 39088 32312 39088 0 _0971_
rlabel metal2 32872 39480 32872 39480 0 _0972_
rlabel metal2 33096 39088 33096 39088 0 _0973_
rlabel metal2 45976 43232 45976 43232 0 _0974_
rlabel metal2 26712 35504 26712 35504 0 _0975_
rlabel metal2 27272 39200 27272 39200 0 _0976_
rlabel metal3 22512 21336 22512 21336 0 _0977_
rlabel metal2 27720 39256 27720 39256 0 _0978_
rlabel metal2 19544 39704 19544 39704 0 _0979_
rlabel metal2 33936 15848 33936 15848 0 _0980_
rlabel metal2 24472 38920 24472 38920 0 _0981_
rlabel metal2 11032 38920 11032 38920 0 _0982_
rlabel metal2 10416 39592 10416 39592 0 _0983_
rlabel metal2 8904 38752 8904 38752 0 _0984_
rlabel metal2 10136 39144 10136 39144 0 _0985_
rlabel metal2 25816 17696 25816 17696 0 _0986_
rlabel metal3 24696 38696 24696 38696 0 _0987_
rlabel metal2 33992 42896 33992 42896 0 _0988_
rlabel metal2 47656 45528 47656 45528 0 _0989_
rlabel metal2 34776 15232 34776 15232 0 _0990_
rlabel metal2 28448 19992 28448 19992 0 _0991_
rlabel metal2 27720 41160 27720 41160 0 _0992_
rlabel metal2 26824 41384 26824 41384 0 _0993_
rlabel metal2 29512 42000 29512 42000 0 _0994_
rlabel metal2 31416 43120 31416 43120 0 _0995_
rlabel metal3 31752 44520 31752 44520 0 _0996_
rlabel metal2 33152 43736 33152 43736 0 _0997_
rlabel metal3 33040 45080 33040 45080 0 _0998_
rlabel metal2 31472 45080 31472 45080 0 _0999_
rlabel metal3 33208 45304 33208 45304 0 _1000_
rlabel metal2 33880 44744 33880 44744 0 _1001_
rlabel metal3 32816 44296 32816 44296 0 _1002_
rlabel metal3 37800 44296 37800 44296 0 _1003_
rlabel metal2 37128 43904 37128 43904 0 _1004_
rlabel metal2 35000 43456 35000 43456 0 _1005_
rlabel metal3 47208 42952 47208 42952 0 _1006_
rlabel metal2 46536 45584 46536 45584 0 _1007_
rlabel metal2 37968 44408 37968 44408 0 _1008_
rlabel metal3 40936 43848 40936 43848 0 _1009_
rlabel metal3 41328 43624 41328 43624 0 _1010_
rlabel metal2 39424 44184 39424 44184 0 _1011_
rlabel metal2 39368 42896 39368 42896 0 _1012_
rlabel metal2 40936 41664 40936 41664 0 _1013_
rlabel metal2 38808 40712 38808 40712 0 _1014_
rlabel metal2 40712 42616 40712 42616 0 _1015_
rlabel metal2 40712 41664 40712 41664 0 _1016_
rlabel metal2 41160 43708 41160 43708 0 _1017_
rlabel metal3 42056 41720 42056 41720 0 _1018_
rlabel metal2 40320 44184 40320 44184 0 _1019_
rlabel metal2 45752 43120 45752 43120 0 _1020_
rlabel metal2 44464 43400 44464 43400 0 _1021_
rlabel metal2 46760 42616 46760 42616 0 _1022_
rlabel metal2 46256 42504 46256 42504 0 _1023_
rlabel metal3 22848 19992 22848 19992 0 clknet_0_wb_clk_i
rlabel metal2 11200 7000 11200 7000 0 clknet_2_0__leaf_wb_clk_i
rlabel metal2 11368 40656 11368 40656 0 clknet_2_1__leaf_wb_clk_i
rlabel metal2 43400 20272 43400 20272 0 clknet_2_2__leaf_wb_clk_i
rlabel metal3 42336 44968 42336 44968 0 clknet_2_3__leaf_wb_clk_i
rlabel metal2 1736 21560 1736 21560 0 clknet_leaf_0_wb_clk_i
rlabel metal2 13664 45080 13664 45080 0 clknet_leaf_10_wb_clk_i
rlabel metal2 24584 43736 24584 43736 0 clknet_leaf_11_wb_clk_i
rlabel metal2 23128 39116 23128 39116 0 clknet_leaf_12_wb_clk_i
rlabel metal2 16408 33376 16408 33376 0 clknet_leaf_13_wb_clk_i
rlabel metal2 26768 26264 26768 26264 0 clknet_leaf_14_wb_clk_i
rlabel metal2 29064 33992 29064 33992 0 clknet_leaf_15_wb_clk_i
rlabel via2 25816 41944 25816 41944 0 clknet_leaf_16_wb_clk_i
rlabel metal2 36568 42784 36568 42784 0 clknet_leaf_17_wb_clk_i
rlabel metal2 44856 44632 44856 44632 0 clknet_leaf_18_wb_clk_i
rlabel metal2 47992 42784 47992 42784 0 clknet_leaf_19_wb_clk_i
rlabel metal2 12824 22008 12824 22008 0 clknet_leaf_1_wb_clk_i
rlabel metal2 47992 30576 47992 30576 0 clknet_leaf_20_wb_clk_i
rlabel metal2 45360 27048 45360 27048 0 clknet_leaf_21_wb_clk_i
rlabel metal2 39592 30632 39592 30632 0 clknet_leaf_22_wb_clk_i
rlabel metal2 30296 23296 30296 23296 0 clknet_leaf_23_wb_clk_i
rlabel metal2 40936 18088 40936 18088 0 clknet_leaf_24_wb_clk_i
rlabel metal2 48104 15680 48104 15680 0 clknet_leaf_25_wb_clk_i
rlabel metal2 44296 16408 44296 16408 0 clknet_leaf_26_wb_clk_i
rlabel metal2 48104 12936 48104 12936 0 clknet_leaf_27_wb_clk_i
rlabel metal2 45416 4368 45416 4368 0 clknet_leaf_28_wb_clk_i
rlabel metal2 35672 9800 35672 9800 0 clknet_leaf_29_wb_clk_i
rlabel metal2 18088 22792 18088 22792 0 clknet_leaf_2_wb_clk_i
rlabel metal2 25816 5880 25816 5880 0 clknet_leaf_30_wb_clk_i
rlabel metal2 26152 10472 26152 10472 0 clknet_leaf_31_wb_clk_i
rlabel metal2 35112 16520 35112 16520 0 clknet_leaf_32_wb_clk_i
rlabel metal2 24920 19992 24920 19992 0 clknet_leaf_33_wb_clk_i
rlabel metal2 16408 15204 16408 15204 0 clknet_leaf_34_wb_clk_i
rlabel metal2 24136 9408 24136 9408 0 clknet_leaf_35_wb_clk_i
rlabel metal2 13608 5488 13608 5488 0 clknet_leaf_36_wb_clk_i
rlabel metal2 8232 6720 8232 6720 0 clknet_leaf_37_wb_clk_i
rlabel metal3 3696 8232 3696 8232 0 clknet_leaf_38_wb_clk_i
rlabel metal2 1848 12936 1848 12936 0 clknet_leaf_39_wb_clk_i
rlabel metal2 20216 25088 20216 25088 0 clknet_leaf_3_wb_clk_i
rlabel metal2 17416 29848 17416 29848 0 clknet_leaf_4_wb_clk_i
rlabel metal2 1848 28224 1848 28224 0 clknet_leaf_5_wb_clk_i
rlabel metal2 1848 30744 1848 30744 0 clknet_leaf_6_wb_clk_i
rlabel metal2 9800 35224 9800 35224 0 clknet_leaf_7_wb_clk_i
rlabel metal2 6104 41608 6104 41608 0 clknet_leaf_8_wb_clk_i
rlabel metal2 10248 44296 10248 44296 0 clknet_leaf_9_wb_clk_i
rlabel metal3 47656 44072 47656 44072 0 custom_settings[0]
rlabel metal2 45304 46480 45304 46480 0 custom_settings[1]
rlabel metal3 48762 2744 48762 2744 0 io_in_1[0]
rlabel metal2 48216 7168 48216 7168 0 io_in_1[1]
rlabel metal2 48216 12656 48216 12656 0 io_in_1[2]
rlabel metal3 48762 17528 48762 17528 0 io_in_1[3]
rlabel metal2 48216 22792 48216 22792 0 io_in_1[4]
rlabel metal2 48216 28000 48216 28000 0 io_in_1[5]
rlabel metal3 44968 35896 44968 35896 0 io_in_1[6]
rlabel metal2 43848 39256 43848 39256 0 io_in_1[7]
rlabel metal2 32648 46144 32648 46144 0 io_in_2[0]
rlabel metal3 43764 45864 43764 45864 0 io_in_2[1]
rlabel metal2 19320 2086 19320 2086 0 io_out[10]
rlabel metal3 21504 3640 21504 3640 0 io_out[11]
rlabel metal2 30296 2198 30296 2198 0 io_out[17]
rlabel metal3 34440 3640 34440 3640 0 io_out[18]
rlabel metal3 33656 5992 33656 5992 0 io_out[19]
rlabel metal3 36512 4872 36512 4872 0 io_out[20]
rlabel metal2 36568 2254 36568 2254 0 io_out[21]
rlabel metal2 16184 854 16184 854 0 io_out[8]
rlabel metal2 17752 1806 17752 1806 0 io_out[9]
rlabel metal3 45696 44968 45696 44968 0 net1
rlabel metal2 48104 33264 48104 33264 0 net10
rlabel metal3 31696 40152 31696 40152 0 net11
rlabel metal2 39312 43960 39312 43960 0 net12
rlabel metal2 21336 18760 21336 18760 0 net13
rlabel metal2 13160 3864 13160 3864 0 net14
rlabel metal2 12936 4760 12936 4760 0 net15
rlabel metal2 24696 3472 24696 3472 0 net16
rlabel metal2 32200 3864 32200 3864 0 net17
rlabel metal2 35112 4256 35112 4256 0 net18
rlabel metal2 23128 16576 23128 16576 0 net19
rlabel metal2 45696 45752 45696 45752 0 net2
rlabel metal2 23912 8232 23912 8232 0 net20
rlabel metal2 16408 3752 16408 3752 0 net21
rlabel metal2 9688 5544 9688 5544 0 net22
rlabel metal2 3640 2030 3640 2030 0 net23
rlabel metal2 5208 2030 5208 2030 0 net24
rlabel metal2 6776 2030 6776 2030 0 net25
rlabel metal2 8344 2030 8344 2030 0 net26
rlabel metal2 9912 2030 9912 2030 0 net27
rlabel metal2 11480 2030 11480 2030 0 net28
rlabel metal2 13048 2030 13048 2030 0 net29
rlabel metal2 31192 19880 31192 19880 0 net3
rlabel metal2 14616 1246 14616 1246 0 net30
rlabel metal3 23856 4424 23856 4424 0 net31
rlabel metal2 24024 2030 24024 2030 0 net32
rlabel metal2 25592 2030 25592 2030 0 net33
rlabel metal2 27160 2030 27160 2030 0 net34
rlabel metal2 28728 1582 28728 1582 0 net35
rlabel metal3 40656 3864 40656 3864 0 net36
rlabel metal2 41272 1246 41272 1246 0 net37
rlabel metal2 42840 2030 42840 2030 0 net38
rlabel metal2 44408 854 44408 854 0 net39
rlabel metal2 47880 6664 47880 6664 0 net4
rlabel metal2 45976 2030 45976 2030 0 net40
rlabel metal2 38136 2030 38136 2030 0 net41
rlabel metal2 34832 17640 34832 17640 0 net5
rlabel metal2 47880 17808 47880 17808 0 net6
rlabel metal2 47880 24248 47880 24248 0 net7
rlabel metal2 44968 32312 44968 32312 0 net8
rlabel metal3 46536 33320 46536 33320 0 net9
rlabel metal2 18592 45976 18592 45976 0 rst_n
rlabel metal3 25872 31864 25872 31864 0 tt_um_rejunity_ay8913.active
rlabel metal2 21280 27832 21280 27832 0 tt_um_rejunity_ay8913.amplitude_A\[0\]
rlabel metal2 20720 24584 20720 24584 0 tt_um_rejunity_ay8913.amplitude_B\[0\]
rlabel metal2 21392 19320 21392 19320 0 tt_um_rejunity_ay8913.amplitude_C\[0\]
rlabel metal3 15736 28784 15736 28784 0 tt_um_rejunity_ay8913.clk_counter\[0\]
rlabel metal3 17080 29288 17080 29288 0 tt_um_rejunity_ay8913.clk_counter\[1\]
rlabel metal2 15904 27832 15904 27832 0 tt_um_rejunity_ay8913.clk_counter\[2\]
rlabel metal2 15512 22904 15512 22904 0 tt_um_rejunity_ay8913.clk_counter\[3\]
rlabel metal3 15148 20776 15148 20776 0 tt_um_rejunity_ay8913.clk_counter\[4\]
rlabel metal2 16856 20384 16856 20384 0 tt_um_rejunity_ay8913.clk_counter\[5\]
rlabel metal2 15288 19936 15288 19936 0 tt_um_rejunity_ay8913.clk_counter\[6\]
rlabel metal2 20664 25928 20664 25928 0 tt_um_rejunity_ay8913.envelope_A
rlabel metal2 18984 21896 18984 21896 0 tt_um_rejunity_ay8913.envelope_B
rlabel metal2 20440 23128 20440 23128 0 tt_um_rejunity_ay8913.envelope_C
rlabel metal3 11984 33432 11984 33432 0 tt_um_rejunity_ay8913.envelope_alternate
rlabel metal2 10920 35392 10920 35392 0 tt_um_rejunity_ay8913.envelope_attack
rlabel metal3 12432 32424 12432 32424 0 tt_um_rejunity_ay8913.envelope_continue
rlabel metal2 5992 34608 5992 34608 0 tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[0\]
rlabel metal2 1736 36176 1736 36176 0 tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[1\]
rlabel metal2 4144 39368 4144 39368 0 tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[2\]
rlabel metal2 1736 38360 1736 38360 0 tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[3\]
rlabel metal2 9912 33992 9912 33992 0 tt_um_rejunity_ay8913.envelope_generator.hold
rlabel metal2 7952 34776 7952 34776 0 tt_um_rejunity_ay8913.envelope_generator.invert_output
rlabel metal3 29680 39592 29680 39592 0 tt_um_rejunity_ay8913.envelope_generator.period\[0\]
rlabel metal2 39480 35616 39480 35616 0 tt_um_rejunity_ay8913.envelope_generator.period\[10\]
rlabel metal2 42616 35168 42616 35168 0 tt_um_rejunity_ay8913.envelope_generator.period\[11\]
rlabel metal2 43736 32984 43736 32984 0 tt_um_rejunity_ay8913.envelope_generator.period\[12\]
rlabel metal2 44968 37296 44968 37296 0 tt_um_rejunity_ay8913.envelope_generator.period\[13\]
rlabel metal2 47432 35896 47432 35896 0 tt_um_rejunity_ay8913.envelope_generator.period\[14\]
rlabel metal2 47880 37968 47880 37968 0 tt_um_rejunity_ay8913.envelope_generator.period\[15\]
rlabel metal2 29288 36512 29288 36512 0 tt_um_rejunity_ay8913.envelope_generator.period\[1\]
rlabel metal2 31024 36456 31024 36456 0 tt_um_rejunity_ay8913.envelope_generator.period\[2\]
rlabel metal3 31640 35672 31640 35672 0 tt_um_rejunity_ay8913.envelope_generator.period\[3\]
rlabel metal2 32984 40880 32984 40880 0 tt_um_rejunity_ay8913.envelope_generator.period\[4\]
rlabel metal3 35112 41048 35112 41048 0 tt_um_rejunity_ay8913.envelope_generator.period\[5\]
rlabel metal2 35112 40096 35112 40096 0 tt_um_rejunity_ay8913.envelope_generator.period\[6\]
rlabel metal2 37688 40656 37688 40656 0 tt_um_rejunity_ay8913.envelope_generator.period\[7\]
rlabel metal2 39816 33656 39816 33656 0 tt_um_rejunity_ay8913.envelope_generator.period\[8\]
rlabel metal3 40488 37128 40488 37128 0 tt_um_rejunity_ay8913.envelope_generator.period\[9\]
rlabel metal2 8176 38696 8176 38696 0 tt_um_rejunity_ay8913.envelope_generator.signal_edge.previous_signal_state_0
rlabel metal3 10080 38920 10080 38920 0 tt_um_rejunity_ay8913.envelope_generator.signal_edge.signal
rlabel metal2 7896 36904 7896 36904 0 tt_um_rejunity_ay8913.envelope_generator.stop
rlabel metal2 26152 40040 26152 40040 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[0\]
rlabel metal2 41384 41496 41384 41496 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[10\]
rlabel metal2 43848 44464 43848 44464 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[11\]
rlabel metal2 46928 42728 46928 42728 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[12\]
rlabel metal2 47040 42616 47040 42616 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[13\]
rlabel metal2 45584 40376 45584 40376 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[14\]
rlabel metal3 46368 39032 46368 39032 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[15\]
rlabel metal2 28952 40936 28952 40936 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[1\]
rlabel metal2 29176 42336 29176 42336 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[2\]
rlabel metal2 30296 43344 30296 43344 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[3\]
rlabel metal2 30632 45360 30632 45360 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[4\]
rlabel metal3 34048 44968 34048 44968 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[5\]
rlabel metal2 36456 43792 36456 43792 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[6\]
rlabel metal3 39032 43736 39032 43736 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[7\]
rlabel metal2 45080 41608 45080 41608 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[8\]
rlabel metal2 40936 39984 40936 39984 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[9\]
rlabel metal2 26152 28672 26152 28672 0 tt_um_rejunity_ay8913.latched_register\[0\]
rlabel metal2 28616 28448 28616 28448 0 tt_um_rejunity_ay8913.latched_register\[1\]
rlabel metal2 30408 30016 30408 30016 0 tt_um_rejunity_ay8913.latched_register\[2\]
rlabel metal2 31640 31472 31640 31472 0 tt_um_rejunity_ay8913.latched_register\[3\]
rlabel metal2 19040 27160 19040 27160 0 tt_um_rejunity_ay8913.noise_disable_A
rlabel metal3 28672 23912 28672 23912 0 tt_um_rejunity_ay8913.noise_disable_B
rlabel metal2 26712 23128 26712 23128 0 tt_um_rejunity_ay8913.noise_disable_C
rlabel metal2 24584 26320 24584 26320 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[0\]
rlabel metal2 3192 28952 3192 28952 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[10\]
rlabel metal2 7728 29960 7728 29960 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[11\]
rlabel metal2 6216 29792 6216 29792 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[12\]
rlabel metal2 6552 31080 6552 31080 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[13\]
rlabel metal2 7784 32256 7784 32256 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[14\]
rlabel metal2 8456 30128 8456 30128 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[15\]
rlabel metal2 7784 26684 7784 26684 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[16\]
rlabel metal3 10584 25256 10584 25256 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[1\]
rlabel metal2 10024 24752 10024 24752 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[2\]
rlabel metal3 9800 23240 9800 23240 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[3\]
rlabel metal2 7560 22400 7560 22400 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[4\]
rlabel metal2 3304 21336 3304 21336 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[5\]
rlabel metal2 4648 22512 4648 22512 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[6\]
rlabel metal2 4200 23352 4200 23352 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[7\]
rlabel metal2 1736 25704 1736 25704 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[8\]
rlabel metal2 4648 25536 4648 25536 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[9\]
rlabel metal2 30856 17360 30856 17360 0 tt_um_rejunity_ay8913.noise_generator.period\[0\]
rlabel metal2 30744 16072 30744 16072 0 tt_um_rejunity_ay8913.noise_generator.period\[1\]
rlabel metal3 30800 13720 30800 13720 0 tt_um_rejunity_ay8913.noise_generator.period\[2\]
rlabel metal3 29512 12712 29512 12712 0 tt_um_rejunity_ay8913.noise_generator.period\[3\]
rlabel metal2 27384 16856 27384 16856 0 tt_um_rejunity_ay8913.noise_generator.period\[4\]
rlabel metal2 8232 18648 8232 18648 0 tt_um_rejunity_ay8913.noise_generator.signal_edge.previous_signal_state_0
rlabel metal3 7336 13720 7336 13720 0 tt_um_rejunity_ay8913.noise_generator.signal_edge.signal
rlabel metal2 26376 17584 26376 17584 0 tt_um_rejunity_ay8913.noise_generator.tone.counter\[0\]
rlabel metal2 27160 16520 27160 16520 0 tt_um_rejunity_ay8913.noise_generator.tone.counter\[1\]
rlabel metal2 26488 14168 26488 14168 0 tt_um_rejunity_ay8913.noise_generator.tone.counter\[2\]
rlabel metal3 25928 12768 25928 12768 0 tt_um_rejunity_ay8913.noise_generator.tone.counter\[3\]
rlabel metal2 28616 11760 28616 11760 0 tt_um_rejunity_ay8913.noise_generator.tone.counter\[4\]
rlabel metal2 15736 17696 15736 17696 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[2\]
rlabel metal2 12712 17696 12712 17696 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[3\]
rlabel metal2 9016 16800 9016 16800 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[4\]
rlabel metal2 9856 15512 9856 15512 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[5\]
rlabel metal2 11592 13776 11592 13776 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[6\]
rlabel metal2 15064 14448 15064 14448 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[7\]
rlabel metal2 14112 12936 14112 12936 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[8\]
rlabel metal3 4872 16856 4872 16856 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[2\]
rlabel metal2 4088 14868 4088 14868 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[3\]
rlabel metal2 3528 11368 3528 11368 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[4\]
rlabel metal2 4648 8372 4648 8372 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[5\]
rlabel metal2 4648 6328 4648 6328 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[6\]
rlabel metal2 6664 6384 6664 6384 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[7\]
rlabel metal3 7224 5880 7224 5880 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[8\]
rlabel metal2 19992 21168 19992 21168 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[2\]
rlabel metal2 11088 19320 11088 19320 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[3\]
rlabel metal2 4424 18984 4424 18984 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[4\]
rlabel metal2 4648 13944 4648 13944 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[5\]
rlabel metal2 5432 12320 5432 12320 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[6\]
rlabel metal2 5992 12096 5992 12096 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[7\]
rlabel metal2 7224 9520 7224 9520 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[8\]
rlabel metal3 22176 16744 22176 16744 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[2\]
rlabel metal2 18760 14896 18760 14896 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[3\]
rlabel metal3 20440 12936 20440 12936 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[4\]
rlabel metal3 18816 12936 18816 12936 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[5\]
rlabel metal2 10192 11480 10192 11480 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[6\]
rlabel metal2 14504 9464 14504 9464 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[7\]
rlabel metal2 11088 6776 11088 6776 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[8\]
rlabel metal2 12488 7784 12488 7784 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[9\]
rlabel metal2 12712 36120 12712 36120 0 tt_um_rejunity_ay8913.restart_envelope
rlabel metal2 28616 4200 28616 4200 0 tt_um_rejunity_ay8913.spi_dac_i_2.counter\[0\]
rlabel metal2 26040 9912 26040 9912 0 tt_um_rejunity_ay8913.spi_dac_i_2.counter\[1\]
rlabel metal2 29624 8624 29624 8624 0 tt_um_rejunity_ay8913.spi_dac_i_2.counter\[2\]
rlabel metal2 28504 8176 28504 8176 0 tt_um_rejunity_ay8913.spi_dac_i_2.counter\[3\]
rlabel metal2 29064 7728 29064 7728 0 tt_um_rejunity_ay8913.spi_dac_i_2.counter\[4\]
rlabel metal3 18704 5208 18704 5208 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[10\]
rlabel metal3 23688 4200 23688 4200 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[11\]
rlabel metal2 24584 5936 24584 5936 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[2\]
rlabel metal2 22008 8568 22008 8568 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[3\]
rlabel metal3 21448 9800 21448 9800 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[4\]
rlabel metal2 20328 9184 20328 9184 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[5\]
rlabel metal3 18816 8120 18816 8120 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[6\]
rlabel metal2 16800 7336 16800 7336 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[7\]
rlabel metal2 16240 6776 16240 6776 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[8\]
rlabel metal2 16408 4312 16408 4312 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[9\]
rlabel metal2 20328 28560 20328 28560 0 tt_um_rejunity_ay8913.tone_A
rlabel metal2 17080 36512 17080 36512 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[0\]
rlabel metal2 12824 41272 12824 41272 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[10\]
rlabel metal2 15680 39480 15680 39480 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[11\]
rlabel metal2 17752 37408 17752 37408 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[1\]
rlabel metal2 20104 39480 20104 39480 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[2\]
rlabel metal3 17248 43624 17248 43624 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[3\]
rlabel metal3 19992 44408 19992 44408 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[4\]
rlabel metal2 16688 44968 16688 44968 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[5\]
rlabel metal2 11480 43960 11480 43960 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[6\]
rlabel metal2 11592 44352 11592 44352 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[7\]
rlabel metal2 12600 43456 12600 43456 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[8\]
rlabel metal2 11928 41832 11928 41832 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[9\]
rlabel metal2 18032 35000 18032 35000 0 tt_um_rejunity_ay8913.tone_A_generator.period\[0\]
rlabel metal2 20440 39144 20440 39144 0 tt_um_rejunity_ay8913.tone_A_generator.period\[10\]
rlabel metal2 22008 37912 22008 37912 0 tt_um_rejunity_ay8913.tone_A_generator.period\[11\]
rlabel metal2 17920 34216 17920 34216 0 tt_um_rejunity_ay8913.tone_A_generator.period\[1\]
rlabel metal2 20440 33656 20440 33656 0 tt_um_rejunity_ay8913.tone_A_generator.period\[2\]
rlabel metal2 18648 42112 18648 42112 0 tt_um_rejunity_ay8913.tone_A_generator.period\[3\]
rlabel metal2 21784 41160 21784 41160 0 tt_um_rejunity_ay8913.tone_A_generator.period\[4\]
rlabel metal2 23912 44800 23912 44800 0 tt_um_rejunity_ay8913.tone_A_generator.period\[5\]
rlabel metal2 23240 44800 23240 44800 0 tt_um_rejunity_ay8913.tone_A_generator.period\[6\]
rlabel metal2 25200 43624 25200 43624 0 tt_um_rejunity_ay8913.tone_A_generator.period\[7\]
rlabel metal2 25984 39928 25984 39928 0 tt_um_rejunity_ay8913.tone_A_generator.period\[8\]
rlabel metal2 25368 36904 25368 36904 0 tt_um_rejunity_ay8913.tone_A_generator.period\[9\]
rlabel metal2 19096 26208 19096 26208 0 tt_um_rejunity_ay8913.tone_B
rlabel metal2 39928 25312 39928 25312 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[0\]
rlabel metal2 44968 19488 44968 19488 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[10\]
rlabel metal2 47656 18928 47656 18928 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[11\]
rlabel metal2 39256 24248 39256 24248 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[1\]
rlabel metal2 39312 27720 39312 27720 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[2\]
rlabel metal2 40320 29512 40320 29512 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[3\]
rlabel metal3 45136 28056 45136 28056 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[4\]
rlabel metal2 47656 26628 47656 26628 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[5\]
rlabel metal2 45192 23352 45192 23352 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[6\]
rlabel metal2 45360 24024 45360 24024 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[7\]
rlabel metal2 44520 23408 44520 23408 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[8\]
rlabel metal3 43344 20888 43344 20888 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[9\]
rlabel metal3 33096 25592 33096 25592 0 tt_um_rejunity_ay8913.tone_B_generator.period\[0\]
rlabel metal3 40600 19992 40600 19992 0 tt_um_rejunity_ay8913.tone_B_generator.period\[10\]
rlabel metal2 39368 19208 39368 19208 0 tt_um_rejunity_ay8913.tone_B_generator.period\[11\]
rlabel metal3 35056 24584 35056 24584 0 tt_um_rejunity_ay8913.tone_B_generator.period\[1\]
rlabel metal3 39872 27048 39872 27048 0 tt_um_rejunity_ay8913.tone_B_generator.period\[2\]
rlabel metal2 39704 26852 39704 26852 0 tt_um_rejunity_ay8913.tone_B_generator.period\[3\]
rlabel metal2 41720 28840 41720 28840 0 tt_um_rejunity_ay8913.tone_B_generator.period\[4\]
rlabel metal2 48160 26376 48160 26376 0 tt_um_rejunity_ay8913.tone_B_generator.period\[5\]
rlabel metal3 44632 25480 44632 25480 0 tt_um_rejunity_ay8913.tone_B_generator.period\[6\]
rlabel metal2 43400 31472 43400 31472 0 tt_um_rejunity_ay8913.tone_B_generator.period\[7\]
rlabel metal2 41944 21840 41944 21840 0 tt_um_rejunity_ay8913.tone_B_generator.period\[8\]
rlabel metal2 41048 20328 41048 20328 0 tt_um_rejunity_ay8913.tone_B_generator.period\[9\]
rlabel metal2 26488 22344 26488 22344 0 tt_um_rejunity_ay8913.tone_C
rlabel via1 39928 16197 39928 16197 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[0\]
rlabel metal2 42168 4872 42168 4872 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[10\]
rlabel metal2 39928 7056 39928 7056 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[11\]
rlabel metal2 38472 13272 38472 13272 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[1\]
rlabel metal3 40264 15176 40264 15176 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[2\]
rlabel metal2 41944 13048 41944 13048 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[3\]
rlabel metal2 42952 12376 42952 12376 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[4\]
rlabel metal2 43400 9856 43400 9856 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[5\]
rlabel metal2 45304 7672 45304 7672 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[6\]
rlabel metal2 42280 8960 42280 8960 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[7\]
rlabel metal2 44072 6608 44072 6608 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[8\]
rlabel metal2 40768 5880 40768 5880 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[9\]
rlabel metal2 37688 11312 37688 11312 0 tt_um_rejunity_ay8913.tone_C_generator.period\[0\]
rlabel metal2 39592 5768 39592 5768 0 tt_um_rejunity_ay8913.tone_C_generator.period\[10\]
rlabel metal3 39592 5880 39592 5880 0 tt_um_rejunity_ay8913.tone_C_generator.period\[11\]
rlabel metal2 36232 12432 36232 12432 0 tt_um_rejunity_ay8913.tone_C_generator.period\[1\]
rlabel metal2 39032 11312 39032 11312 0 tt_um_rejunity_ay8913.tone_C_generator.period\[2\]
rlabel metal3 39088 12152 39088 12152 0 tt_um_rejunity_ay8913.tone_C_generator.period\[3\]
rlabel metal2 41608 17304 41608 17304 0 tt_um_rejunity_ay8913.tone_C_generator.period\[4\]
rlabel metal2 42952 14560 42952 14560 0 tt_um_rejunity_ay8913.tone_C_generator.period\[5\]
rlabel metal2 44744 15148 44744 15148 0 tt_um_rejunity_ay8913.tone_C_generator.period\[6\]
rlabel metal2 45304 16912 45304 16912 0 tt_um_rejunity_ay8913.tone_C_generator.period\[7\]
rlabel metal2 35224 8288 35224 8288 0 tt_um_rejunity_ay8913.tone_C_generator.period\[8\]
rlabel metal3 34552 5880 34552 5880 0 tt_um_rejunity_ay8913.tone_C_generator.period\[9\]
rlabel metal2 20216 29736 20216 29736 0 tt_um_rejunity_ay8913.tone_disable_A
rlabel metal3 17752 26264 17752 26264 0 tt_um_rejunity_ay8913.tone_disable_B
rlabel metal2 26712 24304 26712 24304 0 tt_um_rejunity_ay8913.tone_disable_C
rlabel metal3 25592 24696 25592 24696 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
