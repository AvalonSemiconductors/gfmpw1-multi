VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_sn76489
  CLASS BLOCK ;
  FOREIGN wrapped_sn76489 ;
  ORIGIN 0.000 0.000 ;
  SIZE 250.000 BY 250.000 ;
  PIN custom_settings[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 210.560 250.000 211.120 ;
    END
  END custom_settings[0]
  PIN custom_settings[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 235.200 250.000 235.760 ;
    END
  END custom_settings[1]
  PIN io_in_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    ANTENNADIFFAREA 0.877000 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 13.440 250.000 14.000 ;
    END
  END io_in_1[0]
  PIN io_in_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 38.080 250.000 38.640 ;
    END
  END io_in_1[1]
  PIN io_in_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 62.720 250.000 63.280 ;
    END
  END io_in_1[2]
  PIN io_in_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 87.360 250.000 87.920 ;
    END
  END io_in_1[3]
  PIN io_in_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 112.000 250.000 112.560 ;
    END
  END io_in_1[4]
  PIN io_in_1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 136.640 250.000 137.200 ;
    END
  END io_in_1[5]
  PIN io_in_1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 161.280 250.000 161.840 ;
    END
  END io_in_1[6]
  PIN io_in_1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 185.920 250.000 186.480 ;
    END
  END io_in_1[7]
  PIN io_in_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 207.200 4.000 207.760 ;
    END
  END io_in_2
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal2 ;
        RECT 17.920 246.000 18.480 250.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 96.320 246.000 96.880 250.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 246.000 104.720 250.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 112.000 246.000 112.560 250.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal2 ;
        RECT 119.840 246.000 120.400 250.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 246.000 128.240 250.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal2 ;
        RECT 135.520 246.000 136.080 250.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal2 ;
        RECT 143.360 246.000 143.920 250.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 246.000 151.760 250.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 159.040 246.000 159.600 250.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 166.880 246.000 167.440 250.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal2 ;
        RECT 25.760 246.000 26.320 250.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 174.720 246.000 175.280 250.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 182.560 246.000 183.120 250.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 190.400 246.000 190.960 250.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 198.240 246.000 198.800 250.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 206.080 246.000 206.640 250.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 213.920 246.000 214.480 250.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 246.000 222.320 250.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 229.600 246.000 230.160 250.000 ;
    END
  END io_out[27]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 246.000 34.160 250.000 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal2 ;
        RECT 41.440 246.000 42.000 250.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal2 ;
        RECT 49.280 246.000 49.840 250.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 246.000 57.680 250.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal2 ;
        RECT 64.960 246.000 65.520 250.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal2 ;
        RECT 72.800 246.000 73.360 250.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 246.000 81.200 250.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 88.480 246.000 89.040 250.000 ;
    END
  END io_out[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 124.320 4.000 124.880 ;
    END
  END rst_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 231.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 231.580 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 231.580 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.352000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 41.440 4.000 42.000 ;
    END
  END wb_clk_i
  OBS
      LAYER Nwell ;
        RECT 6.290 15.250 243.470 231.710 ;
      LAYER Metal1 ;
        RECT 6.720 15.380 243.040 231.580 ;
      LAYER Metal2 ;
        RECT 0.140 245.700 17.620 246.820 ;
        RECT 18.780 245.700 25.460 246.820 ;
        RECT 26.620 245.700 33.300 246.820 ;
        RECT 34.460 245.700 41.140 246.820 ;
        RECT 42.300 245.700 48.980 246.820 ;
        RECT 50.140 245.700 56.820 246.820 ;
        RECT 57.980 245.700 64.660 246.820 ;
        RECT 65.820 245.700 72.500 246.820 ;
        RECT 73.660 245.700 80.340 246.820 ;
        RECT 81.500 245.700 88.180 246.820 ;
        RECT 89.340 245.700 96.020 246.820 ;
        RECT 97.180 245.700 103.860 246.820 ;
        RECT 105.020 245.700 111.700 246.820 ;
        RECT 112.860 245.700 119.540 246.820 ;
        RECT 120.700 245.700 127.380 246.820 ;
        RECT 128.540 245.700 135.220 246.820 ;
        RECT 136.380 245.700 143.060 246.820 ;
        RECT 144.220 245.700 150.900 246.820 ;
        RECT 152.060 245.700 158.740 246.820 ;
        RECT 159.900 245.700 166.580 246.820 ;
        RECT 167.740 245.700 174.420 246.820 ;
        RECT 175.580 245.700 182.260 246.820 ;
        RECT 183.420 245.700 190.100 246.820 ;
        RECT 191.260 245.700 197.940 246.820 ;
        RECT 199.100 245.700 205.780 246.820 ;
        RECT 206.940 245.700 213.620 246.820 ;
        RECT 214.780 245.700 221.460 246.820 ;
        RECT 222.620 245.700 229.300 246.820 ;
        RECT 230.460 245.700 244.020 246.820 ;
        RECT 0.140 13.530 244.020 245.700 ;
      LAYER Metal3 ;
        RECT 0.090 234.900 245.700 235.620 ;
        RECT 0.090 211.420 246.820 234.900 ;
        RECT 0.090 210.260 245.700 211.420 ;
        RECT 0.090 208.060 246.820 210.260 ;
        RECT 4.300 206.900 246.820 208.060 ;
        RECT 0.090 186.780 246.820 206.900 ;
        RECT 0.090 185.620 245.700 186.780 ;
        RECT 0.090 162.140 246.820 185.620 ;
        RECT 0.090 160.980 245.700 162.140 ;
        RECT 0.090 137.500 246.820 160.980 ;
        RECT 0.090 136.340 245.700 137.500 ;
        RECT 0.090 125.180 246.820 136.340 ;
        RECT 4.300 124.020 246.820 125.180 ;
        RECT 0.090 112.860 246.820 124.020 ;
        RECT 0.090 111.700 245.700 112.860 ;
        RECT 0.090 88.220 246.820 111.700 ;
        RECT 0.090 87.060 245.700 88.220 ;
        RECT 0.090 63.580 246.820 87.060 ;
        RECT 0.090 62.420 245.700 63.580 ;
        RECT 0.090 42.300 246.820 62.420 ;
        RECT 4.300 41.140 246.820 42.300 ;
        RECT 0.090 38.940 246.820 41.140 ;
        RECT 0.090 37.780 245.700 38.940 ;
        RECT 0.090 14.300 246.820 37.780 ;
        RECT 0.090 13.580 245.700 14.300 ;
      LAYER Metal4 ;
        RECT 32.060 16.330 98.740 227.830 ;
        RECT 100.940 16.330 175.540 227.830 ;
        RECT 177.740 16.330 234.500 227.830 ;
  END
END wrapped_sn76489
END LIBRARY

