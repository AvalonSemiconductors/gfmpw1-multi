magic
tech gf180mcuD
magscale 1 10
timestamp 1702253718
<< metal1 >>
rect 1344 33738 35616 33772
rect 1344 33686 5498 33738
rect 5550 33686 5602 33738
rect 5654 33686 5706 33738
rect 5758 33686 14066 33738
rect 14118 33686 14170 33738
rect 14222 33686 14274 33738
rect 14326 33686 22634 33738
rect 22686 33686 22738 33738
rect 22790 33686 22842 33738
rect 22894 33686 31202 33738
rect 31254 33686 31306 33738
rect 31358 33686 31410 33738
rect 31462 33686 35616 33738
rect 1344 33652 35616 33686
rect 12350 33570 12402 33582
rect 12350 33506 12402 33518
rect 25566 33570 25618 33582
rect 25566 33506 25618 33518
rect 30046 33570 30098 33582
rect 30046 33506 30098 33518
rect 23774 33458 23826 33470
rect 8194 33406 8206 33458
rect 8258 33406 8270 33458
rect 16034 33406 16046 33458
rect 16098 33406 16110 33458
rect 19842 33406 19854 33458
rect 19906 33406 19918 33458
rect 35074 33406 35086 33458
rect 35138 33406 35150 33458
rect 23774 33394 23826 33406
rect 6402 33294 6414 33346
rect 6466 33294 6478 33346
rect 9986 33294 9998 33346
rect 10050 33294 10062 33346
rect 13234 33294 13246 33346
rect 13298 33294 13310 33346
rect 17042 33294 17054 33346
rect 17106 33294 17118 33346
rect 20962 33294 20974 33346
rect 21026 33294 21038 33346
rect 24770 33294 24782 33346
rect 24834 33294 24846 33346
rect 29026 33294 29038 33346
rect 29090 33294 29102 33346
rect 32162 33294 32174 33346
rect 32226 33294 32238 33346
rect 1822 33234 1874 33246
rect 1822 33170 1874 33182
rect 2942 33234 2994 33246
rect 2942 33170 2994 33182
rect 4062 33234 4114 33246
rect 4062 33170 4114 33182
rect 4958 33234 5010 33246
rect 4958 33170 5010 33182
rect 5854 33234 5906 33246
rect 5854 33170 5906 33182
rect 9550 33234 9602 33246
rect 13906 33182 13918 33234
rect 13970 33182 13982 33234
rect 17714 33182 17726 33234
rect 17778 33182 17790 33234
rect 21634 33182 21646 33234
rect 21698 33182 21710 33234
rect 32946 33182 32958 33234
rect 33010 33182 33022 33234
rect 9550 33170 9602 33182
rect 27582 33122 27634 33134
rect 27582 33058 27634 33070
rect 28702 33122 28754 33134
rect 28702 33058 28754 33070
rect 1344 32954 35776 32988
rect 1344 32902 9782 32954
rect 9834 32902 9886 32954
rect 9938 32902 9990 32954
rect 10042 32902 18350 32954
rect 18402 32902 18454 32954
rect 18506 32902 18558 32954
rect 18610 32902 26918 32954
rect 26970 32902 27022 32954
rect 27074 32902 27126 32954
rect 27178 32902 35486 32954
rect 35538 32902 35590 32954
rect 35642 32902 35694 32954
rect 35746 32902 35776 32954
rect 1344 32868 35776 32902
rect 9550 32786 9602 32798
rect 9550 32722 9602 32734
rect 15822 32786 15874 32798
rect 15822 32722 15874 32734
rect 18622 32786 18674 32798
rect 18622 32722 18674 32734
rect 33742 32786 33794 32798
rect 33742 32722 33794 32734
rect 16830 32674 16882 32686
rect 16146 32622 16158 32674
rect 16210 32622 16222 32674
rect 16830 32610 16882 32622
rect 31726 32674 31778 32686
rect 31726 32610 31778 32622
rect 34862 32674 34914 32686
rect 34862 32610 34914 32622
rect 35198 32674 35250 32686
rect 35198 32610 35250 32622
rect 16494 32562 16546 32574
rect 24110 32562 24162 32574
rect 6178 32510 6190 32562
rect 6242 32510 6254 32562
rect 12450 32510 12462 32562
rect 12514 32510 12526 32562
rect 17602 32510 17614 32562
rect 17666 32510 17678 32562
rect 20514 32510 20526 32562
rect 20578 32510 20590 32562
rect 16494 32498 16546 32510
rect 24110 32498 24162 32510
rect 24558 32562 24610 32574
rect 31838 32562 31890 32574
rect 25218 32510 25230 32562
rect 25282 32510 25294 32562
rect 28466 32510 28478 32562
rect 28530 32510 28542 32562
rect 24558 32498 24610 32510
rect 31838 32498 31890 32510
rect 10222 32450 10274 32462
rect 23438 32450 23490 32462
rect 6850 32398 6862 32450
rect 6914 32398 6926 32450
rect 8978 32398 8990 32450
rect 9042 32398 9054 32450
rect 13122 32398 13134 32450
rect 13186 32398 13198 32450
rect 15362 32398 15374 32450
rect 15426 32398 15438 32450
rect 21298 32398 21310 32450
rect 21362 32398 21374 32450
rect 10222 32386 10274 32398
rect 23438 32386 23490 32398
rect 26238 32450 26290 32462
rect 34190 32450 34242 32462
rect 29138 32398 29150 32450
rect 29202 32398 29214 32450
rect 31266 32398 31278 32450
rect 31330 32398 31342 32450
rect 26238 32386 26290 32398
rect 34190 32386 34242 32398
rect 34638 32450 34690 32462
rect 34638 32386 34690 32398
rect 31726 32338 31778 32350
rect 33618 32286 33630 32338
rect 33682 32335 33694 32338
rect 34514 32335 34526 32338
rect 33682 32289 34526 32335
rect 33682 32286 33694 32289
rect 34514 32286 34526 32289
rect 34578 32286 34590 32338
rect 31726 32274 31778 32286
rect 1344 32170 35616 32204
rect 1344 32118 5498 32170
rect 5550 32118 5602 32170
rect 5654 32118 5706 32170
rect 5758 32118 14066 32170
rect 14118 32118 14170 32170
rect 14222 32118 14274 32170
rect 14326 32118 22634 32170
rect 22686 32118 22738 32170
rect 22790 32118 22842 32170
rect 22894 32118 31202 32170
rect 31254 32118 31306 32170
rect 31358 32118 31410 32170
rect 31462 32118 35616 32170
rect 1344 32084 35616 32118
rect 8094 32002 8146 32014
rect 8094 31938 8146 31950
rect 11902 31890 11954 31902
rect 22430 31890 22482 31902
rect 11442 31838 11454 31890
rect 11506 31838 11518 31890
rect 16034 31838 16046 31890
rect 16098 31838 16110 31890
rect 18274 31838 18286 31890
rect 18338 31838 18350 31890
rect 20402 31838 20414 31890
rect 20466 31838 20478 31890
rect 11902 31826 11954 31838
rect 22430 31826 22482 31838
rect 27358 31890 27410 31902
rect 28018 31838 28030 31890
rect 28082 31838 28094 31890
rect 32050 31838 32062 31890
rect 32114 31838 32126 31890
rect 27358 31826 27410 31838
rect 21422 31778 21474 31790
rect 8642 31726 8654 31778
rect 8706 31726 8718 31778
rect 14578 31726 14590 31778
rect 14642 31726 14654 31778
rect 17490 31726 17502 31778
rect 17554 31726 17566 31778
rect 21422 31714 21474 31726
rect 21758 31778 21810 31790
rect 21758 31714 21810 31726
rect 22654 31778 22706 31790
rect 26910 31778 26962 31790
rect 23314 31726 23326 31778
rect 23378 31726 23390 31778
rect 22654 31714 22706 31726
rect 26910 31714 26962 31726
rect 27806 31778 27858 31790
rect 29250 31726 29262 31778
rect 29314 31726 29326 31778
rect 32386 31726 32398 31778
rect 32450 31726 32462 31778
rect 27806 31714 27858 31726
rect 7422 31666 7474 31678
rect 7422 31602 7474 31614
rect 8206 31666 8258 31678
rect 22094 31666 22146 31678
rect 28142 31666 28194 31678
rect 9314 31614 9326 31666
rect 9378 31614 9390 31666
rect 24098 31614 24110 31666
rect 24162 31614 24174 31666
rect 28242 31614 28254 31666
rect 28306 31614 28318 31666
rect 29922 31614 29934 31666
rect 29986 31614 29998 31666
rect 8206 31602 8258 31614
rect 22094 31602 22146 31614
rect 28142 31602 28194 31614
rect 13806 31554 13858 31566
rect 13806 31490 13858 31502
rect 14254 31554 14306 31566
rect 14254 31490 14306 31502
rect 21758 31554 21810 31566
rect 26798 31554 26850 31566
rect 22978 31502 22990 31554
rect 23042 31502 23054 31554
rect 26338 31502 26350 31554
rect 26402 31502 26414 31554
rect 21758 31490 21810 31502
rect 26798 31490 26850 31502
rect 28030 31554 28082 31566
rect 28030 31490 28082 31502
rect 33406 31554 33458 31566
rect 33406 31490 33458 31502
rect 1344 31386 35776 31420
rect 1344 31334 9782 31386
rect 9834 31334 9886 31386
rect 9938 31334 9990 31386
rect 10042 31334 18350 31386
rect 18402 31334 18454 31386
rect 18506 31334 18558 31386
rect 18610 31334 26918 31386
rect 26970 31334 27022 31386
rect 27074 31334 27126 31386
rect 27178 31334 35486 31386
rect 35538 31334 35590 31386
rect 35642 31334 35694 31386
rect 35746 31334 35776 31386
rect 1344 31300 35776 31334
rect 8430 31218 8482 31230
rect 8430 31154 8482 31166
rect 9550 31218 9602 31230
rect 9550 31154 9602 31166
rect 15374 31218 15426 31230
rect 15374 31154 15426 31166
rect 20750 31218 20802 31230
rect 20750 31154 20802 31166
rect 25342 31218 25394 31230
rect 25342 31154 25394 31166
rect 30830 31218 30882 31230
rect 30830 31154 30882 31166
rect 33518 31218 33570 31230
rect 33518 31154 33570 31166
rect 33630 31218 33682 31230
rect 33630 31154 33682 31166
rect 16718 31106 16770 31118
rect 7634 31054 7646 31106
rect 7698 31054 7710 31106
rect 10210 31054 10222 31106
rect 10274 31054 10286 31106
rect 11330 31054 11342 31106
rect 11394 31054 11406 31106
rect 16258 31054 16270 31106
rect 16322 31054 16334 31106
rect 16718 31042 16770 31054
rect 17614 31106 17666 31118
rect 17614 31042 17666 31054
rect 18734 31106 18786 31118
rect 25454 31106 25506 31118
rect 19058 31054 19070 31106
rect 19122 31054 19134 31106
rect 23538 31054 23550 31106
rect 23602 31054 23614 31106
rect 18734 31042 18786 31054
rect 25454 31042 25506 31054
rect 31726 31106 31778 31118
rect 31726 31042 31778 31054
rect 31838 31106 31890 31118
rect 31838 31042 31890 31054
rect 32398 31106 32450 31118
rect 33954 31054 33966 31106
rect 34018 31054 34030 31106
rect 32398 31042 32450 31054
rect 7982 30994 8034 31006
rect 4386 30942 4398 30994
rect 4450 30942 4462 30994
rect 7982 30930 8034 30942
rect 10110 30994 10162 31006
rect 10110 30930 10162 30942
rect 10446 30994 10498 31006
rect 15598 30994 15650 31006
rect 10658 30942 10670 30994
rect 10722 30942 10734 30994
rect 11554 30942 11566 30994
rect 11618 30942 11630 30994
rect 12114 30942 12126 30994
rect 12178 30942 12190 30994
rect 10446 30930 10498 30942
rect 15598 30930 15650 30942
rect 16046 30994 16098 31006
rect 16046 30930 16098 30942
rect 16382 30994 16434 31006
rect 16382 30930 16434 30942
rect 17390 30994 17442 31006
rect 17390 30930 17442 30942
rect 17726 30994 17778 31006
rect 18398 30994 18450 31006
rect 17938 30942 17950 30994
rect 18002 30942 18014 30994
rect 17726 30930 17778 30942
rect 18398 30930 18450 30942
rect 19406 30994 19458 31006
rect 22766 30994 22818 31006
rect 30606 30994 30658 31006
rect 32062 30994 32114 31006
rect 19842 30942 19854 30994
rect 19906 30942 19918 30994
rect 23426 30942 23438 30994
rect 23490 30942 23502 30994
rect 24546 30942 24558 30994
rect 24610 30942 24622 30994
rect 27458 30942 27470 30994
rect 27522 30942 27534 30994
rect 31042 30942 31054 30994
rect 31106 30942 31118 30994
rect 31378 30942 31390 30994
rect 31442 30942 31454 30994
rect 19406 30930 19458 30942
rect 22766 30930 22818 30942
rect 30606 30930 30658 30942
rect 32062 30930 32114 30942
rect 32510 30994 32562 31006
rect 32510 30930 32562 30942
rect 32958 30994 33010 31006
rect 32958 30930 33010 30942
rect 33406 30994 33458 31006
rect 33406 30930 33458 30942
rect 34302 30994 34354 31006
rect 34302 30930 34354 30942
rect 34638 30994 34690 31006
rect 34638 30930 34690 30942
rect 35198 30994 35250 31006
rect 35198 30930 35250 30942
rect 9662 30882 9714 30894
rect 14926 30882 14978 30894
rect 5170 30830 5182 30882
rect 5234 30830 5246 30882
rect 7298 30830 7310 30882
rect 7362 30830 7374 30882
rect 12786 30830 12798 30882
rect 12850 30830 12862 30882
rect 9662 30818 9714 30830
rect 14926 30818 14978 30830
rect 22654 30882 22706 30894
rect 25902 30882 25954 30894
rect 34750 30882 34802 30894
rect 23538 30830 23550 30882
rect 23602 30830 23614 30882
rect 28130 30830 28142 30882
rect 28194 30830 28206 30882
rect 30258 30830 30270 30882
rect 30322 30830 30334 30882
rect 30818 30830 30830 30882
rect 30882 30830 30894 30882
rect 22654 30818 22706 30830
rect 25902 30818 25954 30830
rect 34750 30818 34802 30830
rect 11118 30770 11170 30782
rect 11118 30706 11170 30718
rect 16830 30770 16882 30782
rect 16830 30706 16882 30718
rect 18622 30770 18674 30782
rect 18622 30706 18674 30718
rect 25342 30770 25394 30782
rect 25342 30706 25394 30718
rect 32398 30770 32450 30782
rect 32398 30706 32450 30718
rect 1344 30602 35616 30636
rect 1344 30550 5498 30602
rect 5550 30550 5602 30602
rect 5654 30550 5706 30602
rect 5758 30550 14066 30602
rect 14118 30550 14170 30602
rect 14222 30550 14274 30602
rect 14326 30550 22634 30602
rect 22686 30550 22738 30602
rect 22790 30550 22842 30602
rect 22894 30550 31202 30602
rect 31254 30550 31306 30602
rect 31358 30550 31410 30602
rect 31462 30550 35616 30602
rect 1344 30516 35616 30550
rect 15598 30434 15650 30446
rect 11778 30382 11790 30434
rect 11842 30382 11854 30434
rect 15598 30370 15650 30382
rect 20750 30434 20802 30446
rect 20750 30370 20802 30382
rect 21758 30434 21810 30446
rect 33618 30382 33630 30434
rect 33682 30431 33694 30434
rect 34290 30431 34302 30434
rect 33682 30385 34302 30431
rect 33682 30382 33694 30385
rect 34290 30382 34302 30385
rect 34354 30382 34366 30434
rect 21758 30370 21810 30382
rect 20414 30322 20466 30334
rect 9202 30270 9214 30322
rect 9266 30270 9278 30322
rect 18834 30270 18846 30322
rect 18898 30270 18910 30322
rect 20414 30258 20466 30270
rect 27694 30322 27746 30334
rect 32498 30270 32510 30322
rect 32562 30270 32574 30322
rect 27694 30258 27746 30270
rect 6414 30210 6466 30222
rect 13582 30210 13634 30222
rect 23326 30210 23378 30222
rect 28590 30210 28642 30222
rect 7074 30158 7086 30210
rect 7138 30158 7150 30210
rect 9314 30158 9326 30210
rect 9378 30158 9390 30210
rect 9538 30158 9550 30210
rect 9602 30158 9614 30210
rect 10434 30158 10446 30210
rect 10498 30158 10510 30210
rect 14578 30158 14590 30210
rect 14642 30158 14654 30210
rect 17490 30158 17502 30210
rect 17554 30158 17566 30210
rect 20738 30158 20750 30210
rect 20802 30158 20814 30210
rect 21858 30158 21870 30210
rect 21922 30158 21934 30210
rect 24210 30158 24222 30210
rect 24274 30158 24286 30210
rect 6414 30146 6466 30158
rect 13582 30146 13634 30158
rect 23326 30146 23378 30158
rect 28590 30146 28642 30158
rect 29262 30210 29314 30222
rect 29698 30158 29710 30210
rect 29762 30158 29774 30210
rect 30370 30158 30382 30210
rect 30434 30158 30446 30210
rect 29262 30146 29314 30158
rect 5742 30098 5794 30110
rect 5742 30034 5794 30046
rect 8206 30098 8258 30110
rect 8206 30034 8258 30046
rect 9774 30098 9826 30110
rect 9774 30034 9826 30046
rect 13470 30098 13522 30110
rect 13470 30034 13522 30046
rect 21310 30098 21362 30110
rect 23102 30098 23154 30110
rect 21522 30046 21534 30098
rect 21586 30046 21598 30098
rect 21310 30034 21362 30046
rect 23102 30034 23154 30046
rect 23662 30098 23714 30110
rect 34862 30098 34914 30110
rect 24882 30046 24894 30098
rect 24946 30046 24958 30098
rect 23662 30034 23714 30046
rect 34862 30034 34914 30046
rect 5630 29986 5682 29998
rect 5630 29922 5682 29934
rect 6526 29986 6578 29998
rect 6526 29922 6578 29934
rect 6750 29986 6802 29998
rect 8990 29986 9042 29998
rect 7298 29934 7310 29986
rect 7362 29934 7374 29986
rect 7858 29934 7870 29986
rect 7922 29934 7934 29986
rect 6750 29922 6802 29934
rect 8990 29922 9042 29934
rect 9998 29986 10050 29998
rect 9998 29922 10050 29934
rect 14254 29986 14306 29998
rect 22654 29986 22706 29998
rect 21746 29934 21758 29986
rect 21810 29934 21822 29986
rect 14254 29922 14306 29934
rect 22654 29922 22706 29934
rect 23214 29986 23266 29998
rect 33182 29986 33234 29998
rect 27122 29934 27134 29986
rect 27186 29934 27198 29986
rect 23214 29922 23266 29934
rect 33182 29922 33234 29934
rect 33630 29986 33682 29998
rect 33630 29922 33682 29934
rect 34078 29986 34130 29998
rect 34078 29922 34130 29934
rect 34638 29986 34690 29998
rect 34638 29922 34690 29934
rect 35198 29986 35250 29998
rect 35198 29922 35250 29934
rect 1344 29818 35776 29852
rect 1344 29766 9782 29818
rect 9834 29766 9886 29818
rect 9938 29766 9990 29818
rect 10042 29766 18350 29818
rect 18402 29766 18454 29818
rect 18506 29766 18558 29818
rect 18610 29766 26918 29818
rect 26970 29766 27022 29818
rect 27074 29766 27126 29818
rect 27178 29766 35486 29818
rect 35538 29766 35590 29818
rect 35642 29766 35694 29818
rect 35746 29766 35776 29818
rect 1344 29732 35776 29766
rect 8878 29650 8930 29662
rect 8878 29586 8930 29598
rect 10110 29650 10162 29662
rect 10110 29586 10162 29598
rect 10334 29650 10386 29662
rect 10334 29586 10386 29598
rect 12574 29650 12626 29662
rect 12574 29586 12626 29598
rect 14030 29650 14082 29662
rect 14030 29586 14082 29598
rect 16382 29650 16434 29662
rect 16382 29586 16434 29598
rect 17838 29650 17890 29662
rect 17838 29586 17890 29598
rect 19070 29650 19122 29662
rect 19070 29586 19122 29598
rect 24110 29650 24162 29662
rect 24110 29586 24162 29598
rect 26238 29650 26290 29662
rect 26238 29586 26290 29598
rect 34190 29650 34242 29662
rect 34190 29586 34242 29598
rect 34414 29650 34466 29662
rect 34414 29586 34466 29598
rect 8430 29538 8482 29550
rect 4610 29486 4622 29538
rect 4674 29486 4686 29538
rect 8430 29474 8482 29486
rect 11454 29538 11506 29550
rect 18286 29538 18338 29550
rect 12226 29486 12238 29538
rect 12290 29486 12302 29538
rect 11454 29474 11506 29486
rect 18286 29474 18338 29486
rect 18846 29538 18898 29550
rect 34526 29538 34578 29550
rect 20178 29486 20190 29538
rect 20242 29486 20254 29538
rect 21186 29486 21198 29538
rect 21250 29486 21262 29538
rect 34850 29486 34862 29538
rect 34914 29486 34926 29538
rect 18846 29474 18898 29486
rect 34526 29474 34578 29486
rect 7198 29426 7250 29438
rect 11230 29426 11282 29438
rect 3938 29374 3950 29426
rect 4002 29374 4014 29426
rect 7634 29374 7646 29426
rect 7698 29374 7710 29426
rect 8642 29374 8654 29426
rect 8706 29374 8718 29426
rect 9538 29374 9550 29426
rect 9602 29374 9614 29426
rect 9874 29374 9886 29426
rect 9938 29374 9950 29426
rect 7198 29362 7250 29374
rect 11230 29362 11282 29374
rect 11342 29426 11394 29438
rect 16158 29426 16210 29438
rect 13010 29374 13022 29426
rect 13074 29374 13086 29426
rect 11342 29362 11394 29374
rect 16158 29362 16210 29374
rect 16270 29426 16322 29438
rect 16270 29362 16322 29374
rect 16830 29426 16882 29438
rect 16830 29362 16882 29374
rect 17278 29426 17330 29438
rect 18622 29426 18674 29438
rect 17602 29374 17614 29426
rect 17666 29374 17678 29426
rect 20626 29374 20638 29426
rect 20690 29374 20702 29426
rect 22754 29374 22766 29426
rect 22818 29374 22830 29426
rect 25218 29374 25230 29426
rect 25282 29374 25294 29426
rect 29250 29374 29262 29426
rect 29314 29374 29326 29426
rect 33730 29374 33742 29426
rect 33794 29374 33806 29426
rect 35074 29374 35086 29426
rect 35138 29374 35150 29426
rect 17278 29362 17330 29374
rect 18622 29362 18674 29374
rect 8094 29314 8146 29326
rect 10894 29314 10946 29326
rect 6738 29262 6750 29314
rect 6802 29262 6814 29314
rect 9986 29262 9998 29314
rect 10050 29262 10062 29314
rect 8094 29250 8146 29262
rect 10894 29250 10946 29262
rect 16606 29314 16658 29326
rect 16606 29250 16658 29262
rect 18062 29314 18114 29326
rect 18062 29250 18114 29262
rect 18734 29314 18786 29326
rect 18734 29250 18786 29262
rect 23214 29314 23266 29326
rect 23214 29250 23266 29262
rect 23774 29314 23826 29326
rect 23774 29250 23826 29262
rect 28926 29314 28978 29326
rect 32510 29314 32562 29326
rect 29922 29262 29934 29314
rect 29986 29262 29998 29314
rect 32050 29262 32062 29314
rect 32114 29262 32126 29314
rect 33842 29262 33854 29314
rect 33906 29262 33918 29314
rect 28926 29250 28978 29262
rect 32510 29250 32562 29262
rect 8990 29202 9042 29214
rect 17838 29202 17890 29214
rect 11890 29150 11902 29202
rect 11954 29150 11966 29202
rect 8990 29138 9042 29150
rect 17838 29138 17890 29150
rect 20862 29202 20914 29214
rect 33282 29150 33294 29202
rect 33346 29150 33358 29202
rect 20862 29138 20914 29150
rect 1344 29034 35616 29068
rect 1344 28982 5498 29034
rect 5550 28982 5602 29034
rect 5654 28982 5706 29034
rect 5758 28982 14066 29034
rect 14118 28982 14170 29034
rect 14222 28982 14274 29034
rect 14326 28982 22634 29034
rect 22686 28982 22738 29034
rect 22790 28982 22842 29034
rect 22894 28982 31202 29034
rect 31254 28982 31306 29034
rect 31358 28982 31410 29034
rect 31462 28982 35616 29034
rect 1344 28948 35616 28982
rect 6862 28866 6914 28878
rect 6862 28802 6914 28814
rect 7198 28866 7250 28878
rect 7198 28802 7250 28814
rect 15598 28866 15650 28878
rect 16482 28814 16494 28866
rect 16546 28814 16558 28866
rect 21858 28814 21870 28866
rect 21922 28814 21934 28866
rect 15598 28802 15650 28814
rect 6526 28754 6578 28766
rect 6526 28690 6578 28702
rect 7646 28754 7698 28766
rect 11006 28754 11058 28766
rect 9090 28702 9102 28754
rect 9154 28702 9166 28754
rect 9874 28702 9886 28754
rect 9938 28702 9950 28754
rect 7646 28690 7698 28702
rect 11006 28690 11058 28702
rect 11566 28754 11618 28766
rect 11566 28690 11618 28702
rect 12798 28754 12850 28766
rect 12798 28690 12850 28702
rect 13582 28754 13634 28766
rect 13582 28690 13634 28702
rect 15374 28754 15426 28766
rect 17726 28754 17778 28766
rect 28478 28754 28530 28766
rect 15922 28702 15934 28754
rect 15986 28702 15998 28754
rect 19394 28702 19406 28754
rect 19458 28702 19470 28754
rect 25890 28702 25902 28754
rect 25954 28702 25966 28754
rect 32162 28702 32174 28754
rect 32226 28702 32238 28754
rect 15374 28690 15426 28702
rect 17726 28690 17778 28702
rect 28478 28690 28530 28702
rect 8318 28642 8370 28654
rect 10222 28642 10274 28654
rect 6850 28590 6862 28642
rect 6914 28590 6926 28642
rect 8978 28590 8990 28642
rect 9042 28590 9054 28642
rect 9426 28590 9438 28642
rect 9490 28590 9502 28642
rect 8318 28578 8370 28590
rect 10222 28578 10274 28590
rect 10782 28642 10834 28654
rect 10782 28578 10834 28590
rect 11230 28642 11282 28654
rect 15038 28642 15090 28654
rect 14242 28590 14254 28642
rect 14306 28590 14318 28642
rect 11230 28578 11282 28590
rect 15038 28578 15090 28590
rect 17054 28642 17106 28654
rect 17054 28578 17106 28590
rect 17166 28642 17218 28654
rect 17166 28578 17218 28590
rect 17502 28642 17554 28654
rect 17502 28578 17554 28590
rect 17838 28642 17890 28654
rect 17838 28578 17890 28590
rect 18062 28642 18114 28654
rect 18062 28578 18114 28590
rect 18958 28642 19010 28654
rect 20078 28642 20130 28654
rect 19506 28590 19518 28642
rect 19570 28590 19582 28642
rect 18958 28578 19010 28590
rect 20078 28578 20130 28590
rect 20190 28642 20242 28654
rect 20514 28590 20526 28642
rect 20578 28590 20590 28642
rect 21522 28590 21534 28642
rect 21586 28590 21598 28642
rect 21970 28590 21982 28642
rect 22034 28590 22046 28642
rect 23762 28590 23774 28642
rect 23826 28590 23838 28642
rect 29138 28590 29150 28642
rect 29202 28590 29214 28642
rect 34962 28590 34974 28642
rect 35026 28590 35038 28642
rect 20190 28578 20242 28590
rect 8654 28530 8706 28542
rect 8654 28466 8706 28478
rect 9886 28530 9938 28542
rect 9886 28466 9938 28478
rect 9998 28530 10050 28542
rect 9998 28466 10050 28478
rect 10558 28530 10610 28542
rect 10558 28466 10610 28478
rect 12686 28530 12738 28542
rect 12686 28466 12738 28478
rect 12910 28530 12962 28542
rect 12910 28466 12962 28478
rect 13806 28530 13858 28542
rect 13806 28466 13858 28478
rect 16942 28530 16994 28542
rect 16942 28466 16994 28478
rect 19854 28530 19906 28542
rect 19854 28466 19906 28478
rect 21310 28530 21362 28542
rect 21310 28466 21362 28478
rect 8542 28418 8594 28430
rect 8542 28354 8594 28366
rect 13470 28418 13522 28430
rect 13470 28354 13522 28366
rect 13694 28418 13746 28430
rect 19070 28418 19122 28430
rect 14690 28366 14702 28418
rect 14754 28366 14766 28418
rect 13694 28354 13746 28366
rect 19070 28354 19122 28366
rect 19294 28418 19346 28430
rect 19294 28354 19346 28366
rect 20302 28418 20354 28430
rect 20302 28354 20354 28366
rect 22094 28418 22146 28430
rect 22094 28354 22146 28366
rect 28366 28418 28418 28430
rect 34738 28366 34750 28418
rect 34802 28366 34814 28418
rect 28366 28354 28418 28366
rect 1344 28250 35776 28284
rect 1344 28198 9782 28250
rect 9834 28198 9886 28250
rect 9938 28198 9990 28250
rect 10042 28198 18350 28250
rect 18402 28198 18454 28250
rect 18506 28198 18558 28250
rect 18610 28198 26918 28250
rect 26970 28198 27022 28250
rect 27074 28198 27126 28250
rect 27178 28198 35486 28250
rect 35538 28198 35590 28250
rect 35642 28198 35694 28250
rect 35746 28198 35776 28250
rect 1344 28164 35776 28198
rect 7086 28082 7138 28094
rect 7086 28018 7138 28030
rect 8542 28082 8594 28094
rect 12686 28082 12738 28094
rect 10658 28030 10670 28082
rect 10722 28030 10734 28082
rect 8542 28018 8594 28030
rect 12686 28018 12738 28030
rect 13582 28082 13634 28094
rect 19406 28082 19458 28094
rect 21646 28082 21698 28094
rect 13582 28018 13634 28030
rect 17726 28026 17778 28038
rect 8094 27970 8146 27982
rect 8094 27906 8146 27918
rect 9774 27970 9826 27982
rect 9774 27906 9826 27918
rect 11902 27970 11954 27982
rect 11902 27906 11954 27918
rect 12014 27970 12066 27982
rect 12014 27906 12066 27918
rect 14254 27970 14306 27982
rect 15038 27970 15090 27982
rect 14914 27918 14926 27970
rect 14978 27918 14990 27970
rect 14254 27906 14306 27918
rect 15038 27906 15090 27918
rect 15150 27970 15202 27982
rect 15150 27906 15202 27918
rect 16046 27970 16098 27982
rect 17390 27970 17442 27982
rect 16370 27918 16382 27970
rect 16434 27918 16446 27970
rect 16046 27906 16098 27918
rect 17390 27906 17442 27918
rect 17614 27970 17666 27982
rect 19730 28030 19742 28082
rect 19794 28030 19806 28082
rect 19406 28018 19458 28030
rect 21646 28018 21698 28030
rect 23102 28082 23154 28094
rect 23102 28018 23154 28030
rect 30382 28082 30434 28094
rect 34738 28030 34750 28082
rect 34802 28030 34814 28082
rect 30382 28018 30434 28030
rect 17726 27962 17778 27974
rect 18734 27970 18786 27982
rect 17614 27906 17666 27918
rect 18734 27906 18786 27918
rect 20078 27970 20130 27982
rect 20078 27906 20130 27918
rect 21758 27970 21810 27982
rect 32062 27970 32114 27982
rect 29250 27918 29262 27970
rect 29314 27918 29326 27970
rect 21758 27906 21810 27918
rect 32062 27906 32114 27918
rect 32174 27970 32226 27982
rect 32174 27906 32226 27918
rect 33070 27970 33122 27982
rect 33070 27906 33122 27918
rect 6862 27858 6914 27870
rect 9550 27858 9602 27870
rect 13358 27858 13410 27870
rect 3602 27806 3614 27858
rect 3666 27806 3678 27858
rect 7410 27806 7422 27858
rect 7474 27806 7486 27858
rect 7858 27806 7870 27858
rect 7922 27806 7934 27858
rect 9986 27806 9998 27858
rect 10050 27806 10062 27858
rect 10322 27806 10334 27858
rect 10386 27806 10398 27858
rect 10882 27806 10894 27858
rect 10946 27806 10958 27858
rect 12450 27806 12462 27858
rect 12514 27806 12526 27858
rect 13122 27806 13134 27858
rect 13186 27806 13198 27858
rect 6862 27794 6914 27806
rect 9550 27794 9602 27806
rect 13358 27794 13410 27806
rect 13694 27858 13746 27870
rect 13694 27794 13746 27806
rect 15374 27858 15426 27870
rect 15374 27794 15426 27806
rect 15822 27858 15874 27870
rect 18174 27858 18226 27870
rect 16258 27806 16270 27858
rect 16322 27806 16334 27858
rect 15822 27794 15874 27806
rect 18174 27794 18226 27806
rect 20414 27858 20466 27870
rect 20414 27794 20466 27806
rect 20638 27858 20690 27870
rect 21422 27858 21474 27870
rect 30494 27858 30546 27870
rect 20962 27806 20974 27858
rect 21026 27806 21038 27858
rect 22306 27806 22318 27858
rect 22370 27806 22382 27858
rect 25218 27806 25230 27858
rect 25282 27806 25294 27858
rect 26226 27806 26238 27858
rect 26290 27806 26302 27858
rect 29922 27806 29934 27858
rect 29986 27806 29998 27858
rect 20638 27794 20690 27806
rect 21422 27794 21474 27806
rect 30494 27794 30546 27806
rect 31054 27858 31106 27870
rect 32398 27858 32450 27870
rect 35086 27858 35138 27870
rect 31602 27806 31614 27858
rect 31666 27806 31678 27858
rect 33394 27806 33406 27858
rect 33458 27806 33470 27858
rect 34290 27806 34302 27858
rect 34354 27806 34366 27858
rect 31054 27794 31106 27806
rect 32398 27794 32450 27806
rect 35086 27794 35138 27806
rect 6974 27746 7026 27758
rect 20526 27746 20578 27758
rect 4274 27694 4286 27746
rect 4338 27694 4350 27746
rect 6402 27694 6414 27746
rect 6466 27694 6478 27746
rect 9874 27694 9886 27746
rect 9938 27694 9950 27746
rect 13234 27694 13246 27746
rect 13298 27694 13310 27746
rect 14578 27694 14590 27746
rect 14642 27694 14654 27746
rect 16594 27694 16606 27746
rect 16658 27694 16670 27746
rect 6974 27682 7026 27694
rect 20526 27682 20578 27694
rect 21310 27746 21362 27758
rect 31278 27746 31330 27758
rect 25554 27694 25566 27746
rect 25618 27694 25630 27746
rect 25778 27694 25790 27746
rect 25842 27694 25854 27746
rect 27122 27694 27134 27746
rect 27186 27694 27198 27746
rect 32050 27694 32062 27746
rect 32114 27694 32126 27746
rect 33282 27694 33294 27746
rect 33346 27694 33358 27746
rect 33954 27694 33966 27746
rect 34018 27694 34030 27746
rect 21310 27682 21362 27694
rect 31278 27682 31330 27694
rect 12014 27634 12066 27646
rect 12014 27570 12066 27582
rect 12798 27634 12850 27646
rect 12798 27570 12850 27582
rect 18398 27634 18450 27646
rect 18398 27570 18450 27582
rect 18846 27634 18898 27646
rect 18846 27570 18898 27582
rect 18958 27634 19010 27646
rect 18958 27570 19010 27582
rect 30718 27634 30770 27646
rect 30718 27570 30770 27582
rect 1344 27466 35616 27500
rect 1344 27414 5498 27466
rect 5550 27414 5602 27466
rect 5654 27414 5706 27466
rect 5758 27414 14066 27466
rect 14118 27414 14170 27466
rect 14222 27414 14274 27466
rect 14326 27414 22634 27466
rect 22686 27414 22738 27466
rect 22790 27414 22842 27466
rect 22894 27414 31202 27466
rect 31254 27414 31306 27466
rect 31358 27414 31410 27466
rect 31462 27414 35616 27466
rect 1344 27380 35616 27414
rect 5630 27298 5682 27310
rect 5630 27234 5682 27246
rect 5966 27298 6018 27310
rect 15486 27298 15538 27310
rect 9538 27246 9550 27298
rect 9602 27246 9614 27298
rect 5966 27234 6018 27246
rect 15486 27234 15538 27246
rect 19742 27298 19794 27310
rect 30594 27246 30606 27298
rect 30658 27246 30670 27298
rect 19742 27234 19794 27246
rect 7534 27186 7586 27198
rect 13806 27186 13858 27198
rect 9874 27134 9886 27186
rect 9938 27134 9950 27186
rect 7534 27122 7586 27134
rect 13806 27122 13858 27134
rect 15374 27186 15426 27198
rect 15374 27122 15426 27134
rect 16158 27186 16210 27198
rect 26562 27134 26574 27186
rect 26626 27134 26638 27186
rect 27458 27134 27470 27186
rect 27522 27134 27534 27186
rect 28018 27134 28030 27186
rect 28082 27134 28094 27186
rect 35186 27134 35198 27186
rect 35250 27134 35262 27186
rect 16158 27122 16210 27134
rect 6302 27074 6354 27086
rect 6302 27010 6354 27022
rect 6526 27074 6578 27086
rect 6526 27010 6578 27022
rect 6974 27074 7026 27086
rect 8542 27074 8594 27086
rect 7186 27022 7198 27074
rect 7250 27022 7262 27074
rect 6974 27010 7026 27022
rect 8542 27010 8594 27022
rect 8990 27074 9042 27086
rect 10894 27074 10946 27086
rect 10098 27022 10110 27074
rect 10162 27022 10174 27074
rect 8990 27010 9042 27022
rect 10894 27010 10946 27022
rect 11006 27074 11058 27086
rect 11006 27010 11058 27022
rect 11454 27074 11506 27086
rect 11454 27010 11506 27022
rect 12238 27074 12290 27086
rect 12238 27010 12290 27022
rect 12574 27074 12626 27086
rect 12574 27010 12626 27022
rect 14030 27074 14082 27086
rect 14030 27010 14082 27022
rect 14366 27074 14418 27086
rect 14366 27010 14418 27022
rect 18174 27074 18226 27086
rect 18174 27010 18226 27022
rect 18510 27074 18562 27086
rect 18510 27010 18562 27022
rect 18622 27074 18674 27086
rect 18622 27010 18674 27022
rect 18958 27074 19010 27086
rect 18958 27010 19010 27022
rect 19630 27074 19682 27086
rect 19630 27010 19682 27022
rect 20526 27074 20578 27086
rect 20526 27010 20578 27022
rect 20750 27074 20802 27086
rect 22206 27074 22258 27086
rect 22654 27074 22706 27086
rect 21858 27022 21870 27074
rect 21922 27022 21934 27074
rect 22418 27022 22430 27074
rect 22482 27022 22494 27074
rect 20750 27010 20802 27022
rect 22206 27010 22258 27022
rect 22654 27010 22706 27022
rect 23326 27074 23378 27086
rect 23762 27022 23774 27074
rect 23826 27022 23838 27074
rect 28354 27022 28366 27074
rect 28418 27022 28430 27074
rect 29138 27022 29150 27074
rect 29202 27022 29214 27074
rect 32274 27022 32286 27074
rect 32338 27022 32350 27074
rect 23326 27010 23378 27022
rect 8430 26962 8482 26974
rect 13470 26962 13522 26974
rect 11890 26910 11902 26962
rect 11954 26910 11966 26962
rect 12898 26910 12910 26962
rect 12962 26910 12974 26962
rect 8430 26898 8482 26910
rect 13470 26898 13522 26910
rect 14590 26962 14642 26974
rect 14590 26898 14642 26910
rect 14702 26962 14754 26974
rect 14702 26898 14754 26910
rect 15262 26962 15314 26974
rect 15262 26898 15314 26910
rect 16830 26962 16882 26974
rect 16830 26898 16882 26910
rect 17166 26962 17218 26974
rect 17166 26898 17218 26910
rect 18286 26962 18338 26974
rect 5742 26850 5794 26862
rect 5742 26786 5794 26798
rect 6414 26850 6466 26862
rect 6414 26786 6466 26798
rect 7422 26850 7474 26862
rect 7422 26786 7474 26798
rect 7646 26850 7698 26862
rect 7646 26786 7698 26798
rect 7758 26850 7810 26862
rect 7758 26786 7810 26798
rect 8318 26850 8370 26862
rect 8318 26786 8370 26798
rect 11230 26850 11282 26862
rect 11230 26786 11282 26798
rect 13694 26850 13746 26862
rect 13694 26786 13746 26798
rect 13918 26850 13970 26862
rect 13918 26786 13970 26798
rect 17502 26850 17554 26862
rect 17826 26854 17838 26906
rect 17890 26854 17902 26906
rect 18286 26898 18338 26910
rect 18846 26962 18898 26974
rect 18846 26898 18898 26910
rect 19742 26962 19794 26974
rect 19742 26898 19794 26910
rect 20190 26962 20242 26974
rect 20190 26898 20242 26910
rect 21310 26962 21362 26974
rect 21310 26898 21362 26910
rect 22542 26962 22594 26974
rect 27022 26962 27074 26974
rect 24434 26910 24446 26962
rect 24498 26910 24510 26962
rect 33058 26910 33070 26962
rect 33122 26910 33134 26962
rect 22542 26898 22594 26910
rect 27022 26898 27074 26910
rect 17502 26786 17554 26798
rect 20414 26850 20466 26862
rect 20414 26786 20466 26798
rect 21422 26850 21474 26862
rect 21422 26786 21474 26798
rect 21646 26850 21698 26862
rect 21646 26786 21698 26798
rect 1344 26682 35776 26716
rect 1344 26630 9782 26682
rect 9834 26630 9886 26682
rect 9938 26630 9990 26682
rect 10042 26630 18350 26682
rect 18402 26630 18454 26682
rect 18506 26630 18558 26682
rect 18610 26630 26918 26682
rect 26970 26630 27022 26682
rect 27074 26630 27126 26682
rect 27178 26630 35486 26682
rect 35538 26630 35590 26682
rect 35642 26630 35694 26682
rect 35746 26630 35776 26682
rect 1344 26596 35776 26630
rect 8430 26514 8482 26526
rect 8430 26450 8482 26462
rect 9550 26514 9602 26526
rect 9550 26450 9602 26462
rect 9662 26514 9714 26526
rect 9662 26450 9714 26462
rect 9774 26514 9826 26526
rect 22542 26514 22594 26526
rect 17378 26462 17390 26514
rect 17442 26462 17454 26514
rect 18386 26462 18398 26514
rect 18450 26462 18462 26514
rect 18722 26462 18734 26514
rect 18786 26462 18798 26514
rect 20850 26462 20862 26514
rect 20914 26462 20926 26514
rect 9774 26450 9826 26462
rect 22542 26450 22594 26462
rect 22654 26514 22706 26526
rect 22654 26450 22706 26462
rect 24670 26514 24722 26526
rect 24670 26450 24722 26462
rect 25566 26514 25618 26526
rect 25566 26450 25618 26462
rect 27582 26514 27634 26526
rect 27582 26450 27634 26462
rect 33070 26514 33122 26526
rect 33070 26450 33122 26462
rect 7422 26402 7474 26414
rect 7422 26338 7474 26350
rect 7534 26402 7586 26414
rect 7534 26338 7586 26350
rect 7646 26402 7698 26414
rect 7646 26338 7698 26350
rect 7982 26402 8034 26414
rect 7982 26338 8034 26350
rect 9886 26402 9938 26414
rect 9886 26338 9938 26350
rect 12462 26402 12514 26414
rect 12462 26338 12514 26350
rect 12686 26402 12738 26414
rect 12686 26338 12738 26350
rect 13582 26402 13634 26414
rect 19742 26402 19794 26414
rect 16482 26350 16494 26402
rect 16546 26350 16558 26402
rect 13582 26338 13634 26350
rect 19742 26338 19794 26350
rect 20078 26402 20130 26414
rect 20078 26338 20130 26350
rect 23886 26402 23938 26414
rect 23886 26338 23938 26350
rect 25678 26402 25730 26414
rect 33966 26402 34018 26414
rect 29922 26350 29934 26402
rect 29986 26350 29998 26402
rect 25678 26338 25730 26350
rect 33966 26338 34018 26350
rect 34414 26402 34466 26414
rect 34414 26338 34466 26350
rect 34526 26402 34578 26414
rect 34850 26350 34862 26402
rect 34914 26350 34926 26402
rect 34526 26338 34578 26350
rect 8318 26290 8370 26302
rect 3602 26238 3614 26290
rect 3666 26238 3678 26290
rect 7074 26238 7086 26290
rect 7138 26238 7150 26290
rect 8318 26226 8370 26238
rect 8542 26290 8594 26302
rect 11566 26290 11618 26302
rect 10322 26238 10334 26290
rect 10386 26238 10398 26290
rect 11330 26238 11342 26290
rect 11394 26238 11406 26290
rect 8542 26226 8594 26238
rect 11566 26226 11618 26238
rect 12126 26290 12178 26302
rect 12126 26226 12178 26238
rect 13358 26290 13410 26302
rect 13358 26226 13410 26238
rect 13806 26290 13858 26302
rect 13806 26226 13858 26238
rect 15262 26290 15314 26302
rect 15262 26226 15314 26238
rect 16158 26290 16210 26302
rect 17726 26290 17778 26302
rect 19070 26290 19122 26302
rect 16706 26238 16718 26290
rect 16770 26238 16782 26290
rect 18162 26238 18174 26290
rect 18226 26238 18238 26290
rect 16158 26226 16210 26238
rect 17726 26226 17778 26238
rect 19070 26226 19122 26238
rect 20414 26290 20466 26302
rect 20862 26290 20914 26302
rect 22766 26290 22818 26302
rect 20626 26238 20638 26290
rect 20690 26238 20702 26290
rect 20962 26238 20974 26290
rect 21026 26238 21038 26290
rect 20414 26226 20466 26238
rect 20862 26226 20914 26238
rect 22766 26226 22818 26238
rect 23214 26290 23266 26302
rect 23214 26226 23266 26238
rect 23326 26290 23378 26302
rect 25342 26290 25394 26302
rect 33742 26290 33794 26302
rect 23650 26238 23662 26290
rect 23714 26238 23726 26290
rect 28130 26238 28142 26290
rect 28194 26238 28206 26290
rect 31490 26238 31502 26290
rect 31554 26238 31566 26290
rect 23326 26226 23378 26238
rect 25342 26226 25394 26238
rect 33742 26226 33794 26238
rect 34302 26290 34354 26302
rect 34738 26238 34750 26290
rect 34802 26238 34814 26290
rect 34302 26226 34354 26238
rect 13134 26178 13186 26190
rect 4386 26126 4398 26178
rect 4450 26126 4462 26178
rect 6514 26126 6526 26178
rect 6578 26126 6590 26178
rect 12674 26126 12686 26178
rect 12738 26126 12750 26178
rect 13134 26114 13186 26126
rect 14702 26178 14754 26190
rect 21758 26178 21810 26190
rect 32286 26178 32338 26190
rect 15698 26126 15710 26178
rect 15762 26126 15774 26178
rect 31938 26126 31950 26178
rect 32002 26126 32014 26178
rect 14702 26114 14754 26126
rect 21758 26114 21810 26126
rect 32286 26114 32338 26126
rect 11790 26066 11842 26078
rect 11790 26002 11842 26014
rect 11902 26066 11954 26078
rect 11902 26002 11954 26014
rect 13918 26066 13970 26078
rect 13918 26002 13970 26014
rect 21870 26066 21922 26078
rect 21870 26002 21922 26014
rect 22094 26066 22146 26078
rect 22094 26002 22146 26014
rect 22206 26066 22258 26078
rect 22206 26002 22258 26014
rect 23550 26066 23602 26078
rect 23550 26002 23602 26014
rect 33182 26066 33234 26078
rect 33182 26002 33234 26014
rect 33406 26066 33458 26078
rect 33406 26002 33458 26014
rect 1344 25898 35616 25932
rect 1344 25846 5498 25898
rect 5550 25846 5602 25898
rect 5654 25846 5706 25898
rect 5758 25846 14066 25898
rect 14118 25846 14170 25898
rect 14222 25846 14274 25898
rect 14326 25846 22634 25898
rect 22686 25846 22738 25898
rect 22790 25846 22842 25898
rect 22894 25846 31202 25898
rect 31254 25846 31306 25898
rect 31358 25846 31410 25898
rect 31462 25846 35616 25898
rect 1344 25812 35616 25846
rect 6190 25730 6242 25742
rect 6190 25666 6242 25678
rect 6526 25730 6578 25742
rect 12238 25730 12290 25742
rect 6962 25678 6974 25730
rect 7026 25727 7038 25730
rect 7410 25727 7422 25730
rect 7026 25681 7422 25727
rect 7026 25678 7038 25681
rect 7410 25678 7422 25681
rect 7474 25678 7486 25730
rect 10434 25678 10446 25730
rect 10498 25678 10510 25730
rect 6526 25666 6578 25678
rect 12238 25666 12290 25678
rect 13582 25730 13634 25742
rect 13582 25666 13634 25678
rect 19630 25730 19682 25742
rect 19630 25666 19682 25678
rect 21422 25730 21474 25742
rect 21422 25666 21474 25678
rect 21534 25730 21586 25742
rect 21534 25666 21586 25678
rect 28030 25730 28082 25742
rect 28030 25666 28082 25678
rect 29598 25730 29650 25742
rect 29598 25666 29650 25678
rect 30942 25730 30994 25742
rect 30942 25666 30994 25678
rect 7422 25618 7474 25630
rect 7422 25554 7474 25566
rect 17950 25618 18002 25630
rect 17950 25554 18002 25566
rect 18734 25618 18786 25630
rect 18734 25554 18786 25566
rect 19182 25618 19234 25630
rect 33406 25618 33458 25630
rect 22418 25566 22430 25618
rect 22482 25566 22494 25618
rect 26450 25566 26462 25618
rect 26514 25566 26526 25618
rect 28242 25566 28254 25618
rect 28306 25566 28318 25618
rect 34962 25566 34974 25618
rect 35026 25566 35038 25618
rect 19182 25554 19234 25566
rect 33406 25554 33458 25566
rect 7758 25506 7810 25518
rect 7758 25442 7810 25454
rect 9886 25506 9938 25518
rect 12126 25506 12178 25518
rect 10658 25454 10670 25506
rect 10722 25454 10734 25506
rect 9886 25442 9938 25454
rect 12126 25442 12178 25454
rect 12686 25506 12738 25518
rect 12686 25442 12738 25454
rect 13022 25506 13074 25518
rect 13022 25442 13074 25454
rect 13694 25506 13746 25518
rect 13694 25442 13746 25454
rect 14590 25506 14642 25518
rect 14590 25442 14642 25454
rect 14926 25506 14978 25518
rect 14926 25442 14978 25454
rect 15262 25506 15314 25518
rect 15262 25442 15314 25454
rect 17390 25506 17442 25518
rect 17390 25442 17442 25454
rect 17614 25506 17666 25518
rect 17614 25442 17666 25454
rect 18174 25506 18226 25518
rect 18174 25442 18226 25454
rect 19406 25506 19458 25518
rect 27806 25506 27858 25518
rect 23426 25454 23438 25506
rect 23490 25454 23502 25506
rect 27122 25454 27134 25506
rect 27186 25454 27198 25506
rect 19406 25442 19458 25454
rect 27806 25442 27858 25454
rect 29486 25506 29538 25518
rect 33630 25506 33682 25518
rect 29922 25454 29934 25506
rect 29986 25454 29998 25506
rect 29486 25442 29538 25454
rect 33630 25442 33682 25454
rect 6302 25394 6354 25406
rect 6302 25330 6354 25342
rect 7982 25394 8034 25406
rect 7982 25330 8034 25342
rect 8094 25394 8146 25406
rect 18846 25394 18898 25406
rect 21758 25394 21810 25406
rect 22318 25394 22370 25406
rect 28366 25394 28418 25406
rect 10098 25342 10110 25394
rect 10162 25342 10174 25394
rect 20402 25342 20414 25394
rect 20466 25342 20478 25394
rect 22082 25342 22094 25394
rect 22146 25342 22158 25394
rect 24210 25342 24222 25394
rect 24274 25342 24286 25394
rect 27346 25342 27358 25394
rect 27410 25342 27422 25394
rect 8094 25330 8146 25342
rect 18846 25330 18898 25342
rect 21758 25330 21810 25342
rect 22318 25330 22370 25342
rect 28366 25330 28418 25342
rect 28590 25394 28642 25406
rect 28590 25330 28642 25342
rect 32846 25394 32898 25406
rect 32846 25330 32898 25342
rect 33070 25394 33122 25406
rect 33070 25330 33122 25342
rect 33182 25394 33234 25406
rect 33182 25330 33234 25342
rect 6974 25282 7026 25294
rect 12238 25282 12290 25294
rect 10210 25230 10222 25282
rect 10274 25230 10286 25282
rect 6974 25218 7026 25230
rect 12238 25218 12290 25230
rect 12798 25282 12850 25294
rect 12798 25218 12850 25230
rect 13582 25282 13634 25294
rect 15038 25282 15090 25294
rect 14242 25230 14254 25282
rect 14306 25230 14318 25282
rect 13582 25218 13634 25230
rect 15038 25218 15090 25230
rect 17054 25282 17106 25294
rect 17054 25218 17106 25230
rect 18622 25282 18674 25294
rect 18622 25218 18674 25230
rect 20078 25282 20130 25294
rect 20078 25218 20130 25230
rect 20750 25282 20802 25294
rect 20750 25218 20802 25230
rect 23102 25282 23154 25294
rect 23102 25218 23154 25230
rect 29374 25282 29426 25294
rect 29374 25218 29426 25230
rect 34190 25282 34242 25294
rect 34190 25218 34242 25230
rect 34526 25282 34578 25294
rect 34526 25218 34578 25230
rect 1344 25114 35776 25148
rect 1344 25062 9782 25114
rect 9834 25062 9886 25114
rect 9938 25062 9990 25114
rect 10042 25062 18350 25114
rect 18402 25062 18454 25114
rect 18506 25062 18558 25114
rect 18610 25062 26918 25114
rect 26970 25062 27022 25114
rect 27074 25062 27126 25114
rect 27178 25062 35486 25114
rect 35538 25062 35590 25114
rect 35642 25062 35694 25114
rect 35746 25062 35776 25114
rect 1344 25028 35776 25062
rect 6974 24946 7026 24958
rect 6974 24882 7026 24894
rect 7534 24946 7586 24958
rect 7534 24882 7586 24894
rect 8094 24946 8146 24958
rect 8094 24882 8146 24894
rect 8654 24946 8706 24958
rect 8654 24882 8706 24894
rect 12574 24946 12626 24958
rect 12574 24882 12626 24894
rect 12798 24946 12850 24958
rect 12798 24882 12850 24894
rect 15262 24946 15314 24958
rect 19630 24946 19682 24958
rect 17378 24894 17390 24946
rect 17442 24894 17454 24946
rect 15262 24882 15314 24894
rect 19630 24882 19682 24894
rect 19742 24946 19794 24958
rect 19742 24882 19794 24894
rect 20078 24946 20130 24958
rect 20078 24882 20130 24894
rect 22990 24946 23042 24958
rect 22990 24882 23042 24894
rect 33070 24946 33122 24958
rect 33070 24882 33122 24894
rect 34302 24946 34354 24958
rect 34302 24882 34354 24894
rect 6750 24834 6802 24846
rect 6750 24770 6802 24782
rect 7310 24834 7362 24846
rect 7310 24770 7362 24782
rect 7870 24834 7922 24846
rect 7870 24770 7922 24782
rect 8430 24834 8482 24846
rect 8430 24770 8482 24782
rect 9550 24834 9602 24846
rect 9550 24770 9602 24782
rect 10446 24834 10498 24846
rect 10446 24770 10498 24782
rect 11566 24834 11618 24846
rect 11566 24770 11618 24782
rect 12238 24834 12290 24846
rect 12238 24770 12290 24782
rect 12350 24834 12402 24846
rect 12350 24770 12402 24782
rect 14814 24834 14866 24846
rect 14814 24770 14866 24782
rect 14926 24834 14978 24846
rect 14926 24770 14978 24782
rect 15486 24834 15538 24846
rect 15486 24770 15538 24782
rect 22878 24834 22930 24846
rect 29374 24834 29426 24846
rect 26002 24782 26014 24834
rect 26066 24782 26078 24834
rect 22878 24770 22930 24782
rect 29374 24770 29426 24782
rect 34526 24834 34578 24846
rect 34526 24770 34578 24782
rect 6638 24722 6690 24734
rect 6638 24658 6690 24670
rect 7198 24722 7250 24734
rect 7198 24658 7250 24670
rect 7758 24722 7810 24734
rect 7758 24658 7810 24670
rect 8318 24722 8370 24734
rect 8318 24658 8370 24670
rect 9886 24722 9938 24734
rect 9886 24658 9938 24670
rect 10334 24722 10386 24734
rect 10334 24658 10386 24670
rect 10670 24722 10722 24734
rect 10670 24658 10722 24670
rect 11342 24722 11394 24734
rect 11342 24658 11394 24670
rect 11678 24722 11730 24734
rect 11678 24658 11730 24670
rect 13134 24722 13186 24734
rect 14030 24722 14082 24734
rect 13570 24670 13582 24722
rect 13634 24670 13646 24722
rect 13134 24658 13186 24670
rect 14030 24658 14082 24670
rect 15150 24722 15202 24734
rect 15150 24658 15202 24670
rect 15598 24722 15650 24734
rect 15598 24658 15650 24670
rect 16158 24722 16210 24734
rect 16158 24658 16210 24670
rect 16718 24722 16770 24734
rect 16718 24658 16770 24670
rect 17726 24722 17778 24734
rect 17726 24658 17778 24670
rect 19854 24722 19906 24734
rect 22654 24722 22706 24734
rect 21074 24670 21086 24722
rect 21138 24670 21150 24722
rect 19854 24658 19906 24670
rect 22654 24658 22706 24670
rect 23326 24722 23378 24734
rect 29038 24722 29090 24734
rect 33182 24722 33234 24734
rect 25218 24670 25230 24722
rect 25282 24670 25294 24722
rect 32050 24670 32062 24722
rect 32114 24670 32126 24722
rect 23326 24658 23378 24670
rect 29038 24658 29090 24670
rect 33182 24658 33234 24670
rect 33742 24722 33794 24734
rect 34738 24670 34750 24722
rect 34802 24670 34814 24722
rect 35074 24670 35086 24722
rect 35138 24670 35150 24722
rect 33742 24658 33794 24670
rect 9102 24610 9154 24622
rect 9102 24546 9154 24558
rect 11118 24610 11170 24622
rect 11118 24546 11170 24558
rect 14478 24610 14530 24622
rect 14478 24546 14530 24558
rect 18174 24610 18226 24622
rect 23774 24610 23826 24622
rect 21970 24558 21982 24610
rect 22034 24558 22046 24610
rect 18174 24546 18226 24558
rect 23774 24546 23826 24558
rect 24334 24610 24386 24622
rect 24334 24546 24386 24558
rect 24782 24610 24834 24622
rect 33406 24610 33458 24622
rect 28130 24558 28142 24610
rect 28194 24558 28206 24610
rect 29362 24558 29374 24610
rect 29426 24558 29438 24610
rect 30258 24558 30270 24610
rect 30322 24558 30334 24610
rect 34626 24558 34638 24610
rect 34690 24558 34702 24610
rect 24782 24546 24834 24558
rect 33406 24546 33458 24558
rect 28814 24498 28866 24510
rect 28814 24434 28866 24446
rect 29598 24498 29650 24510
rect 29598 24434 29650 24446
rect 33966 24498 34018 24510
rect 33966 24434 34018 24446
rect 1344 24330 35616 24364
rect 1344 24278 5498 24330
rect 5550 24278 5602 24330
rect 5654 24278 5706 24330
rect 5758 24278 14066 24330
rect 14118 24278 14170 24330
rect 14222 24278 14274 24330
rect 14326 24278 22634 24330
rect 22686 24278 22738 24330
rect 22790 24278 22842 24330
rect 22894 24278 31202 24330
rect 31254 24278 31306 24330
rect 31358 24278 31410 24330
rect 31462 24278 35616 24330
rect 1344 24244 35616 24278
rect 23998 24162 24050 24174
rect 30818 24110 30830 24162
rect 30882 24110 30894 24162
rect 23998 24098 24050 24110
rect 28478 24050 28530 24062
rect 25554 23998 25566 24050
rect 25618 23998 25630 24050
rect 33058 23998 33070 24050
rect 33122 23998 33134 24050
rect 35186 23998 35198 24050
rect 35250 23998 35262 24050
rect 28478 23986 28530 23998
rect 23550 23938 23602 23950
rect 12898 23886 12910 23938
rect 12962 23886 12974 23938
rect 13570 23886 13582 23938
rect 13634 23886 13646 23938
rect 21522 23886 21534 23938
rect 21586 23886 21598 23938
rect 23550 23874 23602 23886
rect 23886 23938 23938 23950
rect 27134 23938 27186 23950
rect 25442 23886 25454 23938
rect 25506 23886 25518 23938
rect 23886 23874 23938 23886
rect 27134 23874 27186 23886
rect 28590 23938 28642 23950
rect 29362 23886 29374 23938
rect 29426 23886 29438 23938
rect 32386 23886 32398 23938
rect 32450 23886 32462 23938
rect 28590 23874 28642 23886
rect 7198 23826 7250 23838
rect 7198 23762 7250 23774
rect 7310 23826 7362 23838
rect 18958 23826 19010 23838
rect 7858 23774 7870 23826
rect 7922 23774 7934 23826
rect 15698 23774 15710 23826
rect 15762 23774 15774 23826
rect 7310 23762 7362 23774
rect 18958 23762 19010 23774
rect 19182 23826 19234 23838
rect 19182 23762 19234 23774
rect 19294 23826 19346 23838
rect 19294 23762 19346 23774
rect 21310 23826 21362 23838
rect 21310 23762 21362 23774
rect 21758 23826 21810 23838
rect 21758 23762 21810 23774
rect 24334 23826 24386 23838
rect 26126 23826 26178 23838
rect 28254 23826 28306 23838
rect 25106 23774 25118 23826
rect 25170 23774 25182 23826
rect 26786 23774 26798 23826
rect 26850 23774 26862 23826
rect 27458 23774 27470 23826
rect 27522 23774 27534 23826
rect 28130 23774 28142 23826
rect 28194 23774 28206 23826
rect 24334 23762 24386 23774
rect 26126 23762 26178 23774
rect 28254 23762 28306 23774
rect 6750 23714 6802 23726
rect 6750 23650 6802 23662
rect 6974 23714 7026 23726
rect 6974 23650 7026 23662
rect 19742 23714 19794 23726
rect 19742 23650 19794 23662
rect 21870 23714 21922 23726
rect 21870 23650 21922 23662
rect 22318 23714 22370 23726
rect 22318 23650 22370 23662
rect 24446 23714 24498 23726
rect 24446 23650 24498 23662
rect 24670 23714 24722 23726
rect 24670 23650 24722 23662
rect 25790 23714 25842 23726
rect 25790 23650 25842 23662
rect 26014 23714 26066 23726
rect 26014 23650 26066 23662
rect 26462 23714 26514 23726
rect 26462 23650 26514 23662
rect 28366 23714 28418 23726
rect 28366 23650 28418 23662
rect 1344 23546 35776 23580
rect 1344 23494 9782 23546
rect 9834 23494 9886 23546
rect 9938 23494 9990 23546
rect 10042 23494 18350 23546
rect 18402 23494 18454 23546
rect 18506 23494 18558 23546
rect 18610 23494 26918 23546
rect 26970 23494 27022 23546
rect 27074 23494 27126 23546
rect 27178 23494 35486 23546
rect 35538 23494 35590 23546
rect 35642 23494 35694 23546
rect 35746 23494 35776 23546
rect 1344 23460 35776 23494
rect 8206 23378 8258 23390
rect 8206 23314 8258 23326
rect 9102 23378 9154 23390
rect 9102 23314 9154 23326
rect 13806 23378 13858 23390
rect 13806 23314 13858 23326
rect 14254 23378 14306 23390
rect 14254 23314 14306 23326
rect 17726 23378 17778 23390
rect 17726 23314 17778 23326
rect 18398 23378 18450 23390
rect 18398 23314 18450 23326
rect 19406 23378 19458 23390
rect 19406 23314 19458 23326
rect 24334 23378 24386 23390
rect 24334 23314 24386 23326
rect 26350 23378 26402 23390
rect 28926 23378 28978 23390
rect 27346 23326 27358 23378
rect 27410 23326 27422 23378
rect 26350 23314 26402 23326
rect 28926 23314 28978 23326
rect 30942 23378 30994 23390
rect 30942 23314 30994 23326
rect 8094 23266 8146 23278
rect 8094 23202 8146 23214
rect 8878 23266 8930 23278
rect 8878 23202 8930 23214
rect 24558 23266 24610 23278
rect 24558 23202 24610 23214
rect 25454 23266 25506 23278
rect 25454 23202 25506 23214
rect 26574 23266 26626 23278
rect 26574 23202 26626 23214
rect 28030 23266 28082 23278
rect 28030 23202 28082 23214
rect 28254 23266 28306 23278
rect 28254 23202 28306 23214
rect 28478 23266 28530 23278
rect 28478 23202 28530 23214
rect 29038 23266 29090 23278
rect 33282 23214 33294 23266
rect 33346 23214 33358 23266
rect 29038 23202 29090 23214
rect 7086 23154 7138 23166
rect 3938 23102 3950 23154
rect 4002 23102 4014 23154
rect 7086 23090 7138 23102
rect 7534 23154 7586 23166
rect 7534 23090 7586 23102
rect 7758 23154 7810 23166
rect 7758 23090 7810 23102
rect 8430 23154 8482 23166
rect 8430 23090 8482 23102
rect 8766 23154 8818 23166
rect 8766 23090 8818 23102
rect 9438 23154 9490 23166
rect 9438 23090 9490 23102
rect 9774 23154 9826 23166
rect 9774 23090 9826 23102
rect 10110 23154 10162 23166
rect 17502 23154 17554 23166
rect 10546 23102 10558 23154
rect 10610 23102 10622 23154
rect 10110 23090 10162 23102
rect 17502 23090 17554 23102
rect 17726 23154 17778 23166
rect 17726 23090 17778 23102
rect 18062 23154 18114 23166
rect 18062 23090 18114 23102
rect 18174 23154 18226 23166
rect 18174 23090 18226 23102
rect 18510 23154 18562 23166
rect 18510 23090 18562 23102
rect 19294 23154 19346 23166
rect 23214 23154 23266 23166
rect 19954 23102 19966 23154
rect 20018 23102 20030 23154
rect 19294 23090 19346 23102
rect 23214 23090 23266 23102
rect 24670 23154 24722 23166
rect 24670 23090 24722 23102
rect 25566 23154 25618 23166
rect 25566 23090 25618 23102
rect 26126 23154 26178 23166
rect 26126 23090 26178 23102
rect 26238 23154 26290 23166
rect 26238 23090 26290 23102
rect 27022 23154 27074 23166
rect 27022 23090 27074 23102
rect 28814 23154 28866 23166
rect 29250 23102 29262 23154
rect 29314 23102 29326 23154
rect 29586 23102 29598 23154
rect 29650 23102 29662 23154
rect 29922 23102 29934 23154
rect 29986 23102 29998 23154
rect 33170 23102 33182 23154
rect 33234 23102 33246 23154
rect 34178 23102 34190 23154
rect 34242 23102 34254 23154
rect 28814 23090 28866 23102
rect 7310 23042 7362 23054
rect 4722 22990 4734 23042
rect 4786 22990 4798 23042
rect 6850 22990 6862 23042
rect 6914 22990 6926 23042
rect 7310 22978 7362 22990
rect 9662 23042 9714 23054
rect 23662 23042 23714 23054
rect 11218 22990 11230 23042
rect 11282 22990 11294 23042
rect 13346 22990 13358 23042
rect 13410 22990 13422 23042
rect 20626 22990 20638 23042
rect 20690 22990 20702 23042
rect 22754 22990 22766 23042
rect 22818 22990 22830 23042
rect 9662 22978 9714 22990
rect 23662 22978 23714 22990
rect 24110 23042 24162 23054
rect 33966 23042 34018 23054
rect 33618 22990 33630 23042
rect 33682 22990 33694 23042
rect 24110 22978 24162 22990
rect 33966 22978 34018 22990
rect 35198 23042 35250 23054
rect 35198 22978 35250 22990
rect 19406 22930 19458 22942
rect 19406 22866 19458 22878
rect 25454 22930 25506 22942
rect 25454 22866 25506 22878
rect 28366 22930 28418 22942
rect 28366 22866 28418 22878
rect 35086 22930 35138 22942
rect 35086 22866 35138 22878
rect 1344 22762 35616 22796
rect 1344 22710 5498 22762
rect 5550 22710 5602 22762
rect 5654 22710 5706 22762
rect 5758 22710 14066 22762
rect 14118 22710 14170 22762
rect 14222 22710 14274 22762
rect 14326 22710 22634 22762
rect 22686 22710 22738 22762
rect 22790 22710 22842 22762
rect 22894 22710 31202 22762
rect 31254 22710 31306 22762
rect 31358 22710 31410 22762
rect 31462 22710 35616 22762
rect 1344 22676 35616 22710
rect 19406 22594 19458 22606
rect 34974 22594 35026 22606
rect 26114 22542 26126 22594
rect 26178 22591 26190 22594
rect 26338 22591 26350 22594
rect 26178 22545 26350 22591
rect 26178 22542 26190 22545
rect 26338 22542 26350 22545
rect 26402 22542 26414 22594
rect 19406 22530 19458 22542
rect 34974 22530 35026 22542
rect 15710 22482 15762 22494
rect 30718 22482 30770 22494
rect 8194 22430 8206 22482
rect 8258 22430 8270 22482
rect 10322 22430 10334 22482
rect 10386 22430 10398 22482
rect 16818 22430 16830 22482
rect 16882 22430 16894 22482
rect 18946 22430 18958 22482
rect 19010 22430 19022 22482
rect 25778 22430 25790 22482
rect 25842 22430 25854 22482
rect 15710 22418 15762 22430
rect 30718 22418 30770 22430
rect 7086 22370 7138 22382
rect 10894 22370 10946 22382
rect 7522 22318 7534 22370
rect 7586 22318 7598 22370
rect 7086 22306 7138 22318
rect 10894 22306 10946 22318
rect 11342 22370 11394 22382
rect 21534 22370 21586 22382
rect 16034 22318 16046 22370
rect 16098 22318 16110 22370
rect 11342 22306 11394 22318
rect 21534 22306 21586 22318
rect 21870 22370 21922 22382
rect 30606 22370 30658 22382
rect 31614 22370 31666 22382
rect 22866 22318 22878 22370
rect 22930 22318 22942 22370
rect 27122 22318 27134 22370
rect 27186 22318 27198 22370
rect 27458 22318 27470 22370
rect 27522 22318 27534 22370
rect 27682 22318 27694 22370
rect 27746 22318 27758 22370
rect 28130 22318 28142 22370
rect 28194 22318 28206 22370
rect 29138 22318 29150 22370
rect 29202 22318 29214 22370
rect 31378 22318 31390 22370
rect 31442 22318 31454 22370
rect 31938 22318 31950 22370
rect 32002 22318 32014 22370
rect 33058 22318 33070 22370
rect 33122 22318 33134 22370
rect 21870 22306 21922 22318
rect 30606 22306 30658 22318
rect 31614 22306 31666 22318
rect 6526 22258 6578 22270
rect 6526 22194 6578 22206
rect 6862 22258 6914 22270
rect 6862 22194 6914 22206
rect 11566 22258 11618 22270
rect 11566 22194 11618 22206
rect 11902 22258 11954 22270
rect 11902 22194 11954 22206
rect 12014 22258 12066 22270
rect 12014 22194 12066 22206
rect 12462 22258 12514 22270
rect 12462 22194 12514 22206
rect 12798 22258 12850 22270
rect 12798 22194 12850 22206
rect 19294 22258 19346 22270
rect 19294 22194 19346 22206
rect 19406 22258 19458 22270
rect 19406 22194 19458 22206
rect 19966 22258 20018 22270
rect 19966 22194 20018 22206
rect 20302 22258 20354 22270
rect 20302 22194 20354 22206
rect 20750 22258 20802 22270
rect 20750 22194 20802 22206
rect 21310 22258 21362 22270
rect 30830 22258 30882 22270
rect 23650 22206 23662 22258
rect 23714 22206 23726 22258
rect 29474 22206 29486 22258
rect 29538 22206 29550 22258
rect 29922 22206 29934 22258
rect 29986 22206 29998 22258
rect 21310 22194 21362 22206
rect 30830 22194 30882 22206
rect 30942 22258 30994 22270
rect 30942 22194 30994 22206
rect 6638 22146 6690 22158
rect 6638 22082 6690 22094
rect 11230 22146 11282 22158
rect 11230 22082 11282 22094
rect 12238 22146 12290 22158
rect 12238 22082 12290 22094
rect 21646 22146 21698 22158
rect 21646 22082 21698 22094
rect 26238 22146 26290 22158
rect 26238 22082 26290 22094
rect 26462 22146 26514 22158
rect 26462 22082 26514 22094
rect 28366 22146 28418 22158
rect 28366 22082 28418 22094
rect 28590 22146 28642 22158
rect 28590 22082 28642 22094
rect 28702 22146 28754 22158
rect 32174 22146 32226 22158
rect 29698 22094 29710 22146
rect 29762 22094 29774 22146
rect 28702 22082 28754 22094
rect 32174 22082 32226 22094
rect 32286 22146 32338 22158
rect 32286 22082 32338 22094
rect 1344 21978 35776 22012
rect 1344 21926 9782 21978
rect 9834 21926 9886 21978
rect 9938 21926 9990 21978
rect 10042 21926 18350 21978
rect 18402 21926 18454 21978
rect 18506 21926 18558 21978
rect 18610 21926 26918 21978
rect 26970 21926 27022 21978
rect 27074 21926 27126 21978
rect 27178 21926 35486 21978
rect 35538 21926 35590 21978
rect 35642 21926 35694 21978
rect 35746 21926 35776 21978
rect 1344 21892 35776 21926
rect 7086 21810 7138 21822
rect 7086 21746 7138 21758
rect 7310 21810 7362 21822
rect 7310 21746 7362 21758
rect 7646 21810 7698 21822
rect 7646 21746 7698 21758
rect 7870 21810 7922 21822
rect 11902 21810 11954 21822
rect 17502 21810 17554 21822
rect 25230 21810 25282 21822
rect 10098 21758 10110 21810
rect 10162 21758 10174 21810
rect 12898 21758 12910 21810
rect 12962 21758 12974 21810
rect 21074 21758 21086 21810
rect 21138 21758 21150 21810
rect 7870 21746 7922 21758
rect 11902 21746 11954 21758
rect 17502 21746 17554 21758
rect 25230 21746 25282 21758
rect 25342 21810 25394 21822
rect 25342 21746 25394 21758
rect 25454 21810 25506 21822
rect 25454 21746 25506 21758
rect 34862 21810 34914 21822
rect 34862 21746 34914 21758
rect 11790 21698 11842 21710
rect 4386 21646 4398 21698
rect 4450 21646 4462 21698
rect 11790 21634 11842 21646
rect 13246 21698 13298 21710
rect 13246 21634 13298 21646
rect 13582 21698 13634 21710
rect 13582 21634 13634 21646
rect 24782 21698 24834 21710
rect 32062 21698 32114 21710
rect 28802 21646 28814 21698
rect 28866 21646 28878 21698
rect 29586 21646 29598 21698
rect 29650 21646 29662 21698
rect 24782 21634 24834 21646
rect 32062 21634 32114 21646
rect 32398 21698 32450 21710
rect 35086 21698 35138 21710
rect 34402 21646 34414 21698
rect 34466 21646 34478 21698
rect 32398 21634 32450 21646
rect 35086 21634 35138 21646
rect 35198 21698 35250 21710
rect 35198 21634 35250 21646
rect 7422 21586 7474 21598
rect 3714 21534 3726 21586
rect 3778 21534 3790 21586
rect 7422 21522 7474 21534
rect 7982 21586 8034 21598
rect 7982 21522 8034 21534
rect 8430 21586 8482 21598
rect 8430 21522 8482 21534
rect 10446 21586 10498 21598
rect 21422 21586 21474 21598
rect 12674 21534 12686 21586
rect 12738 21534 12750 21586
rect 13906 21534 13918 21586
rect 13970 21534 13982 21586
rect 20738 21534 20750 21586
rect 20802 21534 20814 21586
rect 10446 21522 10498 21534
rect 21422 21522 21474 21534
rect 25902 21586 25954 21598
rect 31502 21586 31554 21598
rect 26114 21534 26126 21586
rect 26178 21534 26190 21586
rect 27010 21534 27022 21586
rect 27074 21534 27086 21586
rect 27234 21534 27246 21586
rect 27298 21534 27310 21586
rect 27458 21534 27470 21586
rect 27522 21534 27534 21586
rect 29250 21534 29262 21586
rect 29314 21534 29326 21586
rect 31154 21534 31166 21586
rect 31218 21534 31230 21586
rect 33058 21534 33070 21586
rect 33122 21534 33134 21586
rect 33618 21534 33630 21586
rect 33682 21534 33694 21586
rect 34626 21534 34638 21586
rect 34690 21534 34702 21586
rect 25902 21522 25954 21534
rect 8878 21474 8930 21486
rect 6514 21422 6526 21474
rect 6578 21422 6590 21474
rect 8878 21410 8930 21422
rect 10894 21474 10946 21486
rect 21870 21474 21922 21486
rect 14690 21422 14702 21474
rect 14754 21422 14766 21474
rect 16818 21422 16830 21474
rect 16882 21422 16894 21474
rect 17826 21422 17838 21474
rect 17890 21422 17902 21474
rect 19954 21422 19966 21474
rect 20018 21422 20030 21474
rect 10894 21410 10946 21422
rect 21870 21410 21922 21422
rect 22542 21474 22594 21486
rect 22542 21410 22594 21422
rect 22990 21474 23042 21486
rect 22990 21410 23042 21422
rect 23326 21474 23378 21486
rect 23326 21410 23378 21422
rect 23774 21474 23826 21486
rect 23774 21410 23826 21422
rect 24222 21474 24274 21486
rect 25778 21422 25790 21474
rect 25842 21471 25854 21474
rect 26129 21471 26175 21534
rect 31502 21522 31554 21534
rect 33966 21474 34018 21486
rect 25842 21425 26175 21471
rect 25842 21422 25854 21425
rect 30034 21422 30046 21474
rect 30098 21422 30110 21474
rect 24222 21410 24274 21422
rect 33966 21410 34018 21422
rect 11902 21362 11954 21374
rect 32510 21362 32562 21374
rect 21634 21310 21646 21362
rect 21698 21359 21710 21362
rect 22978 21359 22990 21362
rect 21698 21313 22990 21359
rect 21698 21310 21710 21313
rect 22978 21310 22990 21313
rect 23042 21310 23054 21362
rect 23314 21310 23326 21362
rect 23378 21359 23390 21362
rect 23762 21359 23774 21362
rect 23378 21313 23774 21359
rect 23378 21310 23390 21313
rect 23762 21310 23774 21313
rect 23826 21310 23838 21362
rect 26450 21310 26462 21362
rect 26514 21310 26526 21362
rect 11902 21298 11954 21310
rect 32510 21298 32562 21310
rect 1344 21194 35616 21228
rect 1344 21142 5498 21194
rect 5550 21142 5602 21194
rect 5654 21142 5706 21194
rect 5758 21142 14066 21194
rect 14118 21142 14170 21194
rect 14222 21142 14274 21194
rect 14326 21142 22634 21194
rect 22686 21142 22738 21194
rect 22790 21142 22842 21194
rect 22894 21142 31202 21194
rect 31254 21142 31306 21194
rect 31358 21142 31410 21194
rect 31462 21142 35616 21194
rect 1344 21108 35616 21142
rect 34750 21026 34802 21038
rect 29698 20974 29710 21026
rect 29762 20974 29774 21026
rect 31826 20974 31838 21026
rect 31890 20974 31902 21026
rect 34750 20962 34802 20974
rect 14254 20914 14306 20926
rect 12786 20862 12798 20914
rect 12850 20862 12862 20914
rect 14254 20850 14306 20862
rect 16606 20914 16658 20926
rect 27246 20914 27298 20926
rect 22754 20862 22766 20914
rect 22818 20862 22830 20914
rect 23426 20862 23438 20914
rect 23490 20862 23502 20914
rect 25554 20862 25566 20914
rect 25618 20862 25630 20914
rect 16606 20850 16658 20862
rect 27246 20850 27298 20862
rect 28590 20914 28642 20926
rect 31714 20862 31726 20914
rect 31778 20862 31790 20914
rect 28590 20850 28642 20862
rect 6638 20802 6690 20814
rect 6638 20738 6690 20750
rect 8542 20802 8594 20814
rect 13806 20802 13858 20814
rect 9314 20750 9326 20802
rect 9378 20750 9390 20802
rect 9986 20750 9998 20802
rect 10050 20750 10062 20802
rect 8542 20738 8594 20750
rect 13806 20738 13858 20750
rect 14590 20802 14642 20814
rect 14590 20738 14642 20750
rect 16270 20802 16322 20814
rect 16270 20738 16322 20750
rect 16494 20802 16546 20814
rect 16494 20738 16546 20750
rect 16718 20802 16770 20814
rect 16718 20738 16770 20750
rect 16942 20802 16994 20814
rect 16942 20738 16994 20750
rect 18398 20802 18450 20814
rect 18398 20738 18450 20750
rect 18958 20802 19010 20814
rect 26910 20802 26962 20814
rect 26226 20750 26238 20802
rect 26290 20750 26302 20802
rect 18958 20738 19010 20750
rect 26910 20738 26962 20750
rect 27806 20802 27858 20814
rect 27806 20738 27858 20750
rect 28254 20802 28306 20814
rect 28254 20738 28306 20750
rect 28366 20802 28418 20814
rect 28366 20738 28418 20750
rect 29150 20802 29202 20814
rect 29150 20738 29202 20750
rect 29374 20802 29426 20814
rect 29374 20738 29426 20750
rect 30494 20802 30546 20814
rect 32722 20750 32734 20802
rect 32786 20750 32798 20802
rect 30494 20738 30546 20750
rect 6974 20690 7026 20702
rect 6974 20626 7026 20638
rect 7310 20690 7362 20702
rect 7310 20626 7362 20638
rect 7646 20690 7698 20702
rect 7646 20626 7698 20638
rect 7870 20690 7922 20702
rect 14926 20690 14978 20702
rect 9538 20638 9550 20690
rect 9602 20638 9614 20690
rect 10658 20638 10670 20690
rect 10722 20638 10734 20690
rect 7870 20626 7922 20638
rect 14926 20626 14978 20638
rect 15934 20690 15986 20702
rect 15934 20626 15986 20638
rect 17838 20690 17890 20702
rect 17838 20626 17890 20638
rect 18062 20690 18114 20702
rect 18062 20626 18114 20638
rect 18622 20690 18674 20702
rect 27022 20690 27074 20702
rect 21858 20638 21870 20690
rect 21922 20638 21934 20690
rect 18622 20626 18674 20638
rect 27022 20626 27074 20638
rect 27358 20690 27410 20702
rect 27358 20626 27410 20638
rect 30606 20690 30658 20702
rect 31938 20638 31950 20690
rect 32002 20638 32014 20690
rect 30606 20626 30658 20638
rect 6414 20578 6466 20590
rect 6414 20514 6466 20526
rect 6862 20578 6914 20590
rect 6862 20514 6914 20526
rect 7422 20578 7474 20590
rect 7422 20514 7474 20526
rect 8206 20578 8258 20590
rect 8206 20514 8258 20526
rect 13470 20578 13522 20590
rect 13470 20514 13522 20526
rect 16046 20578 16098 20590
rect 16046 20514 16098 20526
rect 18286 20578 18338 20590
rect 18286 20514 18338 20526
rect 18846 20578 18898 20590
rect 18846 20514 18898 20526
rect 21534 20578 21586 20590
rect 21534 20514 21586 20526
rect 27582 20578 27634 20590
rect 27582 20514 27634 20526
rect 1344 20410 35776 20444
rect 1344 20358 9782 20410
rect 9834 20358 9886 20410
rect 9938 20358 9990 20410
rect 10042 20358 18350 20410
rect 18402 20358 18454 20410
rect 18506 20358 18558 20410
rect 18610 20358 26918 20410
rect 26970 20358 27022 20410
rect 27074 20358 27126 20410
rect 27178 20358 35486 20410
rect 35538 20358 35590 20410
rect 35642 20358 35694 20410
rect 35746 20358 35776 20410
rect 1344 20324 35776 20358
rect 11566 20242 11618 20254
rect 11566 20178 11618 20190
rect 17950 20242 18002 20254
rect 23538 20190 23550 20242
rect 23602 20190 23614 20242
rect 17950 20178 18002 20190
rect 8206 20130 8258 20142
rect 8206 20066 8258 20078
rect 9662 20130 9714 20142
rect 9662 20066 9714 20078
rect 9774 20130 9826 20142
rect 9774 20066 9826 20078
rect 10334 20130 10386 20142
rect 10334 20066 10386 20078
rect 10894 20130 10946 20142
rect 10894 20066 10946 20078
rect 11006 20130 11058 20142
rect 11006 20066 11058 20078
rect 11454 20130 11506 20142
rect 11454 20066 11506 20078
rect 13134 20130 13186 20142
rect 13134 20066 13186 20078
rect 13358 20130 13410 20142
rect 13358 20066 13410 20078
rect 14926 20130 14978 20142
rect 14926 20066 14978 20078
rect 15262 20130 15314 20142
rect 15262 20066 15314 20078
rect 15934 20130 15986 20142
rect 15934 20066 15986 20078
rect 16606 20130 16658 20142
rect 16606 20066 16658 20078
rect 16718 20130 16770 20142
rect 18174 20130 18226 20142
rect 17378 20078 17390 20130
rect 17442 20078 17454 20130
rect 16718 20066 16770 20078
rect 18174 20066 18226 20078
rect 18286 20130 18338 20142
rect 26126 20130 26178 20142
rect 19730 20078 19742 20130
rect 19794 20078 19806 20130
rect 23986 20078 23998 20130
rect 24050 20078 24062 20130
rect 24434 20078 24446 20130
rect 24498 20078 24510 20130
rect 18286 20066 18338 20078
rect 26126 20066 26178 20078
rect 26238 20130 26290 20142
rect 26238 20066 26290 20078
rect 26462 20130 26514 20142
rect 26462 20066 26514 20078
rect 27134 20130 27186 20142
rect 27134 20066 27186 20078
rect 27358 20130 27410 20142
rect 31614 20130 31666 20142
rect 29250 20078 29262 20130
rect 29314 20078 29326 20130
rect 30258 20078 30270 20130
rect 30322 20078 30334 20130
rect 27358 20066 27410 20078
rect 31614 20066 31666 20078
rect 33070 20130 33122 20142
rect 33070 20066 33122 20078
rect 33182 20130 33234 20142
rect 33182 20066 33234 20078
rect 8542 20018 8594 20030
rect 5058 19966 5070 20018
rect 5122 19966 5134 20018
rect 8542 19954 8594 19966
rect 8766 20018 8818 20030
rect 8766 19954 8818 19966
rect 9438 20018 9490 20030
rect 9438 19954 9490 19966
rect 11230 20018 11282 20030
rect 11230 19954 11282 19966
rect 11678 20018 11730 20030
rect 11678 19954 11730 19966
rect 12014 20018 12066 20030
rect 12014 19954 12066 19966
rect 12462 20018 12514 20030
rect 12462 19954 12514 19966
rect 12574 20018 12626 20030
rect 12574 19954 12626 19966
rect 13022 20018 13074 20030
rect 13022 19954 13074 19966
rect 13470 20018 13522 20030
rect 13470 19954 13522 19966
rect 15710 20018 15762 20030
rect 15710 19954 15762 19966
rect 16046 20018 16098 20030
rect 16046 19954 16098 19966
rect 16942 20018 16994 20030
rect 16942 19954 16994 19966
rect 17726 20018 17778 20030
rect 21086 20018 21138 20030
rect 22094 20018 22146 20030
rect 25342 20018 25394 20030
rect 19954 19966 19966 20018
rect 20018 19966 20030 20018
rect 21634 19966 21646 20018
rect 21698 19966 21710 20018
rect 22866 19966 22878 20018
rect 22930 19966 22942 20018
rect 24546 19966 24558 20018
rect 24610 19966 24622 20018
rect 17726 19954 17778 19966
rect 21086 19954 21138 19966
rect 22094 19954 22146 19966
rect 25342 19954 25394 19966
rect 25566 20018 25618 20030
rect 25566 19954 25618 19966
rect 25790 20018 25842 20030
rect 25790 19954 25842 19966
rect 26798 20018 26850 20030
rect 31838 20018 31890 20030
rect 33742 20018 33794 20030
rect 34638 20018 34690 20030
rect 29474 19966 29486 20018
rect 29538 19966 29550 20018
rect 29698 19966 29710 20018
rect 29762 19966 29774 20018
rect 31938 19966 31950 20018
rect 32002 19966 32014 20018
rect 34066 19966 34078 20018
rect 34130 19966 34142 20018
rect 26798 19954 26850 19966
rect 31838 19954 31890 19966
rect 33742 19954 33794 19966
rect 34638 19954 34690 19966
rect 8654 19906 8706 19918
rect 5730 19854 5742 19906
rect 5794 19854 5806 19906
rect 7858 19854 7870 19906
rect 7922 19854 7934 19906
rect 8654 19842 8706 19854
rect 12798 19906 12850 19918
rect 25678 19906 25730 19918
rect 20626 19854 20638 19906
rect 20690 19854 20702 19906
rect 21746 19854 21758 19906
rect 21810 19854 21822 19906
rect 22978 19854 22990 19906
rect 23042 19854 23054 19906
rect 27458 19854 27470 19906
rect 27522 19854 27534 19906
rect 27906 19854 27918 19906
rect 27970 19854 27982 19906
rect 31714 19854 31726 19906
rect 31778 19854 31790 19906
rect 35074 19854 35086 19906
rect 35138 19854 35150 19906
rect 12798 19842 12850 19854
rect 25678 19842 25730 19854
rect 26686 19794 26738 19806
rect 26686 19730 26738 19742
rect 32286 19794 32338 19806
rect 32286 19730 32338 19742
rect 32510 19794 32562 19806
rect 33618 19742 33630 19794
rect 33682 19742 33694 19794
rect 32510 19730 32562 19742
rect 1344 19626 35616 19660
rect 1344 19574 5498 19626
rect 5550 19574 5602 19626
rect 5654 19574 5706 19626
rect 5758 19574 14066 19626
rect 14118 19574 14170 19626
rect 14222 19574 14274 19626
rect 14326 19574 22634 19626
rect 22686 19574 22738 19626
rect 22790 19574 22842 19626
rect 22894 19574 31202 19626
rect 31254 19574 31306 19626
rect 31358 19574 31410 19626
rect 31462 19574 35616 19626
rect 1344 19540 35616 19574
rect 25342 19458 25394 19470
rect 25342 19394 25394 19406
rect 25790 19458 25842 19470
rect 31490 19406 31502 19458
rect 31554 19406 31566 19458
rect 34290 19406 34302 19458
rect 34354 19406 34366 19458
rect 25790 19394 25842 19406
rect 27022 19346 27074 19358
rect 6402 19294 6414 19346
rect 6466 19294 6478 19346
rect 8530 19294 8542 19346
rect 8594 19294 8606 19346
rect 10210 19294 10222 19346
rect 10274 19294 10286 19346
rect 12338 19294 12350 19346
rect 12402 19294 12414 19346
rect 19394 19294 19406 19346
rect 19458 19294 19470 19346
rect 30034 19294 30046 19346
rect 30098 19294 30110 19346
rect 32274 19294 32286 19346
rect 32338 19294 32350 19346
rect 27022 19282 27074 19294
rect 8766 19234 8818 19246
rect 12686 19234 12738 19246
rect 5730 19182 5742 19234
rect 5794 19182 5806 19234
rect 9538 19182 9550 19234
rect 9602 19182 9614 19234
rect 8766 19170 8818 19182
rect 12686 19170 12738 19182
rect 14142 19234 14194 19246
rect 14142 19170 14194 19182
rect 14478 19234 14530 19246
rect 14478 19170 14530 19182
rect 14926 19234 14978 19246
rect 14926 19170 14978 19182
rect 15374 19234 15426 19246
rect 15374 19170 15426 19182
rect 15598 19234 15650 19246
rect 15598 19170 15650 19182
rect 15934 19234 15986 19246
rect 23214 19234 23266 19246
rect 16482 19182 16494 19234
rect 16546 19182 16558 19234
rect 20066 19182 20078 19234
rect 20130 19182 20142 19234
rect 20514 19182 20526 19234
rect 20578 19182 20590 19234
rect 15934 19170 15986 19182
rect 23214 19170 23266 19182
rect 25566 19234 25618 19246
rect 25566 19170 25618 19182
rect 26014 19234 26066 19246
rect 26014 19170 26066 19182
rect 27582 19234 27634 19246
rect 34526 19234 34578 19246
rect 28466 19182 28478 19234
rect 28530 19182 28542 19234
rect 30146 19182 30158 19234
rect 30210 19182 30222 19234
rect 30706 19182 30718 19234
rect 30770 19182 30782 19234
rect 32386 19182 32398 19234
rect 32450 19182 32462 19234
rect 27582 19170 27634 19182
rect 34526 19170 34578 19182
rect 34974 19234 35026 19246
rect 34974 19170 35026 19182
rect 8990 19122 9042 19134
rect 8990 19058 9042 19070
rect 9102 19122 9154 19134
rect 9102 19058 9154 19070
rect 12798 19122 12850 19134
rect 12798 19058 12850 19070
rect 13694 19122 13746 19134
rect 13694 19058 13746 19070
rect 13806 19122 13858 19134
rect 13806 19058 13858 19070
rect 14254 19122 14306 19134
rect 21422 19122 21474 19134
rect 26350 19122 26402 19134
rect 17266 19070 17278 19122
rect 17330 19070 17342 19122
rect 22418 19070 22430 19122
rect 22482 19070 22494 19122
rect 22754 19070 22766 19122
rect 22818 19070 22830 19122
rect 24770 19070 24782 19122
rect 24834 19070 24846 19122
rect 14254 19058 14306 19070
rect 21422 19058 21474 19070
rect 26350 19058 26402 19070
rect 26574 19122 26626 19134
rect 28578 19070 28590 19122
rect 28642 19070 28654 19122
rect 29922 19070 29934 19122
rect 29986 19070 29998 19122
rect 31378 19070 31390 19122
rect 31442 19070 31454 19122
rect 26574 19058 26626 19070
rect 13022 19010 13074 19022
rect 13022 18946 13074 18958
rect 13470 19010 13522 19022
rect 13470 18946 13522 18958
rect 15150 19010 15202 19022
rect 15150 18946 15202 18958
rect 16046 19010 16098 19022
rect 16046 18946 16098 18958
rect 16270 19010 16322 19022
rect 16270 18946 16322 18958
rect 20638 19010 20690 19022
rect 23662 19010 23714 19022
rect 22642 18958 22654 19010
rect 22706 18958 22718 19010
rect 20638 18946 20690 18958
rect 23662 18946 23714 18958
rect 24110 19010 24162 19022
rect 24110 18946 24162 18958
rect 26462 19010 26514 19022
rect 28018 18958 28030 19010
rect 28082 18958 28094 19010
rect 26462 18946 26514 18958
rect 1344 18842 35776 18876
rect 1344 18790 9782 18842
rect 9834 18790 9886 18842
rect 9938 18790 9990 18842
rect 10042 18790 18350 18842
rect 18402 18790 18454 18842
rect 18506 18790 18558 18842
rect 18610 18790 26918 18842
rect 26970 18790 27022 18842
rect 27074 18790 27126 18842
rect 27178 18790 35486 18842
rect 35538 18790 35590 18842
rect 35642 18790 35694 18842
rect 35746 18790 35776 18842
rect 1344 18756 35776 18790
rect 8094 18674 8146 18686
rect 12350 18674 12402 18686
rect 8642 18622 8654 18674
rect 8706 18622 8718 18674
rect 10098 18622 10110 18674
rect 10162 18622 10174 18674
rect 8094 18610 8146 18622
rect 12350 18610 12402 18622
rect 12798 18674 12850 18686
rect 12798 18610 12850 18622
rect 17502 18674 17554 18686
rect 17502 18610 17554 18622
rect 28030 18674 28082 18686
rect 28030 18610 28082 18622
rect 29598 18674 29650 18686
rect 29598 18610 29650 18622
rect 30270 18674 30322 18686
rect 34290 18622 34302 18674
rect 34354 18622 34366 18674
rect 30270 18610 30322 18622
rect 7422 18562 7474 18574
rect 7422 18498 7474 18510
rect 7534 18562 7586 18574
rect 7534 18498 7586 18510
rect 8206 18562 8258 18574
rect 8206 18498 8258 18510
rect 12462 18562 12514 18574
rect 27806 18562 27858 18574
rect 34862 18562 34914 18574
rect 25442 18510 25454 18562
rect 25506 18510 25518 18562
rect 26002 18510 26014 18562
rect 26066 18510 26078 18562
rect 30594 18510 30606 18562
rect 30658 18510 30670 18562
rect 31378 18510 31390 18562
rect 31442 18510 31454 18562
rect 33170 18510 33182 18562
rect 33234 18510 33246 18562
rect 12462 18498 12514 18510
rect 27806 18498 27858 18510
rect 34862 18498 34914 18510
rect 7758 18450 7810 18462
rect 7758 18386 7810 18398
rect 7870 18450 7922 18462
rect 7870 18386 7922 18398
rect 8990 18450 9042 18462
rect 10558 18450 10610 18462
rect 9874 18398 9886 18450
rect 9938 18398 9950 18450
rect 8990 18386 9042 18398
rect 10558 18386 10610 18398
rect 13134 18450 13186 18462
rect 13134 18386 13186 18398
rect 13582 18450 13634 18462
rect 17278 18450 17330 18462
rect 13906 18398 13918 18450
rect 13970 18398 13982 18450
rect 14690 18398 14702 18450
rect 14754 18398 14766 18450
rect 13582 18386 13634 18398
rect 17278 18386 17330 18398
rect 17614 18450 17666 18462
rect 17614 18386 17666 18398
rect 17838 18450 17890 18462
rect 26798 18450 26850 18462
rect 23426 18398 23438 18450
rect 23490 18398 23502 18450
rect 26338 18398 26350 18450
rect 26402 18398 26414 18450
rect 17838 18386 17890 18398
rect 26798 18386 26850 18398
rect 26910 18450 26962 18462
rect 26910 18386 26962 18398
rect 27022 18450 27074 18462
rect 27022 18386 27074 18398
rect 28366 18450 28418 18462
rect 28366 18386 28418 18398
rect 28702 18450 28754 18462
rect 33406 18450 33458 18462
rect 29138 18398 29150 18450
rect 29202 18398 29214 18450
rect 29810 18398 29822 18450
rect 29874 18398 29886 18450
rect 31826 18398 31838 18450
rect 31890 18398 31902 18450
rect 32162 18398 32174 18450
rect 32226 18398 32238 18450
rect 28702 18386 28754 18398
rect 33406 18386 33458 18398
rect 33854 18450 33906 18462
rect 33854 18386 33906 18398
rect 34078 18450 34130 18462
rect 34078 18386 34130 18398
rect 18846 18338 18898 18350
rect 25118 18338 25170 18350
rect 33070 18338 33122 18350
rect 16818 18286 16830 18338
rect 16882 18286 16894 18338
rect 21634 18286 21646 18338
rect 21698 18286 21710 18338
rect 27458 18286 27470 18338
rect 27522 18286 27534 18338
rect 31714 18286 31726 18338
rect 31778 18286 31790 18338
rect 18846 18274 18898 18286
rect 25118 18274 25170 18286
rect 33070 18274 33122 18286
rect 12350 18226 12402 18238
rect 12350 18162 12402 18174
rect 28142 18226 28194 18238
rect 28142 18162 28194 18174
rect 34638 18226 34690 18238
rect 34638 18162 34690 18174
rect 1344 18058 35616 18092
rect 1344 18006 5498 18058
rect 5550 18006 5602 18058
rect 5654 18006 5706 18058
rect 5758 18006 14066 18058
rect 14118 18006 14170 18058
rect 14222 18006 14274 18058
rect 14326 18006 22634 18058
rect 22686 18006 22738 18058
rect 22790 18006 22842 18058
rect 22894 18006 31202 18058
rect 31254 18006 31306 18058
rect 31358 18006 31410 18058
rect 31462 18006 35616 18058
rect 1344 17972 35616 18006
rect 20638 17890 20690 17902
rect 28478 17890 28530 17902
rect 23538 17838 23550 17890
rect 23602 17838 23614 17890
rect 24770 17838 24782 17890
rect 24834 17887 24846 17890
rect 25106 17887 25118 17890
rect 24834 17841 25118 17887
rect 24834 17838 24846 17841
rect 25106 17838 25118 17841
rect 25170 17838 25182 17890
rect 20638 17826 20690 17838
rect 28478 17826 28530 17838
rect 30942 17890 30994 17902
rect 30942 17826 30994 17838
rect 10782 17778 10834 17790
rect 10210 17726 10222 17778
rect 10274 17726 10286 17778
rect 10782 17714 10834 17726
rect 16158 17778 16210 17790
rect 16158 17714 16210 17726
rect 17054 17778 17106 17790
rect 17054 17714 17106 17726
rect 21422 17778 21474 17790
rect 29262 17778 29314 17790
rect 24546 17726 24558 17778
rect 24610 17726 24622 17778
rect 21422 17714 21474 17726
rect 29262 17714 29314 17726
rect 30830 17778 30882 17790
rect 30830 17714 30882 17726
rect 31278 17778 31330 17790
rect 32274 17726 32286 17778
rect 32338 17726 32350 17778
rect 31278 17714 31330 17726
rect 12350 17666 12402 17678
rect 7298 17614 7310 17666
rect 7362 17614 7374 17666
rect 12350 17602 12402 17614
rect 12686 17666 12738 17678
rect 12686 17602 12738 17614
rect 12910 17666 12962 17678
rect 12910 17602 12962 17614
rect 13470 17666 13522 17678
rect 13470 17602 13522 17614
rect 14030 17666 14082 17678
rect 14030 17602 14082 17614
rect 14590 17666 14642 17678
rect 14590 17602 14642 17614
rect 18062 17666 18114 17678
rect 18062 17602 18114 17614
rect 18286 17666 18338 17678
rect 22318 17666 22370 17678
rect 19618 17614 19630 17666
rect 19682 17614 19694 17666
rect 20290 17614 20302 17666
rect 20354 17614 20366 17666
rect 18286 17602 18338 17614
rect 22318 17602 22370 17614
rect 22990 17666 23042 17678
rect 26798 17666 26850 17678
rect 23986 17614 23998 17666
rect 24050 17614 24062 17666
rect 24322 17614 24334 17666
rect 24386 17614 24398 17666
rect 25442 17614 25454 17666
rect 25506 17614 25518 17666
rect 26562 17614 26574 17666
rect 26626 17614 26638 17666
rect 22990 17602 23042 17614
rect 26798 17602 26850 17614
rect 27022 17666 27074 17678
rect 27022 17602 27074 17614
rect 28590 17666 28642 17678
rect 31714 17614 31726 17666
rect 31778 17614 31790 17666
rect 35074 17614 35086 17666
rect 35138 17614 35150 17666
rect 28590 17602 28642 17614
rect 13806 17554 13858 17566
rect 8082 17502 8094 17554
rect 8146 17502 8158 17554
rect 13806 17490 13858 17502
rect 14254 17554 14306 17566
rect 14254 17490 14306 17502
rect 14478 17554 14530 17566
rect 14478 17490 14530 17502
rect 17838 17554 17890 17566
rect 22430 17554 22482 17566
rect 18610 17502 18622 17554
rect 18674 17502 18686 17554
rect 19394 17502 19406 17554
rect 19458 17502 19470 17554
rect 20738 17502 20750 17554
rect 20802 17502 20814 17554
rect 17838 17490 17890 17502
rect 22430 17490 22482 17502
rect 22654 17554 22706 17566
rect 30158 17554 30210 17566
rect 26226 17502 26238 17554
rect 26290 17502 26302 17554
rect 27458 17502 27470 17554
rect 27522 17502 27534 17554
rect 27906 17502 27918 17554
rect 27970 17502 27982 17554
rect 34402 17502 34414 17554
rect 34466 17502 34478 17554
rect 22654 17490 22706 17502
rect 30158 17490 30210 17502
rect 12462 17442 12514 17454
rect 12462 17378 12514 17390
rect 13582 17442 13634 17454
rect 25118 17442 25170 17454
rect 28478 17442 28530 17454
rect 19506 17390 19518 17442
rect 19570 17390 19582 17442
rect 21858 17390 21870 17442
rect 21922 17390 21934 17442
rect 25554 17390 25566 17442
rect 25618 17390 25630 17442
rect 13582 17378 13634 17390
rect 25118 17378 25170 17390
rect 28478 17378 28530 17390
rect 29822 17442 29874 17454
rect 29822 17378 29874 17390
rect 30270 17442 30322 17454
rect 30270 17378 30322 17390
rect 30382 17442 30434 17454
rect 30382 17378 30434 17390
rect 1344 17274 35776 17308
rect 1344 17222 9782 17274
rect 9834 17222 9886 17274
rect 9938 17222 9990 17274
rect 10042 17222 18350 17274
rect 18402 17222 18454 17274
rect 18506 17222 18558 17274
rect 18610 17222 26918 17274
rect 26970 17222 27022 17274
rect 27074 17222 27126 17274
rect 27178 17222 35486 17274
rect 35538 17222 35590 17274
rect 35642 17222 35694 17274
rect 35746 17222 35776 17274
rect 1344 17188 35776 17222
rect 8542 17106 8594 17118
rect 8542 17042 8594 17054
rect 9886 17106 9938 17118
rect 9886 17042 9938 17054
rect 9998 17106 10050 17118
rect 9998 17042 10050 17054
rect 10782 17106 10834 17118
rect 10782 17042 10834 17054
rect 15262 17106 15314 17118
rect 15262 17042 15314 17054
rect 16830 17106 16882 17118
rect 16830 17042 16882 17054
rect 18846 17106 18898 17118
rect 20862 17106 20914 17118
rect 19394 17054 19406 17106
rect 19458 17054 19470 17106
rect 18846 17042 18898 17054
rect 20862 17042 20914 17054
rect 23102 17106 23154 17118
rect 27582 17106 27634 17118
rect 25666 17054 25678 17106
rect 25730 17054 25742 17106
rect 23102 17042 23154 17054
rect 27582 17042 27634 17054
rect 27918 17106 27970 17118
rect 27918 17042 27970 17054
rect 28590 17106 28642 17118
rect 28590 17042 28642 17054
rect 30718 17106 30770 17118
rect 34638 17106 34690 17118
rect 33954 17054 33966 17106
rect 34018 17054 34030 17106
rect 30718 17042 30770 17054
rect 34638 17042 34690 17054
rect 8990 16994 9042 17006
rect 17838 16994 17890 17006
rect 12674 16942 12686 16994
rect 12738 16942 12750 16994
rect 17602 16942 17614 16994
rect 17666 16942 17678 16994
rect 8990 16930 9042 16942
rect 17838 16930 17890 16942
rect 17950 16994 18002 17006
rect 21982 16994 22034 17006
rect 26686 16994 26738 17006
rect 19730 16942 19742 16994
rect 19794 16942 19806 16994
rect 24210 16942 24222 16994
rect 24274 16942 24286 16994
rect 25442 16942 25454 16994
rect 25506 16942 25518 16994
rect 26002 16942 26014 16994
rect 26066 16942 26078 16994
rect 17950 16930 18002 16942
rect 21982 16930 22034 16942
rect 26686 16930 26738 16942
rect 28366 16994 28418 17006
rect 29486 16994 29538 17006
rect 28914 16942 28926 16994
rect 28978 16942 28990 16994
rect 28366 16930 28418 16942
rect 29486 16930 29538 16942
rect 32174 16994 32226 17006
rect 32174 16930 32226 16942
rect 8430 16882 8482 16894
rect 8430 16818 8482 16830
rect 8766 16882 8818 16894
rect 8766 16818 8818 16830
rect 9774 16882 9826 16894
rect 18174 16882 18226 16894
rect 21758 16882 21810 16894
rect 10322 16830 10334 16882
rect 10386 16830 10398 16882
rect 12002 16830 12014 16882
rect 12066 16830 12078 16882
rect 19842 16830 19854 16882
rect 19906 16830 19918 16882
rect 21410 16830 21422 16882
rect 21474 16830 21486 16882
rect 9774 16818 9826 16830
rect 18174 16818 18226 16830
rect 21758 16818 21810 16830
rect 22206 16882 22258 16894
rect 25230 16882 25282 16894
rect 22530 16830 22542 16882
rect 22594 16830 22606 16882
rect 23426 16830 23438 16882
rect 23490 16830 23502 16882
rect 22206 16818 22258 16830
rect 25230 16818 25282 16830
rect 26910 16882 26962 16894
rect 30046 16882 30098 16894
rect 33070 16882 33122 16894
rect 35198 16882 35250 16894
rect 28802 16830 28814 16882
rect 28866 16830 28878 16882
rect 31714 16830 31726 16882
rect 31778 16830 31790 16882
rect 32386 16830 32398 16882
rect 32450 16830 32462 16882
rect 33506 16830 33518 16882
rect 33570 16830 33582 16882
rect 34178 16830 34190 16882
rect 34242 16830 34254 16882
rect 26910 16818 26962 16830
rect 30046 16818 30098 16830
rect 33070 16818 33122 16830
rect 35198 16818 35250 16830
rect 28030 16770 28082 16782
rect 30830 16770 30882 16782
rect 14802 16718 14814 16770
rect 14866 16718 14878 16770
rect 17938 16718 17950 16770
rect 18002 16718 18014 16770
rect 29138 16718 29150 16770
rect 29202 16718 29214 16770
rect 28030 16706 28082 16718
rect 30830 16706 30882 16718
rect 30942 16770 30994 16782
rect 30942 16706 30994 16718
rect 31278 16770 31330 16782
rect 31278 16706 31330 16718
rect 27246 16658 27298 16670
rect 27246 16594 27298 16606
rect 27470 16658 27522 16670
rect 27470 16594 27522 16606
rect 1344 16490 35616 16524
rect 1344 16438 5498 16490
rect 5550 16438 5602 16490
rect 5654 16438 5706 16490
rect 5758 16438 14066 16490
rect 14118 16438 14170 16490
rect 14222 16438 14274 16490
rect 14326 16438 22634 16490
rect 22686 16438 22738 16490
rect 22790 16438 22842 16490
rect 22894 16438 31202 16490
rect 31254 16438 31306 16490
rect 31358 16438 31410 16490
rect 31462 16438 35616 16490
rect 1344 16404 35616 16438
rect 33070 16322 33122 16334
rect 21410 16270 21422 16322
rect 21474 16270 21486 16322
rect 25106 16270 25118 16322
rect 25170 16270 25182 16322
rect 33070 16258 33122 16270
rect 35086 16322 35138 16334
rect 35086 16258 35138 16270
rect 9214 16210 9266 16222
rect 15374 16210 15426 16222
rect 19854 16210 19906 16222
rect 22878 16210 22930 16222
rect 10770 16158 10782 16210
rect 10834 16158 10846 16210
rect 12898 16158 12910 16210
rect 12962 16158 12974 16210
rect 16818 16158 16830 16210
rect 16882 16158 16894 16210
rect 20290 16158 20302 16210
rect 20354 16158 20366 16210
rect 28018 16158 28030 16210
rect 28082 16158 28094 16210
rect 29250 16158 29262 16210
rect 29314 16158 29326 16210
rect 9214 16146 9266 16158
rect 15374 16146 15426 16158
rect 19854 16146 19906 16158
rect 22878 16146 22930 16158
rect 18734 16098 18786 16110
rect 10098 16046 10110 16098
rect 10162 16046 10174 16098
rect 16482 16046 16494 16098
rect 16546 16046 16558 16098
rect 17826 16046 17838 16098
rect 17890 16046 17902 16098
rect 18734 16034 18786 16046
rect 20750 16098 20802 16110
rect 20750 16034 20802 16046
rect 21758 16098 21810 16110
rect 24222 16098 24274 16110
rect 23874 16046 23886 16098
rect 23938 16046 23950 16098
rect 21758 16034 21810 16046
rect 24222 16034 24274 16046
rect 24446 16098 24498 16110
rect 24446 16034 24498 16046
rect 25454 16098 25506 16110
rect 27918 16098 27970 16110
rect 28590 16098 28642 16110
rect 32734 16098 32786 16110
rect 26450 16046 26462 16098
rect 26514 16046 26526 16098
rect 27458 16046 27470 16098
rect 27522 16046 27534 16098
rect 28130 16046 28142 16098
rect 28194 16046 28206 16098
rect 32162 16046 32174 16098
rect 32226 16046 32238 16098
rect 25454 16034 25506 16046
rect 27918 16034 27970 16046
rect 28590 16034 28642 16046
rect 32734 16034 32786 16046
rect 34638 16098 34690 16110
rect 34638 16034 34690 16046
rect 35198 16098 35250 16110
rect 35198 16034 35250 16046
rect 15262 15986 15314 15998
rect 21982 15986 22034 15998
rect 13570 15934 13582 15986
rect 13634 15934 13646 15986
rect 16370 15934 16382 15986
rect 16434 15934 16446 15986
rect 15262 15922 15314 15934
rect 21982 15922 22034 15934
rect 23438 15986 23490 15998
rect 23438 15922 23490 15934
rect 24670 15986 24722 15998
rect 24670 15922 24722 15934
rect 25678 15986 25730 15998
rect 25678 15922 25730 15934
rect 26798 15986 26850 15998
rect 26798 15922 26850 15934
rect 26910 15986 26962 15998
rect 35086 15986 35138 15998
rect 31490 15934 31502 15986
rect 31554 15934 31566 15986
rect 33282 15934 33294 15986
rect 33346 15934 33358 15986
rect 33618 15934 33630 15986
rect 33682 15934 33694 15986
rect 34290 15934 34302 15986
rect 34354 15934 34366 15986
rect 26910 15922 26962 15934
rect 35086 15922 35138 15934
rect 13918 15874 13970 15886
rect 13918 15810 13970 15822
rect 14926 15874 14978 15886
rect 23102 15874 23154 15886
rect 19058 15822 19070 15874
rect 19122 15822 19134 15874
rect 14926 15810 14978 15822
rect 23102 15810 23154 15822
rect 27022 15874 27074 15886
rect 27022 15810 27074 15822
rect 27134 15874 27186 15886
rect 27134 15810 27186 15822
rect 27694 15874 27746 15886
rect 27694 15810 27746 15822
rect 28478 15874 28530 15886
rect 28478 15810 28530 15822
rect 1344 15706 35776 15740
rect 1344 15654 9782 15706
rect 9834 15654 9886 15706
rect 9938 15654 9990 15706
rect 10042 15654 18350 15706
rect 18402 15654 18454 15706
rect 18506 15654 18558 15706
rect 18610 15654 26918 15706
rect 26970 15654 27022 15706
rect 27074 15654 27126 15706
rect 27178 15654 35486 15706
rect 35538 15654 35590 15706
rect 35642 15654 35694 15706
rect 35746 15654 35776 15706
rect 1344 15620 35776 15654
rect 13246 15538 13298 15550
rect 13806 15538 13858 15550
rect 13458 15486 13470 15538
rect 13522 15486 13534 15538
rect 13246 15474 13298 15486
rect 13806 15474 13858 15486
rect 15598 15538 15650 15550
rect 15598 15474 15650 15486
rect 21198 15538 21250 15550
rect 35086 15538 35138 15550
rect 34738 15486 34750 15538
rect 34802 15486 34814 15538
rect 21198 15474 21250 15486
rect 35086 15474 35138 15486
rect 14814 15426 14866 15438
rect 14130 15374 14142 15426
rect 14194 15374 14206 15426
rect 14814 15362 14866 15374
rect 25790 15426 25842 15438
rect 25790 15362 25842 15374
rect 25902 15426 25954 15438
rect 25902 15362 25954 15374
rect 33182 15426 33234 15438
rect 33730 15374 33742 15426
rect 33794 15374 33806 15426
rect 34290 15374 34302 15426
rect 34354 15374 34366 15426
rect 33182 15362 33234 15374
rect 21758 15314 21810 15326
rect 25678 15314 25730 15326
rect 14354 15262 14366 15314
rect 14418 15262 14430 15314
rect 15138 15262 15150 15314
rect 15202 15262 15214 15314
rect 17490 15262 17502 15314
rect 17554 15262 17566 15314
rect 17938 15262 17950 15314
rect 18002 15262 18014 15314
rect 21970 15262 21982 15314
rect 22034 15262 22046 15314
rect 24210 15262 24222 15314
rect 24274 15262 24286 15314
rect 21758 15250 21810 15262
rect 25678 15250 25730 15262
rect 26910 15314 26962 15326
rect 26910 15250 26962 15262
rect 27134 15314 27186 15326
rect 27134 15250 27186 15262
rect 27582 15314 27634 15326
rect 27582 15250 27634 15262
rect 27806 15314 27858 15326
rect 27806 15250 27858 15262
rect 28702 15314 28754 15326
rect 30482 15262 30494 15314
rect 30546 15262 30558 15314
rect 31826 15262 31838 15314
rect 31890 15262 31902 15314
rect 28702 15250 28754 15262
rect 14926 15202 14978 15214
rect 26350 15202 26402 15214
rect 20402 15150 20414 15202
rect 20466 15150 20478 15202
rect 22306 15150 22318 15202
rect 22370 15150 22382 15202
rect 24546 15150 24558 15202
rect 24610 15150 24622 15202
rect 14926 15138 14978 15150
rect 26350 15138 26402 15150
rect 27358 15202 27410 15214
rect 31502 15202 31554 15214
rect 29810 15150 29822 15202
rect 29874 15150 29886 15202
rect 27358 15138 27410 15150
rect 31502 15138 31554 15150
rect 32510 15202 32562 15214
rect 32510 15138 32562 15150
rect 28478 15090 28530 15102
rect 25218 15038 25230 15090
rect 25282 15038 25294 15090
rect 28130 15038 28142 15090
rect 28194 15038 28206 15090
rect 28478 15026 28530 15038
rect 32398 15090 32450 15102
rect 32398 15026 32450 15038
rect 33518 15090 33570 15102
rect 33518 15026 33570 15038
rect 1344 14922 35616 14956
rect 1344 14870 5498 14922
rect 5550 14870 5602 14922
rect 5654 14870 5706 14922
rect 5758 14870 14066 14922
rect 14118 14870 14170 14922
rect 14222 14870 14274 14922
rect 14326 14870 22634 14922
rect 22686 14870 22738 14922
rect 22790 14870 22842 14922
rect 22894 14870 31202 14922
rect 31254 14870 31306 14922
rect 31358 14870 31410 14922
rect 31462 14870 35616 14922
rect 1344 14836 35616 14870
rect 20750 14754 20802 14766
rect 20750 14690 20802 14702
rect 28478 14754 28530 14766
rect 28478 14690 28530 14702
rect 31726 14754 31778 14766
rect 31726 14690 31778 14702
rect 8318 14642 8370 14654
rect 8318 14578 8370 14590
rect 9214 14642 9266 14654
rect 9214 14578 9266 14590
rect 11790 14642 11842 14654
rect 20638 14642 20690 14654
rect 14466 14590 14478 14642
rect 14530 14590 14542 14642
rect 16594 14590 16606 14642
rect 16658 14590 16670 14642
rect 16930 14590 16942 14642
rect 16994 14590 17006 14642
rect 19058 14590 19070 14642
rect 19122 14590 19134 14642
rect 25330 14590 25342 14642
rect 25394 14590 25406 14642
rect 32274 14590 32286 14642
rect 32338 14590 32350 14642
rect 11790 14578 11842 14590
rect 20638 14578 20690 14590
rect 10222 14530 10274 14542
rect 10222 14466 10274 14478
rect 10446 14530 10498 14542
rect 10446 14466 10498 14478
rect 10670 14530 10722 14542
rect 10670 14466 10722 14478
rect 11006 14530 11058 14542
rect 13794 14478 13806 14530
rect 13858 14478 13870 14530
rect 19842 14478 19854 14530
rect 19906 14478 19918 14530
rect 20402 14478 20414 14530
rect 20466 14478 20478 14530
rect 23202 14478 23214 14530
rect 23266 14478 23278 14530
rect 27458 14478 27470 14530
rect 27522 14478 27534 14530
rect 30930 14478 30942 14530
rect 30994 14478 31006 14530
rect 35074 14478 35086 14530
rect 35138 14478 35150 14530
rect 11006 14466 11058 14478
rect 11230 14418 11282 14430
rect 11230 14354 11282 14366
rect 11342 14418 11394 14430
rect 11342 14354 11394 14366
rect 27918 14418 27970 14430
rect 27918 14354 27970 14366
rect 28590 14418 28642 14430
rect 29138 14366 29150 14418
rect 29202 14366 29214 14418
rect 29922 14366 29934 14418
rect 29986 14366 29998 14418
rect 34402 14366 34414 14418
rect 34466 14366 34478 14418
rect 28590 14354 28642 14366
rect 10334 14306 10386 14318
rect 10334 14242 10386 14254
rect 21422 14306 21474 14318
rect 21422 14242 21474 14254
rect 28478 14306 28530 14318
rect 28478 14242 28530 14254
rect 1344 14138 35776 14172
rect 1344 14086 9782 14138
rect 9834 14086 9886 14138
rect 9938 14086 9990 14138
rect 10042 14086 18350 14138
rect 18402 14086 18454 14138
rect 18506 14086 18558 14138
rect 18610 14086 26918 14138
rect 26970 14086 27022 14138
rect 27074 14086 27126 14138
rect 27178 14086 35486 14138
rect 35538 14086 35590 14138
rect 35642 14086 35694 14138
rect 35746 14086 35776 14138
rect 1344 14052 35776 14086
rect 7086 13970 7138 13982
rect 7086 13906 7138 13918
rect 8094 13970 8146 13982
rect 8094 13906 8146 13918
rect 8990 13970 9042 13982
rect 8990 13906 9042 13918
rect 14926 13970 14978 13982
rect 14926 13906 14978 13918
rect 17390 13970 17442 13982
rect 17390 13906 17442 13918
rect 19518 13970 19570 13982
rect 19518 13906 19570 13918
rect 19742 13970 19794 13982
rect 20750 13970 20802 13982
rect 33182 13970 33234 13982
rect 20402 13918 20414 13970
rect 20466 13918 20478 13970
rect 25218 13918 25230 13970
rect 25282 13918 25294 13970
rect 19742 13906 19794 13918
rect 20750 13906 20802 13918
rect 33182 13906 33234 13918
rect 35086 13970 35138 13982
rect 35086 13906 35138 13918
rect 17950 13858 18002 13870
rect 10322 13806 10334 13858
rect 10386 13806 10398 13858
rect 15586 13806 15598 13858
rect 15650 13806 15662 13858
rect 17950 13794 18002 13806
rect 19406 13858 19458 13870
rect 19406 13794 19458 13806
rect 19966 13858 20018 13870
rect 19966 13794 20018 13806
rect 20078 13858 20130 13870
rect 25790 13858 25842 13870
rect 34750 13858 34802 13870
rect 22306 13806 22318 13858
rect 22370 13806 22382 13858
rect 23090 13806 23102 13858
rect 23154 13806 23166 13858
rect 27346 13806 27358 13858
rect 27410 13806 27422 13858
rect 28130 13806 28142 13858
rect 28194 13806 28206 13858
rect 33730 13806 33742 13858
rect 33794 13806 33806 13858
rect 34178 13806 34190 13858
rect 34242 13806 34254 13858
rect 20078 13794 20130 13806
rect 25790 13794 25842 13806
rect 34750 13794 34802 13806
rect 6862 13746 6914 13758
rect 6862 13682 6914 13694
rect 7198 13746 7250 13758
rect 7198 13682 7250 13694
rect 7422 13746 7474 13758
rect 13358 13746 13410 13758
rect 9538 13694 9550 13746
rect 9602 13694 9614 13746
rect 7422 13682 7474 13694
rect 13358 13682 13410 13694
rect 14366 13746 14418 13758
rect 24558 13746 24610 13758
rect 14690 13694 14702 13746
rect 14754 13694 14766 13746
rect 15362 13694 15374 13746
rect 15426 13694 15438 13746
rect 22754 13694 22766 13746
rect 22818 13694 22830 13746
rect 14366 13682 14418 13694
rect 24558 13682 24610 13694
rect 25566 13746 25618 13758
rect 28814 13746 28866 13758
rect 27122 13694 27134 13746
rect 27186 13694 27198 13746
rect 28018 13694 28030 13746
rect 28082 13694 28094 13746
rect 29698 13694 29710 13746
rect 29762 13694 29774 13746
rect 25566 13682 25618 13694
rect 28814 13682 28866 13694
rect 8430 13634 8482 13646
rect 12798 13634 12850 13646
rect 12450 13582 12462 13634
rect 12514 13582 12526 13634
rect 8430 13570 8482 13582
rect 12798 13570 12850 13582
rect 13806 13634 13858 13646
rect 13806 13570 13858 13582
rect 16158 13634 16210 13646
rect 16158 13570 16210 13582
rect 18622 13634 18674 13646
rect 21858 13582 21870 13634
rect 21922 13582 21934 13634
rect 30370 13582 30382 13634
rect 30434 13582 30446 13634
rect 32498 13582 32510 13634
rect 32562 13582 32574 13634
rect 18622 13570 18674 13582
rect 26350 13522 26402 13534
rect 26350 13458 26402 13470
rect 26686 13522 26738 13534
rect 26686 13458 26738 13470
rect 29150 13522 29202 13534
rect 29150 13458 29202 13470
rect 33518 13522 33570 13534
rect 33518 13458 33570 13470
rect 1344 13354 35616 13388
rect 1344 13302 5498 13354
rect 5550 13302 5602 13354
rect 5654 13302 5706 13354
rect 5758 13302 14066 13354
rect 14118 13302 14170 13354
rect 14222 13302 14274 13354
rect 14326 13302 22634 13354
rect 22686 13302 22738 13354
rect 22790 13302 22842 13354
rect 22894 13302 31202 13354
rect 31254 13302 31306 13354
rect 31358 13302 31410 13354
rect 31462 13302 35616 13354
rect 1344 13268 35616 13302
rect 6190 13186 6242 13198
rect 6190 13122 6242 13134
rect 27918 13186 27970 13198
rect 27918 13122 27970 13134
rect 28254 13186 28306 13198
rect 28254 13122 28306 13134
rect 31726 13186 31778 13198
rect 31726 13122 31778 13134
rect 8542 13074 8594 13086
rect 8542 13010 8594 13022
rect 10670 13074 10722 13086
rect 10670 13010 10722 13022
rect 12798 13074 12850 13086
rect 28478 13074 28530 13086
rect 22418 13022 22430 13074
rect 22482 13022 22494 13074
rect 24322 13022 24334 13074
rect 24386 13022 24398 13074
rect 24658 13022 24670 13074
rect 24722 13022 24734 13074
rect 26786 13022 26798 13074
rect 26850 13022 26862 13074
rect 12798 13010 12850 13022
rect 28478 13010 28530 13022
rect 30494 13074 30546 13086
rect 32274 13022 32286 13074
rect 32338 13022 32350 13074
rect 30494 13010 30546 13022
rect 6526 12962 6578 12974
rect 6526 12898 6578 12910
rect 7198 12962 7250 12974
rect 7198 12898 7250 12910
rect 7646 12962 7698 12974
rect 9998 12962 10050 12974
rect 8082 12910 8094 12962
rect 8146 12910 8158 12962
rect 7646 12898 7698 12910
rect 9998 12898 10050 12910
rect 10334 12962 10386 12974
rect 12126 12962 12178 12974
rect 11554 12910 11566 12962
rect 11618 12910 11630 12962
rect 10334 12898 10386 12910
rect 12126 12898 12178 12910
rect 12462 12962 12514 12974
rect 22990 12962 23042 12974
rect 20514 12910 20526 12962
rect 20578 12910 20590 12962
rect 21858 12910 21870 12962
rect 21922 12910 21934 12962
rect 22530 12910 22542 12962
rect 22594 12910 22606 12962
rect 12462 12898 12514 12910
rect 22990 12898 23042 12910
rect 23326 12962 23378 12974
rect 29150 12962 29202 12974
rect 24210 12910 24222 12962
rect 24274 12910 24286 12962
rect 27570 12910 27582 12962
rect 27634 12910 27646 12962
rect 23326 12898 23378 12910
rect 29150 12898 29202 12910
rect 29374 12962 29426 12974
rect 29374 12898 29426 12910
rect 29710 12962 29762 12974
rect 29710 12898 29762 12910
rect 30046 12962 30098 12974
rect 30046 12898 30098 12910
rect 30270 12962 30322 12974
rect 30270 12898 30322 12910
rect 30606 12962 30658 12974
rect 31154 12910 31166 12962
rect 31218 12910 31230 12962
rect 35074 12910 35086 12962
rect 35138 12910 35150 12962
rect 30606 12898 30658 12910
rect 6302 12850 6354 12862
rect 6302 12786 6354 12798
rect 6974 12850 7026 12862
rect 6974 12786 7026 12798
rect 8878 12850 8930 12862
rect 8878 12786 8930 12798
rect 9662 12850 9714 12862
rect 9662 12786 9714 12798
rect 10782 12850 10834 12862
rect 12238 12850 12290 12862
rect 11778 12798 11790 12850
rect 11842 12798 11854 12850
rect 10782 12786 10834 12798
rect 12238 12786 12290 12798
rect 19406 12850 19458 12862
rect 19406 12786 19458 12798
rect 19742 12850 19794 12862
rect 19742 12786 19794 12798
rect 19966 12850 20018 12862
rect 23214 12850 23266 12862
rect 31838 12850 31890 12862
rect 22754 12798 22766 12850
rect 22818 12798 22830 12850
rect 23986 12798 23998 12850
rect 24050 12798 24062 12850
rect 34402 12798 34414 12850
rect 34466 12798 34478 12850
rect 19966 12786 20018 12798
rect 23214 12786 23266 12798
rect 31838 12786 31890 12798
rect 6190 12738 6242 12750
rect 6190 12674 6242 12686
rect 6862 12738 6914 12750
rect 6862 12674 6914 12686
rect 7534 12738 7586 12750
rect 7534 12674 7586 12686
rect 7758 12738 7810 12750
rect 7758 12674 7810 12686
rect 8430 12738 8482 12750
rect 8430 12674 8482 12686
rect 8654 12738 8706 12750
rect 8654 12674 8706 12686
rect 10110 12738 10162 12750
rect 10110 12674 10162 12686
rect 10558 12738 10610 12750
rect 10558 12674 10610 12686
rect 11006 12738 11058 12750
rect 11006 12674 11058 12686
rect 15150 12738 15202 12750
rect 16494 12738 16546 12750
rect 15474 12686 15486 12738
rect 15538 12686 15550 12738
rect 16146 12686 16158 12738
rect 16210 12686 16222 12738
rect 15150 12674 15202 12686
rect 16494 12674 16546 12686
rect 19518 12738 19570 12750
rect 29486 12738 29538 12750
rect 20290 12686 20302 12738
rect 20354 12686 20366 12738
rect 19518 12674 19570 12686
rect 29486 12674 29538 12686
rect 30942 12738 30994 12750
rect 30942 12674 30994 12686
rect 31726 12738 31778 12750
rect 31726 12674 31778 12686
rect 1344 12570 35776 12604
rect 1344 12518 9782 12570
rect 9834 12518 9886 12570
rect 9938 12518 9990 12570
rect 10042 12518 18350 12570
rect 18402 12518 18454 12570
rect 18506 12518 18558 12570
rect 18610 12518 26918 12570
rect 26970 12518 27022 12570
rect 27074 12518 27126 12570
rect 27178 12518 35486 12570
rect 35538 12518 35590 12570
rect 35642 12518 35694 12570
rect 35746 12518 35776 12570
rect 1344 12484 35776 12518
rect 7982 12402 8034 12414
rect 8990 12402 9042 12414
rect 8642 12350 8654 12402
rect 8706 12350 8718 12402
rect 7982 12338 8034 12350
rect 8990 12338 9042 12350
rect 13582 12402 13634 12414
rect 13582 12338 13634 12350
rect 21198 12402 21250 12414
rect 21198 12338 21250 12350
rect 22206 12402 22258 12414
rect 22206 12338 22258 12350
rect 23662 12402 23714 12414
rect 23662 12338 23714 12350
rect 32062 12402 32114 12414
rect 32062 12338 32114 12350
rect 32286 12402 32338 12414
rect 32286 12338 32338 12350
rect 33182 12402 33234 12414
rect 33182 12338 33234 12350
rect 34862 12402 34914 12414
rect 34862 12338 34914 12350
rect 8206 12290 8258 12302
rect 6962 12238 6974 12290
rect 7026 12238 7038 12290
rect 8206 12226 8258 12238
rect 8318 12290 8370 12302
rect 22318 12290 22370 12302
rect 13234 12238 13246 12290
rect 13298 12238 13310 12290
rect 18722 12238 18734 12290
rect 18786 12238 18798 12290
rect 8318 12226 8370 12238
rect 22318 12226 22370 12238
rect 22654 12290 22706 12302
rect 24098 12238 24110 12290
rect 24162 12238 24174 12290
rect 33730 12238 33742 12290
rect 33794 12238 33806 12290
rect 34066 12238 34078 12290
rect 34130 12238 34142 12290
rect 22654 12226 22706 12238
rect 22990 12178 23042 12190
rect 7634 12126 7646 12178
rect 7698 12126 7710 12178
rect 11666 12126 11678 12178
rect 11730 12126 11742 12178
rect 12450 12126 12462 12178
rect 12514 12126 12526 12178
rect 13906 12126 13918 12178
rect 13970 12126 13982 12178
rect 17938 12126 17950 12178
rect 18002 12126 18014 12178
rect 22990 12114 23042 12126
rect 23214 12178 23266 12190
rect 32398 12178 32450 12190
rect 24546 12126 24558 12178
rect 24610 12126 24622 12178
rect 25442 12126 25454 12178
rect 25506 12126 25518 12178
rect 25890 12126 25902 12178
rect 25954 12126 25966 12178
rect 27234 12126 27246 12178
rect 27298 12126 27310 12178
rect 35074 12126 35086 12178
rect 35138 12126 35150 12178
rect 23214 12114 23266 12126
rect 32398 12114 32450 12126
rect 21758 12066 21810 12078
rect 4834 12014 4846 12066
rect 4898 12014 4910 12066
rect 9538 12014 9550 12066
rect 9602 12014 9614 12066
rect 14690 12014 14702 12066
rect 14754 12014 14766 12066
rect 16818 12014 16830 12066
rect 16882 12014 16894 12066
rect 20850 12014 20862 12066
rect 20914 12014 20926 12066
rect 21758 12002 21810 12014
rect 22766 12066 22818 12078
rect 24658 12014 24670 12066
rect 24722 12014 24734 12066
rect 30034 12014 30046 12066
rect 30098 12014 30110 12066
rect 22766 12002 22818 12014
rect 33518 11954 33570 11966
rect 25890 11902 25902 11954
rect 25954 11902 25966 11954
rect 33518 11890 33570 11902
rect 1344 11786 35616 11820
rect 1344 11734 5498 11786
rect 5550 11734 5602 11786
rect 5654 11734 5706 11786
rect 5758 11734 14066 11786
rect 14118 11734 14170 11786
rect 14222 11734 14274 11786
rect 14326 11734 22634 11786
rect 22686 11734 22738 11786
rect 22790 11734 22842 11786
rect 22894 11734 31202 11786
rect 31254 11734 31306 11786
rect 31358 11734 31410 11786
rect 31462 11734 35616 11786
rect 1344 11700 35616 11734
rect 27918 11618 27970 11630
rect 27918 11554 27970 11566
rect 28478 11618 28530 11630
rect 28478 11554 28530 11566
rect 9886 11506 9938 11518
rect 5618 11454 5630 11506
rect 5682 11454 5694 11506
rect 7746 11454 7758 11506
rect 7810 11454 7822 11506
rect 9886 11442 9938 11454
rect 10558 11506 10610 11518
rect 10558 11442 10610 11454
rect 14926 11506 14978 11518
rect 14926 11442 14978 11454
rect 19406 11506 19458 11518
rect 19406 11442 19458 11454
rect 20638 11506 20690 11518
rect 26798 11506 26850 11518
rect 33518 11506 33570 11518
rect 22418 11454 22430 11506
rect 22482 11454 22494 11506
rect 24546 11454 24558 11506
rect 24610 11454 24622 11506
rect 29586 11454 29598 11506
rect 29650 11454 29662 11506
rect 32946 11454 32958 11506
rect 33010 11454 33022 11506
rect 34626 11454 34638 11506
rect 34690 11454 34702 11506
rect 20638 11442 20690 11454
rect 26798 11442 26850 11454
rect 33518 11442 33570 11454
rect 10446 11394 10498 11406
rect 11454 11394 11506 11406
rect 8530 11342 8542 11394
rect 8594 11342 8606 11394
rect 10994 11342 11006 11394
rect 11058 11342 11070 11394
rect 10446 11330 10498 11342
rect 11454 11330 11506 11342
rect 11902 11394 11954 11406
rect 11902 11330 11954 11342
rect 15038 11394 15090 11406
rect 15038 11330 15090 11342
rect 15374 11394 15426 11406
rect 15374 11330 15426 11342
rect 15822 11394 15874 11406
rect 15822 11330 15874 11342
rect 15934 11394 15986 11406
rect 15934 11330 15986 11342
rect 17166 11394 17218 11406
rect 17166 11330 17218 11342
rect 19518 11394 19570 11406
rect 29150 11394 29202 11406
rect 33854 11394 33906 11406
rect 20178 11342 20190 11394
rect 20242 11342 20254 11394
rect 21634 11342 21646 11394
rect 21698 11342 21710 11394
rect 25442 11342 25454 11394
rect 25506 11342 25518 11394
rect 26002 11342 26014 11394
rect 26066 11342 26078 11394
rect 27346 11342 27358 11394
rect 27410 11342 27422 11394
rect 27570 11342 27582 11394
rect 27634 11342 27646 11394
rect 30034 11342 30046 11394
rect 30098 11342 30110 11394
rect 19518 11330 19570 11342
rect 29150 11330 29202 11342
rect 33854 11330 33906 11342
rect 35086 11394 35138 11406
rect 35086 11330 35138 11342
rect 10670 11282 10722 11294
rect 10670 11218 10722 11230
rect 14814 11282 14866 11294
rect 14814 11218 14866 11230
rect 16606 11282 16658 11294
rect 16606 11218 16658 11230
rect 26238 11282 26290 11294
rect 26238 11218 26290 11230
rect 27806 11282 27858 11294
rect 27806 11218 27858 11230
rect 28366 11282 28418 11294
rect 34190 11282 34242 11294
rect 30818 11230 30830 11282
rect 30882 11230 30894 11282
rect 28366 11218 28418 11230
rect 34190 11218 34242 11230
rect 9438 11170 9490 11182
rect 9090 11118 9102 11170
rect 9154 11118 9166 11170
rect 9438 11106 9490 11118
rect 15710 11170 15762 11182
rect 15710 11106 15762 11118
rect 16158 11170 16210 11182
rect 16158 11106 16210 11118
rect 19294 11170 19346 11182
rect 19294 11106 19346 11118
rect 19742 11170 19794 11182
rect 19742 11106 19794 11118
rect 20526 11170 20578 11182
rect 20526 11106 20578 11118
rect 20750 11170 20802 11182
rect 20750 11106 20802 11118
rect 24894 11170 24946 11182
rect 24894 11106 24946 11118
rect 25006 11170 25058 11182
rect 25006 11106 25058 11118
rect 25118 11170 25170 11182
rect 25118 11106 25170 11118
rect 1344 11002 35776 11036
rect 1344 10950 9782 11002
rect 9834 10950 9886 11002
rect 9938 10950 9990 11002
rect 10042 10950 18350 11002
rect 18402 10950 18454 11002
rect 18506 10950 18558 11002
rect 18610 10950 26918 11002
rect 26970 10950 27022 11002
rect 27074 10950 27126 11002
rect 27178 10950 35486 11002
rect 35538 10950 35590 11002
rect 35642 10950 35694 11002
rect 35746 10950 35776 11002
rect 1344 10916 35776 10950
rect 7982 10834 8034 10846
rect 7982 10770 8034 10782
rect 9662 10834 9714 10846
rect 9662 10770 9714 10782
rect 10334 10834 10386 10846
rect 10334 10770 10386 10782
rect 12014 10834 12066 10846
rect 12014 10770 12066 10782
rect 21422 10834 21474 10846
rect 21422 10770 21474 10782
rect 21646 10834 21698 10846
rect 21646 10770 21698 10782
rect 22318 10834 22370 10846
rect 22318 10770 22370 10782
rect 22766 10834 22818 10846
rect 22766 10770 22818 10782
rect 23326 10834 23378 10846
rect 23326 10770 23378 10782
rect 23662 10834 23714 10846
rect 23662 10770 23714 10782
rect 23774 10834 23826 10846
rect 23774 10770 23826 10782
rect 24334 10834 24386 10846
rect 24334 10770 24386 10782
rect 26574 10834 26626 10846
rect 26574 10770 26626 10782
rect 27358 10834 27410 10846
rect 27358 10770 27410 10782
rect 31054 10834 31106 10846
rect 31054 10770 31106 10782
rect 31278 10834 31330 10846
rect 31278 10770 31330 10782
rect 32286 10834 32338 10846
rect 32286 10770 32338 10782
rect 33518 10834 33570 10846
rect 33518 10770 33570 10782
rect 33854 10834 33906 10846
rect 33854 10770 33906 10782
rect 20862 10722 20914 10734
rect 20862 10658 20914 10670
rect 21086 10722 21138 10734
rect 21086 10658 21138 10670
rect 22430 10722 22482 10734
rect 22430 10658 22482 10670
rect 25566 10722 25618 10734
rect 30830 10722 30882 10734
rect 29698 10670 29710 10722
rect 29762 10670 29774 10722
rect 25566 10658 25618 10670
rect 30830 10658 30882 10670
rect 31838 10722 31890 10734
rect 31838 10658 31890 10670
rect 9774 10610 9826 10622
rect 15598 10610 15650 10622
rect 12450 10558 12462 10610
rect 12514 10558 12526 10610
rect 9774 10546 9826 10558
rect 15598 10546 15650 10558
rect 15822 10610 15874 10622
rect 20526 10610 20578 10622
rect 16146 10558 16158 10610
rect 16210 10558 16222 10610
rect 15822 10546 15874 10558
rect 20526 10546 20578 10558
rect 21534 10610 21586 10622
rect 21534 10546 21586 10558
rect 22094 10610 22146 10622
rect 22094 10546 22146 10558
rect 22542 10610 22594 10622
rect 22542 10546 22594 10558
rect 23550 10610 23602 10622
rect 23550 10546 23602 10558
rect 24110 10610 24162 10622
rect 24110 10546 24162 10558
rect 24222 10610 24274 10622
rect 25230 10610 25282 10622
rect 24658 10558 24670 10610
rect 24722 10558 24734 10610
rect 24222 10546 24274 10558
rect 25230 10546 25282 10558
rect 25678 10610 25730 10622
rect 34190 10610 34242 10622
rect 35086 10610 35138 10622
rect 30482 10558 30494 10610
rect 30546 10558 30558 10610
rect 34626 10558 34638 10610
rect 34690 10558 34702 10610
rect 25678 10546 25730 10558
rect 34190 10546 34242 10558
rect 35086 10546 35138 10558
rect 10894 10498 10946 10510
rect 15710 10498 15762 10510
rect 13122 10446 13134 10498
rect 13186 10446 13198 10498
rect 15250 10446 15262 10498
rect 15314 10446 15326 10498
rect 10894 10434 10946 10446
rect 15710 10434 15762 10446
rect 20638 10498 20690 10510
rect 20638 10434 20690 10446
rect 25342 10498 25394 10510
rect 30942 10498 30994 10510
rect 27570 10446 27582 10498
rect 27634 10446 27646 10498
rect 25342 10434 25394 10446
rect 30942 10434 30994 10446
rect 9662 10386 9714 10398
rect 9662 10322 9714 10334
rect 1344 10218 35616 10252
rect 1344 10166 5498 10218
rect 5550 10166 5602 10218
rect 5654 10166 5706 10218
rect 5758 10166 14066 10218
rect 14118 10166 14170 10218
rect 14222 10166 14274 10218
rect 14326 10166 22634 10218
rect 22686 10166 22738 10218
rect 22790 10166 22842 10218
rect 22894 10166 31202 10218
rect 31254 10166 31306 10218
rect 31358 10166 31410 10218
rect 31462 10166 35616 10218
rect 1344 10132 35616 10166
rect 29250 9998 29262 10050
rect 29314 10047 29326 10050
rect 29474 10047 29486 10050
rect 29314 10001 29486 10047
rect 29314 9998 29326 10001
rect 29474 9998 29486 10001
rect 29538 9998 29550 10050
rect 14142 9938 14194 9950
rect 9874 9886 9886 9938
rect 9938 9886 9950 9938
rect 14142 9874 14194 9886
rect 18286 9938 18338 9950
rect 18286 9874 18338 9886
rect 22654 9938 22706 9950
rect 27358 9938 27410 9950
rect 24770 9886 24782 9938
rect 24834 9886 24846 9938
rect 26898 9886 26910 9938
rect 26962 9886 26974 9938
rect 22654 9874 22706 9886
rect 27358 9874 27410 9886
rect 29486 9938 29538 9950
rect 29486 9874 29538 9886
rect 30158 9938 30210 9950
rect 30158 9874 30210 9886
rect 32734 9938 32786 9950
rect 32734 9874 32786 9886
rect 33182 9938 33234 9950
rect 33182 9874 33234 9886
rect 33630 9938 33682 9950
rect 33630 9874 33682 9886
rect 34078 9938 34130 9950
rect 34078 9874 34130 9886
rect 10670 9826 10722 9838
rect 7074 9774 7086 9826
rect 7138 9774 7150 9826
rect 10670 9762 10722 9774
rect 11118 9826 11170 9838
rect 11118 9762 11170 9774
rect 11566 9826 11618 9838
rect 11566 9762 11618 9774
rect 11790 9826 11842 9838
rect 11790 9762 11842 9774
rect 12350 9826 12402 9838
rect 12350 9762 12402 9774
rect 12910 9826 12962 9838
rect 12910 9762 12962 9774
rect 14590 9826 14642 9838
rect 16046 9826 16098 9838
rect 14914 9774 14926 9826
rect 14978 9774 14990 9826
rect 14590 9762 14642 9774
rect 16046 9762 16098 9774
rect 16942 9826 16994 9838
rect 22542 9826 22594 9838
rect 20290 9774 20302 9826
rect 20354 9774 20366 9826
rect 16942 9762 16994 9774
rect 22542 9762 22594 9774
rect 23214 9826 23266 9838
rect 28254 9826 28306 9838
rect 24098 9774 24110 9826
rect 24162 9774 24174 9826
rect 23214 9762 23266 9774
rect 28254 9762 28306 9774
rect 29822 9826 29874 9838
rect 29822 9762 29874 9774
rect 30382 9826 30434 9838
rect 30382 9762 30434 9774
rect 30830 9826 30882 9838
rect 30830 9762 30882 9774
rect 34638 9826 34690 9838
rect 34638 9762 34690 9774
rect 35198 9826 35250 9838
rect 35198 9762 35250 9774
rect 14030 9714 14082 9726
rect 7746 9662 7758 9714
rect 7810 9662 7822 9714
rect 14030 9650 14082 9662
rect 14366 9714 14418 9726
rect 14366 9650 14418 9662
rect 16718 9714 16770 9726
rect 16718 9650 16770 9662
rect 17278 9714 17330 9726
rect 17278 9650 17330 9662
rect 17502 9714 17554 9726
rect 17502 9650 17554 9662
rect 17838 9714 17890 9726
rect 29934 9714 29986 9726
rect 20514 9662 20526 9714
rect 20578 9662 20590 9714
rect 22082 9662 22094 9714
rect 22146 9662 22158 9714
rect 28578 9662 28590 9714
rect 28642 9662 28654 9714
rect 17838 9650 17890 9662
rect 11454 9602 11506 9614
rect 10322 9550 10334 9602
rect 10386 9550 10398 9602
rect 11454 9538 11506 9550
rect 12238 9602 12290 9614
rect 12238 9538 12290 9550
rect 12462 9602 12514 9614
rect 12462 9538 12514 9550
rect 13582 9602 13634 9614
rect 13582 9538 13634 9550
rect 15262 9602 15314 9614
rect 15262 9538 15314 9550
rect 15374 9602 15426 9614
rect 15374 9538 15426 9550
rect 15486 9602 15538 9614
rect 15486 9538 15538 9550
rect 15822 9602 15874 9614
rect 15822 9538 15874 9550
rect 15934 9602 15986 9614
rect 15934 9538 15986 9550
rect 16270 9602 16322 9614
rect 16270 9538 16322 9550
rect 17166 9602 17218 9614
rect 17166 9538 17218 9550
rect 17726 9602 17778 9614
rect 22097 9599 22143 9662
rect 29934 9650 29986 9662
rect 30606 9714 30658 9726
rect 30606 9650 30658 9662
rect 31166 9714 31218 9726
rect 31166 9650 31218 9662
rect 34862 9714 34914 9726
rect 34862 9650 34914 9662
rect 22766 9602 22818 9614
rect 22306 9599 22318 9602
rect 22097 9553 22318 9599
rect 22306 9550 22318 9553
rect 22370 9550 22382 9602
rect 17726 9538 17778 9550
rect 22766 9538 22818 9550
rect 30718 9602 30770 9614
rect 30718 9538 30770 9550
rect 1344 9434 35776 9468
rect 1344 9382 9782 9434
rect 9834 9382 9886 9434
rect 9938 9382 9990 9434
rect 10042 9382 18350 9434
rect 18402 9382 18454 9434
rect 18506 9382 18558 9434
rect 18610 9382 26918 9434
rect 26970 9382 27022 9434
rect 27074 9382 27126 9434
rect 27178 9382 35486 9434
rect 35538 9382 35590 9434
rect 35642 9382 35694 9434
rect 35746 9382 35776 9434
rect 1344 9348 35776 9382
rect 8206 9266 8258 9278
rect 8206 9202 8258 9214
rect 16158 9266 16210 9278
rect 16158 9202 16210 9214
rect 16606 9266 16658 9278
rect 16606 9202 16658 9214
rect 22430 9266 22482 9278
rect 22430 9202 22482 9214
rect 23774 9266 23826 9278
rect 23774 9202 23826 9214
rect 24782 9266 24834 9278
rect 24782 9202 24834 9214
rect 25230 9266 25282 9278
rect 26014 9266 26066 9278
rect 25554 9214 25566 9266
rect 25618 9214 25630 9266
rect 25230 9202 25282 9214
rect 26014 9202 26066 9214
rect 26350 9266 26402 9278
rect 26350 9202 26402 9214
rect 30606 9266 30658 9278
rect 30606 9202 30658 9214
rect 31390 9266 31442 9278
rect 31390 9202 31442 9214
rect 31502 9266 31554 9278
rect 31502 9202 31554 9214
rect 33966 9266 34018 9278
rect 33966 9202 34018 9214
rect 34414 9266 34466 9278
rect 34414 9202 34466 9214
rect 34862 9266 34914 9278
rect 34862 9202 34914 9214
rect 35198 9266 35250 9278
rect 35198 9202 35250 9214
rect 17390 9154 17442 9166
rect 22654 9154 22706 9166
rect 7410 9102 7422 9154
rect 7474 9102 7486 9154
rect 18274 9102 18286 9154
rect 18338 9102 18350 9154
rect 20066 9102 20078 9154
rect 20130 9102 20142 9154
rect 17390 9090 17442 9102
rect 22654 9090 22706 9102
rect 23998 9154 24050 9166
rect 23998 9090 24050 9102
rect 24110 9154 24162 9166
rect 24110 9090 24162 9102
rect 24558 9154 24610 9166
rect 32398 9154 32450 9166
rect 26674 9102 26686 9154
rect 26738 9102 26750 9154
rect 28018 9102 28030 9154
rect 28082 9102 28094 9154
rect 24558 9090 24610 9102
rect 32398 9090 32450 9102
rect 8094 9042 8146 9054
rect 7074 8990 7086 9042
rect 7138 8990 7150 9042
rect 7634 8990 7646 9042
rect 7698 8990 7710 9042
rect 8094 8978 8146 8990
rect 8430 9042 8482 9054
rect 8430 8978 8482 8990
rect 8654 9042 8706 9054
rect 16382 9042 16434 9054
rect 14802 8990 14814 9042
rect 14866 8990 14878 9042
rect 8654 8978 8706 8990
rect 16382 8978 16434 8990
rect 16494 9042 16546 9054
rect 16494 8978 16546 8990
rect 17614 9042 17666 9054
rect 17614 8978 17666 8990
rect 18062 9042 18114 9054
rect 18062 8978 18114 8990
rect 18622 9042 18674 9054
rect 22766 9042 22818 9054
rect 19282 8990 19294 9042
rect 19346 8990 19358 9042
rect 18622 8978 18674 8990
rect 22766 8978 22818 8990
rect 24446 9042 24498 9054
rect 30494 9042 30546 9054
rect 27346 8990 27358 9042
rect 27410 8990 27422 9042
rect 24446 8978 24498 8990
rect 30494 8978 30546 8990
rect 30718 9042 30770 9054
rect 30718 8978 30770 8990
rect 31166 9042 31218 9054
rect 31166 8978 31218 8990
rect 31614 9042 31666 9054
rect 32286 9042 32338 9054
rect 31938 8990 31950 9042
rect 32002 8990 32014 9042
rect 31614 8978 31666 8990
rect 32286 8978 32338 8990
rect 15262 8930 15314 8942
rect 4162 8878 4174 8930
rect 4226 8878 4238 8930
rect 6290 8878 6302 8930
rect 6354 8878 6366 8930
rect 12114 8878 12126 8930
rect 12178 8878 12190 8930
rect 15262 8866 15314 8878
rect 15710 8930 15762 8942
rect 15710 8866 15762 8878
rect 17502 8930 17554 8942
rect 22194 8878 22206 8930
rect 22258 8878 22270 8930
rect 30146 8878 30158 8930
rect 30210 8878 30222 8930
rect 17502 8866 17554 8878
rect 32398 8818 32450 8830
rect 32398 8754 32450 8766
rect 1344 8650 35616 8684
rect 1344 8598 5498 8650
rect 5550 8598 5602 8650
rect 5654 8598 5706 8650
rect 5758 8598 14066 8650
rect 14118 8598 14170 8650
rect 14222 8598 14274 8650
rect 14326 8598 22634 8650
rect 22686 8598 22738 8650
rect 22790 8598 22842 8650
rect 22894 8598 31202 8650
rect 31254 8598 31306 8650
rect 31358 8598 31410 8650
rect 31462 8598 35616 8650
rect 1344 8564 35616 8598
rect 6638 8370 6690 8382
rect 6638 8306 6690 8318
rect 8542 8370 8594 8382
rect 8542 8306 8594 8318
rect 9438 8370 9490 8382
rect 21534 8370 21586 8382
rect 9762 8318 9774 8370
rect 9826 8318 9838 8370
rect 11890 8318 11902 8370
rect 11954 8318 11966 8370
rect 19282 8318 19294 8370
rect 19346 8318 19358 8370
rect 9438 8306 9490 8318
rect 21534 8306 21586 8318
rect 25006 8370 25058 8382
rect 25006 8306 25058 8318
rect 29934 8370 29986 8382
rect 34178 8318 34190 8370
rect 34242 8318 34254 8370
rect 29934 8306 29986 8318
rect 6862 8258 6914 8270
rect 6862 8194 6914 8206
rect 7086 8258 7138 8270
rect 7086 8194 7138 8206
rect 7534 8258 7586 8270
rect 7534 8194 7586 8206
rect 7646 8258 7698 8270
rect 7646 8194 7698 8206
rect 8094 8258 8146 8270
rect 8094 8194 8146 8206
rect 9102 8258 9154 8270
rect 14142 8258 14194 8270
rect 12562 8206 12574 8258
rect 12626 8206 12638 8258
rect 9102 8194 9154 8206
rect 14142 8194 14194 8206
rect 14478 8258 14530 8270
rect 14478 8194 14530 8206
rect 14702 8258 14754 8270
rect 29822 8258 29874 8270
rect 16706 8206 16718 8258
rect 16770 8206 16782 8258
rect 27234 8206 27246 8258
rect 27298 8206 27310 8258
rect 14702 8194 14754 8206
rect 29822 8194 29874 8206
rect 30718 8258 30770 8270
rect 31266 8206 31278 8258
rect 31330 8206 31342 8258
rect 30718 8194 30770 8206
rect 5966 8146 6018 8158
rect 5966 8082 6018 8094
rect 6302 8146 6354 8158
rect 6302 8082 6354 8094
rect 6526 8146 6578 8158
rect 6526 8082 6578 8094
rect 13582 8146 13634 8158
rect 13582 8082 13634 8094
rect 13694 8146 13746 8158
rect 13694 8082 13746 8094
rect 28030 8146 28082 8158
rect 28030 8082 28082 8094
rect 30046 8146 30098 8158
rect 34862 8146 34914 8158
rect 32050 8094 32062 8146
rect 32114 8094 32126 8146
rect 30046 8082 30098 8094
rect 34862 8082 34914 8094
rect 35198 8146 35250 8158
rect 35198 8082 35250 8094
rect 6078 8034 6130 8046
rect 6078 7970 6130 7982
rect 7422 8034 7474 8046
rect 7422 7970 7474 7982
rect 8430 8034 8482 8046
rect 8430 7970 8482 7982
rect 8654 8034 8706 8046
rect 8654 7970 8706 7982
rect 13918 8034 13970 8046
rect 13918 7970 13970 7982
rect 14254 8034 14306 8046
rect 14254 7970 14306 7982
rect 27470 8034 27522 8046
rect 29598 8034 29650 8046
rect 28354 7982 28366 8034
rect 28418 7982 28430 8034
rect 27470 7970 27522 7982
rect 29598 7970 29650 7982
rect 30494 8034 30546 8046
rect 30494 7970 30546 7982
rect 30830 8034 30882 8046
rect 30830 7970 30882 7982
rect 30942 8034 30994 8046
rect 30942 7970 30994 7982
rect 1344 7866 35776 7900
rect 1344 7814 9782 7866
rect 9834 7814 9886 7866
rect 9938 7814 9990 7866
rect 10042 7814 18350 7866
rect 18402 7814 18454 7866
rect 18506 7814 18558 7866
rect 18610 7814 26918 7866
rect 26970 7814 27022 7866
rect 27074 7814 27126 7866
rect 27178 7814 35486 7866
rect 35538 7814 35590 7866
rect 35642 7814 35694 7866
rect 35746 7814 35776 7866
rect 1344 7780 35776 7814
rect 7086 7698 7138 7710
rect 7086 7634 7138 7646
rect 9102 7698 9154 7710
rect 9102 7634 9154 7646
rect 10782 7698 10834 7710
rect 15598 7698 15650 7710
rect 11106 7646 11118 7698
rect 11170 7646 11182 7698
rect 10782 7634 10834 7646
rect 15598 7634 15650 7646
rect 15710 7698 15762 7710
rect 15710 7634 15762 7646
rect 15822 7698 15874 7710
rect 17726 7698 17778 7710
rect 17378 7646 17390 7698
rect 17442 7646 17454 7698
rect 15822 7634 15874 7646
rect 17726 7634 17778 7646
rect 18398 7698 18450 7710
rect 18398 7634 18450 7646
rect 20190 7698 20242 7710
rect 20190 7634 20242 7646
rect 20750 7698 20802 7710
rect 20750 7634 20802 7646
rect 24446 7698 24498 7710
rect 24446 7634 24498 7646
rect 25902 7698 25954 7710
rect 25902 7634 25954 7646
rect 29374 7698 29426 7710
rect 29374 7634 29426 7646
rect 29598 7698 29650 7710
rect 29598 7634 29650 7646
rect 29822 7698 29874 7710
rect 29822 7634 29874 7646
rect 31166 7698 31218 7710
rect 31166 7634 31218 7646
rect 31614 7698 31666 7710
rect 31614 7634 31666 7646
rect 32062 7698 32114 7710
rect 32062 7634 32114 7646
rect 33966 7698 34018 7710
rect 33966 7634 34018 7646
rect 35310 7698 35362 7710
rect 35310 7634 35362 7646
rect 6414 7586 6466 7598
rect 6414 7522 6466 7534
rect 7982 7586 8034 7598
rect 7982 7522 8034 7534
rect 9550 7586 9602 7598
rect 9550 7522 9602 7534
rect 11566 7586 11618 7598
rect 18510 7586 18562 7598
rect 12898 7534 12910 7586
rect 12962 7534 12974 7586
rect 16482 7534 16494 7586
rect 16546 7534 16558 7586
rect 11566 7522 11618 7534
rect 18510 7522 18562 7534
rect 18846 7586 18898 7598
rect 18846 7522 18898 7534
rect 19182 7586 19234 7598
rect 19182 7522 19234 7534
rect 19518 7586 19570 7598
rect 19518 7522 19570 7534
rect 19854 7586 19906 7598
rect 19854 7522 19906 7534
rect 20974 7586 21026 7598
rect 20974 7522 21026 7534
rect 21086 7586 21138 7598
rect 21086 7522 21138 7534
rect 21422 7586 21474 7598
rect 21422 7522 21474 7534
rect 21534 7586 21586 7598
rect 21534 7522 21586 7534
rect 25342 7586 25394 7598
rect 25342 7522 25394 7534
rect 26574 7586 26626 7598
rect 27582 7586 27634 7598
rect 27234 7534 27246 7586
rect 27298 7534 27310 7586
rect 26574 7522 26626 7534
rect 27582 7522 27634 7534
rect 28030 7586 28082 7598
rect 28030 7522 28082 7534
rect 28590 7586 28642 7598
rect 28590 7522 28642 7534
rect 30046 7586 30098 7598
rect 30046 7522 30098 7534
rect 30270 7586 30322 7598
rect 30270 7522 30322 7534
rect 31838 7586 31890 7598
rect 31838 7522 31890 7534
rect 6302 7474 6354 7486
rect 6302 7410 6354 7422
rect 6862 7474 6914 7486
rect 6862 7410 6914 7422
rect 7198 7474 7250 7486
rect 7198 7410 7250 7422
rect 7310 7474 7362 7486
rect 7310 7410 7362 7422
rect 7758 7474 7810 7486
rect 7758 7410 7810 7422
rect 8206 7474 8258 7486
rect 11454 7474 11506 7486
rect 16270 7474 16322 7486
rect 18174 7474 18226 7486
rect 23438 7474 23490 7486
rect 8530 7422 8542 7474
rect 8594 7422 8606 7474
rect 9986 7422 9998 7474
rect 10050 7422 10062 7474
rect 12114 7422 12126 7474
rect 12178 7422 12190 7474
rect 16706 7422 16718 7474
rect 16770 7422 16782 7474
rect 20402 7422 20414 7474
rect 20466 7422 20478 7474
rect 8206 7410 8258 7422
rect 11454 7410 11506 7422
rect 16270 7410 16322 7422
rect 18174 7410 18226 7422
rect 23438 7410 23490 7422
rect 23774 7474 23826 7486
rect 23774 7410 23826 7422
rect 23998 7474 24050 7486
rect 23998 7410 24050 7422
rect 24222 7474 24274 7486
rect 24222 7410 24274 7422
rect 24558 7474 24610 7486
rect 24558 7410 24610 7422
rect 25118 7474 25170 7486
rect 25118 7410 25170 7422
rect 25454 7474 25506 7486
rect 25454 7410 25506 7422
rect 25790 7474 25842 7486
rect 25790 7410 25842 7422
rect 26126 7474 26178 7486
rect 27806 7474 27858 7486
rect 26786 7422 26798 7474
rect 26850 7422 26862 7474
rect 26126 7410 26178 7422
rect 27806 7410 27858 7422
rect 28142 7474 28194 7486
rect 28142 7410 28194 7422
rect 28478 7474 28530 7486
rect 28478 7410 28530 7422
rect 28814 7474 28866 7486
rect 28814 7410 28866 7422
rect 29262 7474 29314 7486
rect 29262 7410 29314 7422
rect 29934 7474 29986 7486
rect 29934 7410 29986 7422
rect 30830 7474 30882 7486
rect 30830 7410 30882 7422
rect 31054 7474 31106 7486
rect 31054 7410 31106 7422
rect 31278 7474 31330 7486
rect 31278 7410 31330 7422
rect 6638 7362 6690 7374
rect 6638 7298 6690 7310
rect 8094 7362 8146 7374
rect 23550 7362 23602 7374
rect 15026 7310 15038 7362
rect 15090 7310 15102 7362
rect 8094 7298 8146 7310
rect 23550 7298 23602 7310
rect 31726 7362 31778 7374
rect 31726 7298 31778 7310
rect 34078 7362 34130 7374
rect 34078 7298 34130 7310
rect 11566 7250 11618 7262
rect 11566 7186 11618 7198
rect 21534 7250 21586 7262
rect 21534 7186 21586 7198
rect 1344 7082 35616 7116
rect 1344 7030 5498 7082
rect 5550 7030 5602 7082
rect 5654 7030 5706 7082
rect 5758 7030 14066 7082
rect 14118 7030 14170 7082
rect 14222 7030 14274 7082
rect 14326 7030 22634 7082
rect 22686 7030 22738 7082
rect 22790 7030 22842 7082
rect 22894 7030 31202 7082
rect 31254 7030 31306 7082
rect 31358 7030 31410 7082
rect 31462 7030 35616 7082
rect 1344 6996 35616 7030
rect 15026 6750 15038 6802
rect 15090 6750 15102 6802
rect 24210 6750 24222 6802
rect 24274 6750 24286 6802
rect 6526 6690 6578 6702
rect 6526 6626 6578 6638
rect 6750 6690 6802 6702
rect 6750 6626 6802 6638
rect 7198 6690 7250 6702
rect 13918 6690 13970 6702
rect 18734 6690 18786 6702
rect 9650 6638 9662 6690
rect 9714 6638 9726 6690
rect 12450 6638 12462 6690
rect 12514 6638 12526 6690
rect 17154 6638 17166 6690
rect 17218 6638 17230 6690
rect 17938 6638 17950 6690
rect 18002 6638 18014 6690
rect 7198 6626 7250 6638
rect 13918 6626 13970 6638
rect 18734 6626 18786 6638
rect 19294 6690 19346 6702
rect 19294 6626 19346 6638
rect 19630 6690 19682 6702
rect 19630 6626 19682 6638
rect 20302 6690 20354 6702
rect 20302 6626 20354 6638
rect 20862 6690 20914 6702
rect 25566 6690 25618 6702
rect 21298 6638 21310 6690
rect 21362 6638 21374 6690
rect 22082 6638 22094 6690
rect 22146 6638 22158 6690
rect 25106 6638 25118 6690
rect 25170 6638 25182 6690
rect 20862 6626 20914 6638
rect 25566 6626 25618 6638
rect 25678 6690 25730 6702
rect 25678 6626 25730 6638
rect 26462 6690 26514 6702
rect 26462 6626 26514 6638
rect 26910 6690 26962 6702
rect 26910 6626 26962 6638
rect 27470 6690 27522 6702
rect 27470 6626 27522 6638
rect 28142 6690 28194 6702
rect 28142 6626 28194 6638
rect 29038 6690 29090 6702
rect 29038 6626 29090 6638
rect 29598 6690 29650 6702
rect 29598 6626 29650 6638
rect 29934 6690 29986 6702
rect 29934 6626 29986 6638
rect 30382 6690 30434 6702
rect 30382 6626 30434 6638
rect 30606 6690 30658 6702
rect 30606 6626 30658 6638
rect 31166 6690 31218 6702
rect 31166 6626 31218 6638
rect 14478 6578 14530 6590
rect 8306 6526 8318 6578
rect 8370 6526 8382 6578
rect 11218 6526 11230 6578
rect 11282 6526 11294 6578
rect 14478 6514 14530 6526
rect 18286 6578 18338 6590
rect 18286 6514 18338 6526
rect 18622 6578 18674 6590
rect 18622 6514 18674 6526
rect 19182 6578 19234 6590
rect 19182 6514 19234 6526
rect 20078 6578 20130 6590
rect 20078 6514 20130 6526
rect 24558 6578 24610 6590
rect 24558 6514 24610 6526
rect 26014 6578 26066 6590
rect 26014 6514 26066 6526
rect 6862 6466 6914 6478
rect 6862 6402 6914 6414
rect 14030 6466 14082 6478
rect 14030 6402 14082 6414
rect 14254 6466 14306 6478
rect 14254 6402 14306 6414
rect 14590 6466 14642 6478
rect 14590 6402 14642 6414
rect 14814 6466 14866 6478
rect 14814 6402 14866 6414
rect 18398 6466 18450 6478
rect 18398 6402 18450 6414
rect 18958 6466 19010 6478
rect 18958 6402 19010 6414
rect 19966 6466 20018 6478
rect 19966 6402 20018 6414
rect 24670 6466 24722 6478
rect 24670 6402 24722 6414
rect 24782 6466 24834 6478
rect 24782 6402 24834 6414
rect 25902 6466 25954 6478
rect 29486 6466 29538 6478
rect 27794 6414 27806 6466
rect 27858 6414 27870 6466
rect 25902 6402 25954 6414
rect 29486 6402 29538 6414
rect 29710 6466 29762 6478
rect 29710 6402 29762 6414
rect 30158 6466 30210 6478
rect 30158 6402 30210 6414
rect 30830 6466 30882 6478
rect 30830 6402 30882 6414
rect 31054 6466 31106 6478
rect 31054 6402 31106 6414
rect 1344 6298 35776 6332
rect 1344 6246 9782 6298
rect 9834 6246 9886 6298
rect 9938 6246 9990 6298
rect 10042 6246 18350 6298
rect 18402 6246 18454 6298
rect 18506 6246 18558 6298
rect 18610 6246 26918 6298
rect 26970 6246 27022 6298
rect 27074 6246 27126 6298
rect 27178 6246 35486 6298
rect 35538 6246 35590 6298
rect 35642 6246 35694 6298
rect 35746 6246 35776 6298
rect 1344 6212 35776 6246
rect 5742 6130 5794 6142
rect 5742 6066 5794 6078
rect 20190 6130 20242 6142
rect 20190 6066 20242 6078
rect 24222 6130 24274 6142
rect 24222 6066 24274 6078
rect 24334 6130 24386 6142
rect 24334 6066 24386 6078
rect 24558 6130 24610 6142
rect 24558 6066 24610 6078
rect 26686 6130 26738 6142
rect 26686 6066 26738 6078
rect 27022 6130 27074 6142
rect 27022 6066 27074 6078
rect 28142 6130 28194 6142
rect 28142 6066 28194 6078
rect 5966 6018 6018 6030
rect 5966 5954 6018 5966
rect 9774 6018 9826 6030
rect 9774 5954 9826 5966
rect 9886 6018 9938 6030
rect 9886 5954 9938 5966
rect 10334 6018 10386 6030
rect 10334 5954 10386 5966
rect 10782 6018 10834 6030
rect 10782 5954 10834 5966
rect 11342 6018 11394 6030
rect 11342 5954 11394 5966
rect 15486 6018 15538 6030
rect 15486 5954 15538 5966
rect 20414 6018 20466 6030
rect 20414 5954 20466 5966
rect 20526 6018 20578 6030
rect 20526 5954 20578 5966
rect 25230 6018 25282 6030
rect 25230 5954 25282 5966
rect 27918 6018 27970 6030
rect 29810 5966 29822 6018
rect 29874 5966 29886 6018
rect 27918 5954 27970 5966
rect 5630 5906 5682 5918
rect 9550 5906 9602 5918
rect 8754 5854 8766 5906
rect 8818 5854 8830 5906
rect 5630 5842 5682 5854
rect 9550 5842 9602 5854
rect 10110 5906 10162 5918
rect 10110 5842 10162 5854
rect 10446 5906 10498 5918
rect 10446 5842 10498 5854
rect 11006 5906 11058 5918
rect 15150 5906 15202 5918
rect 11778 5854 11790 5906
rect 11842 5854 11854 5906
rect 11006 5842 11058 5854
rect 15150 5842 15202 5854
rect 15374 5906 15426 5918
rect 15374 5842 15426 5854
rect 15710 5906 15762 5918
rect 15710 5842 15762 5854
rect 15822 5906 15874 5918
rect 15822 5842 15874 5854
rect 16158 5906 16210 5918
rect 16158 5842 16210 5854
rect 16494 5906 16546 5918
rect 24110 5906 24162 5918
rect 17378 5854 17390 5906
rect 17442 5854 17454 5906
rect 20850 5854 20862 5906
rect 20914 5854 20926 5906
rect 16494 5842 16546 5854
rect 24110 5842 24162 5854
rect 25454 5906 25506 5918
rect 25454 5842 25506 5854
rect 25678 5906 25730 5918
rect 26462 5906 26514 5918
rect 26114 5854 26126 5906
rect 26178 5854 26190 5906
rect 25678 5842 25730 5854
rect 26462 5842 26514 5854
rect 27246 5906 27298 5918
rect 27246 5842 27298 5854
rect 27694 5906 27746 5918
rect 28466 5854 28478 5906
rect 28530 5854 28542 5906
rect 29026 5854 29038 5906
rect 29090 5854 29102 5906
rect 27694 5842 27746 5854
rect 10894 5794 10946 5806
rect 16046 5794 16098 5806
rect 25342 5794 25394 5806
rect 12450 5742 12462 5794
rect 12514 5742 12526 5794
rect 14578 5742 14590 5794
rect 14642 5742 14654 5794
rect 19058 5742 19070 5794
rect 19122 5742 19134 5794
rect 10894 5730 10946 5742
rect 16046 5730 16098 5742
rect 25342 5730 25394 5742
rect 26574 5794 26626 5806
rect 26574 5730 26626 5742
rect 27134 5794 27186 5806
rect 27134 5730 27186 5742
rect 28030 5794 28082 5806
rect 31938 5742 31950 5794
rect 32002 5742 32014 5794
rect 28030 5730 28082 5742
rect 6638 5682 6690 5694
rect 6638 5618 6690 5630
rect 21870 5682 21922 5694
rect 21870 5618 21922 5630
rect 1344 5514 35616 5548
rect 1344 5462 5498 5514
rect 5550 5462 5602 5514
rect 5654 5462 5706 5514
rect 5758 5462 14066 5514
rect 14118 5462 14170 5514
rect 14222 5462 14274 5514
rect 14326 5462 22634 5514
rect 22686 5462 22738 5514
rect 22790 5462 22842 5514
rect 22894 5462 31202 5514
rect 31254 5462 31306 5514
rect 31358 5462 31410 5514
rect 31462 5462 35616 5514
rect 1344 5428 35616 5462
rect 28030 5346 28082 5358
rect 28030 5282 28082 5294
rect 29262 5346 29314 5358
rect 29262 5282 29314 5294
rect 2270 5234 2322 5246
rect 13582 5234 13634 5246
rect 25454 5234 25506 5246
rect 6850 5182 6862 5234
rect 6914 5182 6926 5234
rect 8978 5182 8990 5234
rect 9042 5182 9054 5234
rect 10658 5182 10670 5234
rect 10722 5182 10734 5234
rect 12786 5182 12798 5234
rect 12850 5182 12862 5234
rect 14578 5182 14590 5234
rect 14642 5182 14654 5234
rect 18610 5182 18622 5234
rect 18674 5182 18686 5234
rect 20738 5182 20750 5234
rect 20802 5182 20814 5234
rect 22530 5182 22542 5234
rect 22594 5182 22606 5234
rect 24658 5182 24670 5234
rect 24722 5182 24734 5234
rect 2270 5170 2322 5182
rect 13582 5170 13634 5182
rect 25454 5170 25506 5182
rect 26350 5234 26402 5246
rect 26350 5170 26402 5182
rect 28590 5234 28642 5246
rect 28590 5170 28642 5182
rect 13470 5122 13522 5134
rect 4610 5070 4622 5122
rect 4674 5070 4686 5122
rect 6066 5070 6078 5122
rect 6130 5070 6142 5122
rect 9874 5070 9886 5122
rect 9938 5070 9950 5122
rect 13470 5058 13522 5070
rect 13806 5122 13858 5134
rect 13806 5058 13858 5070
rect 14030 5122 14082 5134
rect 24894 5122 24946 5134
rect 17490 5070 17502 5122
rect 17554 5070 17566 5122
rect 17938 5070 17950 5122
rect 18002 5070 18014 5122
rect 21746 5070 21758 5122
rect 21810 5070 21822 5122
rect 14030 5058 14082 5070
rect 24894 5058 24946 5070
rect 25790 5122 25842 5134
rect 25790 5058 25842 5070
rect 27134 5122 27186 5134
rect 27134 5058 27186 5070
rect 27470 5122 27522 5134
rect 27470 5058 27522 5070
rect 27694 5122 27746 5134
rect 27694 5058 27746 5070
rect 34638 5122 34690 5134
rect 34638 5058 34690 5070
rect 35198 5122 35250 5134
rect 35198 5058 35250 5070
rect 9326 5010 9378 5022
rect 9326 4946 9378 4958
rect 9438 5010 9490 5022
rect 25342 5010 25394 5022
rect 16706 4958 16718 5010
rect 16770 4958 16782 5010
rect 9438 4946 9490 4958
rect 25342 4946 25394 4958
rect 25566 5010 25618 5022
rect 25566 4946 25618 4958
rect 26462 5010 26514 5022
rect 26462 4946 26514 4958
rect 28142 5010 28194 5022
rect 28142 4946 28194 4958
rect 29374 5010 29426 5022
rect 29374 4946 29426 4958
rect 34862 5010 34914 5022
rect 34862 4946 34914 4958
rect 9662 4898 9714 4910
rect 9662 4834 9714 4846
rect 26238 4898 26290 4910
rect 26238 4834 26290 4846
rect 27358 4898 27410 4910
rect 27358 4834 27410 4846
rect 29822 4898 29874 4910
rect 29822 4834 29874 4846
rect 1344 4730 35776 4764
rect 1344 4678 9782 4730
rect 9834 4678 9886 4730
rect 9938 4678 9990 4730
rect 10042 4678 18350 4730
rect 18402 4678 18454 4730
rect 18506 4678 18558 4730
rect 18610 4678 26918 4730
rect 26970 4678 27022 4730
rect 27074 4678 27126 4730
rect 27178 4678 35486 4730
rect 35538 4678 35590 4730
rect 35642 4678 35694 4730
rect 35746 4678 35776 4730
rect 1344 4644 35776 4678
rect 17502 4562 17554 4574
rect 17502 4498 17554 4510
rect 18622 4562 18674 4574
rect 18622 4498 18674 4510
rect 18958 4562 19010 4574
rect 18958 4498 19010 4510
rect 23214 4562 23266 4574
rect 23214 4498 23266 4510
rect 24110 4562 24162 4574
rect 24110 4498 24162 4510
rect 24558 4562 24610 4574
rect 24558 4498 24610 4510
rect 31726 4562 31778 4574
rect 31726 4498 31778 4510
rect 32174 4562 32226 4574
rect 32174 4498 32226 4510
rect 13358 4450 13410 4462
rect 17950 4450 18002 4462
rect 6626 4398 6638 4450
rect 6690 4398 6702 4450
rect 16034 4398 16046 4450
rect 16098 4398 16110 4450
rect 13358 4386 13410 4398
rect 17950 4386 18002 4398
rect 18286 4450 18338 4462
rect 18286 4386 18338 4398
rect 18398 4450 18450 4462
rect 22654 4450 22706 4462
rect 20066 4398 20078 4450
rect 20130 4398 20142 4450
rect 18398 4386 18450 4398
rect 22654 4386 22706 4398
rect 22766 4450 22818 4462
rect 26002 4398 26014 4450
rect 26066 4398 26078 4450
rect 30594 4398 30606 4450
rect 30658 4398 30670 4450
rect 22766 4386 22818 4398
rect 12686 4338 12738 4350
rect 5282 4286 5294 4338
rect 5346 4286 5358 4338
rect 5954 4286 5966 4338
rect 6018 4286 6030 4338
rect 12450 4286 12462 4338
rect 12514 4286 12526 4338
rect 12686 4274 12738 4286
rect 13022 4338 13074 4350
rect 17278 4338 17330 4350
rect 16818 4286 16830 4338
rect 16882 4286 16894 4338
rect 13022 4274 13074 4286
rect 17278 4274 17330 4286
rect 17614 4338 17666 4350
rect 19282 4286 19294 4338
rect 19346 4286 19358 4338
rect 25330 4286 25342 4338
rect 25394 4286 25406 4338
rect 31266 4286 31278 4338
rect 31330 4286 31342 4338
rect 17614 4274 17666 4286
rect 12910 4226 12962 4238
rect 23774 4226 23826 4238
rect 3378 4174 3390 4226
rect 3442 4174 3454 4226
rect 8754 4174 8766 4226
rect 8818 4174 8830 4226
rect 9538 4174 9550 4226
rect 9602 4174 9614 4226
rect 11666 4174 11678 4226
rect 11730 4174 11742 4226
rect 13906 4174 13918 4226
rect 13970 4174 13982 4226
rect 22194 4174 22206 4226
rect 22258 4174 22270 4226
rect 12910 4162 12962 4174
rect 23774 4162 23826 4174
rect 24222 4226 24274 4238
rect 24222 4162 24274 4174
rect 24670 4226 24722 4238
rect 31838 4226 31890 4238
rect 28130 4174 28142 4226
rect 28194 4174 28206 4226
rect 28466 4174 28478 4226
rect 28530 4174 28542 4226
rect 24670 4162 24722 4174
rect 31838 4162 31890 4174
rect 32286 4226 32338 4238
rect 32286 4162 32338 4174
rect 33294 4226 33346 4238
rect 33294 4162 33346 4174
rect 22654 4114 22706 4126
rect 22654 4050 22706 4062
rect 1344 3946 35616 3980
rect 1344 3894 5498 3946
rect 5550 3894 5602 3946
rect 5654 3894 5706 3946
rect 5758 3894 14066 3946
rect 14118 3894 14170 3946
rect 14222 3894 14274 3946
rect 14326 3894 22634 3946
rect 22686 3894 22738 3946
rect 22790 3894 22842 3946
rect 22894 3894 31202 3946
rect 31254 3894 31306 3946
rect 31358 3894 31410 3946
rect 31462 3894 35616 3946
rect 1344 3860 35616 3894
rect 12350 3666 12402 3678
rect 18622 3666 18674 3678
rect 25566 3666 25618 3678
rect 15922 3614 15934 3666
rect 15986 3614 15998 3666
rect 21858 3614 21870 3666
rect 21922 3614 21934 3666
rect 12350 3602 12402 3614
rect 18622 3602 18674 3614
rect 25566 3602 25618 3614
rect 5630 3554 5682 3566
rect 4498 3502 4510 3554
rect 4562 3502 4574 3554
rect 5630 3490 5682 3502
rect 5966 3554 6018 3566
rect 9214 3554 9266 3566
rect 8754 3502 8766 3554
rect 8818 3502 8830 3554
rect 5966 3490 6018 3502
rect 9214 3490 9266 3502
rect 9550 3554 9602 3566
rect 13246 3554 13298 3566
rect 10434 3502 10446 3554
rect 10498 3502 10510 3554
rect 9550 3490 9602 3502
rect 13246 3490 13298 3502
rect 13582 3554 13634 3566
rect 17054 3554 17106 3566
rect 14242 3502 14254 3554
rect 14306 3502 14318 3554
rect 13582 3490 13634 3502
rect 17054 3490 17106 3502
rect 17390 3554 17442 3566
rect 28702 3554 28754 3566
rect 17602 3502 17614 3554
rect 17666 3502 17678 3554
rect 20738 3502 20750 3554
rect 20802 3502 20814 3554
rect 23762 3502 23774 3554
rect 23826 3502 23838 3554
rect 24770 3502 24782 3554
rect 24834 3502 24846 3554
rect 17390 3490 17442 3502
rect 28702 3490 28754 3502
rect 29374 3554 29426 3566
rect 29374 3490 29426 3502
rect 31054 3554 31106 3566
rect 32958 3554 33010 3566
rect 32386 3502 32398 3554
rect 32450 3502 32462 3554
rect 33618 3502 33630 3554
rect 33682 3502 33694 3554
rect 35074 3502 35086 3554
rect 35138 3502 35150 3554
rect 31054 3490 31106 3502
rect 32958 3490 33010 3502
rect 5742 3442 5794 3454
rect 5742 3378 5794 3390
rect 9438 3442 9490 3454
rect 9438 3378 9490 3390
rect 13358 3442 13410 3454
rect 13358 3378 13410 3390
rect 17166 3442 17218 3454
rect 17166 3378 17218 3390
rect 23998 3442 24050 3454
rect 23998 3378 24050 3390
rect 27470 3442 27522 3454
rect 27470 3378 27522 3390
rect 27806 3442 27858 3454
rect 27806 3378 27858 3390
rect 28366 3442 28418 3454
rect 28366 3378 28418 3390
rect 29038 3442 29090 3454
rect 29038 3378 29090 3390
rect 29822 3442 29874 3454
rect 29822 3378 29874 3390
rect 30270 3442 30322 3454
rect 30270 3378 30322 3390
rect 30606 3442 30658 3454
rect 30606 3378 30658 3390
rect 31502 3442 31554 3454
rect 31502 3378 31554 3390
rect 32174 3442 32226 3454
rect 32174 3378 32226 3390
rect 34638 3442 34690 3454
rect 34638 3378 34690 3390
rect 3950 3330 4002 3342
rect 3950 3266 4002 3278
rect 7758 3330 7810 3342
rect 7758 3266 7810 3278
rect 33406 3330 33458 3342
rect 33406 3266 33458 3278
rect 34862 3330 34914 3342
rect 34862 3266 34914 3278
rect 1344 3162 35776 3196
rect 1344 3110 9782 3162
rect 9834 3110 9886 3162
rect 9938 3110 9990 3162
rect 10042 3110 18350 3162
rect 18402 3110 18454 3162
rect 18506 3110 18558 3162
rect 18610 3110 26918 3162
rect 26970 3110 27022 3162
rect 27074 3110 27126 3162
rect 27178 3110 35486 3162
rect 35538 3110 35590 3162
rect 35642 3110 35694 3162
rect 35746 3110 35776 3162
rect 1344 3076 35776 3110
<< via1 >>
rect 5498 33686 5550 33738
rect 5602 33686 5654 33738
rect 5706 33686 5758 33738
rect 14066 33686 14118 33738
rect 14170 33686 14222 33738
rect 14274 33686 14326 33738
rect 22634 33686 22686 33738
rect 22738 33686 22790 33738
rect 22842 33686 22894 33738
rect 31202 33686 31254 33738
rect 31306 33686 31358 33738
rect 31410 33686 31462 33738
rect 12350 33518 12402 33570
rect 25566 33518 25618 33570
rect 30046 33518 30098 33570
rect 8206 33406 8258 33458
rect 16046 33406 16098 33458
rect 19854 33406 19906 33458
rect 23774 33406 23826 33458
rect 35086 33406 35138 33458
rect 6414 33294 6466 33346
rect 9998 33294 10050 33346
rect 13246 33294 13298 33346
rect 17054 33294 17106 33346
rect 20974 33294 21026 33346
rect 24782 33294 24834 33346
rect 29038 33294 29090 33346
rect 32174 33294 32226 33346
rect 1822 33182 1874 33234
rect 2942 33182 2994 33234
rect 4062 33182 4114 33234
rect 4958 33182 5010 33234
rect 5854 33182 5906 33234
rect 9550 33182 9602 33234
rect 13918 33182 13970 33234
rect 17726 33182 17778 33234
rect 21646 33182 21698 33234
rect 32958 33182 33010 33234
rect 27582 33070 27634 33122
rect 28702 33070 28754 33122
rect 9782 32902 9834 32954
rect 9886 32902 9938 32954
rect 9990 32902 10042 32954
rect 18350 32902 18402 32954
rect 18454 32902 18506 32954
rect 18558 32902 18610 32954
rect 26918 32902 26970 32954
rect 27022 32902 27074 32954
rect 27126 32902 27178 32954
rect 35486 32902 35538 32954
rect 35590 32902 35642 32954
rect 35694 32902 35746 32954
rect 9550 32734 9602 32786
rect 15822 32734 15874 32786
rect 18622 32734 18674 32786
rect 33742 32734 33794 32786
rect 16158 32622 16210 32674
rect 16830 32622 16882 32674
rect 31726 32622 31778 32674
rect 34862 32622 34914 32674
rect 35198 32622 35250 32674
rect 6190 32510 6242 32562
rect 12462 32510 12514 32562
rect 16494 32510 16546 32562
rect 17614 32510 17666 32562
rect 20526 32510 20578 32562
rect 24110 32510 24162 32562
rect 24558 32510 24610 32562
rect 25230 32510 25282 32562
rect 28478 32510 28530 32562
rect 31838 32510 31890 32562
rect 6862 32398 6914 32450
rect 8990 32398 9042 32450
rect 10222 32398 10274 32450
rect 13134 32398 13186 32450
rect 15374 32398 15426 32450
rect 21310 32398 21362 32450
rect 23438 32398 23490 32450
rect 26238 32398 26290 32450
rect 29150 32398 29202 32450
rect 31278 32398 31330 32450
rect 34190 32398 34242 32450
rect 34638 32398 34690 32450
rect 31726 32286 31778 32338
rect 33630 32286 33682 32338
rect 34526 32286 34578 32338
rect 5498 32118 5550 32170
rect 5602 32118 5654 32170
rect 5706 32118 5758 32170
rect 14066 32118 14118 32170
rect 14170 32118 14222 32170
rect 14274 32118 14326 32170
rect 22634 32118 22686 32170
rect 22738 32118 22790 32170
rect 22842 32118 22894 32170
rect 31202 32118 31254 32170
rect 31306 32118 31358 32170
rect 31410 32118 31462 32170
rect 8094 31950 8146 32002
rect 11454 31838 11506 31890
rect 11902 31838 11954 31890
rect 16046 31838 16098 31890
rect 18286 31838 18338 31890
rect 20414 31838 20466 31890
rect 22430 31838 22482 31890
rect 27358 31838 27410 31890
rect 28030 31838 28082 31890
rect 32062 31838 32114 31890
rect 8654 31726 8706 31778
rect 14590 31726 14642 31778
rect 17502 31726 17554 31778
rect 21422 31726 21474 31778
rect 21758 31726 21810 31778
rect 22654 31726 22706 31778
rect 23326 31726 23378 31778
rect 26910 31726 26962 31778
rect 27806 31726 27858 31778
rect 29262 31726 29314 31778
rect 32398 31726 32450 31778
rect 7422 31614 7474 31666
rect 8206 31614 8258 31666
rect 9326 31614 9378 31666
rect 22094 31614 22146 31666
rect 24110 31614 24162 31666
rect 28142 31614 28194 31666
rect 28254 31614 28306 31666
rect 29934 31614 29986 31666
rect 13806 31502 13858 31554
rect 14254 31502 14306 31554
rect 21758 31502 21810 31554
rect 22990 31502 23042 31554
rect 26350 31502 26402 31554
rect 26798 31502 26850 31554
rect 28030 31502 28082 31554
rect 33406 31502 33458 31554
rect 9782 31334 9834 31386
rect 9886 31334 9938 31386
rect 9990 31334 10042 31386
rect 18350 31334 18402 31386
rect 18454 31334 18506 31386
rect 18558 31334 18610 31386
rect 26918 31334 26970 31386
rect 27022 31334 27074 31386
rect 27126 31334 27178 31386
rect 35486 31334 35538 31386
rect 35590 31334 35642 31386
rect 35694 31334 35746 31386
rect 8430 31166 8482 31218
rect 9550 31166 9602 31218
rect 15374 31166 15426 31218
rect 20750 31166 20802 31218
rect 25342 31166 25394 31218
rect 30830 31166 30882 31218
rect 33518 31166 33570 31218
rect 33630 31166 33682 31218
rect 7646 31054 7698 31106
rect 10222 31054 10274 31106
rect 11342 31054 11394 31106
rect 16270 31054 16322 31106
rect 16718 31054 16770 31106
rect 17614 31054 17666 31106
rect 18734 31054 18786 31106
rect 19070 31054 19122 31106
rect 23550 31054 23602 31106
rect 25454 31054 25506 31106
rect 31726 31054 31778 31106
rect 31838 31054 31890 31106
rect 32398 31054 32450 31106
rect 33966 31054 34018 31106
rect 4398 30942 4450 30994
rect 7982 30942 8034 30994
rect 10110 30942 10162 30994
rect 10446 30942 10498 30994
rect 10670 30942 10722 30994
rect 11566 30942 11618 30994
rect 12126 30942 12178 30994
rect 15598 30942 15650 30994
rect 16046 30942 16098 30994
rect 16382 30942 16434 30994
rect 17390 30942 17442 30994
rect 17726 30942 17778 30994
rect 17950 30942 18002 30994
rect 18398 30942 18450 30994
rect 19406 30942 19458 30994
rect 19854 30942 19906 30994
rect 22766 30942 22818 30994
rect 23438 30942 23490 30994
rect 24558 30942 24610 30994
rect 27470 30942 27522 30994
rect 30606 30942 30658 30994
rect 31054 30942 31106 30994
rect 31390 30942 31442 30994
rect 32062 30942 32114 30994
rect 32510 30942 32562 30994
rect 32958 30942 33010 30994
rect 33406 30942 33458 30994
rect 34302 30942 34354 30994
rect 34638 30942 34690 30994
rect 35198 30942 35250 30994
rect 5182 30830 5234 30882
rect 7310 30830 7362 30882
rect 9662 30830 9714 30882
rect 12798 30830 12850 30882
rect 14926 30830 14978 30882
rect 22654 30830 22706 30882
rect 23550 30830 23602 30882
rect 25902 30830 25954 30882
rect 28142 30830 28194 30882
rect 30270 30830 30322 30882
rect 30830 30830 30882 30882
rect 34750 30830 34802 30882
rect 11118 30718 11170 30770
rect 16830 30718 16882 30770
rect 18622 30718 18674 30770
rect 25342 30718 25394 30770
rect 32398 30718 32450 30770
rect 5498 30550 5550 30602
rect 5602 30550 5654 30602
rect 5706 30550 5758 30602
rect 14066 30550 14118 30602
rect 14170 30550 14222 30602
rect 14274 30550 14326 30602
rect 22634 30550 22686 30602
rect 22738 30550 22790 30602
rect 22842 30550 22894 30602
rect 31202 30550 31254 30602
rect 31306 30550 31358 30602
rect 31410 30550 31462 30602
rect 11790 30382 11842 30434
rect 15598 30382 15650 30434
rect 20750 30382 20802 30434
rect 21758 30382 21810 30434
rect 33630 30382 33682 30434
rect 34302 30382 34354 30434
rect 9214 30270 9266 30322
rect 18846 30270 18898 30322
rect 20414 30270 20466 30322
rect 27694 30270 27746 30322
rect 32510 30270 32562 30322
rect 6414 30158 6466 30210
rect 7086 30158 7138 30210
rect 9326 30158 9378 30210
rect 9550 30158 9602 30210
rect 10446 30158 10498 30210
rect 13582 30158 13634 30210
rect 14590 30158 14642 30210
rect 17502 30158 17554 30210
rect 20750 30158 20802 30210
rect 21870 30158 21922 30210
rect 23326 30158 23378 30210
rect 24222 30158 24274 30210
rect 28590 30158 28642 30210
rect 29262 30158 29314 30210
rect 29710 30158 29762 30210
rect 30382 30158 30434 30210
rect 5742 30046 5794 30098
rect 8206 30046 8258 30098
rect 9774 30046 9826 30098
rect 13470 30046 13522 30098
rect 21310 30046 21362 30098
rect 21534 30046 21586 30098
rect 23102 30046 23154 30098
rect 23662 30046 23714 30098
rect 24894 30046 24946 30098
rect 34862 30046 34914 30098
rect 5630 29934 5682 29986
rect 6526 29934 6578 29986
rect 6750 29934 6802 29986
rect 7310 29934 7362 29986
rect 7870 29934 7922 29986
rect 8990 29934 9042 29986
rect 9998 29934 10050 29986
rect 14254 29934 14306 29986
rect 21758 29934 21810 29986
rect 22654 29934 22706 29986
rect 23214 29934 23266 29986
rect 27134 29934 27186 29986
rect 33182 29934 33234 29986
rect 33630 29934 33682 29986
rect 34078 29934 34130 29986
rect 34638 29934 34690 29986
rect 35198 29934 35250 29986
rect 9782 29766 9834 29818
rect 9886 29766 9938 29818
rect 9990 29766 10042 29818
rect 18350 29766 18402 29818
rect 18454 29766 18506 29818
rect 18558 29766 18610 29818
rect 26918 29766 26970 29818
rect 27022 29766 27074 29818
rect 27126 29766 27178 29818
rect 35486 29766 35538 29818
rect 35590 29766 35642 29818
rect 35694 29766 35746 29818
rect 8878 29598 8930 29650
rect 10110 29598 10162 29650
rect 10334 29598 10386 29650
rect 12574 29598 12626 29650
rect 14030 29598 14082 29650
rect 16382 29598 16434 29650
rect 17838 29598 17890 29650
rect 19070 29598 19122 29650
rect 24110 29598 24162 29650
rect 26238 29598 26290 29650
rect 34190 29598 34242 29650
rect 34414 29598 34466 29650
rect 4622 29486 4674 29538
rect 8430 29486 8482 29538
rect 11454 29486 11506 29538
rect 12238 29486 12290 29538
rect 18286 29486 18338 29538
rect 18846 29486 18898 29538
rect 20190 29486 20242 29538
rect 21198 29486 21250 29538
rect 34526 29486 34578 29538
rect 34862 29486 34914 29538
rect 3950 29374 4002 29426
rect 7198 29374 7250 29426
rect 7646 29374 7698 29426
rect 8654 29374 8706 29426
rect 9550 29374 9602 29426
rect 9886 29374 9938 29426
rect 11230 29374 11282 29426
rect 11342 29374 11394 29426
rect 13022 29374 13074 29426
rect 16158 29374 16210 29426
rect 16270 29374 16322 29426
rect 16830 29374 16882 29426
rect 17278 29374 17330 29426
rect 17614 29374 17666 29426
rect 18622 29374 18674 29426
rect 20638 29374 20690 29426
rect 22766 29374 22818 29426
rect 25230 29374 25282 29426
rect 29262 29374 29314 29426
rect 33742 29374 33794 29426
rect 35086 29374 35138 29426
rect 6750 29262 6802 29314
rect 8094 29262 8146 29314
rect 9998 29262 10050 29314
rect 10894 29262 10946 29314
rect 16606 29262 16658 29314
rect 18062 29262 18114 29314
rect 18734 29262 18786 29314
rect 23214 29262 23266 29314
rect 23774 29262 23826 29314
rect 28926 29262 28978 29314
rect 29934 29262 29986 29314
rect 32062 29262 32114 29314
rect 32510 29262 32562 29314
rect 33854 29262 33906 29314
rect 8990 29150 9042 29202
rect 11902 29150 11954 29202
rect 17838 29150 17890 29202
rect 20862 29150 20914 29202
rect 33294 29150 33346 29202
rect 5498 28982 5550 29034
rect 5602 28982 5654 29034
rect 5706 28982 5758 29034
rect 14066 28982 14118 29034
rect 14170 28982 14222 29034
rect 14274 28982 14326 29034
rect 22634 28982 22686 29034
rect 22738 28982 22790 29034
rect 22842 28982 22894 29034
rect 31202 28982 31254 29034
rect 31306 28982 31358 29034
rect 31410 28982 31462 29034
rect 6862 28814 6914 28866
rect 7198 28814 7250 28866
rect 15598 28814 15650 28866
rect 16494 28814 16546 28866
rect 21870 28814 21922 28866
rect 6526 28702 6578 28754
rect 7646 28702 7698 28754
rect 9102 28702 9154 28754
rect 9886 28702 9938 28754
rect 11006 28702 11058 28754
rect 11566 28702 11618 28754
rect 12798 28702 12850 28754
rect 13582 28702 13634 28754
rect 15374 28702 15426 28754
rect 15934 28702 15986 28754
rect 17726 28702 17778 28754
rect 19406 28702 19458 28754
rect 25902 28702 25954 28754
rect 28478 28702 28530 28754
rect 32174 28702 32226 28754
rect 6862 28590 6914 28642
rect 8318 28590 8370 28642
rect 8990 28590 9042 28642
rect 9438 28590 9490 28642
rect 10222 28590 10274 28642
rect 10782 28590 10834 28642
rect 11230 28590 11282 28642
rect 14254 28590 14306 28642
rect 15038 28590 15090 28642
rect 17054 28590 17106 28642
rect 17166 28590 17218 28642
rect 17502 28590 17554 28642
rect 17838 28590 17890 28642
rect 18062 28590 18114 28642
rect 18958 28590 19010 28642
rect 19518 28590 19570 28642
rect 20078 28590 20130 28642
rect 20190 28590 20242 28642
rect 20526 28590 20578 28642
rect 21534 28590 21586 28642
rect 21982 28590 22034 28642
rect 23774 28590 23826 28642
rect 29150 28590 29202 28642
rect 34974 28590 35026 28642
rect 8654 28478 8706 28530
rect 9886 28478 9938 28530
rect 9998 28478 10050 28530
rect 10558 28478 10610 28530
rect 12686 28478 12738 28530
rect 12910 28478 12962 28530
rect 13806 28478 13858 28530
rect 16942 28478 16994 28530
rect 19854 28478 19906 28530
rect 21310 28478 21362 28530
rect 8542 28366 8594 28418
rect 13470 28366 13522 28418
rect 13694 28366 13746 28418
rect 14702 28366 14754 28418
rect 19070 28366 19122 28418
rect 19294 28366 19346 28418
rect 20302 28366 20354 28418
rect 22094 28366 22146 28418
rect 28366 28366 28418 28418
rect 34750 28366 34802 28418
rect 9782 28198 9834 28250
rect 9886 28198 9938 28250
rect 9990 28198 10042 28250
rect 18350 28198 18402 28250
rect 18454 28198 18506 28250
rect 18558 28198 18610 28250
rect 26918 28198 26970 28250
rect 27022 28198 27074 28250
rect 27126 28198 27178 28250
rect 35486 28198 35538 28250
rect 35590 28198 35642 28250
rect 35694 28198 35746 28250
rect 7086 28030 7138 28082
rect 8542 28030 8594 28082
rect 10670 28030 10722 28082
rect 12686 28030 12738 28082
rect 13582 28030 13634 28082
rect 8094 27918 8146 27970
rect 9774 27918 9826 27970
rect 11902 27918 11954 27970
rect 12014 27918 12066 27970
rect 14254 27918 14306 27970
rect 14926 27918 14978 27970
rect 15038 27918 15090 27970
rect 15150 27918 15202 27970
rect 16046 27918 16098 27970
rect 16382 27918 16434 27970
rect 17390 27918 17442 27970
rect 17614 27918 17666 27970
rect 17726 27974 17778 28026
rect 19406 28030 19458 28082
rect 19742 28030 19794 28082
rect 21646 28030 21698 28082
rect 23102 28030 23154 28082
rect 30382 28030 30434 28082
rect 34750 28030 34802 28082
rect 18734 27918 18786 27970
rect 20078 27918 20130 27970
rect 21758 27918 21810 27970
rect 29262 27918 29314 27970
rect 32062 27918 32114 27970
rect 32174 27918 32226 27970
rect 33070 27918 33122 27970
rect 3614 27806 3666 27858
rect 6862 27806 6914 27858
rect 7422 27806 7474 27858
rect 7870 27806 7922 27858
rect 9550 27806 9602 27858
rect 9998 27806 10050 27858
rect 10334 27806 10386 27858
rect 10894 27806 10946 27858
rect 12462 27806 12514 27858
rect 13134 27806 13186 27858
rect 13358 27806 13410 27858
rect 13694 27806 13746 27858
rect 15374 27806 15426 27858
rect 15822 27806 15874 27858
rect 16270 27806 16322 27858
rect 18174 27806 18226 27858
rect 20414 27806 20466 27858
rect 20638 27806 20690 27858
rect 20974 27806 21026 27858
rect 21422 27806 21474 27858
rect 22318 27806 22370 27858
rect 25230 27806 25282 27858
rect 26238 27806 26290 27858
rect 29934 27806 29986 27858
rect 30494 27806 30546 27858
rect 31054 27806 31106 27858
rect 31614 27806 31666 27858
rect 32398 27806 32450 27858
rect 33406 27806 33458 27858
rect 34302 27806 34354 27858
rect 35086 27806 35138 27858
rect 4286 27694 4338 27746
rect 6414 27694 6466 27746
rect 6974 27694 7026 27746
rect 9886 27694 9938 27746
rect 13246 27694 13298 27746
rect 14590 27694 14642 27746
rect 16606 27694 16658 27746
rect 20526 27694 20578 27746
rect 21310 27694 21362 27746
rect 25566 27694 25618 27746
rect 25790 27694 25842 27746
rect 27134 27694 27186 27746
rect 31278 27694 31330 27746
rect 32062 27694 32114 27746
rect 33294 27694 33346 27746
rect 33966 27694 34018 27746
rect 12014 27582 12066 27634
rect 12798 27582 12850 27634
rect 18398 27582 18450 27634
rect 18846 27582 18898 27634
rect 18958 27582 19010 27634
rect 30718 27582 30770 27634
rect 5498 27414 5550 27466
rect 5602 27414 5654 27466
rect 5706 27414 5758 27466
rect 14066 27414 14118 27466
rect 14170 27414 14222 27466
rect 14274 27414 14326 27466
rect 22634 27414 22686 27466
rect 22738 27414 22790 27466
rect 22842 27414 22894 27466
rect 31202 27414 31254 27466
rect 31306 27414 31358 27466
rect 31410 27414 31462 27466
rect 5630 27246 5682 27298
rect 5966 27246 6018 27298
rect 9550 27246 9602 27298
rect 15486 27246 15538 27298
rect 19742 27246 19794 27298
rect 30606 27246 30658 27298
rect 7534 27134 7586 27186
rect 9886 27134 9938 27186
rect 13806 27134 13858 27186
rect 15374 27134 15426 27186
rect 16158 27134 16210 27186
rect 26574 27134 26626 27186
rect 27470 27134 27522 27186
rect 28030 27134 28082 27186
rect 35198 27134 35250 27186
rect 6302 27022 6354 27074
rect 6526 27022 6578 27074
rect 6974 27022 7026 27074
rect 7198 27022 7250 27074
rect 8542 27022 8594 27074
rect 8990 27022 9042 27074
rect 10110 27022 10162 27074
rect 10894 27022 10946 27074
rect 11006 27022 11058 27074
rect 11454 27022 11506 27074
rect 12238 27022 12290 27074
rect 12574 27022 12626 27074
rect 14030 27022 14082 27074
rect 14366 27022 14418 27074
rect 18174 27022 18226 27074
rect 18510 27022 18562 27074
rect 18622 27022 18674 27074
rect 18958 27022 19010 27074
rect 19630 27022 19682 27074
rect 20526 27022 20578 27074
rect 20750 27022 20802 27074
rect 21870 27022 21922 27074
rect 22206 27022 22258 27074
rect 22430 27022 22482 27074
rect 22654 27022 22706 27074
rect 23326 27022 23378 27074
rect 23774 27022 23826 27074
rect 28366 27022 28418 27074
rect 29150 27022 29202 27074
rect 32286 27022 32338 27074
rect 8430 26910 8482 26962
rect 11902 26910 11954 26962
rect 12910 26910 12962 26962
rect 13470 26910 13522 26962
rect 14590 26910 14642 26962
rect 14702 26910 14754 26962
rect 15262 26910 15314 26962
rect 16830 26910 16882 26962
rect 17166 26910 17218 26962
rect 18286 26910 18338 26962
rect 5742 26798 5794 26850
rect 6414 26798 6466 26850
rect 7422 26798 7474 26850
rect 7646 26798 7698 26850
rect 7758 26798 7810 26850
rect 8318 26798 8370 26850
rect 11230 26798 11282 26850
rect 13694 26798 13746 26850
rect 13918 26798 13970 26850
rect 17838 26854 17890 26906
rect 18846 26910 18898 26962
rect 19742 26910 19794 26962
rect 20190 26910 20242 26962
rect 21310 26910 21362 26962
rect 22542 26910 22594 26962
rect 24446 26910 24498 26962
rect 27022 26910 27074 26962
rect 33070 26910 33122 26962
rect 17502 26798 17554 26850
rect 20414 26798 20466 26850
rect 21422 26798 21474 26850
rect 21646 26798 21698 26850
rect 9782 26630 9834 26682
rect 9886 26630 9938 26682
rect 9990 26630 10042 26682
rect 18350 26630 18402 26682
rect 18454 26630 18506 26682
rect 18558 26630 18610 26682
rect 26918 26630 26970 26682
rect 27022 26630 27074 26682
rect 27126 26630 27178 26682
rect 35486 26630 35538 26682
rect 35590 26630 35642 26682
rect 35694 26630 35746 26682
rect 8430 26462 8482 26514
rect 9550 26462 9602 26514
rect 9662 26462 9714 26514
rect 9774 26462 9826 26514
rect 17390 26462 17442 26514
rect 18398 26462 18450 26514
rect 18734 26462 18786 26514
rect 20862 26462 20914 26514
rect 22542 26462 22594 26514
rect 22654 26462 22706 26514
rect 24670 26462 24722 26514
rect 25566 26462 25618 26514
rect 27582 26462 27634 26514
rect 33070 26462 33122 26514
rect 7422 26350 7474 26402
rect 7534 26350 7586 26402
rect 7646 26350 7698 26402
rect 7982 26350 8034 26402
rect 9886 26350 9938 26402
rect 12462 26350 12514 26402
rect 12686 26350 12738 26402
rect 13582 26350 13634 26402
rect 16494 26350 16546 26402
rect 19742 26350 19794 26402
rect 20078 26350 20130 26402
rect 23886 26350 23938 26402
rect 25678 26350 25730 26402
rect 29934 26350 29986 26402
rect 33966 26350 34018 26402
rect 34414 26350 34466 26402
rect 34526 26350 34578 26402
rect 34862 26350 34914 26402
rect 3614 26238 3666 26290
rect 7086 26238 7138 26290
rect 8318 26238 8370 26290
rect 8542 26238 8594 26290
rect 10334 26238 10386 26290
rect 11342 26238 11394 26290
rect 11566 26238 11618 26290
rect 12126 26238 12178 26290
rect 13358 26238 13410 26290
rect 13806 26238 13858 26290
rect 15262 26238 15314 26290
rect 16158 26238 16210 26290
rect 16718 26238 16770 26290
rect 17726 26238 17778 26290
rect 18174 26238 18226 26290
rect 19070 26238 19122 26290
rect 20414 26238 20466 26290
rect 20638 26238 20690 26290
rect 20862 26238 20914 26290
rect 20974 26238 21026 26290
rect 22766 26238 22818 26290
rect 23214 26238 23266 26290
rect 23326 26238 23378 26290
rect 23662 26238 23714 26290
rect 25342 26238 25394 26290
rect 28142 26238 28194 26290
rect 31502 26238 31554 26290
rect 33742 26238 33794 26290
rect 34302 26238 34354 26290
rect 34750 26238 34802 26290
rect 4398 26126 4450 26178
rect 6526 26126 6578 26178
rect 12686 26126 12738 26178
rect 13134 26126 13186 26178
rect 14702 26126 14754 26178
rect 15710 26126 15762 26178
rect 21758 26126 21810 26178
rect 31950 26126 32002 26178
rect 32286 26126 32338 26178
rect 11790 26014 11842 26066
rect 11902 26014 11954 26066
rect 13918 26014 13970 26066
rect 21870 26014 21922 26066
rect 22094 26014 22146 26066
rect 22206 26014 22258 26066
rect 23550 26014 23602 26066
rect 33182 26014 33234 26066
rect 33406 26014 33458 26066
rect 5498 25846 5550 25898
rect 5602 25846 5654 25898
rect 5706 25846 5758 25898
rect 14066 25846 14118 25898
rect 14170 25846 14222 25898
rect 14274 25846 14326 25898
rect 22634 25846 22686 25898
rect 22738 25846 22790 25898
rect 22842 25846 22894 25898
rect 31202 25846 31254 25898
rect 31306 25846 31358 25898
rect 31410 25846 31462 25898
rect 6190 25678 6242 25730
rect 6526 25678 6578 25730
rect 6974 25678 7026 25730
rect 7422 25678 7474 25730
rect 10446 25678 10498 25730
rect 12238 25678 12290 25730
rect 13582 25678 13634 25730
rect 19630 25678 19682 25730
rect 21422 25678 21474 25730
rect 21534 25678 21586 25730
rect 28030 25678 28082 25730
rect 29598 25678 29650 25730
rect 30942 25678 30994 25730
rect 7422 25566 7474 25618
rect 17950 25566 18002 25618
rect 18734 25566 18786 25618
rect 19182 25566 19234 25618
rect 22430 25566 22482 25618
rect 26462 25566 26514 25618
rect 28254 25566 28306 25618
rect 33406 25566 33458 25618
rect 34974 25566 35026 25618
rect 7758 25454 7810 25506
rect 9886 25454 9938 25506
rect 10670 25454 10722 25506
rect 12126 25454 12178 25506
rect 12686 25454 12738 25506
rect 13022 25454 13074 25506
rect 13694 25454 13746 25506
rect 14590 25454 14642 25506
rect 14926 25454 14978 25506
rect 15262 25454 15314 25506
rect 17390 25454 17442 25506
rect 17614 25454 17666 25506
rect 18174 25454 18226 25506
rect 19406 25454 19458 25506
rect 23438 25454 23490 25506
rect 27134 25454 27186 25506
rect 27806 25454 27858 25506
rect 29486 25454 29538 25506
rect 29934 25454 29986 25506
rect 33630 25454 33682 25506
rect 6302 25342 6354 25394
rect 7982 25342 8034 25394
rect 8094 25342 8146 25394
rect 10110 25342 10162 25394
rect 18846 25342 18898 25394
rect 20414 25342 20466 25394
rect 21758 25342 21810 25394
rect 22094 25342 22146 25394
rect 22318 25342 22370 25394
rect 24222 25342 24274 25394
rect 27358 25342 27410 25394
rect 28366 25342 28418 25394
rect 28590 25342 28642 25394
rect 32846 25342 32898 25394
rect 33070 25342 33122 25394
rect 33182 25342 33234 25394
rect 6974 25230 7026 25282
rect 10222 25230 10274 25282
rect 12238 25230 12290 25282
rect 12798 25230 12850 25282
rect 13582 25230 13634 25282
rect 14254 25230 14306 25282
rect 15038 25230 15090 25282
rect 17054 25230 17106 25282
rect 18622 25230 18674 25282
rect 20078 25230 20130 25282
rect 20750 25230 20802 25282
rect 23102 25230 23154 25282
rect 29374 25230 29426 25282
rect 34190 25230 34242 25282
rect 34526 25230 34578 25282
rect 9782 25062 9834 25114
rect 9886 25062 9938 25114
rect 9990 25062 10042 25114
rect 18350 25062 18402 25114
rect 18454 25062 18506 25114
rect 18558 25062 18610 25114
rect 26918 25062 26970 25114
rect 27022 25062 27074 25114
rect 27126 25062 27178 25114
rect 35486 25062 35538 25114
rect 35590 25062 35642 25114
rect 35694 25062 35746 25114
rect 6974 24894 7026 24946
rect 7534 24894 7586 24946
rect 8094 24894 8146 24946
rect 8654 24894 8706 24946
rect 12574 24894 12626 24946
rect 12798 24894 12850 24946
rect 15262 24894 15314 24946
rect 17390 24894 17442 24946
rect 19630 24894 19682 24946
rect 19742 24894 19794 24946
rect 20078 24894 20130 24946
rect 22990 24894 23042 24946
rect 33070 24894 33122 24946
rect 34302 24894 34354 24946
rect 6750 24782 6802 24834
rect 7310 24782 7362 24834
rect 7870 24782 7922 24834
rect 8430 24782 8482 24834
rect 9550 24782 9602 24834
rect 10446 24782 10498 24834
rect 11566 24782 11618 24834
rect 12238 24782 12290 24834
rect 12350 24782 12402 24834
rect 14814 24782 14866 24834
rect 14926 24782 14978 24834
rect 15486 24782 15538 24834
rect 22878 24782 22930 24834
rect 26014 24782 26066 24834
rect 29374 24782 29426 24834
rect 34526 24782 34578 24834
rect 6638 24670 6690 24722
rect 7198 24670 7250 24722
rect 7758 24670 7810 24722
rect 8318 24670 8370 24722
rect 9886 24670 9938 24722
rect 10334 24670 10386 24722
rect 10670 24670 10722 24722
rect 11342 24670 11394 24722
rect 11678 24670 11730 24722
rect 13134 24670 13186 24722
rect 13582 24670 13634 24722
rect 14030 24670 14082 24722
rect 15150 24670 15202 24722
rect 15598 24670 15650 24722
rect 16158 24670 16210 24722
rect 16718 24670 16770 24722
rect 17726 24670 17778 24722
rect 19854 24670 19906 24722
rect 21086 24670 21138 24722
rect 22654 24670 22706 24722
rect 23326 24670 23378 24722
rect 25230 24670 25282 24722
rect 29038 24670 29090 24722
rect 32062 24670 32114 24722
rect 33182 24670 33234 24722
rect 33742 24670 33794 24722
rect 34750 24670 34802 24722
rect 35086 24670 35138 24722
rect 9102 24558 9154 24610
rect 11118 24558 11170 24610
rect 14478 24558 14530 24610
rect 18174 24558 18226 24610
rect 21982 24558 22034 24610
rect 23774 24558 23826 24610
rect 24334 24558 24386 24610
rect 24782 24558 24834 24610
rect 28142 24558 28194 24610
rect 29374 24558 29426 24610
rect 30270 24558 30322 24610
rect 33406 24558 33458 24610
rect 34638 24558 34690 24610
rect 28814 24446 28866 24498
rect 29598 24446 29650 24498
rect 33966 24446 34018 24498
rect 5498 24278 5550 24330
rect 5602 24278 5654 24330
rect 5706 24278 5758 24330
rect 14066 24278 14118 24330
rect 14170 24278 14222 24330
rect 14274 24278 14326 24330
rect 22634 24278 22686 24330
rect 22738 24278 22790 24330
rect 22842 24278 22894 24330
rect 31202 24278 31254 24330
rect 31306 24278 31358 24330
rect 31410 24278 31462 24330
rect 23998 24110 24050 24162
rect 30830 24110 30882 24162
rect 25566 23998 25618 24050
rect 28478 23998 28530 24050
rect 33070 23998 33122 24050
rect 35198 23998 35250 24050
rect 12910 23886 12962 23938
rect 13582 23886 13634 23938
rect 21534 23886 21586 23938
rect 23550 23886 23602 23938
rect 23886 23886 23938 23938
rect 25454 23886 25506 23938
rect 27134 23886 27186 23938
rect 28590 23886 28642 23938
rect 29374 23886 29426 23938
rect 32398 23886 32450 23938
rect 7198 23774 7250 23826
rect 7310 23774 7362 23826
rect 7870 23774 7922 23826
rect 15710 23774 15762 23826
rect 18958 23774 19010 23826
rect 19182 23774 19234 23826
rect 19294 23774 19346 23826
rect 21310 23774 21362 23826
rect 21758 23774 21810 23826
rect 24334 23774 24386 23826
rect 25118 23774 25170 23826
rect 26126 23774 26178 23826
rect 26798 23774 26850 23826
rect 27470 23774 27522 23826
rect 28142 23774 28194 23826
rect 28254 23774 28306 23826
rect 6750 23662 6802 23714
rect 6974 23662 7026 23714
rect 19742 23662 19794 23714
rect 21870 23662 21922 23714
rect 22318 23662 22370 23714
rect 24446 23662 24498 23714
rect 24670 23662 24722 23714
rect 25790 23662 25842 23714
rect 26014 23662 26066 23714
rect 26462 23662 26514 23714
rect 28366 23662 28418 23714
rect 9782 23494 9834 23546
rect 9886 23494 9938 23546
rect 9990 23494 10042 23546
rect 18350 23494 18402 23546
rect 18454 23494 18506 23546
rect 18558 23494 18610 23546
rect 26918 23494 26970 23546
rect 27022 23494 27074 23546
rect 27126 23494 27178 23546
rect 35486 23494 35538 23546
rect 35590 23494 35642 23546
rect 35694 23494 35746 23546
rect 8206 23326 8258 23378
rect 9102 23326 9154 23378
rect 13806 23326 13858 23378
rect 14254 23326 14306 23378
rect 17726 23326 17778 23378
rect 18398 23326 18450 23378
rect 19406 23326 19458 23378
rect 24334 23326 24386 23378
rect 26350 23326 26402 23378
rect 27358 23326 27410 23378
rect 28926 23326 28978 23378
rect 30942 23326 30994 23378
rect 8094 23214 8146 23266
rect 8878 23214 8930 23266
rect 24558 23214 24610 23266
rect 25454 23214 25506 23266
rect 26574 23214 26626 23266
rect 28030 23214 28082 23266
rect 28254 23214 28306 23266
rect 28478 23214 28530 23266
rect 29038 23214 29090 23266
rect 33294 23214 33346 23266
rect 3950 23102 4002 23154
rect 7086 23102 7138 23154
rect 7534 23102 7586 23154
rect 7758 23102 7810 23154
rect 8430 23102 8482 23154
rect 8766 23102 8818 23154
rect 9438 23102 9490 23154
rect 9774 23102 9826 23154
rect 10110 23102 10162 23154
rect 10558 23102 10610 23154
rect 17502 23102 17554 23154
rect 17726 23102 17778 23154
rect 18062 23102 18114 23154
rect 18174 23102 18226 23154
rect 18510 23102 18562 23154
rect 19294 23102 19346 23154
rect 19966 23102 20018 23154
rect 23214 23102 23266 23154
rect 24670 23102 24722 23154
rect 25566 23102 25618 23154
rect 26126 23102 26178 23154
rect 26238 23102 26290 23154
rect 27022 23102 27074 23154
rect 28814 23102 28866 23154
rect 29262 23102 29314 23154
rect 29598 23102 29650 23154
rect 29934 23102 29986 23154
rect 33182 23102 33234 23154
rect 34190 23102 34242 23154
rect 4734 22990 4786 23042
rect 6862 22990 6914 23042
rect 7310 22990 7362 23042
rect 9662 22990 9714 23042
rect 11230 22990 11282 23042
rect 13358 22990 13410 23042
rect 20638 22990 20690 23042
rect 22766 22990 22818 23042
rect 23662 22990 23714 23042
rect 24110 22990 24162 23042
rect 33630 22990 33682 23042
rect 33966 22990 34018 23042
rect 35198 22990 35250 23042
rect 19406 22878 19458 22930
rect 25454 22878 25506 22930
rect 28366 22878 28418 22930
rect 35086 22878 35138 22930
rect 5498 22710 5550 22762
rect 5602 22710 5654 22762
rect 5706 22710 5758 22762
rect 14066 22710 14118 22762
rect 14170 22710 14222 22762
rect 14274 22710 14326 22762
rect 22634 22710 22686 22762
rect 22738 22710 22790 22762
rect 22842 22710 22894 22762
rect 31202 22710 31254 22762
rect 31306 22710 31358 22762
rect 31410 22710 31462 22762
rect 19406 22542 19458 22594
rect 26126 22542 26178 22594
rect 26350 22542 26402 22594
rect 34974 22542 35026 22594
rect 8206 22430 8258 22482
rect 10334 22430 10386 22482
rect 15710 22430 15762 22482
rect 16830 22430 16882 22482
rect 18958 22430 19010 22482
rect 25790 22430 25842 22482
rect 30718 22430 30770 22482
rect 7086 22318 7138 22370
rect 7534 22318 7586 22370
rect 10894 22318 10946 22370
rect 11342 22318 11394 22370
rect 16046 22318 16098 22370
rect 21534 22318 21586 22370
rect 21870 22318 21922 22370
rect 22878 22318 22930 22370
rect 27134 22318 27186 22370
rect 27470 22318 27522 22370
rect 27694 22318 27746 22370
rect 28142 22318 28194 22370
rect 29150 22318 29202 22370
rect 30606 22318 30658 22370
rect 31390 22318 31442 22370
rect 31614 22318 31666 22370
rect 31950 22318 32002 22370
rect 33070 22318 33122 22370
rect 6526 22206 6578 22258
rect 6862 22206 6914 22258
rect 11566 22206 11618 22258
rect 11902 22206 11954 22258
rect 12014 22206 12066 22258
rect 12462 22206 12514 22258
rect 12798 22206 12850 22258
rect 19294 22206 19346 22258
rect 19406 22206 19458 22258
rect 19966 22206 20018 22258
rect 20302 22206 20354 22258
rect 20750 22206 20802 22258
rect 21310 22206 21362 22258
rect 23662 22206 23714 22258
rect 29486 22206 29538 22258
rect 29934 22206 29986 22258
rect 30830 22206 30882 22258
rect 30942 22206 30994 22258
rect 6638 22094 6690 22146
rect 11230 22094 11282 22146
rect 12238 22094 12290 22146
rect 21646 22094 21698 22146
rect 26238 22094 26290 22146
rect 26462 22094 26514 22146
rect 28366 22094 28418 22146
rect 28590 22094 28642 22146
rect 28702 22094 28754 22146
rect 29710 22094 29762 22146
rect 32174 22094 32226 22146
rect 32286 22094 32338 22146
rect 9782 21926 9834 21978
rect 9886 21926 9938 21978
rect 9990 21926 10042 21978
rect 18350 21926 18402 21978
rect 18454 21926 18506 21978
rect 18558 21926 18610 21978
rect 26918 21926 26970 21978
rect 27022 21926 27074 21978
rect 27126 21926 27178 21978
rect 35486 21926 35538 21978
rect 35590 21926 35642 21978
rect 35694 21926 35746 21978
rect 7086 21758 7138 21810
rect 7310 21758 7362 21810
rect 7646 21758 7698 21810
rect 7870 21758 7922 21810
rect 10110 21758 10162 21810
rect 11902 21758 11954 21810
rect 12910 21758 12962 21810
rect 17502 21758 17554 21810
rect 21086 21758 21138 21810
rect 25230 21758 25282 21810
rect 25342 21758 25394 21810
rect 25454 21758 25506 21810
rect 34862 21758 34914 21810
rect 4398 21646 4450 21698
rect 11790 21646 11842 21698
rect 13246 21646 13298 21698
rect 13582 21646 13634 21698
rect 24782 21646 24834 21698
rect 28814 21646 28866 21698
rect 29598 21646 29650 21698
rect 32062 21646 32114 21698
rect 32398 21646 32450 21698
rect 34414 21646 34466 21698
rect 35086 21646 35138 21698
rect 35198 21646 35250 21698
rect 3726 21534 3778 21586
rect 7422 21534 7474 21586
rect 7982 21534 8034 21586
rect 8430 21534 8482 21586
rect 10446 21534 10498 21586
rect 12686 21534 12738 21586
rect 13918 21534 13970 21586
rect 20750 21534 20802 21586
rect 21422 21534 21474 21586
rect 25902 21534 25954 21586
rect 26126 21534 26178 21586
rect 27022 21534 27074 21586
rect 27246 21534 27298 21586
rect 27470 21534 27522 21586
rect 29262 21534 29314 21586
rect 31166 21534 31218 21586
rect 31502 21534 31554 21586
rect 33070 21534 33122 21586
rect 33630 21534 33682 21586
rect 34638 21534 34690 21586
rect 6526 21422 6578 21474
rect 8878 21422 8930 21474
rect 10894 21422 10946 21474
rect 14702 21422 14754 21474
rect 16830 21422 16882 21474
rect 17838 21422 17890 21474
rect 19966 21422 20018 21474
rect 21870 21422 21922 21474
rect 22542 21422 22594 21474
rect 22990 21422 23042 21474
rect 23326 21422 23378 21474
rect 23774 21422 23826 21474
rect 24222 21422 24274 21474
rect 25790 21422 25842 21474
rect 30046 21422 30098 21474
rect 33966 21422 34018 21474
rect 11902 21310 11954 21362
rect 21646 21310 21698 21362
rect 22990 21310 23042 21362
rect 23326 21310 23378 21362
rect 23774 21310 23826 21362
rect 26462 21310 26514 21362
rect 32510 21310 32562 21362
rect 5498 21142 5550 21194
rect 5602 21142 5654 21194
rect 5706 21142 5758 21194
rect 14066 21142 14118 21194
rect 14170 21142 14222 21194
rect 14274 21142 14326 21194
rect 22634 21142 22686 21194
rect 22738 21142 22790 21194
rect 22842 21142 22894 21194
rect 31202 21142 31254 21194
rect 31306 21142 31358 21194
rect 31410 21142 31462 21194
rect 29710 20974 29762 21026
rect 31838 20974 31890 21026
rect 34750 20974 34802 21026
rect 12798 20862 12850 20914
rect 14254 20862 14306 20914
rect 16606 20862 16658 20914
rect 22766 20862 22818 20914
rect 23438 20862 23490 20914
rect 25566 20862 25618 20914
rect 27246 20862 27298 20914
rect 28590 20862 28642 20914
rect 31726 20862 31778 20914
rect 6638 20750 6690 20802
rect 8542 20750 8594 20802
rect 9326 20750 9378 20802
rect 9998 20750 10050 20802
rect 13806 20750 13858 20802
rect 14590 20750 14642 20802
rect 16270 20750 16322 20802
rect 16494 20750 16546 20802
rect 16718 20750 16770 20802
rect 16942 20750 16994 20802
rect 18398 20750 18450 20802
rect 18958 20750 19010 20802
rect 26238 20750 26290 20802
rect 26910 20750 26962 20802
rect 27806 20750 27858 20802
rect 28254 20750 28306 20802
rect 28366 20750 28418 20802
rect 29150 20750 29202 20802
rect 29374 20750 29426 20802
rect 30494 20750 30546 20802
rect 32734 20750 32786 20802
rect 6974 20638 7026 20690
rect 7310 20638 7362 20690
rect 7646 20638 7698 20690
rect 7870 20638 7922 20690
rect 9550 20638 9602 20690
rect 10670 20638 10722 20690
rect 14926 20638 14978 20690
rect 15934 20638 15986 20690
rect 17838 20638 17890 20690
rect 18062 20638 18114 20690
rect 18622 20638 18674 20690
rect 21870 20638 21922 20690
rect 27022 20638 27074 20690
rect 27358 20638 27410 20690
rect 30606 20638 30658 20690
rect 31950 20638 32002 20690
rect 6414 20526 6466 20578
rect 6862 20526 6914 20578
rect 7422 20526 7474 20578
rect 8206 20526 8258 20578
rect 13470 20526 13522 20578
rect 16046 20526 16098 20578
rect 18286 20526 18338 20578
rect 18846 20526 18898 20578
rect 21534 20526 21586 20578
rect 27582 20526 27634 20578
rect 9782 20358 9834 20410
rect 9886 20358 9938 20410
rect 9990 20358 10042 20410
rect 18350 20358 18402 20410
rect 18454 20358 18506 20410
rect 18558 20358 18610 20410
rect 26918 20358 26970 20410
rect 27022 20358 27074 20410
rect 27126 20358 27178 20410
rect 35486 20358 35538 20410
rect 35590 20358 35642 20410
rect 35694 20358 35746 20410
rect 11566 20190 11618 20242
rect 17950 20190 18002 20242
rect 23550 20190 23602 20242
rect 8206 20078 8258 20130
rect 9662 20078 9714 20130
rect 9774 20078 9826 20130
rect 10334 20078 10386 20130
rect 10894 20078 10946 20130
rect 11006 20078 11058 20130
rect 11454 20078 11506 20130
rect 13134 20078 13186 20130
rect 13358 20078 13410 20130
rect 14926 20078 14978 20130
rect 15262 20078 15314 20130
rect 15934 20078 15986 20130
rect 16606 20078 16658 20130
rect 16718 20078 16770 20130
rect 17390 20078 17442 20130
rect 18174 20078 18226 20130
rect 18286 20078 18338 20130
rect 19742 20078 19794 20130
rect 23998 20078 24050 20130
rect 24446 20078 24498 20130
rect 26126 20078 26178 20130
rect 26238 20078 26290 20130
rect 26462 20078 26514 20130
rect 27134 20078 27186 20130
rect 27358 20078 27410 20130
rect 29262 20078 29314 20130
rect 30270 20078 30322 20130
rect 31614 20078 31666 20130
rect 33070 20078 33122 20130
rect 33182 20078 33234 20130
rect 5070 19966 5122 20018
rect 8542 19966 8594 20018
rect 8766 19966 8818 20018
rect 9438 19966 9490 20018
rect 11230 19966 11282 20018
rect 11678 19966 11730 20018
rect 12014 19966 12066 20018
rect 12462 19966 12514 20018
rect 12574 19966 12626 20018
rect 13022 19966 13074 20018
rect 13470 19966 13522 20018
rect 15710 19966 15762 20018
rect 16046 19966 16098 20018
rect 16942 19966 16994 20018
rect 17726 19966 17778 20018
rect 19966 19966 20018 20018
rect 21086 19966 21138 20018
rect 21646 19966 21698 20018
rect 22094 19966 22146 20018
rect 22878 19966 22930 20018
rect 24558 19966 24610 20018
rect 25342 19966 25394 20018
rect 25566 19966 25618 20018
rect 25790 19966 25842 20018
rect 26798 19966 26850 20018
rect 29486 19966 29538 20018
rect 29710 19966 29762 20018
rect 31838 19966 31890 20018
rect 31950 19966 32002 20018
rect 33742 19966 33794 20018
rect 34078 19966 34130 20018
rect 34638 19966 34690 20018
rect 5742 19854 5794 19906
rect 7870 19854 7922 19906
rect 8654 19854 8706 19906
rect 12798 19854 12850 19906
rect 20638 19854 20690 19906
rect 21758 19854 21810 19906
rect 22990 19854 23042 19906
rect 25678 19854 25730 19906
rect 27470 19854 27522 19906
rect 27918 19854 27970 19906
rect 31726 19854 31778 19906
rect 35086 19854 35138 19906
rect 26686 19742 26738 19794
rect 32286 19742 32338 19794
rect 32510 19742 32562 19794
rect 33630 19742 33682 19794
rect 5498 19574 5550 19626
rect 5602 19574 5654 19626
rect 5706 19574 5758 19626
rect 14066 19574 14118 19626
rect 14170 19574 14222 19626
rect 14274 19574 14326 19626
rect 22634 19574 22686 19626
rect 22738 19574 22790 19626
rect 22842 19574 22894 19626
rect 31202 19574 31254 19626
rect 31306 19574 31358 19626
rect 31410 19574 31462 19626
rect 25342 19406 25394 19458
rect 25790 19406 25842 19458
rect 31502 19406 31554 19458
rect 34302 19406 34354 19458
rect 6414 19294 6466 19346
rect 8542 19294 8594 19346
rect 10222 19294 10274 19346
rect 12350 19294 12402 19346
rect 19406 19294 19458 19346
rect 27022 19294 27074 19346
rect 30046 19294 30098 19346
rect 32286 19294 32338 19346
rect 5742 19182 5794 19234
rect 8766 19182 8818 19234
rect 9550 19182 9602 19234
rect 12686 19182 12738 19234
rect 14142 19182 14194 19234
rect 14478 19182 14530 19234
rect 14926 19182 14978 19234
rect 15374 19182 15426 19234
rect 15598 19182 15650 19234
rect 15934 19182 15986 19234
rect 16494 19182 16546 19234
rect 20078 19182 20130 19234
rect 20526 19182 20578 19234
rect 23214 19182 23266 19234
rect 25566 19182 25618 19234
rect 26014 19182 26066 19234
rect 27582 19182 27634 19234
rect 28478 19182 28530 19234
rect 30158 19182 30210 19234
rect 30718 19182 30770 19234
rect 32398 19182 32450 19234
rect 34526 19182 34578 19234
rect 34974 19182 35026 19234
rect 8990 19070 9042 19122
rect 9102 19070 9154 19122
rect 12798 19070 12850 19122
rect 13694 19070 13746 19122
rect 13806 19070 13858 19122
rect 14254 19070 14306 19122
rect 17278 19070 17330 19122
rect 21422 19070 21474 19122
rect 22430 19070 22482 19122
rect 22766 19070 22818 19122
rect 24782 19070 24834 19122
rect 26350 19070 26402 19122
rect 26574 19070 26626 19122
rect 28590 19070 28642 19122
rect 29934 19070 29986 19122
rect 31390 19070 31442 19122
rect 13022 18958 13074 19010
rect 13470 18958 13522 19010
rect 15150 18958 15202 19010
rect 16046 18958 16098 19010
rect 16270 18958 16322 19010
rect 20638 18958 20690 19010
rect 22654 18958 22706 19010
rect 23662 18958 23714 19010
rect 24110 18958 24162 19010
rect 26462 18958 26514 19010
rect 28030 18958 28082 19010
rect 9782 18790 9834 18842
rect 9886 18790 9938 18842
rect 9990 18790 10042 18842
rect 18350 18790 18402 18842
rect 18454 18790 18506 18842
rect 18558 18790 18610 18842
rect 26918 18790 26970 18842
rect 27022 18790 27074 18842
rect 27126 18790 27178 18842
rect 35486 18790 35538 18842
rect 35590 18790 35642 18842
rect 35694 18790 35746 18842
rect 8094 18622 8146 18674
rect 8654 18622 8706 18674
rect 10110 18622 10162 18674
rect 12350 18622 12402 18674
rect 12798 18622 12850 18674
rect 17502 18622 17554 18674
rect 28030 18622 28082 18674
rect 29598 18622 29650 18674
rect 30270 18622 30322 18674
rect 34302 18622 34354 18674
rect 7422 18510 7474 18562
rect 7534 18510 7586 18562
rect 8206 18510 8258 18562
rect 12462 18510 12514 18562
rect 25454 18510 25506 18562
rect 26014 18510 26066 18562
rect 27806 18510 27858 18562
rect 30606 18510 30658 18562
rect 31390 18510 31442 18562
rect 33182 18510 33234 18562
rect 34862 18510 34914 18562
rect 7758 18398 7810 18450
rect 7870 18398 7922 18450
rect 8990 18398 9042 18450
rect 9886 18398 9938 18450
rect 10558 18398 10610 18450
rect 13134 18398 13186 18450
rect 13582 18398 13634 18450
rect 13918 18398 13970 18450
rect 14702 18398 14754 18450
rect 17278 18398 17330 18450
rect 17614 18398 17666 18450
rect 17838 18398 17890 18450
rect 23438 18398 23490 18450
rect 26350 18398 26402 18450
rect 26798 18398 26850 18450
rect 26910 18398 26962 18450
rect 27022 18398 27074 18450
rect 28366 18398 28418 18450
rect 28702 18398 28754 18450
rect 29150 18398 29202 18450
rect 29822 18398 29874 18450
rect 31838 18398 31890 18450
rect 32174 18398 32226 18450
rect 33406 18398 33458 18450
rect 33854 18398 33906 18450
rect 34078 18398 34130 18450
rect 16830 18286 16882 18338
rect 18846 18286 18898 18338
rect 21646 18286 21698 18338
rect 25118 18286 25170 18338
rect 27470 18286 27522 18338
rect 31726 18286 31778 18338
rect 33070 18286 33122 18338
rect 12350 18174 12402 18226
rect 28142 18174 28194 18226
rect 34638 18174 34690 18226
rect 5498 18006 5550 18058
rect 5602 18006 5654 18058
rect 5706 18006 5758 18058
rect 14066 18006 14118 18058
rect 14170 18006 14222 18058
rect 14274 18006 14326 18058
rect 22634 18006 22686 18058
rect 22738 18006 22790 18058
rect 22842 18006 22894 18058
rect 31202 18006 31254 18058
rect 31306 18006 31358 18058
rect 31410 18006 31462 18058
rect 20638 17838 20690 17890
rect 23550 17838 23602 17890
rect 24782 17838 24834 17890
rect 25118 17838 25170 17890
rect 28478 17838 28530 17890
rect 30942 17838 30994 17890
rect 10222 17726 10274 17778
rect 10782 17726 10834 17778
rect 16158 17726 16210 17778
rect 17054 17726 17106 17778
rect 21422 17726 21474 17778
rect 24558 17726 24610 17778
rect 29262 17726 29314 17778
rect 30830 17726 30882 17778
rect 31278 17726 31330 17778
rect 32286 17726 32338 17778
rect 7310 17614 7362 17666
rect 12350 17614 12402 17666
rect 12686 17614 12738 17666
rect 12910 17614 12962 17666
rect 13470 17614 13522 17666
rect 14030 17614 14082 17666
rect 14590 17614 14642 17666
rect 18062 17614 18114 17666
rect 18286 17614 18338 17666
rect 19630 17614 19682 17666
rect 20302 17614 20354 17666
rect 22318 17614 22370 17666
rect 22990 17614 23042 17666
rect 23998 17614 24050 17666
rect 24334 17614 24386 17666
rect 25454 17614 25506 17666
rect 26574 17614 26626 17666
rect 26798 17614 26850 17666
rect 27022 17614 27074 17666
rect 28590 17614 28642 17666
rect 31726 17614 31778 17666
rect 35086 17614 35138 17666
rect 8094 17502 8146 17554
rect 13806 17502 13858 17554
rect 14254 17502 14306 17554
rect 14478 17502 14530 17554
rect 17838 17502 17890 17554
rect 18622 17502 18674 17554
rect 19406 17502 19458 17554
rect 20750 17502 20802 17554
rect 22430 17502 22482 17554
rect 22654 17502 22706 17554
rect 26238 17502 26290 17554
rect 27470 17502 27522 17554
rect 27918 17502 27970 17554
rect 30158 17502 30210 17554
rect 34414 17502 34466 17554
rect 12462 17390 12514 17442
rect 13582 17390 13634 17442
rect 19518 17390 19570 17442
rect 21870 17390 21922 17442
rect 25118 17390 25170 17442
rect 25566 17390 25618 17442
rect 28478 17390 28530 17442
rect 29822 17390 29874 17442
rect 30270 17390 30322 17442
rect 30382 17390 30434 17442
rect 9782 17222 9834 17274
rect 9886 17222 9938 17274
rect 9990 17222 10042 17274
rect 18350 17222 18402 17274
rect 18454 17222 18506 17274
rect 18558 17222 18610 17274
rect 26918 17222 26970 17274
rect 27022 17222 27074 17274
rect 27126 17222 27178 17274
rect 35486 17222 35538 17274
rect 35590 17222 35642 17274
rect 35694 17222 35746 17274
rect 8542 17054 8594 17106
rect 9886 17054 9938 17106
rect 9998 17054 10050 17106
rect 10782 17054 10834 17106
rect 15262 17054 15314 17106
rect 16830 17054 16882 17106
rect 18846 17054 18898 17106
rect 19406 17054 19458 17106
rect 20862 17054 20914 17106
rect 23102 17054 23154 17106
rect 25678 17054 25730 17106
rect 27582 17054 27634 17106
rect 27918 17054 27970 17106
rect 28590 17054 28642 17106
rect 30718 17054 30770 17106
rect 33966 17054 34018 17106
rect 34638 17054 34690 17106
rect 8990 16942 9042 16994
rect 12686 16942 12738 16994
rect 17614 16942 17666 16994
rect 17838 16942 17890 16994
rect 17950 16942 18002 16994
rect 19742 16942 19794 16994
rect 21982 16942 22034 16994
rect 24222 16942 24274 16994
rect 25454 16942 25506 16994
rect 26014 16942 26066 16994
rect 26686 16942 26738 16994
rect 28366 16942 28418 16994
rect 28926 16942 28978 16994
rect 29486 16942 29538 16994
rect 32174 16942 32226 16994
rect 8430 16830 8482 16882
rect 8766 16830 8818 16882
rect 9774 16830 9826 16882
rect 10334 16830 10386 16882
rect 12014 16830 12066 16882
rect 18174 16830 18226 16882
rect 19854 16830 19906 16882
rect 21422 16830 21474 16882
rect 21758 16830 21810 16882
rect 22206 16830 22258 16882
rect 22542 16830 22594 16882
rect 23438 16830 23490 16882
rect 25230 16830 25282 16882
rect 26910 16830 26962 16882
rect 28814 16830 28866 16882
rect 30046 16830 30098 16882
rect 31726 16830 31778 16882
rect 32398 16830 32450 16882
rect 33070 16830 33122 16882
rect 33518 16830 33570 16882
rect 34190 16830 34242 16882
rect 35198 16830 35250 16882
rect 14814 16718 14866 16770
rect 17950 16718 18002 16770
rect 28030 16718 28082 16770
rect 29150 16718 29202 16770
rect 30830 16718 30882 16770
rect 30942 16718 30994 16770
rect 31278 16718 31330 16770
rect 27246 16606 27298 16658
rect 27470 16606 27522 16658
rect 5498 16438 5550 16490
rect 5602 16438 5654 16490
rect 5706 16438 5758 16490
rect 14066 16438 14118 16490
rect 14170 16438 14222 16490
rect 14274 16438 14326 16490
rect 22634 16438 22686 16490
rect 22738 16438 22790 16490
rect 22842 16438 22894 16490
rect 31202 16438 31254 16490
rect 31306 16438 31358 16490
rect 31410 16438 31462 16490
rect 21422 16270 21474 16322
rect 25118 16270 25170 16322
rect 33070 16270 33122 16322
rect 35086 16270 35138 16322
rect 9214 16158 9266 16210
rect 10782 16158 10834 16210
rect 12910 16158 12962 16210
rect 15374 16158 15426 16210
rect 16830 16158 16882 16210
rect 19854 16158 19906 16210
rect 20302 16158 20354 16210
rect 22878 16158 22930 16210
rect 28030 16158 28082 16210
rect 29262 16158 29314 16210
rect 10110 16046 10162 16098
rect 16494 16046 16546 16098
rect 17838 16046 17890 16098
rect 18734 16046 18786 16098
rect 20750 16046 20802 16098
rect 21758 16046 21810 16098
rect 23886 16046 23938 16098
rect 24222 16046 24274 16098
rect 24446 16046 24498 16098
rect 25454 16046 25506 16098
rect 26462 16046 26514 16098
rect 27470 16046 27522 16098
rect 27918 16046 27970 16098
rect 28142 16046 28194 16098
rect 28590 16046 28642 16098
rect 32174 16046 32226 16098
rect 32734 16046 32786 16098
rect 34638 16046 34690 16098
rect 35198 16046 35250 16098
rect 13582 15934 13634 15986
rect 15262 15934 15314 15986
rect 16382 15934 16434 15986
rect 21982 15934 22034 15986
rect 23438 15934 23490 15986
rect 24670 15934 24722 15986
rect 25678 15934 25730 15986
rect 26798 15934 26850 15986
rect 26910 15934 26962 15986
rect 31502 15934 31554 15986
rect 33294 15934 33346 15986
rect 33630 15934 33682 15986
rect 34302 15934 34354 15986
rect 35086 15934 35138 15986
rect 13918 15822 13970 15874
rect 14926 15822 14978 15874
rect 19070 15822 19122 15874
rect 23102 15822 23154 15874
rect 27022 15822 27074 15874
rect 27134 15822 27186 15874
rect 27694 15822 27746 15874
rect 28478 15822 28530 15874
rect 9782 15654 9834 15706
rect 9886 15654 9938 15706
rect 9990 15654 10042 15706
rect 18350 15654 18402 15706
rect 18454 15654 18506 15706
rect 18558 15654 18610 15706
rect 26918 15654 26970 15706
rect 27022 15654 27074 15706
rect 27126 15654 27178 15706
rect 35486 15654 35538 15706
rect 35590 15654 35642 15706
rect 35694 15654 35746 15706
rect 13246 15486 13298 15538
rect 13470 15486 13522 15538
rect 13806 15486 13858 15538
rect 15598 15486 15650 15538
rect 21198 15486 21250 15538
rect 34750 15486 34802 15538
rect 35086 15486 35138 15538
rect 14142 15374 14194 15426
rect 14814 15374 14866 15426
rect 25790 15374 25842 15426
rect 25902 15374 25954 15426
rect 33182 15374 33234 15426
rect 33742 15374 33794 15426
rect 34302 15374 34354 15426
rect 14366 15262 14418 15314
rect 15150 15262 15202 15314
rect 17502 15262 17554 15314
rect 17950 15262 18002 15314
rect 21758 15262 21810 15314
rect 21982 15262 22034 15314
rect 24222 15262 24274 15314
rect 25678 15262 25730 15314
rect 26910 15262 26962 15314
rect 27134 15262 27186 15314
rect 27582 15262 27634 15314
rect 27806 15262 27858 15314
rect 28702 15262 28754 15314
rect 30494 15262 30546 15314
rect 31838 15262 31890 15314
rect 14926 15150 14978 15202
rect 20414 15150 20466 15202
rect 22318 15150 22370 15202
rect 24558 15150 24610 15202
rect 26350 15150 26402 15202
rect 27358 15150 27410 15202
rect 29822 15150 29874 15202
rect 31502 15150 31554 15202
rect 32510 15150 32562 15202
rect 25230 15038 25282 15090
rect 28142 15038 28194 15090
rect 28478 15038 28530 15090
rect 32398 15038 32450 15090
rect 33518 15038 33570 15090
rect 5498 14870 5550 14922
rect 5602 14870 5654 14922
rect 5706 14870 5758 14922
rect 14066 14870 14118 14922
rect 14170 14870 14222 14922
rect 14274 14870 14326 14922
rect 22634 14870 22686 14922
rect 22738 14870 22790 14922
rect 22842 14870 22894 14922
rect 31202 14870 31254 14922
rect 31306 14870 31358 14922
rect 31410 14870 31462 14922
rect 20750 14702 20802 14754
rect 28478 14702 28530 14754
rect 31726 14702 31778 14754
rect 8318 14590 8370 14642
rect 9214 14590 9266 14642
rect 11790 14590 11842 14642
rect 14478 14590 14530 14642
rect 16606 14590 16658 14642
rect 16942 14590 16994 14642
rect 19070 14590 19122 14642
rect 20638 14590 20690 14642
rect 25342 14590 25394 14642
rect 32286 14590 32338 14642
rect 10222 14478 10274 14530
rect 10446 14478 10498 14530
rect 10670 14478 10722 14530
rect 11006 14478 11058 14530
rect 13806 14478 13858 14530
rect 19854 14478 19906 14530
rect 20414 14478 20466 14530
rect 23214 14478 23266 14530
rect 27470 14478 27522 14530
rect 30942 14478 30994 14530
rect 35086 14478 35138 14530
rect 11230 14366 11282 14418
rect 11342 14366 11394 14418
rect 27918 14366 27970 14418
rect 28590 14366 28642 14418
rect 29150 14366 29202 14418
rect 29934 14366 29986 14418
rect 34414 14366 34466 14418
rect 10334 14254 10386 14306
rect 21422 14254 21474 14306
rect 28478 14254 28530 14306
rect 9782 14086 9834 14138
rect 9886 14086 9938 14138
rect 9990 14086 10042 14138
rect 18350 14086 18402 14138
rect 18454 14086 18506 14138
rect 18558 14086 18610 14138
rect 26918 14086 26970 14138
rect 27022 14086 27074 14138
rect 27126 14086 27178 14138
rect 35486 14086 35538 14138
rect 35590 14086 35642 14138
rect 35694 14086 35746 14138
rect 7086 13918 7138 13970
rect 8094 13918 8146 13970
rect 8990 13918 9042 13970
rect 14926 13918 14978 13970
rect 17390 13918 17442 13970
rect 19518 13918 19570 13970
rect 19742 13918 19794 13970
rect 20414 13918 20466 13970
rect 20750 13918 20802 13970
rect 25230 13918 25282 13970
rect 33182 13918 33234 13970
rect 35086 13918 35138 13970
rect 10334 13806 10386 13858
rect 15598 13806 15650 13858
rect 17950 13806 18002 13858
rect 19406 13806 19458 13858
rect 19966 13806 20018 13858
rect 20078 13806 20130 13858
rect 22318 13806 22370 13858
rect 23102 13806 23154 13858
rect 25790 13806 25842 13858
rect 27358 13806 27410 13858
rect 28142 13806 28194 13858
rect 33742 13806 33794 13858
rect 34190 13806 34242 13858
rect 34750 13806 34802 13858
rect 6862 13694 6914 13746
rect 7198 13694 7250 13746
rect 7422 13694 7474 13746
rect 9550 13694 9602 13746
rect 13358 13694 13410 13746
rect 14366 13694 14418 13746
rect 14702 13694 14754 13746
rect 15374 13694 15426 13746
rect 22766 13694 22818 13746
rect 24558 13694 24610 13746
rect 25566 13694 25618 13746
rect 27134 13694 27186 13746
rect 28030 13694 28082 13746
rect 28814 13694 28866 13746
rect 29710 13694 29762 13746
rect 8430 13582 8482 13634
rect 12462 13582 12514 13634
rect 12798 13582 12850 13634
rect 13806 13582 13858 13634
rect 16158 13582 16210 13634
rect 18622 13582 18674 13634
rect 21870 13582 21922 13634
rect 30382 13582 30434 13634
rect 32510 13582 32562 13634
rect 26350 13470 26402 13522
rect 26686 13470 26738 13522
rect 29150 13470 29202 13522
rect 33518 13470 33570 13522
rect 5498 13302 5550 13354
rect 5602 13302 5654 13354
rect 5706 13302 5758 13354
rect 14066 13302 14118 13354
rect 14170 13302 14222 13354
rect 14274 13302 14326 13354
rect 22634 13302 22686 13354
rect 22738 13302 22790 13354
rect 22842 13302 22894 13354
rect 31202 13302 31254 13354
rect 31306 13302 31358 13354
rect 31410 13302 31462 13354
rect 6190 13134 6242 13186
rect 27918 13134 27970 13186
rect 28254 13134 28306 13186
rect 31726 13134 31778 13186
rect 8542 13022 8594 13074
rect 10670 13022 10722 13074
rect 12798 13022 12850 13074
rect 22430 13022 22482 13074
rect 24334 13022 24386 13074
rect 24670 13022 24722 13074
rect 26798 13022 26850 13074
rect 28478 13022 28530 13074
rect 30494 13022 30546 13074
rect 32286 13022 32338 13074
rect 6526 12910 6578 12962
rect 7198 12910 7250 12962
rect 7646 12910 7698 12962
rect 8094 12910 8146 12962
rect 9998 12910 10050 12962
rect 10334 12910 10386 12962
rect 11566 12910 11618 12962
rect 12126 12910 12178 12962
rect 12462 12910 12514 12962
rect 20526 12910 20578 12962
rect 21870 12910 21922 12962
rect 22542 12910 22594 12962
rect 22990 12910 23042 12962
rect 23326 12910 23378 12962
rect 24222 12910 24274 12962
rect 27582 12910 27634 12962
rect 29150 12910 29202 12962
rect 29374 12910 29426 12962
rect 29710 12910 29762 12962
rect 30046 12910 30098 12962
rect 30270 12910 30322 12962
rect 30606 12910 30658 12962
rect 31166 12910 31218 12962
rect 35086 12910 35138 12962
rect 6302 12798 6354 12850
rect 6974 12798 7026 12850
rect 8878 12798 8930 12850
rect 9662 12798 9714 12850
rect 10782 12798 10834 12850
rect 11790 12798 11842 12850
rect 12238 12798 12290 12850
rect 19406 12798 19458 12850
rect 19742 12798 19794 12850
rect 19966 12798 20018 12850
rect 22766 12798 22818 12850
rect 23214 12798 23266 12850
rect 23998 12798 24050 12850
rect 31838 12798 31890 12850
rect 34414 12798 34466 12850
rect 6190 12686 6242 12738
rect 6862 12686 6914 12738
rect 7534 12686 7586 12738
rect 7758 12686 7810 12738
rect 8430 12686 8482 12738
rect 8654 12686 8706 12738
rect 10110 12686 10162 12738
rect 10558 12686 10610 12738
rect 11006 12686 11058 12738
rect 15150 12686 15202 12738
rect 15486 12686 15538 12738
rect 16158 12686 16210 12738
rect 16494 12686 16546 12738
rect 19518 12686 19570 12738
rect 20302 12686 20354 12738
rect 29486 12686 29538 12738
rect 30942 12686 30994 12738
rect 31726 12686 31778 12738
rect 9782 12518 9834 12570
rect 9886 12518 9938 12570
rect 9990 12518 10042 12570
rect 18350 12518 18402 12570
rect 18454 12518 18506 12570
rect 18558 12518 18610 12570
rect 26918 12518 26970 12570
rect 27022 12518 27074 12570
rect 27126 12518 27178 12570
rect 35486 12518 35538 12570
rect 35590 12518 35642 12570
rect 35694 12518 35746 12570
rect 7982 12350 8034 12402
rect 8654 12350 8706 12402
rect 8990 12350 9042 12402
rect 13582 12350 13634 12402
rect 21198 12350 21250 12402
rect 22206 12350 22258 12402
rect 23662 12350 23714 12402
rect 32062 12350 32114 12402
rect 32286 12350 32338 12402
rect 33182 12350 33234 12402
rect 34862 12350 34914 12402
rect 6974 12238 7026 12290
rect 8206 12238 8258 12290
rect 8318 12238 8370 12290
rect 13246 12238 13298 12290
rect 18734 12238 18786 12290
rect 22318 12238 22370 12290
rect 22654 12238 22706 12290
rect 24110 12238 24162 12290
rect 33742 12238 33794 12290
rect 34078 12238 34130 12290
rect 7646 12126 7698 12178
rect 11678 12126 11730 12178
rect 12462 12126 12514 12178
rect 13918 12126 13970 12178
rect 17950 12126 18002 12178
rect 22990 12126 23042 12178
rect 23214 12126 23266 12178
rect 24558 12126 24610 12178
rect 25454 12126 25506 12178
rect 25902 12126 25954 12178
rect 27246 12126 27298 12178
rect 32398 12126 32450 12178
rect 35086 12126 35138 12178
rect 4846 12014 4898 12066
rect 9550 12014 9602 12066
rect 14702 12014 14754 12066
rect 16830 12014 16882 12066
rect 20862 12014 20914 12066
rect 21758 12014 21810 12066
rect 22766 12014 22818 12066
rect 24670 12014 24722 12066
rect 30046 12014 30098 12066
rect 25902 11902 25954 11954
rect 33518 11902 33570 11954
rect 5498 11734 5550 11786
rect 5602 11734 5654 11786
rect 5706 11734 5758 11786
rect 14066 11734 14118 11786
rect 14170 11734 14222 11786
rect 14274 11734 14326 11786
rect 22634 11734 22686 11786
rect 22738 11734 22790 11786
rect 22842 11734 22894 11786
rect 31202 11734 31254 11786
rect 31306 11734 31358 11786
rect 31410 11734 31462 11786
rect 27918 11566 27970 11618
rect 28478 11566 28530 11618
rect 5630 11454 5682 11506
rect 7758 11454 7810 11506
rect 9886 11454 9938 11506
rect 10558 11454 10610 11506
rect 14926 11454 14978 11506
rect 19406 11454 19458 11506
rect 20638 11454 20690 11506
rect 22430 11454 22482 11506
rect 24558 11454 24610 11506
rect 26798 11454 26850 11506
rect 29598 11454 29650 11506
rect 32958 11454 33010 11506
rect 33518 11454 33570 11506
rect 34638 11454 34690 11506
rect 8542 11342 8594 11394
rect 10446 11342 10498 11394
rect 11006 11342 11058 11394
rect 11454 11342 11506 11394
rect 11902 11342 11954 11394
rect 15038 11342 15090 11394
rect 15374 11342 15426 11394
rect 15822 11342 15874 11394
rect 15934 11342 15986 11394
rect 17166 11342 17218 11394
rect 19518 11342 19570 11394
rect 20190 11342 20242 11394
rect 21646 11342 21698 11394
rect 25454 11342 25506 11394
rect 26014 11342 26066 11394
rect 27358 11342 27410 11394
rect 27582 11342 27634 11394
rect 29150 11342 29202 11394
rect 30046 11342 30098 11394
rect 33854 11342 33906 11394
rect 35086 11342 35138 11394
rect 10670 11230 10722 11282
rect 14814 11230 14866 11282
rect 16606 11230 16658 11282
rect 26238 11230 26290 11282
rect 27806 11230 27858 11282
rect 28366 11230 28418 11282
rect 30830 11230 30882 11282
rect 34190 11230 34242 11282
rect 9102 11118 9154 11170
rect 9438 11118 9490 11170
rect 15710 11118 15762 11170
rect 16158 11118 16210 11170
rect 19294 11118 19346 11170
rect 19742 11118 19794 11170
rect 20526 11118 20578 11170
rect 20750 11118 20802 11170
rect 24894 11118 24946 11170
rect 25006 11118 25058 11170
rect 25118 11118 25170 11170
rect 9782 10950 9834 11002
rect 9886 10950 9938 11002
rect 9990 10950 10042 11002
rect 18350 10950 18402 11002
rect 18454 10950 18506 11002
rect 18558 10950 18610 11002
rect 26918 10950 26970 11002
rect 27022 10950 27074 11002
rect 27126 10950 27178 11002
rect 35486 10950 35538 11002
rect 35590 10950 35642 11002
rect 35694 10950 35746 11002
rect 7982 10782 8034 10834
rect 9662 10782 9714 10834
rect 10334 10782 10386 10834
rect 12014 10782 12066 10834
rect 21422 10782 21474 10834
rect 21646 10782 21698 10834
rect 22318 10782 22370 10834
rect 22766 10782 22818 10834
rect 23326 10782 23378 10834
rect 23662 10782 23714 10834
rect 23774 10782 23826 10834
rect 24334 10782 24386 10834
rect 26574 10782 26626 10834
rect 27358 10782 27410 10834
rect 31054 10782 31106 10834
rect 31278 10782 31330 10834
rect 32286 10782 32338 10834
rect 33518 10782 33570 10834
rect 33854 10782 33906 10834
rect 20862 10670 20914 10722
rect 21086 10670 21138 10722
rect 22430 10670 22482 10722
rect 25566 10670 25618 10722
rect 29710 10670 29762 10722
rect 30830 10670 30882 10722
rect 31838 10670 31890 10722
rect 9774 10558 9826 10610
rect 12462 10558 12514 10610
rect 15598 10558 15650 10610
rect 15822 10558 15874 10610
rect 16158 10558 16210 10610
rect 20526 10558 20578 10610
rect 21534 10558 21586 10610
rect 22094 10558 22146 10610
rect 22542 10558 22594 10610
rect 23550 10558 23602 10610
rect 24110 10558 24162 10610
rect 24222 10558 24274 10610
rect 24670 10558 24722 10610
rect 25230 10558 25282 10610
rect 25678 10558 25730 10610
rect 30494 10558 30546 10610
rect 34190 10558 34242 10610
rect 34638 10558 34690 10610
rect 35086 10558 35138 10610
rect 10894 10446 10946 10498
rect 13134 10446 13186 10498
rect 15262 10446 15314 10498
rect 15710 10446 15762 10498
rect 20638 10446 20690 10498
rect 25342 10446 25394 10498
rect 27582 10446 27634 10498
rect 30942 10446 30994 10498
rect 9662 10334 9714 10386
rect 5498 10166 5550 10218
rect 5602 10166 5654 10218
rect 5706 10166 5758 10218
rect 14066 10166 14118 10218
rect 14170 10166 14222 10218
rect 14274 10166 14326 10218
rect 22634 10166 22686 10218
rect 22738 10166 22790 10218
rect 22842 10166 22894 10218
rect 31202 10166 31254 10218
rect 31306 10166 31358 10218
rect 31410 10166 31462 10218
rect 29262 9998 29314 10050
rect 29486 9998 29538 10050
rect 9886 9886 9938 9938
rect 14142 9886 14194 9938
rect 18286 9886 18338 9938
rect 22654 9886 22706 9938
rect 24782 9886 24834 9938
rect 26910 9886 26962 9938
rect 27358 9886 27410 9938
rect 29486 9886 29538 9938
rect 30158 9886 30210 9938
rect 32734 9886 32786 9938
rect 33182 9886 33234 9938
rect 33630 9886 33682 9938
rect 34078 9886 34130 9938
rect 7086 9774 7138 9826
rect 10670 9774 10722 9826
rect 11118 9774 11170 9826
rect 11566 9774 11618 9826
rect 11790 9774 11842 9826
rect 12350 9774 12402 9826
rect 12910 9774 12962 9826
rect 14590 9774 14642 9826
rect 14926 9774 14978 9826
rect 16046 9774 16098 9826
rect 16942 9774 16994 9826
rect 20302 9774 20354 9826
rect 22542 9774 22594 9826
rect 23214 9774 23266 9826
rect 24110 9774 24162 9826
rect 28254 9774 28306 9826
rect 29822 9774 29874 9826
rect 30382 9774 30434 9826
rect 30830 9774 30882 9826
rect 34638 9774 34690 9826
rect 35198 9774 35250 9826
rect 7758 9662 7810 9714
rect 14030 9662 14082 9714
rect 14366 9662 14418 9714
rect 16718 9662 16770 9714
rect 17278 9662 17330 9714
rect 17502 9662 17554 9714
rect 17838 9662 17890 9714
rect 20526 9662 20578 9714
rect 22094 9662 22146 9714
rect 28590 9662 28642 9714
rect 29934 9662 29986 9714
rect 10334 9550 10386 9602
rect 11454 9550 11506 9602
rect 12238 9550 12290 9602
rect 12462 9550 12514 9602
rect 13582 9550 13634 9602
rect 15262 9550 15314 9602
rect 15374 9550 15426 9602
rect 15486 9550 15538 9602
rect 15822 9550 15874 9602
rect 15934 9550 15986 9602
rect 16270 9550 16322 9602
rect 17166 9550 17218 9602
rect 17726 9550 17778 9602
rect 30606 9662 30658 9714
rect 31166 9662 31218 9714
rect 34862 9662 34914 9714
rect 22318 9550 22370 9602
rect 22766 9550 22818 9602
rect 30718 9550 30770 9602
rect 9782 9382 9834 9434
rect 9886 9382 9938 9434
rect 9990 9382 10042 9434
rect 18350 9382 18402 9434
rect 18454 9382 18506 9434
rect 18558 9382 18610 9434
rect 26918 9382 26970 9434
rect 27022 9382 27074 9434
rect 27126 9382 27178 9434
rect 35486 9382 35538 9434
rect 35590 9382 35642 9434
rect 35694 9382 35746 9434
rect 8206 9214 8258 9266
rect 16158 9214 16210 9266
rect 16606 9214 16658 9266
rect 22430 9214 22482 9266
rect 23774 9214 23826 9266
rect 24782 9214 24834 9266
rect 25230 9214 25282 9266
rect 25566 9214 25618 9266
rect 26014 9214 26066 9266
rect 26350 9214 26402 9266
rect 30606 9214 30658 9266
rect 31390 9214 31442 9266
rect 31502 9214 31554 9266
rect 33966 9214 34018 9266
rect 34414 9214 34466 9266
rect 34862 9214 34914 9266
rect 35198 9214 35250 9266
rect 7422 9102 7474 9154
rect 17390 9102 17442 9154
rect 18286 9102 18338 9154
rect 20078 9102 20130 9154
rect 22654 9102 22706 9154
rect 23998 9102 24050 9154
rect 24110 9102 24162 9154
rect 24558 9102 24610 9154
rect 26686 9102 26738 9154
rect 28030 9102 28082 9154
rect 32398 9102 32450 9154
rect 7086 8990 7138 9042
rect 7646 8990 7698 9042
rect 8094 8990 8146 9042
rect 8430 8990 8482 9042
rect 8654 8990 8706 9042
rect 14814 8990 14866 9042
rect 16382 8990 16434 9042
rect 16494 8990 16546 9042
rect 17614 8990 17666 9042
rect 18062 8990 18114 9042
rect 18622 8990 18674 9042
rect 19294 8990 19346 9042
rect 22766 8990 22818 9042
rect 24446 8990 24498 9042
rect 27358 8990 27410 9042
rect 30494 8990 30546 9042
rect 30718 8990 30770 9042
rect 31166 8990 31218 9042
rect 31614 8990 31666 9042
rect 31950 8990 32002 9042
rect 32286 8990 32338 9042
rect 4174 8878 4226 8930
rect 6302 8878 6354 8930
rect 12126 8878 12178 8930
rect 15262 8878 15314 8930
rect 15710 8878 15762 8930
rect 17502 8878 17554 8930
rect 22206 8878 22258 8930
rect 30158 8878 30210 8930
rect 32398 8766 32450 8818
rect 5498 8598 5550 8650
rect 5602 8598 5654 8650
rect 5706 8598 5758 8650
rect 14066 8598 14118 8650
rect 14170 8598 14222 8650
rect 14274 8598 14326 8650
rect 22634 8598 22686 8650
rect 22738 8598 22790 8650
rect 22842 8598 22894 8650
rect 31202 8598 31254 8650
rect 31306 8598 31358 8650
rect 31410 8598 31462 8650
rect 6638 8318 6690 8370
rect 8542 8318 8594 8370
rect 9438 8318 9490 8370
rect 9774 8318 9826 8370
rect 11902 8318 11954 8370
rect 19294 8318 19346 8370
rect 21534 8318 21586 8370
rect 25006 8318 25058 8370
rect 29934 8318 29986 8370
rect 34190 8318 34242 8370
rect 6862 8206 6914 8258
rect 7086 8206 7138 8258
rect 7534 8206 7586 8258
rect 7646 8206 7698 8258
rect 8094 8206 8146 8258
rect 9102 8206 9154 8258
rect 12574 8206 12626 8258
rect 14142 8206 14194 8258
rect 14478 8206 14530 8258
rect 14702 8206 14754 8258
rect 16718 8206 16770 8258
rect 27246 8206 27298 8258
rect 29822 8206 29874 8258
rect 30718 8206 30770 8258
rect 31278 8206 31330 8258
rect 5966 8094 6018 8146
rect 6302 8094 6354 8146
rect 6526 8094 6578 8146
rect 13582 8094 13634 8146
rect 13694 8094 13746 8146
rect 28030 8094 28082 8146
rect 30046 8094 30098 8146
rect 32062 8094 32114 8146
rect 34862 8094 34914 8146
rect 35198 8094 35250 8146
rect 6078 7982 6130 8034
rect 7422 7982 7474 8034
rect 8430 7982 8482 8034
rect 8654 7982 8706 8034
rect 13918 7982 13970 8034
rect 14254 7982 14306 8034
rect 27470 7982 27522 8034
rect 28366 7982 28418 8034
rect 29598 7982 29650 8034
rect 30494 7982 30546 8034
rect 30830 7982 30882 8034
rect 30942 7982 30994 8034
rect 9782 7814 9834 7866
rect 9886 7814 9938 7866
rect 9990 7814 10042 7866
rect 18350 7814 18402 7866
rect 18454 7814 18506 7866
rect 18558 7814 18610 7866
rect 26918 7814 26970 7866
rect 27022 7814 27074 7866
rect 27126 7814 27178 7866
rect 35486 7814 35538 7866
rect 35590 7814 35642 7866
rect 35694 7814 35746 7866
rect 7086 7646 7138 7698
rect 9102 7646 9154 7698
rect 10782 7646 10834 7698
rect 11118 7646 11170 7698
rect 15598 7646 15650 7698
rect 15710 7646 15762 7698
rect 15822 7646 15874 7698
rect 17390 7646 17442 7698
rect 17726 7646 17778 7698
rect 18398 7646 18450 7698
rect 20190 7646 20242 7698
rect 20750 7646 20802 7698
rect 24446 7646 24498 7698
rect 25902 7646 25954 7698
rect 29374 7646 29426 7698
rect 29598 7646 29650 7698
rect 29822 7646 29874 7698
rect 31166 7646 31218 7698
rect 31614 7646 31666 7698
rect 32062 7646 32114 7698
rect 33966 7646 34018 7698
rect 35310 7646 35362 7698
rect 6414 7534 6466 7586
rect 7982 7534 8034 7586
rect 9550 7534 9602 7586
rect 11566 7534 11618 7586
rect 12910 7534 12962 7586
rect 16494 7534 16546 7586
rect 18510 7534 18562 7586
rect 18846 7534 18898 7586
rect 19182 7534 19234 7586
rect 19518 7534 19570 7586
rect 19854 7534 19906 7586
rect 20974 7534 21026 7586
rect 21086 7534 21138 7586
rect 21422 7534 21474 7586
rect 21534 7534 21586 7586
rect 25342 7534 25394 7586
rect 26574 7534 26626 7586
rect 27246 7534 27298 7586
rect 27582 7534 27634 7586
rect 28030 7534 28082 7586
rect 28590 7534 28642 7586
rect 30046 7534 30098 7586
rect 30270 7534 30322 7586
rect 31838 7534 31890 7586
rect 6302 7422 6354 7474
rect 6862 7422 6914 7474
rect 7198 7422 7250 7474
rect 7310 7422 7362 7474
rect 7758 7422 7810 7474
rect 8206 7422 8258 7474
rect 8542 7422 8594 7474
rect 9998 7422 10050 7474
rect 11454 7422 11506 7474
rect 12126 7422 12178 7474
rect 16270 7422 16322 7474
rect 16718 7422 16770 7474
rect 18174 7422 18226 7474
rect 20414 7422 20466 7474
rect 23438 7422 23490 7474
rect 23774 7422 23826 7474
rect 23998 7422 24050 7474
rect 24222 7422 24274 7474
rect 24558 7422 24610 7474
rect 25118 7422 25170 7474
rect 25454 7422 25506 7474
rect 25790 7422 25842 7474
rect 26126 7422 26178 7474
rect 26798 7422 26850 7474
rect 27806 7422 27858 7474
rect 28142 7422 28194 7474
rect 28478 7422 28530 7474
rect 28814 7422 28866 7474
rect 29262 7422 29314 7474
rect 29934 7422 29986 7474
rect 30830 7422 30882 7474
rect 31054 7422 31106 7474
rect 31278 7422 31330 7474
rect 6638 7310 6690 7362
rect 8094 7310 8146 7362
rect 15038 7310 15090 7362
rect 23550 7310 23602 7362
rect 31726 7310 31778 7362
rect 34078 7310 34130 7362
rect 11566 7198 11618 7250
rect 21534 7198 21586 7250
rect 5498 7030 5550 7082
rect 5602 7030 5654 7082
rect 5706 7030 5758 7082
rect 14066 7030 14118 7082
rect 14170 7030 14222 7082
rect 14274 7030 14326 7082
rect 22634 7030 22686 7082
rect 22738 7030 22790 7082
rect 22842 7030 22894 7082
rect 31202 7030 31254 7082
rect 31306 7030 31358 7082
rect 31410 7030 31462 7082
rect 15038 6750 15090 6802
rect 24222 6750 24274 6802
rect 6526 6638 6578 6690
rect 6750 6638 6802 6690
rect 7198 6638 7250 6690
rect 9662 6638 9714 6690
rect 12462 6638 12514 6690
rect 13918 6638 13970 6690
rect 17166 6638 17218 6690
rect 17950 6638 18002 6690
rect 18734 6638 18786 6690
rect 19294 6638 19346 6690
rect 19630 6638 19682 6690
rect 20302 6638 20354 6690
rect 20862 6638 20914 6690
rect 21310 6638 21362 6690
rect 22094 6638 22146 6690
rect 25118 6638 25170 6690
rect 25566 6638 25618 6690
rect 25678 6638 25730 6690
rect 26462 6638 26514 6690
rect 26910 6638 26962 6690
rect 27470 6638 27522 6690
rect 28142 6638 28194 6690
rect 29038 6638 29090 6690
rect 29598 6638 29650 6690
rect 29934 6638 29986 6690
rect 30382 6638 30434 6690
rect 30606 6638 30658 6690
rect 31166 6638 31218 6690
rect 8318 6526 8370 6578
rect 11230 6526 11282 6578
rect 14478 6526 14530 6578
rect 18286 6526 18338 6578
rect 18622 6526 18674 6578
rect 19182 6526 19234 6578
rect 20078 6526 20130 6578
rect 24558 6526 24610 6578
rect 26014 6526 26066 6578
rect 6862 6414 6914 6466
rect 14030 6414 14082 6466
rect 14254 6414 14306 6466
rect 14590 6414 14642 6466
rect 14814 6414 14866 6466
rect 18398 6414 18450 6466
rect 18958 6414 19010 6466
rect 19966 6414 20018 6466
rect 24670 6414 24722 6466
rect 24782 6414 24834 6466
rect 25902 6414 25954 6466
rect 27806 6414 27858 6466
rect 29486 6414 29538 6466
rect 29710 6414 29762 6466
rect 30158 6414 30210 6466
rect 30830 6414 30882 6466
rect 31054 6414 31106 6466
rect 9782 6246 9834 6298
rect 9886 6246 9938 6298
rect 9990 6246 10042 6298
rect 18350 6246 18402 6298
rect 18454 6246 18506 6298
rect 18558 6246 18610 6298
rect 26918 6246 26970 6298
rect 27022 6246 27074 6298
rect 27126 6246 27178 6298
rect 35486 6246 35538 6298
rect 35590 6246 35642 6298
rect 35694 6246 35746 6298
rect 5742 6078 5794 6130
rect 20190 6078 20242 6130
rect 24222 6078 24274 6130
rect 24334 6078 24386 6130
rect 24558 6078 24610 6130
rect 26686 6078 26738 6130
rect 27022 6078 27074 6130
rect 28142 6078 28194 6130
rect 5966 5966 6018 6018
rect 9774 5966 9826 6018
rect 9886 5966 9938 6018
rect 10334 5966 10386 6018
rect 10782 5966 10834 6018
rect 11342 5966 11394 6018
rect 15486 5966 15538 6018
rect 20414 5966 20466 6018
rect 20526 5966 20578 6018
rect 25230 5966 25282 6018
rect 27918 5966 27970 6018
rect 29822 5966 29874 6018
rect 5630 5854 5682 5906
rect 8766 5854 8818 5906
rect 9550 5854 9602 5906
rect 10110 5854 10162 5906
rect 10446 5854 10498 5906
rect 11006 5854 11058 5906
rect 11790 5854 11842 5906
rect 15150 5854 15202 5906
rect 15374 5854 15426 5906
rect 15710 5854 15762 5906
rect 15822 5854 15874 5906
rect 16158 5854 16210 5906
rect 16494 5854 16546 5906
rect 17390 5854 17442 5906
rect 20862 5854 20914 5906
rect 24110 5854 24162 5906
rect 25454 5854 25506 5906
rect 25678 5854 25730 5906
rect 26126 5854 26178 5906
rect 26462 5854 26514 5906
rect 27246 5854 27298 5906
rect 27694 5854 27746 5906
rect 28478 5854 28530 5906
rect 29038 5854 29090 5906
rect 10894 5742 10946 5794
rect 12462 5742 12514 5794
rect 14590 5742 14642 5794
rect 16046 5742 16098 5794
rect 19070 5742 19122 5794
rect 25342 5742 25394 5794
rect 26574 5742 26626 5794
rect 27134 5742 27186 5794
rect 28030 5742 28082 5794
rect 31950 5742 32002 5794
rect 6638 5630 6690 5682
rect 21870 5630 21922 5682
rect 5498 5462 5550 5514
rect 5602 5462 5654 5514
rect 5706 5462 5758 5514
rect 14066 5462 14118 5514
rect 14170 5462 14222 5514
rect 14274 5462 14326 5514
rect 22634 5462 22686 5514
rect 22738 5462 22790 5514
rect 22842 5462 22894 5514
rect 31202 5462 31254 5514
rect 31306 5462 31358 5514
rect 31410 5462 31462 5514
rect 28030 5294 28082 5346
rect 29262 5294 29314 5346
rect 2270 5182 2322 5234
rect 6862 5182 6914 5234
rect 8990 5182 9042 5234
rect 10670 5182 10722 5234
rect 12798 5182 12850 5234
rect 13582 5182 13634 5234
rect 14590 5182 14642 5234
rect 18622 5182 18674 5234
rect 20750 5182 20802 5234
rect 22542 5182 22594 5234
rect 24670 5182 24722 5234
rect 25454 5182 25506 5234
rect 26350 5182 26402 5234
rect 28590 5182 28642 5234
rect 4622 5070 4674 5122
rect 6078 5070 6130 5122
rect 9886 5070 9938 5122
rect 13470 5070 13522 5122
rect 13806 5070 13858 5122
rect 14030 5070 14082 5122
rect 17502 5070 17554 5122
rect 17950 5070 18002 5122
rect 21758 5070 21810 5122
rect 24894 5070 24946 5122
rect 25790 5070 25842 5122
rect 27134 5070 27186 5122
rect 27470 5070 27522 5122
rect 27694 5070 27746 5122
rect 34638 5070 34690 5122
rect 35198 5070 35250 5122
rect 9326 4958 9378 5010
rect 9438 4958 9490 5010
rect 16718 4958 16770 5010
rect 25342 4958 25394 5010
rect 25566 4958 25618 5010
rect 26462 4958 26514 5010
rect 28142 4958 28194 5010
rect 29374 4958 29426 5010
rect 34862 4958 34914 5010
rect 9662 4846 9714 4898
rect 26238 4846 26290 4898
rect 27358 4846 27410 4898
rect 29822 4846 29874 4898
rect 9782 4678 9834 4730
rect 9886 4678 9938 4730
rect 9990 4678 10042 4730
rect 18350 4678 18402 4730
rect 18454 4678 18506 4730
rect 18558 4678 18610 4730
rect 26918 4678 26970 4730
rect 27022 4678 27074 4730
rect 27126 4678 27178 4730
rect 35486 4678 35538 4730
rect 35590 4678 35642 4730
rect 35694 4678 35746 4730
rect 17502 4510 17554 4562
rect 18622 4510 18674 4562
rect 18958 4510 19010 4562
rect 23214 4510 23266 4562
rect 24110 4510 24162 4562
rect 24558 4510 24610 4562
rect 31726 4510 31778 4562
rect 32174 4510 32226 4562
rect 6638 4398 6690 4450
rect 13358 4398 13410 4450
rect 16046 4398 16098 4450
rect 17950 4398 18002 4450
rect 18286 4398 18338 4450
rect 18398 4398 18450 4450
rect 20078 4398 20130 4450
rect 22654 4398 22706 4450
rect 22766 4398 22818 4450
rect 26014 4398 26066 4450
rect 30606 4398 30658 4450
rect 5294 4286 5346 4338
rect 5966 4286 6018 4338
rect 12462 4286 12514 4338
rect 12686 4286 12738 4338
rect 13022 4286 13074 4338
rect 16830 4286 16882 4338
rect 17278 4286 17330 4338
rect 17614 4286 17666 4338
rect 19294 4286 19346 4338
rect 25342 4286 25394 4338
rect 31278 4286 31330 4338
rect 3390 4174 3442 4226
rect 8766 4174 8818 4226
rect 9550 4174 9602 4226
rect 11678 4174 11730 4226
rect 12910 4174 12962 4226
rect 13918 4174 13970 4226
rect 22206 4174 22258 4226
rect 23774 4174 23826 4226
rect 24222 4174 24274 4226
rect 24670 4174 24722 4226
rect 28142 4174 28194 4226
rect 28478 4174 28530 4226
rect 31838 4174 31890 4226
rect 32286 4174 32338 4226
rect 33294 4174 33346 4226
rect 22654 4062 22706 4114
rect 5498 3894 5550 3946
rect 5602 3894 5654 3946
rect 5706 3894 5758 3946
rect 14066 3894 14118 3946
rect 14170 3894 14222 3946
rect 14274 3894 14326 3946
rect 22634 3894 22686 3946
rect 22738 3894 22790 3946
rect 22842 3894 22894 3946
rect 31202 3894 31254 3946
rect 31306 3894 31358 3946
rect 31410 3894 31462 3946
rect 12350 3614 12402 3666
rect 15934 3614 15986 3666
rect 18622 3614 18674 3666
rect 21870 3614 21922 3666
rect 25566 3614 25618 3666
rect 4510 3502 4562 3554
rect 5630 3502 5682 3554
rect 5966 3502 6018 3554
rect 8766 3502 8818 3554
rect 9214 3502 9266 3554
rect 9550 3502 9602 3554
rect 10446 3502 10498 3554
rect 13246 3502 13298 3554
rect 13582 3502 13634 3554
rect 14254 3502 14306 3554
rect 17054 3502 17106 3554
rect 17390 3502 17442 3554
rect 17614 3502 17666 3554
rect 20750 3502 20802 3554
rect 23774 3502 23826 3554
rect 24782 3502 24834 3554
rect 28702 3502 28754 3554
rect 29374 3502 29426 3554
rect 31054 3502 31106 3554
rect 32398 3502 32450 3554
rect 32958 3502 33010 3554
rect 33630 3502 33682 3554
rect 35086 3502 35138 3554
rect 5742 3390 5794 3442
rect 9438 3390 9490 3442
rect 13358 3390 13410 3442
rect 17166 3390 17218 3442
rect 23998 3390 24050 3442
rect 27470 3390 27522 3442
rect 27806 3390 27858 3442
rect 28366 3390 28418 3442
rect 29038 3390 29090 3442
rect 29822 3390 29874 3442
rect 30270 3390 30322 3442
rect 30606 3390 30658 3442
rect 31502 3390 31554 3442
rect 32174 3390 32226 3442
rect 34638 3390 34690 3442
rect 3950 3278 4002 3330
rect 7758 3278 7810 3330
rect 33406 3278 33458 3330
rect 34862 3278 34914 3330
rect 9782 3110 9834 3162
rect 9886 3110 9938 3162
rect 9990 3110 10042 3162
rect 18350 3110 18402 3162
rect 18454 3110 18506 3162
rect 18558 3110 18610 3162
rect 26918 3110 26970 3162
rect 27022 3110 27074 3162
rect 27126 3110 27178 3162
rect 35486 3110 35538 3162
rect 35590 3110 35642 3162
rect 35694 3110 35746 3162
<< metal2 >>
rect 1568 36200 1680 37000
rect 2688 36200 2800 37000
rect 3808 36200 3920 37000
rect 4928 36200 5040 37000
rect 6048 36200 6160 37000
rect 7168 36200 7280 37000
rect 8288 36200 8400 37000
rect 9408 36200 9520 37000
rect 10528 36200 10640 37000
rect 11648 36200 11760 37000
rect 12768 36200 12880 37000
rect 13888 36200 14000 37000
rect 15008 36200 15120 37000
rect 16128 36200 16240 37000
rect 17248 36200 17360 37000
rect 18368 36200 18480 37000
rect 19488 36200 19600 37000
rect 20608 36200 20720 37000
rect 21728 36200 21840 37000
rect 22848 36200 22960 37000
rect 23968 36200 24080 37000
rect 24332 36204 24724 36260
rect 1596 33236 1652 36200
rect 1820 33236 1876 33246
rect 1596 33234 1876 33236
rect 1596 33182 1822 33234
rect 1874 33182 1876 33234
rect 1596 33180 1876 33182
rect 2716 33236 2772 36200
rect 2940 33236 2996 33246
rect 2716 33234 2996 33236
rect 2716 33182 2942 33234
rect 2994 33182 2996 33234
rect 2716 33180 2996 33182
rect 3836 33236 3892 36200
rect 4060 33236 4116 33246
rect 3836 33234 4116 33236
rect 3836 33182 4062 33234
rect 4114 33182 4116 33234
rect 3836 33180 4116 33182
rect 1820 33170 1876 33180
rect 2940 33170 2996 33180
rect 4060 33170 4116 33180
rect 4956 33234 5012 36200
rect 5496 33740 5760 33750
rect 5552 33684 5600 33740
rect 5656 33684 5704 33740
rect 5496 33674 5760 33684
rect 4956 33182 4958 33234
rect 5010 33182 5012 33234
rect 4956 33170 5012 33182
rect 5852 33236 5908 33246
rect 6076 33236 6132 36200
rect 7196 33908 7252 36200
rect 7196 33852 7476 33908
rect 5852 33234 6132 33236
rect 5852 33182 5854 33234
rect 5906 33182 6132 33234
rect 5852 33180 6132 33182
rect 6412 33346 6468 33358
rect 6412 33294 6414 33346
rect 6466 33294 6468 33346
rect 5852 33170 5908 33180
rect 6188 32564 6244 32574
rect 6188 32562 6356 32564
rect 6188 32510 6190 32562
rect 6242 32510 6356 32562
rect 6188 32508 6356 32510
rect 6188 32498 6244 32508
rect 5496 32172 5760 32182
rect 5552 32116 5600 32172
rect 5656 32116 5704 32172
rect 5496 32106 5760 32116
rect 6300 31892 6356 32508
rect 6300 31826 6356 31836
rect 4396 30996 4452 31006
rect 3948 30994 4452 30996
rect 3948 30942 4398 30994
rect 4450 30942 4452 30994
rect 3948 30940 4452 30942
rect 3948 29428 4004 30940
rect 4396 30930 4452 30940
rect 5180 30882 5236 30894
rect 5180 30830 5182 30882
rect 5234 30830 5236 30882
rect 4620 29988 4676 29998
rect 4620 29538 4676 29932
rect 4620 29486 4622 29538
rect 4674 29486 4676 29538
rect 4620 29474 4676 29486
rect 3612 29426 4004 29428
rect 3612 29374 3950 29426
rect 4002 29374 4004 29426
rect 3612 29372 4004 29374
rect 3612 27858 3668 29372
rect 3948 29362 4004 29372
rect 5180 28868 5236 30830
rect 5496 30604 5760 30614
rect 5552 30548 5600 30604
rect 5656 30548 5704 30604
rect 5496 30538 5760 30548
rect 6412 30212 6468 33294
rect 6860 32452 6916 32462
rect 6860 32358 6916 32396
rect 6524 31892 6580 31902
rect 6580 31836 6692 31892
rect 6524 31826 6580 31836
rect 5740 30098 5796 30110
rect 5740 30046 5742 30098
rect 5794 30046 5796 30098
rect 5628 29988 5684 29998
rect 5628 29894 5684 29932
rect 5740 29540 5796 30046
rect 5740 29474 5796 29484
rect 5496 29036 5760 29046
rect 5552 28980 5600 29036
rect 5656 28980 5704 29036
rect 5496 28970 5760 28980
rect 5180 28802 5236 28812
rect 3612 27806 3614 27858
rect 3666 27806 3668 27858
rect 3612 26290 3668 27806
rect 4284 27746 4340 27758
rect 4284 27694 4286 27746
rect 4338 27694 4340 27746
rect 4284 27300 4340 27694
rect 5964 27748 6020 27758
rect 5496 27468 5760 27478
rect 5552 27412 5600 27468
rect 5656 27412 5704 27468
rect 5496 27402 5760 27412
rect 4284 27234 4340 27244
rect 5628 27300 5684 27310
rect 5628 27206 5684 27244
rect 5964 27298 6020 27692
rect 6412 27746 6468 30156
rect 6524 29986 6580 29998
rect 6524 29934 6526 29986
rect 6578 29934 6580 29986
rect 6524 29428 6580 29934
rect 6524 29362 6580 29372
rect 6524 28756 6580 28766
rect 6636 28756 6692 31836
rect 7420 31666 7476 33852
rect 8204 33572 8260 33582
rect 8204 33458 8260 33516
rect 8204 33406 8206 33458
rect 8258 33406 8260 33458
rect 8204 33394 8260 33406
rect 8316 32788 8372 36200
rect 8316 32722 8372 32732
rect 8988 33348 9044 33358
rect 7868 32452 7924 32462
rect 7924 32396 8148 32452
rect 7868 32386 7924 32396
rect 8092 32002 8148 32396
rect 8988 32450 9044 33292
rect 9436 33236 9492 36200
rect 10556 33572 10612 36200
rect 10556 33506 10612 33516
rect 9996 33348 10052 33358
rect 10052 33292 10164 33348
rect 9996 33254 10052 33292
rect 9548 33236 9604 33246
rect 9436 33234 9604 33236
rect 9436 33182 9550 33234
rect 9602 33182 9604 33234
rect 9436 33180 9604 33182
rect 9548 33170 9604 33180
rect 9780 32956 10044 32966
rect 9836 32900 9884 32956
rect 9940 32900 9988 32956
rect 9780 32890 10044 32900
rect 9548 32788 9604 32798
rect 9548 32694 9604 32732
rect 8988 32398 8990 32450
rect 9042 32398 9044 32450
rect 8988 32386 9044 32398
rect 8092 31950 8094 32002
rect 8146 31950 8148 32002
rect 8092 31938 8148 31950
rect 8652 31892 8708 31902
rect 7420 31614 7422 31666
rect 7474 31614 7476 31666
rect 7420 31602 7476 31614
rect 8092 31780 8148 31790
rect 8652 31780 8708 31836
rect 7644 31108 7700 31118
rect 7532 31106 7700 31108
rect 7532 31054 7646 31106
rect 7698 31054 7700 31106
rect 7532 31052 7700 31054
rect 7308 30996 7364 31006
rect 7308 30882 7364 30940
rect 7308 30830 7310 30882
rect 7362 30830 7364 30882
rect 7308 30818 7364 30830
rect 7084 30212 7140 30222
rect 7084 30118 7140 30156
rect 6748 29988 6804 29998
rect 7308 29988 7364 29998
rect 6748 29986 6916 29988
rect 6748 29934 6750 29986
rect 6802 29934 6916 29986
rect 6748 29932 6916 29934
rect 6748 29922 6804 29932
rect 6748 29764 6804 29774
rect 6748 29314 6804 29708
rect 6860 29428 6916 29932
rect 7196 29428 7252 29438
rect 6860 29426 7252 29428
rect 6860 29374 7198 29426
rect 7250 29374 7252 29426
rect 6860 29372 7252 29374
rect 7196 29362 7252 29372
rect 6748 29262 6750 29314
rect 6802 29262 6804 29314
rect 6748 29250 6804 29262
rect 7308 29092 7364 29932
rect 7532 29428 7588 31052
rect 7644 31042 7700 31052
rect 7980 30996 8036 31006
rect 7980 30902 8036 30940
rect 7868 29986 7924 29998
rect 7868 29934 7870 29986
rect 7922 29934 7924 29986
rect 7868 29652 7924 29934
rect 7532 29362 7588 29372
rect 7644 29596 7868 29652
rect 7644 29426 7700 29596
rect 7868 29586 7924 29596
rect 8092 29540 8148 31724
rect 8428 31778 8708 31780
rect 8428 31726 8654 31778
rect 8706 31726 8708 31778
rect 8428 31724 8708 31726
rect 8204 31668 8260 31678
rect 8204 31574 8260 31612
rect 8428 31218 8484 31724
rect 8652 31714 8708 31724
rect 8428 31166 8430 31218
rect 8482 31166 8484 31218
rect 8428 31154 8484 31166
rect 9212 31668 9268 31678
rect 9212 30322 9268 31612
rect 9324 31668 9380 31678
rect 9324 31666 9604 31668
rect 9324 31614 9326 31666
rect 9378 31614 9604 31666
rect 9324 31612 9604 31614
rect 9324 31602 9380 31612
rect 9548 31218 9604 31612
rect 9780 31388 10044 31398
rect 9836 31332 9884 31388
rect 9940 31332 9988 31388
rect 9780 31322 10044 31332
rect 9548 31166 9550 31218
rect 9602 31166 9604 31218
rect 9548 31154 9604 31166
rect 10108 30996 10164 33292
rect 10220 32450 10276 32462
rect 10220 32398 10222 32450
rect 10274 32398 10276 32450
rect 10220 31892 10276 32398
rect 10220 31826 10276 31836
rect 11452 31892 11508 31902
rect 11452 31890 11620 31892
rect 11452 31838 11454 31890
rect 11506 31838 11620 31890
rect 11452 31836 11620 31838
rect 11452 31826 11508 31836
rect 9772 30994 10164 30996
rect 9772 30942 10110 30994
rect 10162 30942 10164 30994
rect 9772 30940 10164 30942
rect 9660 30882 9716 30894
rect 9660 30830 9662 30882
rect 9714 30830 9716 30882
rect 9212 30270 9214 30322
rect 9266 30270 9268 30322
rect 9212 30258 9268 30270
rect 9548 30324 9604 30334
rect 9324 30210 9380 30222
rect 9324 30158 9326 30210
rect 9378 30158 9380 30210
rect 8204 30100 8260 30110
rect 9324 30100 9380 30158
rect 9548 30210 9604 30268
rect 9548 30158 9550 30210
rect 9602 30158 9604 30210
rect 9548 30146 9604 30158
rect 8204 29764 8260 30044
rect 9212 30044 9380 30100
rect 8204 29698 8260 29708
rect 8316 29988 8372 29998
rect 7980 29484 8148 29540
rect 8316 29540 8372 29932
rect 8988 29988 9044 29998
rect 9212 29988 9268 30044
rect 8988 29986 9268 29988
rect 8988 29934 8990 29986
rect 9042 29934 9268 29986
rect 8988 29932 9268 29934
rect 8988 29922 9044 29932
rect 9212 29764 9268 29932
rect 9212 29698 9268 29708
rect 9548 29764 9604 29774
rect 8876 29652 8932 29662
rect 8876 29558 8932 29596
rect 8428 29540 8484 29550
rect 8316 29538 8484 29540
rect 8316 29486 8430 29538
rect 8482 29486 8484 29538
rect 8316 29484 8484 29486
rect 7644 29374 7646 29426
rect 7698 29374 7700 29426
rect 7644 29362 7700 29374
rect 7756 29428 7812 29438
rect 7084 29036 7364 29092
rect 6860 28868 6916 28878
rect 6860 28774 6916 28812
rect 6524 28754 6636 28756
rect 6524 28702 6526 28754
rect 6578 28702 6636 28754
rect 6524 28700 6636 28702
rect 6524 28690 6580 28700
rect 6636 28662 6692 28700
rect 6860 28644 6916 28654
rect 6860 28550 6916 28588
rect 7084 28082 7140 29036
rect 7196 28924 7588 28980
rect 7196 28866 7252 28924
rect 7196 28814 7198 28866
rect 7250 28814 7252 28866
rect 7196 28802 7252 28814
rect 7084 28030 7086 28082
rect 7138 28030 7140 28082
rect 7084 28018 7140 28030
rect 7308 28756 7364 28766
rect 6412 27694 6414 27746
rect 6466 27694 6468 27746
rect 6412 27682 6468 27694
rect 6860 27858 6916 27870
rect 6860 27806 6862 27858
rect 6914 27806 6916 27858
rect 6524 27636 6580 27646
rect 5964 27246 5966 27298
rect 6018 27246 6020 27298
rect 5964 27234 6020 27246
rect 6300 27412 6356 27422
rect 6300 27074 6356 27356
rect 6300 27022 6302 27074
rect 6354 27022 6356 27074
rect 6300 27010 6356 27022
rect 6524 27074 6580 27580
rect 6860 27412 6916 27806
rect 6972 27748 7028 27758
rect 6972 27654 7028 27692
rect 7196 27412 7252 27422
rect 6860 27356 7196 27412
rect 6972 27188 7028 27198
rect 6524 27022 6526 27074
rect 6578 27022 6580 27074
rect 6524 27010 6580 27022
rect 6860 27076 6916 27086
rect 6860 26908 6916 27020
rect 5740 26850 5796 26862
rect 5740 26798 5742 26850
rect 5794 26798 5796 26850
rect 5740 26516 5796 26798
rect 5740 26450 5796 26460
rect 6412 26850 6468 26862
rect 6412 26798 6414 26850
rect 6466 26798 6468 26850
rect 3612 26238 3614 26290
rect 3666 26238 3668 26290
rect 3612 25284 3668 26238
rect 4396 26180 4452 26190
rect 4396 26086 4452 26124
rect 6188 26180 6244 26190
rect 5496 25900 5760 25910
rect 5552 25844 5600 25900
rect 5656 25844 5704 25900
rect 5496 25834 5760 25844
rect 6188 25730 6244 26124
rect 6188 25678 6190 25730
rect 6242 25678 6244 25730
rect 6188 25666 6244 25678
rect 6412 25732 6468 26798
rect 6524 26852 6916 26908
rect 6972 27074 7028 27132
rect 6972 27022 6974 27074
rect 7026 27022 7028 27074
rect 6524 26178 6580 26852
rect 6524 26126 6526 26178
rect 6578 26126 6580 26178
rect 6524 26114 6580 26126
rect 6860 26628 6916 26638
rect 6524 25732 6580 25742
rect 6412 25730 6580 25732
rect 6412 25678 6526 25730
rect 6578 25678 6580 25730
rect 6412 25676 6580 25678
rect 6524 25666 6580 25676
rect 6300 25396 6356 25406
rect 6300 25302 6356 25340
rect 3612 25218 3668 25228
rect 6860 25284 6916 26572
rect 6972 25730 7028 27022
rect 7196 27074 7252 27356
rect 7196 27022 7198 27074
rect 7250 27022 7252 27074
rect 7196 27010 7252 27022
rect 7308 26628 7364 28700
rect 7420 28084 7476 28094
rect 7420 27858 7476 28028
rect 7420 27806 7422 27858
rect 7474 27806 7476 27858
rect 7420 27188 7476 27806
rect 7420 27122 7476 27132
rect 7532 27186 7588 28924
rect 7644 28756 7700 28766
rect 7644 28662 7700 28700
rect 7756 28532 7812 29372
rect 7532 27134 7534 27186
rect 7586 27134 7588 27186
rect 7532 27122 7588 27134
rect 7644 28476 7812 28532
rect 7420 26852 7476 26862
rect 7420 26850 7588 26852
rect 7420 26798 7422 26850
rect 7474 26798 7588 26850
rect 7420 26796 7588 26798
rect 7420 26786 7476 26796
rect 7308 26562 7364 26572
rect 7420 26404 7476 26414
rect 7420 26310 7476 26348
rect 7532 26402 7588 26796
rect 7644 26850 7700 28476
rect 7868 27860 7924 27870
rect 7980 27860 8036 29484
rect 8092 29316 8148 29326
rect 8092 29314 8372 29316
rect 8092 29262 8094 29314
rect 8146 29262 8372 29314
rect 8092 29260 8372 29262
rect 8092 29250 8148 29260
rect 8316 28642 8372 29260
rect 8316 28590 8318 28642
rect 8370 28590 8372 28642
rect 8316 28578 8372 28590
rect 7868 27858 8036 27860
rect 7868 27806 7870 27858
rect 7922 27806 8036 27858
rect 7868 27804 8036 27806
rect 8092 27970 8148 27982
rect 8092 27918 8094 27970
rect 8146 27918 8148 27970
rect 7868 27076 7924 27804
rect 8092 27636 8148 27918
rect 8092 27570 8148 27580
rect 8428 27524 8484 29484
rect 8652 29428 8708 29438
rect 9324 29428 9380 29438
rect 8652 29334 8708 29372
rect 9100 29372 9324 29428
rect 8988 29204 9044 29214
rect 8988 29110 9044 29148
rect 8764 28980 8820 28990
rect 8652 28530 8708 28542
rect 8652 28478 8654 28530
rect 8706 28478 8708 28530
rect 8540 28418 8596 28430
rect 8540 28366 8542 28418
rect 8594 28366 8596 28418
rect 8540 28308 8596 28366
rect 8540 28242 8596 28252
rect 8540 28084 8596 28094
rect 8540 27990 8596 28028
rect 8428 27468 8596 27524
rect 8540 27076 8596 27468
rect 7868 27010 7924 27020
rect 7980 27020 8484 27076
rect 7980 26908 8036 27020
rect 7644 26798 7646 26850
rect 7698 26798 7700 26850
rect 7644 26628 7700 26798
rect 7756 26852 8036 26908
rect 8428 26962 8484 27020
rect 8540 26982 8596 27020
rect 8428 26910 8430 26962
rect 8482 26910 8484 26962
rect 8428 26898 8484 26910
rect 7756 26850 7812 26852
rect 7756 26798 7758 26850
rect 7810 26798 7812 26850
rect 7756 26786 7812 26798
rect 7644 26562 7700 26572
rect 7868 26740 7924 26750
rect 7532 26350 7534 26402
rect 7586 26350 7588 26402
rect 7532 26338 7588 26350
rect 7644 26404 7700 26414
rect 7644 26402 7812 26404
rect 7644 26350 7646 26402
rect 7698 26350 7812 26402
rect 7644 26348 7812 26350
rect 7644 26338 7700 26348
rect 6972 25678 6974 25730
rect 7026 25678 7028 25730
rect 6972 25666 7028 25678
rect 7084 26290 7140 26302
rect 7084 26238 7086 26290
rect 7138 26238 7140 26290
rect 6972 25284 7028 25294
rect 6916 25282 7028 25284
rect 6916 25230 6974 25282
rect 7026 25230 7028 25282
rect 6916 25228 7028 25230
rect 6748 24834 6804 24846
rect 6748 24782 6750 24834
rect 6802 24782 6804 24834
rect 6636 24724 6692 24734
rect 6636 24630 6692 24668
rect 5496 24332 5760 24342
rect 5552 24276 5600 24332
rect 5656 24276 5704 24332
rect 5496 24266 5760 24276
rect 6748 23940 6804 24782
rect 6636 23884 6804 23940
rect 6636 23492 6692 23884
rect 6748 23716 6804 23726
rect 6860 23716 6916 25228
rect 6972 25218 7028 25228
rect 6972 24948 7028 24958
rect 7084 24948 7140 26238
rect 7420 25730 7476 25742
rect 7420 25678 7422 25730
rect 7474 25678 7476 25730
rect 7420 25618 7476 25678
rect 7420 25566 7422 25618
rect 7474 25566 7476 25618
rect 7420 25554 7476 25566
rect 7756 25506 7812 26348
rect 7756 25454 7758 25506
rect 7810 25454 7812 25506
rect 7756 25442 7812 25454
rect 7868 25284 7924 26684
rect 7980 26402 8036 26852
rect 8316 26850 8372 26862
rect 8316 26798 8318 26850
rect 8370 26798 8372 26850
rect 8316 26740 8372 26798
rect 8316 26684 8596 26740
rect 8204 26628 8260 26638
rect 7980 26350 7982 26402
rect 8034 26350 8036 26402
rect 7980 26338 8036 26350
rect 8092 26572 8204 26628
rect 8092 26068 8148 26572
rect 8204 26562 8260 26572
rect 8540 26628 8596 26684
rect 8540 26562 8596 26572
rect 8428 26516 8484 26526
rect 8428 26422 8484 26460
rect 7980 26012 8148 26068
rect 8204 26404 8260 26414
rect 7980 25394 8036 26012
rect 7980 25342 7982 25394
rect 8034 25342 8036 25394
rect 7980 25330 8036 25342
rect 8092 25394 8148 25406
rect 8092 25342 8094 25394
rect 8146 25342 8148 25394
rect 6972 24946 7140 24948
rect 6972 24894 6974 24946
rect 7026 24894 7140 24946
rect 6972 24892 7140 24894
rect 7532 25228 7924 25284
rect 8092 25284 8148 25342
rect 7532 24946 7588 25228
rect 8092 25218 8148 25228
rect 8204 25060 8260 26348
rect 7532 24894 7534 24946
rect 7586 24894 7588 24946
rect 6972 24882 7028 24892
rect 7532 24882 7588 24894
rect 8092 25004 8260 25060
rect 8316 26290 8372 26302
rect 8316 26238 8318 26290
rect 8370 26238 8372 26290
rect 8092 24946 8148 25004
rect 8316 24948 8372 26238
rect 8540 26290 8596 26302
rect 8540 26238 8542 26290
rect 8594 26238 8596 26290
rect 8540 25956 8596 26238
rect 8540 25890 8596 25900
rect 8092 24894 8094 24946
rect 8146 24894 8148 24946
rect 8092 24882 8148 24894
rect 8204 24892 8372 24948
rect 8652 24946 8708 28478
rect 8764 28084 8820 28924
rect 9100 28754 9156 29372
rect 9324 29362 9380 29372
rect 9548 29426 9604 29708
rect 9548 29374 9550 29426
rect 9602 29374 9604 29426
rect 9548 29316 9604 29374
rect 9548 29250 9604 29260
rect 9660 29204 9716 30830
rect 9772 30098 9828 30940
rect 10108 30930 10164 30940
rect 10220 31106 10276 31118
rect 10220 31054 10222 31106
rect 10274 31054 10276 31106
rect 9772 30046 9774 30098
rect 9826 30046 9828 30098
rect 9772 30034 9828 30046
rect 9996 29988 10052 30026
rect 9996 29922 10052 29932
rect 9780 29820 10044 29830
rect 9836 29764 9884 29820
rect 9940 29764 9988 29820
rect 9780 29754 10044 29764
rect 10108 29652 10164 29662
rect 10220 29652 10276 31054
rect 11340 31106 11396 31118
rect 11340 31054 11342 31106
rect 11394 31054 11396 31106
rect 10444 30996 10500 31006
rect 10444 30210 10500 30940
rect 10444 30158 10446 30210
rect 10498 30158 10500 30210
rect 10444 30146 10500 30158
rect 10668 30994 10724 31006
rect 10668 30942 10670 30994
rect 10722 30942 10724 30994
rect 10668 30212 10724 30942
rect 10668 30146 10724 30156
rect 11116 30770 11172 30782
rect 11116 30718 11118 30770
rect 11170 30718 11172 30770
rect 10892 29988 10948 29998
rect 10948 29932 11060 29988
rect 10892 29922 10948 29932
rect 10164 29596 10276 29652
rect 10332 29876 10388 29886
rect 10332 29650 10388 29820
rect 10332 29598 10334 29650
rect 10386 29598 10388 29650
rect 10108 29558 10164 29596
rect 9996 29540 10052 29550
rect 9884 29428 9940 29438
rect 9884 29334 9940 29372
rect 9996 29314 10052 29484
rect 9996 29262 9998 29314
rect 10050 29262 10052 29314
rect 9996 29250 10052 29262
rect 9660 29148 9940 29204
rect 9100 28702 9102 28754
rect 9154 28702 9156 28754
rect 9100 28690 9156 28702
rect 9324 28980 9380 28990
rect 8988 28642 9044 28654
rect 8988 28590 8990 28642
rect 9042 28590 9044 28642
rect 8988 28532 9044 28590
rect 9324 28532 9380 28924
rect 9884 28754 9940 29148
rect 9884 28702 9886 28754
rect 9938 28702 9940 28754
rect 9884 28690 9940 28702
rect 10332 28756 10388 29598
rect 10892 29314 10948 29326
rect 10892 29262 10894 29314
rect 10946 29262 10948 29314
rect 10780 29204 10836 29214
rect 10332 28700 10724 28756
rect 9436 28642 9492 28654
rect 9436 28590 9438 28642
rect 9490 28590 9492 28642
rect 9436 28532 9492 28590
rect 10220 28644 10276 28654
rect 10332 28644 10388 28700
rect 10220 28642 10388 28644
rect 10220 28590 10222 28642
rect 10274 28590 10388 28642
rect 10220 28588 10388 28590
rect 10220 28578 10276 28588
rect 9884 28532 9940 28542
rect 8988 28476 9156 28532
rect 9324 28476 9492 28532
rect 9772 28530 9940 28532
rect 9772 28478 9886 28530
rect 9938 28478 9940 28530
rect 9772 28476 9940 28478
rect 8764 28018 8820 28028
rect 9100 27972 9156 28476
rect 9772 28420 9828 28476
rect 9884 28466 9940 28476
rect 9996 28532 10052 28542
rect 10052 28476 10164 28532
rect 9996 28438 10052 28476
rect 9660 28364 9828 28420
rect 9324 28308 9380 28318
rect 9380 28252 9492 28308
rect 9324 28242 9380 28252
rect 9100 27906 9156 27916
rect 8988 27860 9044 27870
rect 9436 27860 9492 28252
rect 9548 27860 9604 27870
rect 8988 27074 9044 27804
rect 8988 27022 8990 27074
rect 9042 27022 9044 27074
rect 8988 27010 9044 27022
rect 9324 27858 9604 27860
rect 9324 27806 9550 27858
rect 9602 27806 9604 27858
rect 9324 27804 9604 27806
rect 9324 26908 9380 27804
rect 9548 27794 9604 27804
rect 9548 27298 9604 27310
rect 9548 27246 9550 27298
rect 9602 27246 9604 27298
rect 9324 26852 9492 26908
rect 9436 26292 9492 26852
rect 9548 26514 9604 27246
rect 9548 26462 9550 26514
rect 9602 26462 9604 26514
rect 9548 26450 9604 26462
rect 9660 26514 9716 28364
rect 9780 28252 10044 28262
rect 9836 28196 9884 28252
rect 9940 28196 9988 28252
rect 9780 28186 10044 28196
rect 9772 27970 9828 27982
rect 9772 27918 9774 27970
rect 9826 27918 9828 27970
rect 9772 27188 9828 27918
rect 9996 27858 10052 27870
rect 9996 27806 9998 27858
rect 10050 27806 10052 27858
rect 9884 27748 9940 27758
rect 9884 27654 9940 27692
rect 9884 27188 9940 27198
rect 9772 27132 9884 27188
rect 9884 27094 9940 27132
rect 9996 26908 10052 27806
rect 10108 27076 10164 28476
rect 10556 28530 10612 28542
rect 10556 28478 10558 28530
rect 10610 28478 10612 28530
rect 10108 26982 10164 27020
rect 10332 27972 10388 27982
rect 10332 27858 10388 27916
rect 10332 27806 10334 27858
rect 10386 27806 10388 27858
rect 10332 27300 10388 27806
rect 9884 26852 10052 26908
rect 9884 26786 9940 26796
rect 9780 26684 10044 26694
rect 9836 26628 9884 26684
rect 9940 26628 9988 26684
rect 9780 26618 10044 26628
rect 9660 26462 9662 26514
rect 9714 26462 9716 26514
rect 9660 26450 9716 26462
rect 9772 26516 9828 26526
rect 9772 26422 9828 26460
rect 9884 26404 9940 26414
rect 9884 26310 9940 26348
rect 9436 26226 9492 26236
rect 10332 26290 10388 27244
rect 10556 26908 10612 28478
rect 10668 28082 10724 28700
rect 10780 28642 10836 29148
rect 10892 28980 10948 29262
rect 10892 28914 10948 28924
rect 11004 28754 11060 29932
rect 11116 29652 11172 30718
rect 11116 29586 11172 29596
rect 11228 30772 11284 30782
rect 11228 29428 11284 30716
rect 11004 28702 11006 28754
rect 11058 28702 11060 28754
rect 11004 28690 11060 28702
rect 11116 29426 11284 29428
rect 11116 29374 11230 29426
rect 11282 29374 11284 29426
rect 11116 29372 11284 29374
rect 10780 28590 10782 28642
rect 10834 28590 10836 28642
rect 10780 28578 10836 28590
rect 10668 28030 10670 28082
rect 10722 28030 10724 28082
rect 10668 28018 10724 28030
rect 10892 27860 10948 27870
rect 10892 27766 10948 27804
rect 10892 27636 10948 27646
rect 11116 27636 11172 29372
rect 11228 29362 11284 29372
rect 11340 29426 11396 31054
rect 11564 30996 11620 31836
rect 11676 31556 11732 36200
rect 12348 33572 12404 33582
rect 12348 33478 12404 33516
rect 12796 32788 12852 36200
rect 13916 33572 13972 36200
rect 14064 33740 14328 33750
rect 14120 33684 14168 33740
rect 14224 33684 14272 33740
rect 14064 33674 14328 33684
rect 13916 33506 13972 33516
rect 12572 32732 12852 32788
rect 13244 33346 13300 33358
rect 13244 33294 13246 33346
rect 13298 33294 13300 33346
rect 12460 32562 12516 32574
rect 12460 32510 12462 32562
rect 12514 32510 12516 32562
rect 11900 31892 11956 31902
rect 11900 31798 11956 31836
rect 12124 31556 12180 31566
rect 11676 31500 11844 31556
rect 11564 30902 11620 30940
rect 11788 30434 11844 31500
rect 12124 30994 12180 31500
rect 12460 31556 12516 32510
rect 12460 31490 12516 31500
rect 12124 30942 12126 30994
rect 12178 30942 12180 30994
rect 12124 30930 12180 30942
rect 11788 30382 11790 30434
rect 11842 30382 11844 30434
rect 11788 30370 11844 30382
rect 12572 30436 12628 32732
rect 13132 32452 13188 32462
rect 12572 30370 12628 30380
rect 12684 32450 13188 32452
rect 12684 32398 13134 32450
rect 13186 32398 13188 32450
rect 12684 32396 13188 32398
rect 12572 30212 12628 30222
rect 11452 29652 11508 29662
rect 11452 29538 11508 29596
rect 12572 29652 12628 30156
rect 12572 29558 12628 29596
rect 11452 29486 11454 29538
rect 11506 29486 11508 29538
rect 11452 29474 11508 29486
rect 12236 29538 12292 29550
rect 12236 29486 12238 29538
rect 12290 29486 12292 29538
rect 11340 29374 11342 29426
rect 11394 29374 11396 29426
rect 11228 28868 11284 28878
rect 11228 28642 11284 28812
rect 11228 28590 11230 28642
rect 11282 28590 11284 28642
rect 11228 28578 11284 28590
rect 11340 28532 11396 29374
rect 11564 29204 11620 29214
rect 11564 28754 11620 29148
rect 11900 29202 11956 29214
rect 11900 29150 11902 29202
rect 11954 29150 11956 29202
rect 11564 28702 11566 28754
rect 11618 28702 11620 28754
rect 11564 28690 11620 28702
rect 11788 28756 11844 28766
rect 11340 28466 11396 28476
rect 11788 28084 11844 28700
rect 10948 27580 11172 27636
rect 11452 28028 11844 28084
rect 10892 27074 10948 27580
rect 11452 27188 11508 28028
rect 11900 27972 11956 29150
rect 12236 28756 12292 29486
rect 12684 29204 12740 32396
rect 13132 32386 13188 32396
rect 13244 31556 13300 33294
rect 13916 33236 13972 33246
rect 13244 31490 13300 31500
rect 13580 33234 13972 33236
rect 13580 33182 13918 33234
rect 13970 33182 13972 33234
rect 13580 33180 13972 33182
rect 12236 28690 12292 28700
rect 12572 29148 12740 29204
rect 12796 30882 12852 30894
rect 12796 30830 12798 30882
rect 12850 30830 12852 30882
rect 12460 28644 12516 28654
rect 10892 27022 10894 27074
rect 10946 27022 10948 27074
rect 10892 27010 10948 27022
rect 11004 27076 11060 27086
rect 11004 26982 11060 27020
rect 11452 27074 11508 27132
rect 11452 27022 11454 27074
rect 11506 27022 11508 27074
rect 11452 27010 11508 27022
rect 11788 27970 11956 27972
rect 11788 27918 11902 27970
rect 11954 27918 11956 27970
rect 11788 27916 11956 27918
rect 11788 26908 11844 27916
rect 11900 27906 11956 27916
rect 12012 27970 12068 27982
rect 12012 27918 12014 27970
rect 12066 27918 12068 27970
rect 12012 27860 12068 27918
rect 12012 27794 12068 27804
rect 12460 27858 12516 28588
rect 12572 28196 12628 29148
rect 12796 28754 12852 30830
rect 13580 30210 13636 33180
rect 13916 33170 13972 33180
rect 14064 32172 14328 32182
rect 14120 32116 14168 32172
rect 14224 32116 14272 32172
rect 14064 32106 14328 32116
rect 14588 31780 14644 31790
rect 14588 31686 14644 31724
rect 13804 31556 13860 31566
rect 14252 31556 14308 31566
rect 13860 31554 14532 31556
rect 13860 31502 14254 31554
rect 14306 31502 14532 31554
rect 13860 31500 14532 31502
rect 13804 31462 13860 31500
rect 14252 31490 14308 31500
rect 14064 30604 14328 30614
rect 14120 30548 14168 30604
rect 14224 30548 14272 30604
rect 14064 30538 14328 30548
rect 13580 30158 13582 30210
rect 13634 30158 13636 30210
rect 13580 30146 13636 30158
rect 14028 30436 14084 30446
rect 13020 30100 13076 30110
rect 13020 29426 13076 30044
rect 13020 29374 13022 29426
rect 13074 29374 13076 29426
rect 13020 29362 13076 29374
rect 13468 30098 13524 30110
rect 13468 30046 13470 30098
rect 13522 30046 13524 30098
rect 12796 28702 12798 28754
rect 12850 28702 12852 28754
rect 12796 28690 12852 28702
rect 13468 28756 13524 30046
rect 14028 29650 14084 30380
rect 14252 29986 14308 29998
rect 14252 29934 14254 29986
rect 14306 29934 14308 29986
rect 14252 29876 14308 29934
rect 14476 29876 14532 31500
rect 14588 30996 14644 31006
rect 14588 30210 14644 30940
rect 14924 30884 14980 30894
rect 14588 30158 14590 30210
rect 14642 30158 14644 30210
rect 14588 30146 14644 30158
rect 14812 30828 14924 30884
rect 14252 29820 14532 29876
rect 14028 29598 14030 29650
rect 14082 29598 14084 29650
rect 14028 29586 14084 29598
rect 14064 29036 14328 29046
rect 14120 28980 14168 29036
rect 14224 28980 14272 29036
rect 14064 28970 14328 28980
rect 13580 28756 13636 28766
rect 13468 28754 13636 28756
rect 13468 28702 13582 28754
rect 13634 28702 13636 28754
rect 13468 28700 13636 28702
rect 13580 28690 13636 28700
rect 12684 28644 12740 28654
rect 12684 28530 12740 28588
rect 14252 28642 14308 28654
rect 14252 28590 14254 28642
rect 14306 28590 14308 28642
rect 12684 28478 12686 28530
rect 12738 28478 12740 28530
rect 12684 28466 12740 28478
rect 12908 28532 12964 28542
rect 13804 28532 13860 28542
rect 12908 28530 13300 28532
rect 12908 28478 12910 28530
rect 12962 28478 13300 28530
rect 12908 28476 13300 28478
rect 12908 28466 12964 28476
rect 12572 28140 12740 28196
rect 12684 28082 12740 28140
rect 12684 28030 12686 28082
rect 12738 28030 12740 28082
rect 12684 28018 12740 28030
rect 12460 27806 12462 27858
rect 12514 27806 12516 27858
rect 12460 27794 12516 27806
rect 13132 27858 13188 27870
rect 13132 27806 13134 27858
rect 13186 27806 13188 27858
rect 12012 27634 12068 27646
rect 12012 27582 12014 27634
rect 12066 27582 12068 27634
rect 10556 26852 10836 26908
rect 10780 26628 10836 26852
rect 11228 26852 11284 26862
rect 11564 26852 11844 26908
rect 11900 27300 11956 27310
rect 11900 26962 11956 27244
rect 11900 26910 11902 26962
rect 11954 26910 11956 26962
rect 11900 26898 11956 26910
rect 12012 26908 12068 27582
rect 12796 27636 12852 27646
rect 12796 27542 12852 27580
rect 12908 27412 12964 27422
rect 12236 27132 12628 27188
rect 12236 27074 12292 27132
rect 12236 27022 12238 27074
rect 12290 27022 12292 27074
rect 12236 27010 12292 27022
rect 12572 27076 12628 27132
rect 12572 26982 12628 27020
rect 12348 26964 12404 26974
rect 12012 26852 12180 26908
rect 11228 26850 11396 26852
rect 11228 26798 11230 26850
rect 11282 26798 11396 26850
rect 11228 26796 11396 26798
rect 11228 26786 11284 26796
rect 10332 26238 10334 26290
rect 10386 26238 10388 26290
rect 10332 26226 10388 26238
rect 10668 26572 10780 26628
rect 10444 26068 10500 26078
rect 9884 25956 9940 25966
rect 9884 25506 9940 25900
rect 10444 25730 10500 26012
rect 10444 25678 10446 25730
rect 10498 25678 10500 25730
rect 10444 25666 10500 25678
rect 9884 25454 9886 25506
rect 9938 25454 9940 25506
rect 9884 25442 9940 25454
rect 10668 25506 10724 26572
rect 10780 26562 10836 26572
rect 11340 26290 11396 26796
rect 11340 26238 11342 26290
rect 11394 26238 11396 26290
rect 11340 26226 11396 26238
rect 11564 26404 11620 26852
rect 11564 26290 11620 26348
rect 11564 26238 11566 26290
rect 11618 26238 11620 26290
rect 11564 26226 11620 26238
rect 12124 26290 12180 26852
rect 12124 26238 12126 26290
rect 12178 26238 12180 26290
rect 12124 26180 12180 26238
rect 10668 25454 10670 25506
rect 10722 25454 10724 25506
rect 10668 25442 10724 25454
rect 11788 26066 11844 26078
rect 11788 26014 11790 26066
rect 11842 26014 11844 26066
rect 10108 25394 10164 25406
rect 10108 25342 10110 25394
rect 10162 25342 10164 25394
rect 9780 25116 10044 25126
rect 9836 25060 9884 25116
rect 9940 25060 9988 25116
rect 9780 25050 10044 25060
rect 8652 24894 8654 24946
rect 8706 24894 8708 24946
rect 7308 24836 7364 24846
rect 7868 24836 7924 24846
rect 7308 24834 7476 24836
rect 7308 24782 7310 24834
rect 7362 24782 7476 24834
rect 7308 24780 7476 24782
rect 7308 24770 7364 24780
rect 7196 24724 7252 24734
rect 7196 24630 7252 24668
rect 7420 24052 7476 24780
rect 7868 24834 8036 24836
rect 7868 24782 7870 24834
rect 7922 24782 8036 24834
rect 7868 24780 8036 24782
rect 7868 24770 7924 24780
rect 7756 24724 7812 24734
rect 7756 24630 7812 24668
rect 7196 23996 7476 24052
rect 7196 23826 7252 23996
rect 7196 23774 7198 23826
rect 7250 23774 7252 23826
rect 6804 23660 6916 23716
rect 6972 23716 7028 23726
rect 6972 23714 7140 23716
rect 6972 23662 6974 23714
rect 7026 23662 7140 23714
rect 6972 23660 7140 23662
rect 6748 23622 6804 23660
rect 6972 23650 7028 23660
rect 6972 23492 7028 23502
rect 6636 23436 6804 23492
rect 3948 23154 4004 23166
rect 3948 23102 3950 23154
rect 4002 23102 4004 23154
rect 3724 21588 3780 21598
rect 3948 21588 4004 23102
rect 4732 23044 4788 23054
rect 4732 22950 4788 22988
rect 5496 22764 5760 22774
rect 5552 22708 5600 22764
rect 5656 22708 5704 22764
rect 5496 22698 5760 22708
rect 6524 22258 6580 22270
rect 6524 22206 6526 22258
rect 6578 22206 6580 22258
rect 4396 22148 4452 22158
rect 4396 21698 4452 22092
rect 4396 21646 4398 21698
rect 4450 21646 4452 21698
rect 4396 21634 4452 21646
rect 6524 21700 6580 22206
rect 6636 22148 6692 22158
rect 6636 22054 6692 22092
rect 6748 21812 6804 23436
rect 6860 23436 6972 23492
rect 6860 23042 6916 23436
rect 6972 23426 7028 23436
rect 7084 23154 7140 23660
rect 7084 23102 7086 23154
rect 7138 23102 7140 23154
rect 7084 23090 7140 23102
rect 6860 22990 6862 23042
rect 6914 22990 6916 23042
rect 6860 22978 6916 22990
rect 7084 22596 7140 22606
rect 7084 22370 7140 22540
rect 7084 22318 7086 22370
rect 7138 22318 7140 22370
rect 7084 22306 7140 22318
rect 6860 22260 6916 22270
rect 6860 22258 7028 22260
rect 6860 22206 6862 22258
rect 6914 22206 7028 22258
rect 6860 22204 7028 22206
rect 6860 22194 6916 22204
rect 6972 21812 7028 22204
rect 7084 21812 7140 21822
rect 6748 21756 6916 21812
rect 6972 21810 7140 21812
rect 6972 21758 7086 21810
rect 7138 21758 7140 21810
rect 6972 21756 7140 21758
rect 6860 21700 6916 21756
rect 7084 21746 7140 21756
rect 7196 21812 7252 23774
rect 7308 23828 7364 23838
rect 7308 23734 7364 23772
rect 7756 23828 7812 23838
rect 7420 23716 7476 23726
rect 7308 23044 7364 23054
rect 7308 22950 7364 22988
rect 7420 22372 7476 23660
rect 7756 23380 7812 23772
rect 7868 23826 7924 23838
rect 7868 23774 7870 23826
rect 7922 23774 7924 23826
rect 7868 23716 7924 23774
rect 7868 23650 7924 23660
rect 7980 23492 8036 24780
rect 8204 23604 8260 24892
rect 8652 24882 8708 24894
rect 10108 24948 10164 25342
rect 10220 25396 10276 25406
rect 10220 25282 10276 25340
rect 10220 25230 10222 25282
rect 10274 25230 10276 25282
rect 10220 25218 10276 25230
rect 11788 25060 11844 26014
rect 11900 26068 11956 26078
rect 11900 25974 11956 26012
rect 12124 25506 12180 26124
rect 12236 25732 12292 25742
rect 12348 25732 12404 26908
rect 12908 26962 12964 27356
rect 12908 26910 12910 26962
rect 12962 26910 12964 26962
rect 12908 26898 12964 26910
rect 13132 26908 13188 27806
rect 13244 27746 13300 28476
rect 13804 28438 13860 28476
rect 13468 28418 13524 28430
rect 13468 28366 13470 28418
rect 13522 28366 13524 28418
rect 13244 27694 13246 27746
rect 13298 27694 13300 27746
rect 13244 27682 13300 27694
rect 13356 27858 13412 27870
rect 13356 27806 13358 27858
rect 13410 27806 13412 27858
rect 13020 26852 13188 26908
rect 12460 26404 12516 26414
rect 12684 26404 12740 26414
rect 12460 26310 12516 26348
rect 12572 26402 12740 26404
rect 12572 26350 12686 26402
rect 12738 26350 12740 26402
rect 12572 26348 12740 26350
rect 12572 26180 12628 26348
rect 12684 26338 12740 26348
rect 12236 25730 12404 25732
rect 12236 25678 12238 25730
rect 12290 25678 12404 25730
rect 12236 25676 12404 25678
rect 12460 26124 12628 26180
rect 12684 26178 12740 26190
rect 12684 26126 12686 26178
rect 12738 26126 12740 26178
rect 12236 25666 12292 25676
rect 12124 25454 12126 25506
rect 12178 25454 12180 25506
rect 12124 25442 12180 25454
rect 12236 25284 12292 25294
rect 12460 25284 12516 26124
rect 12684 25506 12740 26126
rect 12684 25454 12686 25506
rect 12738 25454 12740 25506
rect 12684 25442 12740 25454
rect 12908 25508 12964 25518
rect 12796 25284 12852 25294
rect 12292 25228 12516 25284
rect 12572 25282 12852 25284
rect 12572 25230 12798 25282
rect 12850 25230 12852 25282
rect 12572 25228 12852 25230
rect 12236 25190 12292 25228
rect 11788 25004 12292 25060
rect 12236 24948 12292 25004
rect 10108 24892 10500 24948
rect 8428 24836 8484 24846
rect 8428 24834 8596 24836
rect 8428 24782 8430 24834
rect 8482 24782 8596 24834
rect 8428 24780 8596 24782
rect 8428 24770 8484 24780
rect 8316 24724 8372 24734
rect 8316 24630 8372 24668
rect 8204 23548 8372 23604
rect 8036 23436 8260 23492
rect 7980 23426 8036 23436
rect 7756 23324 7924 23380
rect 7868 23268 7924 23324
rect 8204 23378 8260 23436
rect 8204 23326 8206 23378
rect 8258 23326 8260 23378
rect 8092 23268 8148 23278
rect 7868 23266 8148 23268
rect 7868 23214 8094 23266
rect 8146 23214 8148 23266
rect 7868 23212 8148 23214
rect 8092 23202 8148 23212
rect 7532 23156 7588 23166
rect 7532 23154 7700 23156
rect 7532 23102 7534 23154
rect 7586 23102 7700 23154
rect 7532 23100 7700 23102
rect 7532 23090 7588 23100
rect 7532 22372 7588 22382
rect 7420 22370 7588 22372
rect 7420 22318 7534 22370
rect 7586 22318 7588 22370
rect 7420 22316 7588 22318
rect 7308 21812 7364 21822
rect 7196 21810 7364 21812
rect 7196 21758 7310 21810
rect 7362 21758 7364 21810
rect 7196 21756 7364 21758
rect 6524 21644 6692 21700
rect 6860 21644 7028 21700
rect 3724 21586 4004 21588
rect 3724 21534 3726 21586
rect 3778 21534 4004 21586
rect 3724 21532 4004 21534
rect 3724 20244 3780 21532
rect 6524 21476 6580 21486
rect 6524 21382 6580 21420
rect 5496 21196 5760 21206
rect 5552 21140 5600 21196
rect 5656 21140 5704 21196
rect 5496 21130 5760 21140
rect 6636 20802 6692 21644
rect 6972 20916 7028 21644
rect 7196 21476 7252 21756
rect 7308 21746 7364 21756
rect 7196 21410 7252 21420
rect 7420 21586 7476 21598
rect 7420 21534 7422 21586
rect 7474 21534 7476 21586
rect 7420 21252 7476 21534
rect 7532 21476 7588 22316
rect 7644 21810 7700 23100
rect 7756 23154 7812 23166
rect 7756 23102 7758 23154
rect 7810 23102 7812 23154
rect 7756 22596 7812 23102
rect 8204 23044 8260 23326
rect 7756 22530 7812 22540
rect 7868 22988 8260 23044
rect 7644 21758 7646 21810
rect 7698 21758 7700 21810
rect 7644 21746 7700 21758
rect 7868 21810 7924 22988
rect 8204 22708 8260 22718
rect 8204 22482 8260 22652
rect 8204 22430 8206 22482
rect 8258 22430 8260 22482
rect 8204 22418 8260 22430
rect 7868 21758 7870 21810
rect 7922 21758 7924 21810
rect 7868 21746 7924 21758
rect 7532 21410 7588 21420
rect 7980 21586 8036 21598
rect 7980 21534 7982 21586
rect 8034 21534 8036 21586
rect 7980 21252 8036 21534
rect 7420 21196 8036 21252
rect 6972 20860 7588 20916
rect 6636 20750 6638 20802
rect 6690 20750 6692 20802
rect 6636 20738 6692 20750
rect 6972 20690 7028 20702
rect 6972 20638 6974 20690
rect 7026 20638 7028 20690
rect 6412 20580 6468 20590
rect 6300 20578 6468 20580
rect 6300 20526 6414 20578
rect 6466 20526 6468 20578
rect 6300 20524 6468 20526
rect 3724 20178 3780 20188
rect 5068 20244 5124 20254
rect 5068 20018 5124 20188
rect 5068 19966 5070 20018
rect 5122 19966 5124 20018
rect 5068 19954 5124 19966
rect 6300 20244 6356 20524
rect 6412 20514 6468 20524
rect 6524 20580 6580 20590
rect 5740 19908 5796 19918
rect 5740 19814 5796 19852
rect 5496 19628 5760 19638
rect 5552 19572 5600 19628
rect 5656 19572 5704 19628
rect 5496 19562 5760 19572
rect 5740 19234 5796 19246
rect 5740 19182 5742 19234
rect 5794 19182 5796 19234
rect 5740 18564 5796 19182
rect 6076 18564 6132 18574
rect 6300 18564 6356 20188
rect 6412 19348 6468 19358
rect 6524 19348 6580 20524
rect 6860 20578 6916 20590
rect 6860 20526 6862 20578
rect 6914 20526 6916 20578
rect 6860 19796 6916 20526
rect 6860 19730 6916 19740
rect 6412 19346 6580 19348
rect 6412 19294 6414 19346
rect 6466 19294 6580 19346
rect 6412 19292 6580 19294
rect 6412 19282 6468 19292
rect 6972 18788 7028 20638
rect 6972 18722 7028 18732
rect 7308 20690 7364 20702
rect 7308 20638 7310 20690
rect 7362 20638 7364 20690
rect 7308 18676 7364 20638
rect 7420 20580 7476 20590
rect 7420 20486 7476 20524
rect 7308 18610 7364 18620
rect 7532 19348 7588 20860
rect 7644 20692 7700 20702
rect 7644 20690 7812 20692
rect 7644 20638 7646 20690
rect 7698 20638 7812 20690
rect 7644 20636 7812 20638
rect 7644 20626 7700 20636
rect 5740 18508 6076 18564
rect 6132 18508 6356 18564
rect 7420 18564 7476 18574
rect 6076 18498 6132 18508
rect 7420 18470 7476 18508
rect 7532 18562 7588 19292
rect 7532 18510 7534 18562
rect 7586 18510 7588 18562
rect 7532 18498 7588 18510
rect 7308 18452 7364 18462
rect 5496 18060 5760 18070
rect 5552 18004 5600 18060
rect 5656 18004 5704 18060
rect 5496 17994 5760 18004
rect 7308 17666 7364 18396
rect 7756 18450 7812 20636
rect 7868 20690 7924 20702
rect 7868 20638 7870 20690
rect 7922 20638 7924 20690
rect 7868 20244 7924 20638
rect 7868 20178 7924 20188
rect 7980 20468 8036 21196
rect 8204 20578 8260 20590
rect 8204 20526 8206 20578
rect 8258 20526 8260 20578
rect 8204 20468 8260 20526
rect 7980 20412 8260 20468
rect 7980 20132 8036 20412
rect 7868 19906 7924 19918
rect 7868 19854 7870 19906
rect 7922 19854 7924 19906
rect 7868 19796 7924 19854
rect 7868 19730 7924 19740
rect 7756 18398 7758 18450
rect 7810 18398 7812 18450
rect 7756 18386 7812 18398
rect 7868 18676 7924 18686
rect 7868 18450 7924 18620
rect 7980 18564 8036 20076
rect 8204 20244 8260 20254
rect 8204 20130 8260 20188
rect 8204 20078 8206 20130
rect 8258 20078 8260 20130
rect 8204 20066 8260 20078
rect 8316 19908 8372 23548
rect 8428 23156 8484 23166
rect 8428 23062 8484 23100
rect 8428 21588 8484 21598
rect 8428 21494 8484 21532
rect 8540 21252 8596 24780
rect 9548 24834 9604 24846
rect 9548 24782 9550 24834
rect 9602 24782 9604 24834
rect 9548 24724 9604 24782
rect 10444 24834 10500 24892
rect 10444 24782 10446 24834
rect 10498 24782 10500 24834
rect 9548 24658 9604 24668
rect 9884 24722 9940 24734
rect 10332 24724 10388 24734
rect 9884 24670 9886 24722
rect 9938 24670 9940 24722
rect 9100 24610 9156 24622
rect 9100 24558 9102 24610
rect 9154 24558 9156 24610
rect 9100 24500 9156 24558
rect 9100 24434 9156 24444
rect 9884 24500 9940 24670
rect 9884 24434 9940 24444
rect 10220 24722 10388 24724
rect 10220 24670 10334 24722
rect 10386 24670 10388 24722
rect 10220 24668 10388 24670
rect 10220 23828 10276 24668
rect 10332 24658 10388 24668
rect 9780 23548 10044 23558
rect 9836 23492 9884 23548
rect 9940 23492 9988 23548
rect 9780 23482 10044 23492
rect 9100 23380 9156 23390
rect 9100 23378 9828 23380
rect 9100 23326 9102 23378
rect 9154 23326 9828 23378
rect 9100 23324 9828 23326
rect 9100 23314 9156 23324
rect 8876 23266 8932 23278
rect 8876 23214 8878 23266
rect 8930 23214 8932 23266
rect 7980 18498 8036 18508
rect 8092 19852 8372 19908
rect 8428 21196 8596 21252
rect 8764 23154 8820 23166
rect 8764 23102 8766 23154
rect 8818 23102 8820 23154
rect 8092 18674 8148 19852
rect 8428 19796 8484 21196
rect 8540 20804 8596 20814
rect 8540 20710 8596 20748
rect 8764 20692 8820 23102
rect 8876 22484 8932 23214
rect 9436 23156 9492 23166
rect 9436 23062 9492 23100
rect 9772 23154 9828 23324
rect 9772 23102 9774 23154
rect 9826 23102 9828 23154
rect 9772 23090 9828 23102
rect 10108 23154 10164 23166
rect 10108 23102 10110 23154
rect 10162 23102 10164 23154
rect 9660 23042 9716 23054
rect 9660 22990 9662 23042
rect 9714 22990 9716 23042
rect 9660 22708 9716 22990
rect 9660 22642 9716 22652
rect 10108 22596 10164 23102
rect 10108 22530 10164 22540
rect 8876 22418 8932 22428
rect 10220 22372 10276 23772
rect 10332 22484 10388 22494
rect 10444 22484 10500 24782
rect 11564 24836 11620 24846
rect 11564 24742 11620 24780
rect 12012 24836 12068 24846
rect 10668 24724 10724 24734
rect 10668 24722 10948 24724
rect 10668 24670 10670 24722
rect 10722 24670 10948 24722
rect 10668 24668 10948 24670
rect 10668 24658 10724 24668
rect 10388 22428 10500 22484
rect 10556 23156 10612 23166
rect 10332 22390 10388 22428
rect 10108 22316 10276 22372
rect 10108 22148 10164 22316
rect 9780 21980 10044 21990
rect 9836 21924 9884 21980
rect 9940 21924 9988 21980
rect 9780 21914 10044 21924
rect 10108 21810 10164 22092
rect 10556 22036 10612 23100
rect 10892 22370 10948 24668
rect 11340 24722 11396 24734
rect 11340 24670 11342 24722
rect 11394 24670 11396 24722
rect 11116 24610 11172 24622
rect 11116 24558 11118 24610
rect 11170 24558 11172 24610
rect 11116 24500 11172 24558
rect 11116 24434 11172 24444
rect 10892 22318 10894 22370
rect 10946 22318 10948 22370
rect 10892 22306 10948 22318
rect 11228 23042 11284 23054
rect 11228 22990 11230 23042
rect 11282 22990 11284 23042
rect 11228 22146 11284 22990
rect 11340 22370 11396 24670
rect 11676 24722 11732 24734
rect 11676 24670 11678 24722
rect 11730 24670 11732 24722
rect 11340 22318 11342 22370
rect 11394 22318 11396 22370
rect 11340 22306 11396 22318
rect 11564 22596 11620 22606
rect 11564 22260 11620 22540
rect 11564 22166 11620 22204
rect 11228 22094 11230 22146
rect 11282 22094 11284 22146
rect 11228 22082 11284 22094
rect 10108 21758 10110 21810
rect 10162 21758 10164 21810
rect 10108 21746 10164 21758
rect 10220 21980 10612 22036
rect 10220 21588 10276 21980
rect 10444 21812 10500 21822
rect 9996 21532 10276 21588
rect 10332 21756 10444 21812
rect 10332 21588 10388 21756
rect 10444 21746 10500 21756
rect 11676 21700 11732 24670
rect 12012 23604 12068 24780
rect 12236 24834 12292 24892
rect 12572 24946 12628 25228
rect 12796 25218 12852 25228
rect 12572 24894 12574 24946
rect 12626 24894 12628 24946
rect 12572 24882 12628 24894
rect 12796 24948 12852 24958
rect 12796 24854 12852 24892
rect 12236 24782 12238 24834
rect 12290 24782 12292 24834
rect 12236 24770 12292 24782
rect 12348 24836 12404 24846
rect 12348 24742 12404 24780
rect 12908 24164 12964 25452
rect 13020 25506 13076 26852
rect 13356 26740 13412 27806
rect 13468 27412 13524 28366
rect 13692 28420 13748 28430
rect 13692 28326 13748 28364
rect 13580 28084 13636 28094
rect 13580 28082 13972 28084
rect 13580 28030 13582 28082
rect 13634 28030 13972 28082
rect 13580 28028 13972 28030
rect 13580 28018 13636 28028
rect 13692 27860 13748 27870
rect 13692 27766 13748 27804
rect 13468 27346 13524 27356
rect 13804 27636 13860 27646
rect 13804 27186 13860 27580
rect 13804 27134 13806 27186
rect 13858 27134 13860 27186
rect 13804 27122 13860 27134
rect 13916 27076 13972 28028
rect 14252 27972 14308 28590
rect 14252 27878 14308 27916
rect 14064 27468 14328 27478
rect 14120 27412 14168 27468
rect 14224 27412 14272 27468
rect 14064 27402 14328 27412
rect 14028 27076 14084 27086
rect 14364 27076 14420 27086
rect 13916 27074 14420 27076
rect 13916 27022 14030 27074
rect 14082 27022 14366 27074
rect 14418 27022 14420 27074
rect 13916 27020 14420 27022
rect 14028 27010 14084 27020
rect 14364 27010 14420 27020
rect 13468 26962 13524 26974
rect 13468 26910 13470 26962
rect 13522 26910 13524 26962
rect 13468 26740 13524 26910
rect 13692 26852 13748 26862
rect 13244 26684 13524 26740
rect 13580 26850 13748 26852
rect 13580 26798 13694 26850
rect 13746 26798 13748 26850
rect 13580 26796 13748 26798
rect 13132 26180 13188 26190
rect 13132 26086 13188 26124
rect 13020 25454 13022 25506
rect 13074 25454 13076 25506
rect 13020 25442 13076 25454
rect 13244 25060 13300 26684
rect 13356 26516 13412 26526
rect 13356 26290 13412 26460
rect 13580 26402 13636 26796
rect 13692 26786 13748 26796
rect 13916 26852 13972 26862
rect 13580 26350 13582 26402
rect 13634 26350 13636 26402
rect 13580 26338 13636 26350
rect 13356 26238 13358 26290
rect 13410 26238 13412 26290
rect 13356 26226 13412 26238
rect 13804 26292 13860 26302
rect 13916 26292 13972 26796
rect 13804 26290 13972 26292
rect 13804 26238 13806 26290
rect 13858 26238 13972 26290
rect 13804 26236 13972 26238
rect 13804 26226 13860 26236
rect 13916 26068 13972 26078
rect 13580 26066 13972 26068
rect 13580 26014 13918 26066
rect 13970 26014 13972 26066
rect 13580 26012 13972 26014
rect 13580 25730 13636 26012
rect 13916 26002 13972 26012
rect 14064 25900 14328 25910
rect 14120 25844 14168 25900
rect 14224 25844 14272 25900
rect 14064 25834 14328 25844
rect 13580 25678 13582 25730
rect 13634 25678 13636 25730
rect 13580 25666 13636 25678
rect 13692 25620 13748 25630
rect 13692 25506 13748 25564
rect 13692 25454 13694 25506
rect 13746 25454 13748 25506
rect 13692 25442 13748 25454
rect 14028 25620 14084 25630
rect 13244 24994 13300 25004
rect 13580 25282 13636 25294
rect 13580 25230 13582 25282
rect 13634 25230 13636 25282
rect 13580 24948 13636 25230
rect 13468 24892 13636 24948
rect 13692 25172 13748 25182
rect 13132 24722 13188 24734
rect 13132 24670 13134 24722
rect 13186 24670 13188 24722
rect 13132 24500 13188 24670
rect 13132 24434 13188 24444
rect 11900 22258 11956 22270
rect 11900 22206 11902 22258
rect 11954 22206 11956 22258
rect 11900 22148 11956 22206
rect 12012 22258 12068 23548
rect 12012 22206 12014 22258
rect 12066 22206 12068 22258
rect 12012 22194 12068 22206
rect 12124 24108 12964 24164
rect 11900 22082 11956 22092
rect 11900 21924 11956 21934
rect 11900 21810 11956 21868
rect 11900 21758 11902 21810
rect 11954 21758 11956 21810
rect 11900 21746 11956 21758
rect 11788 21700 11844 21710
rect 11564 21698 11844 21700
rect 11564 21646 11790 21698
rect 11842 21646 11844 21698
rect 11564 21644 11844 21646
rect 8764 20626 8820 20636
rect 8876 21476 8932 21486
rect 8540 20020 8596 20030
rect 8540 19926 8596 19964
rect 8764 20018 8820 20030
rect 8764 19966 8766 20018
rect 8818 19966 8820 20018
rect 8652 19908 8708 19918
rect 8652 19814 8708 19852
rect 8428 19730 8484 19740
rect 8540 19348 8596 19358
rect 8540 19254 8596 19292
rect 8764 19234 8820 19966
rect 8764 19182 8766 19234
rect 8818 19182 8820 19234
rect 8764 19170 8820 19182
rect 8092 18622 8094 18674
rect 8146 18622 8148 18674
rect 7868 18398 7870 18450
rect 7922 18398 7924 18450
rect 7868 18386 7924 18398
rect 8092 18340 8148 18622
rect 8204 18788 8260 18798
rect 8204 18676 8260 18732
rect 8652 18676 8708 18686
rect 8204 18674 8708 18676
rect 8204 18622 8654 18674
rect 8706 18622 8708 18674
rect 8204 18620 8708 18622
rect 8204 18562 8260 18620
rect 8204 18510 8206 18562
rect 8258 18510 8260 18562
rect 8204 18498 8260 18510
rect 8092 18274 8148 18284
rect 7308 17614 7310 17666
rect 7362 17614 7364 17666
rect 7308 17602 7364 17614
rect 8092 17556 8148 17566
rect 8092 17554 8596 17556
rect 8092 17502 8094 17554
rect 8146 17502 8596 17554
rect 8092 17500 8596 17502
rect 8092 17490 8148 17500
rect 8540 17106 8596 17500
rect 8540 17054 8542 17106
rect 8594 17054 8596 17106
rect 8540 17042 8596 17054
rect 8428 16884 8484 16894
rect 8652 16884 8708 18620
rect 8876 18452 8932 21420
rect 9324 21364 9380 21374
rect 9324 20804 9380 21308
rect 9324 20710 9380 20748
rect 9996 20802 10052 21532
rect 9996 20750 9998 20802
rect 10050 20750 10052 20802
rect 9996 20738 10052 20750
rect 9548 20692 9604 20702
rect 9548 20598 9604 20636
rect 9780 20412 10044 20422
rect 9836 20356 9884 20412
rect 9940 20356 9988 20412
rect 9780 20346 10044 20356
rect 10332 20244 10388 21532
rect 9660 20130 9716 20142
rect 9660 20078 9662 20130
rect 9714 20078 9716 20130
rect 9436 20020 9492 20030
rect 9436 19926 9492 19964
rect 9660 19796 9716 20078
rect 9772 20132 9828 20142
rect 9772 20038 9828 20076
rect 10332 20130 10388 20188
rect 10332 20078 10334 20130
rect 10386 20078 10388 20130
rect 10332 20066 10388 20078
rect 10444 21588 10500 21598
rect 10780 21588 10836 21598
rect 10444 21586 10780 21588
rect 10444 21534 10446 21586
rect 10498 21534 10780 21586
rect 10444 21532 10780 21534
rect 9660 19730 9716 19740
rect 10220 19908 10276 19918
rect 8988 19348 9044 19358
rect 8988 19122 9044 19292
rect 10220 19346 10276 19852
rect 10220 19294 10222 19346
rect 10274 19294 10276 19346
rect 10220 19282 10276 19294
rect 9548 19234 9604 19246
rect 9548 19182 9550 19234
rect 9602 19182 9604 19234
rect 8988 19070 8990 19122
rect 9042 19070 9044 19122
rect 8988 19058 9044 19070
rect 9100 19122 9156 19134
rect 9100 19070 9102 19122
rect 9154 19070 9156 19122
rect 9100 18788 9156 19070
rect 9100 18722 9156 18732
rect 8876 18386 8932 18396
rect 8988 18450 9044 18462
rect 8988 18398 8990 18450
rect 9042 18398 9044 18450
rect 8988 17892 9044 18398
rect 9548 18452 9604 19182
rect 9780 18844 10044 18854
rect 9836 18788 9884 18844
rect 9940 18788 9988 18844
rect 9780 18778 10044 18788
rect 10108 18676 10164 18686
rect 10444 18676 10500 21532
rect 10780 21522 10836 21532
rect 10892 21476 10948 21486
rect 10892 21382 10948 21420
rect 11564 20916 11620 21644
rect 11788 21634 11844 21644
rect 11900 21364 11956 21374
rect 11564 20850 11620 20860
rect 11676 21362 11956 21364
rect 11676 21310 11902 21362
rect 11954 21310 11956 21362
rect 11676 21308 11956 21310
rect 10668 20692 10724 20702
rect 10668 20690 11620 20692
rect 10668 20638 10670 20690
rect 10722 20638 11620 20690
rect 10668 20636 11620 20638
rect 10668 20626 10724 20636
rect 10892 20468 10948 20478
rect 10892 20130 10948 20412
rect 11452 20468 11508 20478
rect 10892 20078 10894 20130
rect 10946 20078 10948 20130
rect 10892 20066 10948 20078
rect 11004 20130 11060 20142
rect 11004 20078 11006 20130
rect 11058 20078 11060 20130
rect 11004 19796 11060 20078
rect 11452 20130 11508 20412
rect 11564 20242 11620 20636
rect 11564 20190 11566 20242
rect 11618 20190 11620 20242
rect 11564 20178 11620 20190
rect 11452 20078 11454 20130
rect 11506 20078 11508 20130
rect 11452 20066 11508 20078
rect 11228 20020 11284 20030
rect 11228 19926 11284 19964
rect 11676 20018 11732 21308
rect 11900 21298 11956 21308
rect 12124 20244 12180 24108
rect 12908 23940 12964 23950
rect 12908 23846 12964 23884
rect 13356 23604 13412 23614
rect 13356 23042 13412 23548
rect 13356 22990 13358 23042
rect 13410 22990 13412 23042
rect 13356 22978 13412 22990
rect 12460 22260 12516 22270
rect 12460 22166 12516 22204
rect 12796 22258 12852 22270
rect 12796 22206 12798 22258
rect 12850 22206 12852 22258
rect 12236 22146 12292 22158
rect 12236 22094 12238 22146
rect 12290 22094 12292 22146
rect 12236 20468 12292 22094
rect 12684 21586 12740 21598
rect 12684 21534 12686 21586
rect 12738 21534 12740 21586
rect 12684 21476 12740 21534
rect 12796 21476 12852 22206
rect 12908 22260 12964 22270
rect 12908 21812 12964 22204
rect 12908 21718 12964 21756
rect 13356 21924 13412 21934
rect 13468 21924 13524 24892
rect 13580 24722 13636 24734
rect 13580 24670 13582 24722
rect 13634 24670 13636 24722
rect 13580 24500 13636 24670
rect 13580 24434 13636 24444
rect 13580 23940 13636 23950
rect 13580 23846 13636 23884
rect 13412 21868 13524 21924
rect 13580 22148 13636 22158
rect 13244 21698 13300 21710
rect 13244 21646 13246 21698
rect 13298 21646 13300 21698
rect 13244 21476 13300 21646
rect 12684 21420 13300 21476
rect 12796 20914 12852 20926
rect 12796 20862 12798 20914
rect 12850 20862 12852 20914
rect 12796 20580 12852 20862
rect 13244 20804 13300 21420
rect 13244 20738 13300 20748
rect 13356 20580 13412 21868
rect 13580 21698 13636 22092
rect 13580 21646 13582 21698
rect 13634 21646 13636 21698
rect 13580 21634 13636 21646
rect 13692 21364 13748 25116
rect 14028 24722 14084 25564
rect 14252 25282 14308 25294
rect 14252 25230 14254 25282
rect 14306 25230 14308 25282
rect 14252 25060 14308 25230
rect 14252 24994 14308 25004
rect 14476 24836 14532 29820
rect 14588 28532 14644 28542
rect 14588 27746 14644 28476
rect 14588 27694 14590 27746
rect 14642 27694 14644 27746
rect 14588 27682 14644 27694
rect 14700 28420 14756 28430
rect 14588 27300 14644 27310
rect 14588 26962 14644 27244
rect 14700 27188 14756 28364
rect 14812 27860 14868 30828
rect 14924 30790 14980 30828
rect 15036 30436 15092 36200
rect 16044 33460 16100 33470
rect 15932 33404 16044 33460
rect 15820 32788 15876 32798
rect 15820 32694 15876 32732
rect 15372 32452 15428 32462
rect 15372 32358 15428 32396
rect 15372 31220 15428 31230
rect 15372 31126 15428 31164
rect 15708 31220 15764 31230
rect 15596 30996 15652 31006
rect 15596 30902 15652 30940
rect 15596 30436 15652 30446
rect 15036 30434 15652 30436
rect 15036 30382 15598 30434
rect 15650 30382 15652 30434
rect 15036 30380 15652 30382
rect 15596 30370 15652 30380
rect 15596 28868 15652 28878
rect 15708 28868 15764 31164
rect 15932 28980 15988 33404
rect 16044 33366 16100 33404
rect 16156 33236 16212 36200
rect 17276 33460 17332 36200
rect 18396 33572 18452 36200
rect 18396 33516 18788 33572
rect 17276 33404 17668 33460
rect 17052 33348 17108 33358
rect 17052 33346 17556 33348
rect 17052 33294 17054 33346
rect 17106 33294 17556 33346
rect 17052 33292 17556 33294
rect 17052 33282 17108 33292
rect 16044 33180 16212 33236
rect 16044 31890 16100 33180
rect 16044 31838 16046 31890
rect 16098 31838 16100 31890
rect 16044 31826 16100 31838
rect 16156 32674 16212 32686
rect 16156 32622 16158 32674
rect 16210 32622 16212 32674
rect 16156 31332 16212 32622
rect 16828 32676 16884 32686
rect 16828 32582 16884 32620
rect 16492 32562 16548 32574
rect 16492 32510 16494 32562
rect 16546 32510 16548 32562
rect 16268 32452 16324 32462
rect 16324 32396 16436 32452
rect 16268 32386 16324 32396
rect 16044 30996 16100 31006
rect 16044 30902 16100 30940
rect 16156 29764 16212 31276
rect 16268 31106 16324 31118
rect 16268 31054 16270 31106
rect 16322 31054 16324 31106
rect 16268 30996 16324 31054
rect 16268 30930 16324 30940
rect 16380 30994 16436 32396
rect 16380 30942 16382 30994
rect 16434 30942 16436 30994
rect 16380 29876 16436 30942
rect 16380 29810 16436 29820
rect 16156 29708 16324 29764
rect 16268 29652 16324 29708
rect 16380 29652 16436 29662
rect 16268 29650 16436 29652
rect 16268 29598 16382 29650
rect 16434 29598 16436 29650
rect 16268 29596 16436 29598
rect 15596 28866 15764 28868
rect 15596 28814 15598 28866
rect 15650 28814 15764 28866
rect 15596 28812 15764 28814
rect 15820 28924 15988 28980
rect 16156 29426 16212 29438
rect 16156 29374 16158 29426
rect 16210 29374 16212 29426
rect 15596 28802 15652 28812
rect 15372 28756 15428 28766
rect 15372 28662 15428 28700
rect 15036 28644 15092 28654
rect 15036 28550 15092 28588
rect 15820 28644 15876 28924
rect 15932 28756 15988 28766
rect 16156 28756 16212 29374
rect 16268 29428 16324 29438
rect 16268 29334 16324 29372
rect 15988 28700 16212 28756
rect 16268 29204 16324 29214
rect 15932 28662 15988 28700
rect 15820 28578 15876 28588
rect 15596 28196 15652 28206
rect 14812 27794 14868 27804
rect 14924 27970 14980 27982
rect 14924 27918 14926 27970
rect 14978 27918 14980 27970
rect 14700 27122 14756 27132
rect 14588 26910 14590 26962
rect 14642 26910 14644 26962
rect 14588 26898 14644 26910
rect 14700 26964 14756 27002
rect 14924 26964 14980 27918
rect 15036 27970 15092 27982
rect 15036 27918 15038 27970
rect 15090 27918 15092 27970
rect 15036 27748 15092 27918
rect 15148 27972 15204 27982
rect 15148 27878 15204 27916
rect 15036 27682 15092 27692
rect 15372 27858 15428 27870
rect 15372 27806 15374 27858
rect 15426 27806 15428 27858
rect 15260 27188 15316 27198
rect 14924 26908 15204 26964
rect 14700 26898 14756 26908
rect 14812 26852 14868 26862
rect 14700 26178 14756 26190
rect 14700 26126 14702 26178
rect 14754 26126 14756 26178
rect 14700 26068 14756 26126
rect 14700 26002 14756 26012
rect 14588 25508 14644 25518
rect 14812 25508 14868 26796
rect 14588 25506 14868 25508
rect 14588 25454 14590 25506
rect 14642 25454 14868 25506
rect 14588 25452 14868 25454
rect 14924 26404 14980 26414
rect 14924 26068 14980 26348
rect 14924 25506 14980 26012
rect 14924 25454 14926 25506
rect 14978 25454 14980 25506
rect 14588 25442 14644 25452
rect 14924 25442 14980 25454
rect 15036 25956 15092 25966
rect 15036 25508 15092 25900
rect 15036 25442 15092 25452
rect 15036 25284 15092 25294
rect 14028 24670 14030 24722
rect 14082 24670 14084 24722
rect 14028 24658 14084 24670
rect 14364 24780 14532 24836
rect 14588 25282 15092 25284
rect 14588 25230 15038 25282
rect 15090 25230 15092 25282
rect 14588 25228 15092 25230
rect 14364 24500 14420 24780
rect 13804 24444 14420 24500
rect 14476 24610 14532 24622
rect 14476 24558 14478 24610
rect 14530 24558 14532 24610
rect 14476 24500 14532 24558
rect 13804 23378 13860 24444
rect 14476 24434 14532 24444
rect 14064 24332 14328 24342
rect 14120 24276 14168 24332
rect 14224 24276 14272 24332
rect 14064 24266 14328 24276
rect 13804 23326 13806 23378
rect 13858 23326 13860 23378
rect 13804 23156 13860 23326
rect 14252 23940 14308 23950
rect 14252 23378 14308 23884
rect 14252 23326 14254 23378
rect 14306 23326 14308 23378
rect 14252 23314 14308 23326
rect 13804 22484 13860 23100
rect 14064 22764 14328 22774
rect 14120 22708 14168 22764
rect 14224 22708 14272 22764
rect 14064 22698 14328 22708
rect 13804 21588 13860 22428
rect 14476 21812 14532 21822
rect 13916 21588 13972 21598
rect 13804 21586 13972 21588
rect 13804 21534 13918 21586
rect 13970 21534 13972 21586
rect 13804 21532 13972 21534
rect 13580 21308 13748 21364
rect 12796 20524 13412 20580
rect 13468 20578 13524 20590
rect 13468 20526 13470 20578
rect 13522 20526 13524 20578
rect 12236 20402 12292 20412
rect 11676 19966 11678 20018
rect 11730 19966 11732 20018
rect 11676 19954 11732 19966
rect 11788 20188 12180 20244
rect 12908 20244 12964 20254
rect 11004 19730 11060 19740
rect 10108 18674 10500 18676
rect 10108 18622 10110 18674
rect 10162 18622 10500 18674
rect 10108 18620 10500 18622
rect 10108 18610 10164 18620
rect 9548 18386 9604 18396
rect 9884 18450 9940 18462
rect 9884 18398 9886 18450
rect 9938 18398 9940 18450
rect 8988 17826 9044 17836
rect 9884 17892 9940 18398
rect 9884 17826 9940 17836
rect 10220 18340 10276 18350
rect 10220 17780 10276 18284
rect 10108 17778 10276 17780
rect 10108 17726 10222 17778
rect 10274 17726 10276 17778
rect 10108 17724 10276 17726
rect 9780 17276 10044 17286
rect 9836 17220 9884 17276
rect 9940 17220 9988 17276
rect 9780 17210 10044 17220
rect 9884 17108 9940 17118
rect 8988 17106 9940 17108
rect 8988 17054 9886 17106
rect 9938 17054 9940 17106
rect 8988 17052 9940 17054
rect 8988 16994 9044 17052
rect 9884 17042 9940 17052
rect 9996 17108 10052 17118
rect 10108 17108 10164 17724
rect 10220 17714 10276 17724
rect 10444 18340 10500 18620
rect 11004 19348 11060 19358
rect 10556 18452 10612 18462
rect 10612 18396 10836 18452
rect 10556 18358 10612 18396
rect 9996 17106 10164 17108
rect 9996 17054 9998 17106
rect 10050 17054 10164 17106
rect 9996 17052 10164 17054
rect 10332 17108 10388 17118
rect 9996 17042 10052 17052
rect 8988 16942 8990 16994
rect 9042 16942 9044 16994
rect 8988 16930 9044 16942
rect 8428 16882 8708 16884
rect 8428 16830 8430 16882
rect 8482 16830 8708 16882
rect 8428 16828 8708 16830
rect 8764 16882 8820 16894
rect 8764 16830 8766 16882
rect 8818 16830 8820 16882
rect 8428 16818 8484 16828
rect 8316 16660 8372 16670
rect 5496 16492 5760 16502
rect 5552 16436 5600 16492
rect 5656 16436 5704 16492
rect 5496 16426 5760 16436
rect 5496 14924 5760 14934
rect 5552 14868 5600 14924
rect 5656 14868 5704 14924
rect 5496 14858 5760 14868
rect 8316 14644 8372 16604
rect 8764 16212 8820 16830
rect 9772 16884 9828 16894
rect 9772 16790 9828 16828
rect 10332 16882 10388 17052
rect 10332 16830 10334 16882
rect 10386 16830 10388 16882
rect 10332 16818 10388 16830
rect 10444 16884 10500 18284
rect 10780 17778 10836 18396
rect 10780 17726 10782 17778
rect 10834 17726 10836 17778
rect 10780 17714 10836 17726
rect 10892 17444 10948 17454
rect 10780 17108 10836 17118
rect 10780 17014 10836 17052
rect 10444 16818 10500 16828
rect 10108 16772 10164 16782
rect 9212 16212 9268 16222
rect 8764 16156 9212 16212
rect 9212 16118 9268 16156
rect 10108 16098 10164 16716
rect 10780 16212 10836 16222
rect 10892 16212 10948 17388
rect 11004 16660 11060 19292
rect 11788 16772 11844 20188
rect 12012 20020 12068 20030
rect 12460 20020 12516 20030
rect 12012 20018 12516 20020
rect 12012 19966 12014 20018
rect 12066 19966 12462 20018
rect 12514 19966 12516 20018
rect 12012 19964 12516 19966
rect 12012 19954 12068 19964
rect 12348 19796 12404 19806
rect 12348 19346 12404 19740
rect 12460 19460 12516 19964
rect 12572 20020 12628 20030
rect 12572 19926 12628 19964
rect 12796 19908 12852 19918
rect 12796 19814 12852 19852
rect 12908 19460 12964 20188
rect 13132 20130 13188 20142
rect 13132 20078 13134 20130
rect 13186 20078 13188 20130
rect 13020 20020 13076 20030
rect 13132 20020 13188 20078
rect 13244 20132 13300 20524
rect 13468 20244 13524 20526
rect 13468 20178 13524 20188
rect 13356 20132 13412 20142
rect 13244 20130 13412 20132
rect 13244 20078 13358 20130
rect 13410 20078 13412 20130
rect 13244 20076 13412 20078
rect 13356 20066 13412 20076
rect 13020 20018 13188 20020
rect 13020 19966 13022 20018
rect 13074 19966 13188 20018
rect 13020 19964 13188 19966
rect 13468 20018 13524 20030
rect 13468 19966 13470 20018
rect 13522 19966 13524 20018
rect 13020 19954 13076 19964
rect 12460 19404 12964 19460
rect 12348 19294 12350 19346
rect 12402 19294 12404 19346
rect 12348 18674 12404 19294
rect 12684 19236 12740 19246
rect 12684 18788 12740 19180
rect 12796 19124 12852 19134
rect 12796 19030 12852 19068
rect 12348 18622 12350 18674
rect 12402 18622 12404 18674
rect 12348 18610 12404 18622
rect 12460 18732 12852 18788
rect 12460 18562 12516 18732
rect 12796 18674 12852 18732
rect 12796 18622 12798 18674
rect 12850 18622 12852 18674
rect 12796 18610 12852 18622
rect 12460 18510 12462 18562
rect 12514 18510 12516 18562
rect 12460 18498 12516 18510
rect 12684 18564 12740 18574
rect 12348 18226 12404 18238
rect 12348 18174 12350 18226
rect 12402 18174 12404 18226
rect 12348 17666 12404 18174
rect 12348 17614 12350 17666
rect 12402 17614 12404 17666
rect 12348 17602 12404 17614
rect 12684 17666 12740 18508
rect 12684 17614 12686 17666
rect 12738 17614 12740 17666
rect 12684 17602 12740 17614
rect 12908 17668 12964 19404
rect 13468 19236 13524 19966
rect 13468 19170 13524 19180
rect 13020 19012 13076 19022
rect 13020 19010 13412 19012
rect 13020 18958 13022 19010
rect 13074 18958 13412 19010
rect 13020 18956 13412 18958
rect 13020 18946 13076 18956
rect 12908 17574 12964 17612
rect 13020 18788 13076 18798
rect 12460 17444 12516 17454
rect 12460 17350 12516 17388
rect 12796 17108 12852 17118
rect 12684 16996 12740 17006
rect 12684 16902 12740 16940
rect 12012 16884 12068 16894
rect 12012 16790 12068 16828
rect 11004 16594 11060 16604
rect 11676 16716 11844 16772
rect 10780 16210 10948 16212
rect 10780 16158 10782 16210
rect 10834 16158 10948 16210
rect 10780 16156 10948 16158
rect 11676 16212 11732 16716
rect 10780 16146 10836 16156
rect 10108 16046 10110 16098
rect 10162 16046 10164 16098
rect 10108 16034 10164 16046
rect 9780 15708 10044 15718
rect 9836 15652 9884 15708
rect 9940 15652 9988 15708
rect 9780 15642 10044 15652
rect 9212 14756 9268 14766
rect 9212 14644 9268 14700
rect 8092 14642 8372 14644
rect 8092 14590 8318 14642
rect 8370 14590 8372 14642
rect 8092 14588 8372 14590
rect 7084 13970 7140 13982
rect 7084 13918 7086 13970
rect 7138 13918 7140 13970
rect 6860 13748 6916 13758
rect 6860 13654 6916 13692
rect 5496 13356 5760 13366
rect 5552 13300 5600 13356
rect 5656 13300 5704 13356
rect 5496 13290 5760 13300
rect 6188 13186 6244 13198
rect 6188 13134 6190 13186
rect 6242 13134 6244 13186
rect 6188 13076 6244 13134
rect 6188 13020 6468 13076
rect 6412 12964 6468 13020
rect 6524 12964 6580 12974
rect 6412 12962 6580 12964
rect 6412 12910 6526 12962
rect 6578 12910 6580 12962
rect 6412 12908 6580 12910
rect 6524 12898 6580 12908
rect 6300 12850 6356 12862
rect 6300 12798 6302 12850
rect 6354 12798 6356 12850
rect 6188 12738 6244 12750
rect 6188 12686 6190 12738
rect 6242 12686 6244 12738
rect 6188 12516 6244 12686
rect 6300 12628 6356 12798
rect 6972 12852 7028 12862
rect 6972 12758 7028 12796
rect 6300 12562 6356 12572
rect 6860 12738 6916 12750
rect 6860 12686 6862 12738
rect 6914 12686 6916 12738
rect 4844 12404 4900 12414
rect 4844 12066 4900 12348
rect 4844 12014 4846 12066
rect 4898 12014 4900 12066
rect 4172 8930 4228 8942
rect 4172 8878 4174 8930
rect 4226 8878 4228 8930
rect 4172 8484 4228 8878
rect 2268 5236 2324 5246
rect 1820 5234 2324 5236
rect 1820 5182 2270 5234
rect 2322 5182 2324 5234
rect 1820 5180 2324 5182
rect 1820 800 1876 5180
rect 2268 5170 2324 5180
rect 3388 4226 3444 4238
rect 3388 4174 3390 4226
rect 3442 4174 3444 4226
rect 3388 800 3444 4174
rect 4172 3556 4228 8428
rect 4620 5124 4676 5134
rect 4844 5124 4900 12014
rect 5496 11788 5760 11798
rect 5552 11732 5600 11788
rect 5656 11732 5704 11788
rect 5496 11722 5760 11732
rect 5628 11508 5684 11518
rect 6188 11508 6244 12460
rect 6860 12292 6916 12686
rect 6972 12292 7028 12302
rect 6860 12290 7028 12292
rect 6860 12238 6974 12290
rect 7026 12238 7028 12290
rect 6860 12236 7028 12238
rect 6972 12226 7028 12236
rect 7084 11956 7140 13918
rect 8092 13970 8148 14588
rect 8316 14578 8372 14588
rect 8988 14642 9268 14644
rect 8988 14590 9214 14642
rect 9266 14590 9268 14642
rect 8988 14588 9268 14590
rect 8092 13918 8094 13970
rect 8146 13918 8148 13970
rect 7196 13746 7252 13758
rect 7196 13694 7198 13746
rect 7250 13694 7252 13746
rect 7196 13188 7252 13694
rect 7196 13122 7252 13132
rect 7420 13746 7476 13758
rect 7420 13694 7422 13746
rect 7474 13694 7476 13746
rect 7420 13188 7476 13694
rect 7420 13122 7476 13132
rect 7868 13748 7924 13758
rect 7196 12964 7252 12974
rect 7644 12964 7700 12974
rect 7196 12962 7700 12964
rect 7196 12910 7198 12962
rect 7250 12910 7646 12962
rect 7698 12910 7700 12962
rect 7196 12908 7700 12910
rect 7196 12898 7252 12908
rect 7644 12898 7700 12908
rect 7532 12740 7588 12750
rect 7532 12646 7588 12684
rect 7756 12738 7812 12750
rect 7756 12686 7758 12738
rect 7810 12686 7812 12738
rect 7756 12404 7812 12686
rect 7868 12404 7924 13692
rect 8092 12964 8148 13918
rect 8988 13970 9044 14588
rect 9212 14578 9268 14588
rect 10220 14700 11060 14756
rect 10220 14530 10276 14700
rect 10220 14478 10222 14530
rect 10274 14478 10276 14530
rect 10220 14466 10276 14478
rect 10444 14530 10500 14542
rect 10444 14478 10446 14530
rect 10498 14478 10500 14530
rect 10332 14306 10388 14318
rect 10332 14254 10334 14306
rect 10386 14254 10388 14306
rect 9780 14140 10044 14150
rect 9836 14084 9884 14140
rect 9940 14084 9988 14140
rect 9780 14074 10044 14084
rect 8988 13918 8990 13970
rect 9042 13918 9044 13970
rect 8428 13634 8484 13646
rect 8428 13582 8430 13634
rect 8482 13582 8484 13634
rect 8092 12870 8148 12908
rect 8316 13300 8372 13310
rect 8316 12628 8372 13244
rect 8428 12740 8484 13582
rect 8540 13188 8596 13198
rect 8540 13074 8596 13132
rect 8540 13022 8542 13074
rect 8594 13022 8596 13074
rect 8540 13010 8596 13022
rect 8876 12964 8932 12974
rect 8764 12852 8820 12862
rect 8652 12740 8708 12750
rect 8428 12646 8484 12684
rect 8540 12738 8708 12740
rect 8540 12686 8654 12738
rect 8706 12686 8708 12738
rect 8540 12684 8708 12686
rect 7980 12404 8036 12414
rect 7868 12402 8036 12404
rect 7868 12350 7982 12402
rect 8034 12350 8036 12402
rect 7868 12348 8036 12350
rect 7756 12338 7812 12348
rect 7980 12338 8036 12348
rect 8204 12290 8260 12302
rect 8204 12238 8206 12290
rect 8258 12238 8260 12290
rect 7644 12180 7700 12190
rect 7644 12086 7700 12124
rect 7084 11900 7812 11956
rect 5628 11506 6244 11508
rect 5628 11454 5630 11506
rect 5682 11454 6244 11506
rect 5628 11452 6244 11454
rect 7756 11506 7812 11900
rect 7756 11454 7758 11506
rect 7810 11454 7812 11506
rect 5628 10388 5684 11452
rect 7756 11442 7812 11454
rect 7980 11620 8036 11630
rect 7980 10836 8036 11564
rect 4620 5122 4900 5124
rect 4620 5070 4622 5122
rect 4674 5070 4900 5122
rect 4620 5068 4900 5070
rect 5292 10332 5684 10388
rect 7644 10834 8036 10836
rect 7644 10782 7982 10834
rect 8034 10782 8036 10834
rect 7644 10780 8036 10782
rect 4620 5058 4676 5068
rect 5292 4338 5348 10332
rect 5496 10220 5760 10230
rect 5552 10164 5600 10220
rect 5656 10164 5704 10220
rect 5496 10154 5760 10164
rect 7644 10164 7700 10780
rect 7980 10770 8036 10780
rect 6748 9940 6804 9950
rect 6300 8932 6356 8942
rect 6300 8930 6692 8932
rect 6300 8878 6302 8930
rect 6354 8878 6692 8930
rect 6300 8876 6692 8878
rect 6300 8866 6356 8876
rect 5496 8652 5760 8662
rect 5552 8596 5600 8652
rect 5656 8596 5704 8652
rect 5496 8586 5760 8596
rect 6636 8370 6692 8876
rect 6748 8484 6804 9884
rect 7084 9826 7140 9838
rect 7084 9774 7086 9826
rect 7138 9774 7140 9826
rect 7084 9042 7140 9774
rect 7084 8990 7086 9042
rect 7138 8990 7140 9042
rect 7084 8932 7140 8990
rect 7084 8866 7140 8876
rect 7420 9154 7476 9166
rect 7420 9102 7422 9154
rect 7474 9102 7476 9154
rect 7420 8820 7476 9102
rect 7644 9042 7700 10108
rect 8204 9940 8260 12238
rect 8316 12290 8372 12572
rect 8428 12516 8484 12526
rect 8540 12516 8596 12684
rect 8652 12674 8708 12684
rect 8484 12460 8596 12516
rect 8428 12450 8484 12460
rect 8652 12404 8708 12414
rect 8764 12404 8820 12796
rect 8876 12850 8932 12908
rect 8876 12798 8878 12850
rect 8930 12798 8932 12850
rect 8876 12786 8932 12798
rect 8652 12402 8820 12404
rect 8652 12350 8654 12402
rect 8706 12350 8820 12402
rect 8652 12348 8820 12350
rect 8988 12402 9044 13918
rect 10332 13858 10388 14254
rect 10332 13806 10334 13858
rect 10386 13806 10388 13858
rect 10332 13794 10388 13806
rect 9548 13748 9604 13758
rect 8988 12350 8990 12402
rect 9042 12350 9044 12402
rect 8652 12338 8708 12348
rect 8316 12238 8318 12290
rect 8370 12238 8372 12290
rect 8316 12226 8372 12238
rect 8540 12180 8596 12190
rect 8540 11394 8596 12124
rect 8988 11620 9044 12350
rect 9436 13746 9604 13748
rect 9436 13694 9550 13746
rect 9602 13694 9604 13746
rect 9436 13692 9604 13694
rect 9100 12180 9156 12190
rect 9436 12180 9492 13692
rect 9548 13682 9604 13692
rect 10444 13300 10500 14478
rect 9996 13244 10500 13300
rect 10668 14530 10724 14542
rect 10668 14478 10670 14530
rect 10722 14478 10724 14530
rect 9996 12962 10052 13244
rect 10668 13074 10724 14478
rect 11004 14530 11060 14700
rect 11004 14478 11006 14530
rect 11058 14478 11060 14530
rect 11004 14466 11060 14478
rect 11228 14644 11284 14654
rect 11228 14418 11284 14588
rect 11228 14366 11230 14418
rect 11282 14366 11284 14418
rect 11228 14354 11284 14366
rect 11340 14418 11396 14430
rect 11340 14366 11342 14418
rect 11394 14366 11396 14418
rect 11340 13300 11396 14366
rect 11340 13234 11396 13244
rect 10668 13022 10670 13074
rect 10722 13022 10724 13074
rect 10668 13010 10724 13022
rect 11564 13076 11620 13086
rect 9996 12910 9998 12962
rect 10050 12910 10052 12962
rect 9156 12124 9492 12180
rect 9660 12850 9716 12862
rect 9660 12798 9662 12850
rect 9714 12798 9716 12850
rect 9660 12180 9716 12798
rect 9996 12852 10052 12910
rect 10332 12964 10388 12974
rect 10332 12870 10388 12908
rect 11564 12962 11620 13020
rect 11564 12910 11566 12962
rect 11618 12910 11620 12962
rect 9996 12786 10052 12796
rect 10780 12852 10836 12862
rect 10780 12758 10836 12796
rect 10108 12738 10164 12750
rect 10108 12686 10110 12738
rect 10162 12686 10164 12738
rect 9780 12572 10044 12582
rect 9836 12516 9884 12572
rect 9940 12516 9988 12572
rect 9780 12506 10044 12516
rect 9660 12124 9828 12180
rect 9100 12114 9156 12124
rect 9548 12068 9604 12078
rect 9548 12066 9716 12068
rect 9548 12014 9550 12066
rect 9602 12014 9716 12066
rect 9548 12012 9716 12014
rect 9548 12002 9604 12012
rect 8988 11554 9044 11564
rect 8540 11342 8542 11394
rect 8594 11342 8596 11394
rect 8428 10388 8484 10398
rect 8204 9874 8260 9884
rect 8316 10332 8428 10388
rect 7756 9716 7812 9726
rect 7756 9714 8260 9716
rect 7756 9662 7758 9714
rect 7810 9662 8260 9714
rect 7756 9660 8260 9662
rect 7756 9650 7812 9660
rect 8204 9266 8260 9660
rect 8204 9214 8206 9266
rect 8258 9214 8260 9266
rect 8204 9202 8260 9214
rect 7644 8990 7646 9042
rect 7698 8990 7700 9042
rect 7644 8978 7700 8990
rect 8092 9044 8148 9054
rect 8316 9044 8372 10332
rect 8428 10322 8484 10332
rect 8092 9042 8372 9044
rect 8092 8990 8094 9042
rect 8146 8990 8372 9042
rect 8092 8988 8372 8990
rect 8428 9042 8484 9054
rect 8428 8990 8430 9042
rect 8482 8990 8484 9042
rect 8092 8978 8148 8988
rect 8428 8932 8484 8990
rect 8204 8876 8484 8932
rect 8540 8932 8596 11342
rect 9660 11284 9716 12012
rect 9772 11508 9828 12124
rect 10108 12068 10164 12686
rect 10444 12740 10500 12750
rect 10556 12740 10612 12750
rect 10500 12738 10612 12740
rect 10500 12686 10558 12738
rect 10610 12686 10612 12738
rect 10500 12684 10612 12686
rect 10108 12002 10164 12012
rect 10332 12180 10388 12190
rect 9772 11442 9828 11452
rect 9884 11620 9940 11630
rect 9884 11506 9940 11564
rect 9884 11454 9886 11506
rect 9938 11454 9940 11506
rect 9884 11442 9940 11454
rect 9100 11170 9156 11182
rect 9100 11118 9102 11170
rect 9154 11118 9156 11170
rect 9100 10612 9156 11118
rect 9436 11172 9492 11182
rect 9436 11078 9492 11116
rect 9660 10834 9716 11228
rect 10332 11172 10388 12124
rect 10444 11394 10500 12684
rect 10556 12674 10612 12684
rect 11004 12738 11060 12750
rect 11004 12686 11006 12738
rect 11058 12686 11060 12738
rect 10556 11508 10612 11518
rect 10556 11414 10612 11452
rect 10444 11342 10446 11394
rect 10498 11342 10500 11394
rect 10444 11330 10500 11342
rect 11004 11396 11060 12686
rect 11564 12628 11620 12910
rect 11564 12562 11620 12572
rect 11676 12516 11732 16156
rect 11788 14644 11844 14654
rect 11788 14550 11844 14588
rect 12460 13636 12516 13646
rect 12796 13636 12852 17052
rect 12908 16212 12964 16222
rect 13020 16212 13076 18732
rect 13132 18450 13188 18462
rect 13132 18398 13134 18450
rect 13186 18398 13188 18450
rect 13132 18340 13188 18398
rect 13132 18274 13188 18284
rect 13356 17668 13412 18956
rect 13468 19010 13524 19022
rect 13468 18958 13470 19010
rect 13522 18958 13524 19010
rect 13468 18564 13524 18958
rect 13580 18676 13636 21308
rect 13916 21028 13972 21532
rect 14064 21196 14328 21206
rect 14120 21140 14168 21196
rect 14224 21140 14272 21196
rect 14064 21130 14328 21140
rect 13916 20972 14308 21028
rect 13804 20804 13860 20814
rect 13804 20710 13860 20748
rect 13692 19460 13748 19470
rect 13692 19124 13748 19404
rect 13692 19030 13748 19068
rect 13804 19122 13860 19134
rect 13804 19070 13806 19122
rect 13858 19070 13860 19122
rect 13804 18900 13860 19070
rect 13804 18834 13860 18844
rect 13580 18620 13748 18676
rect 13468 18498 13524 18508
rect 13580 18452 13636 18462
rect 13580 18358 13636 18396
rect 13468 17668 13524 17678
rect 13356 17666 13524 17668
rect 13356 17614 13470 17666
rect 13522 17614 13524 17666
rect 13356 17612 13524 17614
rect 13468 17602 13524 17612
rect 13580 17442 13636 17454
rect 13580 17390 13582 17442
rect 13634 17390 13636 17442
rect 13580 16996 13636 17390
rect 13580 16930 13636 16940
rect 12908 16210 13076 16212
rect 12908 16158 12910 16210
rect 12962 16158 13076 16210
rect 12908 16156 13076 16158
rect 13244 16884 13300 16894
rect 12908 16146 12964 16156
rect 13244 15538 13300 16828
rect 13580 15988 13636 15998
rect 13692 15988 13748 18620
rect 13916 18450 13972 20972
rect 14252 20914 14308 20972
rect 14252 20862 14254 20914
rect 14306 20862 14308 20914
rect 14252 20850 14308 20862
rect 14064 19628 14328 19638
rect 14120 19572 14168 19628
rect 14224 19572 14272 19628
rect 14064 19562 14328 19572
rect 14476 19460 14532 21756
rect 14588 21028 14644 25228
rect 15036 25218 15092 25228
rect 14812 24948 14868 24958
rect 15148 24948 15204 26908
rect 15260 26962 15316 27132
rect 15372 27186 15428 27806
rect 15484 27748 15540 27758
rect 15484 27298 15540 27692
rect 15484 27246 15486 27298
rect 15538 27246 15540 27298
rect 15484 27234 15540 27246
rect 15372 27134 15374 27186
rect 15426 27134 15428 27186
rect 15372 27122 15428 27134
rect 15260 26910 15262 26962
rect 15314 26910 15316 26962
rect 15260 26898 15316 26910
rect 15596 26908 15652 28140
rect 16268 28084 16324 29148
rect 16380 28980 16436 29596
rect 16380 28914 16436 28924
rect 16492 28866 16548 32510
rect 17500 32564 17556 33292
rect 17612 33012 17668 33404
rect 17724 33236 17780 33246
rect 17724 33234 17892 33236
rect 17724 33182 17726 33234
rect 17778 33182 17892 33234
rect 17724 33180 17892 33182
rect 17724 33170 17780 33180
rect 17612 32956 17780 33012
rect 17388 31892 17444 31902
rect 16716 31108 16772 31118
rect 16716 31014 16772 31052
rect 17388 31108 17444 31836
rect 17500 31778 17556 32508
rect 17612 32562 17668 32574
rect 17612 32510 17614 32562
rect 17666 32510 17668 32562
rect 17612 32452 17668 32510
rect 17612 32386 17668 32396
rect 17500 31726 17502 31778
rect 17554 31726 17556 31778
rect 17500 31714 17556 31726
rect 17724 31780 17780 32956
rect 17724 31714 17780 31724
rect 17500 31332 17556 31342
rect 17556 31276 17668 31332
rect 17500 31266 17556 31276
rect 17388 30994 17444 31052
rect 17612 31108 17668 31276
rect 17612 31014 17668 31052
rect 17388 30942 17390 30994
rect 17442 30942 17444 30994
rect 17388 30930 17444 30942
rect 17500 30996 17556 31006
rect 16828 30770 16884 30782
rect 16828 30718 16830 30770
rect 16882 30718 16884 30770
rect 16828 29652 16884 30718
rect 17500 30210 17556 30940
rect 17724 30994 17780 31006
rect 17724 30942 17726 30994
rect 17778 30942 17780 30994
rect 17724 30436 17780 30942
rect 17724 30370 17780 30380
rect 17500 30158 17502 30210
rect 17554 30158 17556 30210
rect 17500 30146 17556 30158
rect 16828 29586 16884 29596
rect 17836 29650 17892 33180
rect 18348 32956 18612 32966
rect 18404 32900 18452 32956
rect 18508 32900 18556 32956
rect 18348 32890 18612 32900
rect 18620 32788 18676 32798
rect 18732 32788 18788 33516
rect 18620 32786 18788 32788
rect 18620 32734 18622 32786
rect 18674 32734 18788 32786
rect 18620 32732 18788 32734
rect 18620 32722 18676 32732
rect 18284 32676 18340 32686
rect 18284 31890 18340 32620
rect 18284 31838 18286 31890
rect 18338 31838 18340 31890
rect 18284 31826 18340 31838
rect 18844 31780 18900 31790
rect 18348 31388 18612 31398
rect 18404 31332 18452 31388
rect 18508 31332 18556 31388
rect 18348 31322 18612 31332
rect 17948 31220 18004 31230
rect 17948 30994 18004 31164
rect 18732 31108 18788 31118
rect 18732 31014 18788 31052
rect 17948 30942 17950 30994
rect 18002 30942 18004 30994
rect 17948 30930 18004 30942
rect 18396 30996 18452 31006
rect 18396 30902 18452 30940
rect 18620 30772 18676 30782
rect 18508 30770 18676 30772
rect 18508 30718 18622 30770
rect 18674 30718 18676 30770
rect 18508 30716 18676 30718
rect 18508 30324 18564 30716
rect 18620 30706 18676 30716
rect 17836 29598 17838 29650
rect 17890 29598 17892 29650
rect 17836 29586 17892 29598
rect 18172 30268 18564 30324
rect 18844 30322 18900 31724
rect 19516 31220 19572 36200
rect 20636 33572 20692 36200
rect 20636 33506 20692 33516
rect 19516 31154 19572 31164
rect 19852 33458 19908 33470
rect 19852 33406 19854 33458
rect 19906 33406 19908 33458
rect 19852 32788 19908 33406
rect 19068 31108 19124 31118
rect 18844 30270 18846 30322
rect 18898 30270 18900 30322
rect 16940 29540 16996 29550
rect 18172 29540 18228 30268
rect 18844 30258 18900 30270
rect 18956 31052 19068 31108
rect 18348 29820 18612 29830
rect 18404 29764 18452 29820
rect 18508 29764 18556 29820
rect 18348 29754 18612 29764
rect 18284 29540 18340 29550
rect 18172 29538 18340 29540
rect 18172 29486 18286 29538
rect 18338 29486 18340 29538
rect 18172 29484 18340 29486
rect 16828 29428 16884 29438
rect 16940 29428 16996 29484
rect 18284 29474 18340 29484
rect 18844 29540 18900 29550
rect 18844 29446 18900 29484
rect 16828 29426 16996 29428
rect 16828 29374 16830 29426
rect 16882 29374 16996 29426
rect 16828 29372 16996 29374
rect 17276 29428 17332 29438
rect 16604 29316 16660 29326
rect 16604 29222 16660 29260
rect 16492 28814 16494 28866
rect 16546 28814 16548 28866
rect 16492 28802 16548 28814
rect 16604 29092 16660 29102
rect 16156 28028 16324 28084
rect 16044 27970 16100 27982
rect 16044 27918 16046 27970
rect 16098 27918 16100 27970
rect 15820 27858 15876 27870
rect 15820 27806 15822 27858
rect 15874 27806 15876 27858
rect 15372 26852 15652 26908
rect 15708 27300 15764 27310
rect 15260 26292 15316 26302
rect 15260 26198 15316 26236
rect 15260 25508 15316 25518
rect 15372 25508 15428 26852
rect 15708 26516 15764 27244
rect 15708 26178 15764 26460
rect 15820 26404 15876 27806
rect 16044 27748 16100 27918
rect 16044 27682 16100 27692
rect 16156 27186 16212 28028
rect 16380 27970 16436 27982
rect 16380 27918 16382 27970
rect 16434 27918 16436 27970
rect 16156 27134 16158 27186
rect 16210 27134 16212 27186
rect 16156 26908 16212 27134
rect 15820 26338 15876 26348
rect 16044 26852 16212 26908
rect 16268 27858 16324 27870
rect 16268 27806 16270 27858
rect 16322 27806 16324 27858
rect 15708 26126 15710 26178
rect 15762 26126 15764 26178
rect 15708 26114 15764 26126
rect 15260 25506 15428 25508
rect 15260 25454 15262 25506
rect 15314 25454 15428 25506
rect 15260 25452 15428 25454
rect 15484 25844 15540 25854
rect 15260 25442 15316 25452
rect 15484 25284 15540 25788
rect 15372 25228 15540 25284
rect 15260 24948 15316 24958
rect 15148 24946 15316 24948
rect 15148 24894 15262 24946
rect 15314 24894 15316 24946
rect 15148 24892 15316 24894
rect 14812 24834 14868 24892
rect 15260 24882 15316 24892
rect 14812 24782 14814 24834
rect 14866 24782 14868 24834
rect 14812 24770 14868 24782
rect 14924 24834 14980 24846
rect 14924 24782 14926 24834
rect 14978 24782 14980 24834
rect 14700 21476 14756 21486
rect 14700 21382 14756 21420
rect 14588 20972 14756 21028
rect 14588 20804 14644 20814
rect 14588 20710 14644 20748
rect 14700 19796 14756 20972
rect 14924 20916 14980 24782
rect 15148 24724 15204 24734
rect 15372 24724 15428 25228
rect 15148 24722 15428 24724
rect 15148 24670 15150 24722
rect 15202 24670 15428 24722
rect 15148 24668 15428 24670
rect 15484 24834 15540 24846
rect 15484 24782 15486 24834
rect 15538 24782 15540 24834
rect 15148 24658 15204 24668
rect 15484 21812 15540 24782
rect 15596 24724 15652 24734
rect 15596 24630 15652 24668
rect 15708 23826 15764 23838
rect 15708 23774 15710 23826
rect 15762 23774 15764 23826
rect 15708 22484 15764 23774
rect 16044 22596 16100 26852
rect 16156 26292 16212 26302
rect 16156 24722 16212 26236
rect 16268 25844 16324 27806
rect 16380 27412 16436 27918
rect 16604 27746 16660 29036
rect 16828 28084 16884 29372
rect 17276 29334 17332 29372
rect 17612 29426 17668 29438
rect 17836 29428 17892 29438
rect 17612 29374 17614 29426
rect 17666 29374 17668 29426
rect 17164 29204 17220 29214
rect 17052 29092 17108 29102
rect 17052 28642 17108 29036
rect 17052 28590 17054 28642
rect 17106 28590 17108 28642
rect 17052 28578 17108 28590
rect 17164 28642 17220 29148
rect 17164 28590 17166 28642
rect 17218 28590 17220 28642
rect 17164 28578 17220 28590
rect 17388 29204 17444 29214
rect 16940 28532 16996 28542
rect 16940 28438 16996 28476
rect 17388 28420 17444 29148
rect 17500 28756 17556 28766
rect 17500 28642 17556 28700
rect 17500 28590 17502 28642
rect 17554 28590 17556 28642
rect 17500 28578 17556 28590
rect 17052 28364 17444 28420
rect 16828 28028 16996 28084
rect 16604 27694 16606 27746
rect 16658 27694 16660 27746
rect 16604 27682 16660 27694
rect 16380 27346 16436 27356
rect 16828 26964 16884 27002
rect 16828 26898 16884 26908
rect 16940 26740 16996 28028
rect 16940 26674 16996 26684
rect 16492 26402 16548 26414
rect 16492 26350 16494 26402
rect 16546 26350 16548 26402
rect 16492 26180 16548 26350
rect 16492 26114 16548 26124
rect 16716 26292 16772 26302
rect 16268 25778 16324 25788
rect 16716 25732 16772 26236
rect 16716 25666 16772 25676
rect 17052 25508 17108 28364
rect 17500 28308 17556 28318
rect 17388 27972 17444 27982
rect 17388 27878 17444 27916
rect 17500 27748 17556 28252
rect 17612 28196 17668 29374
rect 17724 29372 17836 29428
rect 17724 29316 17780 29372
rect 17836 29362 17892 29372
rect 18620 29428 18676 29438
rect 18620 29334 18676 29372
rect 17724 28754 17780 29260
rect 18060 29316 18116 29326
rect 17836 29204 17892 29242
rect 18060 29222 18116 29260
rect 18732 29314 18788 29326
rect 18732 29262 18734 29314
rect 18786 29262 18788 29314
rect 17836 29138 17892 29148
rect 17724 28702 17726 28754
rect 17778 28702 17780 28754
rect 17724 28690 17780 28702
rect 17836 28980 17892 28990
rect 17836 28642 17892 28924
rect 17836 28590 17838 28642
rect 17890 28590 17892 28642
rect 17836 28578 17892 28590
rect 18060 28642 18116 28654
rect 18060 28590 18062 28642
rect 18114 28590 18116 28642
rect 17612 28130 17668 28140
rect 17724 28308 17780 28318
rect 17724 28026 17780 28252
rect 17612 27970 17668 27982
rect 17612 27918 17614 27970
rect 17666 27918 17668 27970
rect 17724 27974 17726 28026
rect 17778 27974 17780 28026
rect 17724 27962 17780 27974
rect 17612 27860 17668 27918
rect 17724 27860 17780 27870
rect 17612 27804 17724 27860
rect 17724 27794 17780 27804
rect 17500 27692 17668 27748
rect 17500 27076 17556 27086
rect 17164 26962 17220 26974
rect 17164 26910 17166 26962
rect 17218 26910 17220 26962
rect 17164 26404 17220 26910
rect 17164 26338 17220 26348
rect 17276 26964 17332 26974
rect 17052 25452 17220 25508
rect 17052 25282 17108 25294
rect 17052 25230 17054 25282
rect 17106 25230 17108 25282
rect 16156 24670 16158 24722
rect 16210 24670 16212 24722
rect 16156 24658 16212 24670
rect 16716 24724 16772 24734
rect 16716 24630 16772 24668
rect 17052 24724 17108 25230
rect 17052 24658 17108 24668
rect 17164 24612 17220 25452
rect 17164 24546 17220 24556
rect 17164 23380 17220 23390
rect 16828 23324 17164 23380
rect 16044 22540 16212 22596
rect 15708 22482 16100 22484
rect 15708 22430 15710 22482
rect 15762 22430 16100 22482
rect 15708 22428 16100 22430
rect 15708 22418 15764 22428
rect 16044 22372 16100 22428
rect 16044 22278 16100 22316
rect 15484 21746 15540 21756
rect 14700 19730 14756 19740
rect 14812 20860 14980 20916
rect 15260 21364 15316 21374
rect 14252 19404 14532 19460
rect 14812 19460 14868 20860
rect 14924 20692 14980 20702
rect 14924 20598 14980 20636
rect 15260 20244 15316 21308
rect 15708 20692 15764 20702
rect 15764 20636 15876 20692
rect 15708 20626 15764 20636
rect 14924 20130 14980 20142
rect 14924 20078 14926 20130
rect 14978 20078 14980 20130
rect 14924 19460 14980 20078
rect 15260 20130 15316 20188
rect 15260 20078 15262 20130
rect 15314 20078 15316 20130
rect 15260 20066 15316 20078
rect 15708 20020 15764 20030
rect 15372 20018 15764 20020
rect 15372 19966 15710 20018
rect 15762 19966 15764 20018
rect 15372 19964 15764 19966
rect 14924 19404 15092 19460
rect 14140 19236 14196 19246
rect 14140 19142 14196 19180
rect 14252 19122 14308 19404
rect 14252 19070 14254 19122
rect 14306 19070 14308 19122
rect 14252 19058 14308 19070
rect 14364 18788 14420 19404
rect 14812 19394 14868 19404
rect 14476 19236 14532 19246
rect 14924 19236 14980 19246
rect 14476 19234 14980 19236
rect 14476 19182 14478 19234
rect 14530 19182 14926 19234
rect 14978 19182 14980 19234
rect 14476 19180 14980 19182
rect 14476 19170 14532 19180
rect 14924 19170 14980 19180
rect 15036 19236 15092 19404
rect 14700 19012 14756 19022
rect 14588 18900 14644 18910
rect 14364 18732 14532 18788
rect 13916 18398 13918 18450
rect 13970 18398 13972 18450
rect 13804 17556 13860 17566
rect 13804 17462 13860 17500
rect 13916 16884 13972 18398
rect 14064 18060 14328 18070
rect 14120 18004 14168 18060
rect 14224 18004 14272 18060
rect 14064 17994 14328 18004
rect 14028 17668 14084 17678
rect 14028 17574 14084 17612
rect 14252 17556 14308 17566
rect 14252 17462 14308 17500
rect 14476 17554 14532 18732
rect 14588 17666 14644 18844
rect 14700 18450 14756 18956
rect 14924 18900 14980 18910
rect 15036 18900 15092 19180
rect 15372 19234 15428 19964
rect 15708 19954 15764 19964
rect 15820 19796 15876 20636
rect 15932 20690 15988 20702
rect 15932 20638 15934 20690
rect 15986 20638 15988 20690
rect 15932 20356 15988 20638
rect 16044 20578 16100 20590
rect 16044 20526 16046 20578
rect 16098 20526 16100 20578
rect 16044 20468 16100 20526
rect 16156 20580 16212 22540
rect 16828 22482 16884 23324
rect 17164 23314 17220 23324
rect 16828 22430 16830 22482
rect 16882 22430 16884 22482
rect 16828 22418 16884 22430
rect 16828 22036 16884 22046
rect 16716 21980 16828 22036
rect 16604 21476 16660 21486
rect 16604 20914 16660 21420
rect 16604 20862 16606 20914
rect 16658 20862 16660 20914
rect 16604 20850 16660 20862
rect 16268 20804 16324 20814
rect 16492 20804 16548 20814
rect 16268 20802 16548 20804
rect 16268 20750 16270 20802
rect 16322 20750 16494 20802
rect 16546 20750 16548 20802
rect 16268 20748 16548 20750
rect 16268 20738 16324 20748
rect 16492 20738 16548 20748
rect 16716 20802 16772 21980
rect 16828 21970 16884 21980
rect 16828 21474 16884 21486
rect 16828 21422 16830 21474
rect 16882 21422 16884 21474
rect 16828 21364 16884 21422
rect 17052 21364 17108 21374
rect 16828 21308 17052 21364
rect 17052 21298 17108 21308
rect 16716 20750 16718 20802
rect 16770 20750 16772 20802
rect 16716 20738 16772 20750
rect 16940 20802 16996 20814
rect 16940 20750 16942 20802
rect 16994 20750 16996 20802
rect 16940 20692 16996 20750
rect 16940 20626 16996 20636
rect 16156 20524 16436 20580
rect 16044 20412 16324 20468
rect 15932 20300 16212 20356
rect 15932 20130 15988 20142
rect 15932 20078 15934 20130
rect 15986 20078 15988 20130
rect 15932 20020 15988 20078
rect 16156 20132 16212 20300
rect 16156 20066 16212 20076
rect 15932 19954 15988 19964
rect 16044 20018 16100 20030
rect 16044 19966 16046 20018
rect 16098 19966 16100 20018
rect 15372 19182 15374 19234
rect 15426 19182 15428 19234
rect 15372 19170 15428 19182
rect 15596 19740 15876 19796
rect 15596 19234 15652 19740
rect 15932 19460 15988 19470
rect 15596 19182 15598 19234
rect 15650 19182 15652 19234
rect 15148 19012 15204 19022
rect 15148 18918 15204 18956
rect 14980 18844 15092 18900
rect 14924 18834 14980 18844
rect 14700 18398 14702 18450
rect 14754 18398 14756 18450
rect 14700 18386 14756 18398
rect 15596 18340 15652 19182
rect 15820 19404 15932 19460
rect 15820 19012 15876 19404
rect 15932 19394 15988 19404
rect 15932 19236 15988 19246
rect 16044 19236 16100 19966
rect 16268 19460 16324 20412
rect 16380 19460 16436 20524
rect 17276 20356 17332 26908
rect 17500 26850 17556 27020
rect 17500 26798 17502 26850
rect 17554 26798 17556 26850
rect 17500 26786 17556 26798
rect 17388 26740 17444 26750
rect 17388 26514 17444 26684
rect 17388 26462 17390 26514
rect 17442 26462 17444 26514
rect 17388 26450 17444 26462
rect 17612 25732 17668 27692
rect 18060 27300 18116 28590
rect 18732 28644 18788 29262
rect 18956 28980 19012 31052
rect 19068 31014 19124 31052
rect 19404 30996 19460 31006
rect 19404 30902 19460 30940
rect 19852 30994 19908 32732
rect 20972 33346 21028 33358
rect 20972 33294 20974 33346
rect 21026 33294 21028 33346
rect 20524 32564 20580 32574
rect 20524 32470 20580 32508
rect 20972 32564 21028 33294
rect 21644 33236 21700 33246
rect 20972 32498 21028 32508
rect 21532 33234 21700 33236
rect 21532 33182 21646 33234
rect 21698 33182 21700 33234
rect 21532 33180 21700 33182
rect 21308 32452 21364 32462
rect 21084 32450 21364 32452
rect 21084 32398 21310 32450
rect 21362 32398 21364 32450
rect 21084 32396 21364 32398
rect 20412 31892 20468 31902
rect 20412 31798 20468 31836
rect 19852 30942 19854 30994
rect 19906 30942 19908 30994
rect 19852 30930 19908 30942
rect 20076 31668 20132 31678
rect 19404 30324 19460 30334
rect 19068 29652 19124 29662
rect 19068 29558 19124 29596
rect 18956 28914 19012 28924
rect 19292 28756 19348 28766
rect 19180 28700 19292 28756
rect 18732 28578 18788 28588
rect 18956 28642 19012 28654
rect 18956 28590 18958 28642
rect 19010 28590 19012 28642
rect 18956 28420 19012 28590
rect 18956 28354 19012 28364
rect 19068 28418 19124 28430
rect 19068 28366 19070 28418
rect 19122 28366 19124 28418
rect 18172 28308 18228 28318
rect 18844 28308 18900 28318
rect 18172 27860 18228 28252
rect 18348 28252 18612 28262
rect 18404 28196 18452 28252
rect 18508 28196 18556 28252
rect 18348 28186 18612 28196
rect 18732 28252 18844 28308
rect 18732 27970 18788 28252
rect 18844 28242 18900 28252
rect 19068 28084 19124 28366
rect 18732 27918 18734 27970
rect 18786 27918 18788 27970
rect 18732 27906 18788 27918
rect 18844 28028 19124 28084
rect 18172 27858 18564 27860
rect 18172 27806 18174 27858
rect 18226 27806 18564 27858
rect 18172 27804 18564 27806
rect 18172 27794 18228 27804
rect 18396 27636 18452 27646
rect 17724 27244 18116 27300
rect 17724 26516 17780 27244
rect 17836 27076 17892 27086
rect 18060 27076 18116 27244
rect 18284 27634 18452 27636
rect 18284 27582 18398 27634
rect 18450 27582 18452 27634
rect 18284 27580 18452 27582
rect 18284 27300 18340 27580
rect 18396 27570 18452 27580
rect 18508 27524 18564 27804
rect 18844 27634 18900 28028
rect 19068 27748 19124 27758
rect 18844 27582 18846 27634
rect 18898 27582 18900 27634
rect 18844 27570 18900 27582
rect 18956 27634 19012 27646
rect 18956 27582 18958 27634
rect 19010 27582 19012 27634
rect 18508 27468 18676 27524
rect 18284 27234 18340 27244
rect 18508 27300 18564 27310
rect 18172 27076 18228 27086
rect 18060 27074 18228 27076
rect 18060 27022 18174 27074
rect 18226 27022 18228 27074
rect 18060 27020 18228 27022
rect 17836 26906 17892 27020
rect 18172 27010 18228 27020
rect 18508 27074 18564 27244
rect 18508 27022 18510 27074
rect 18562 27022 18564 27074
rect 18508 27010 18564 27022
rect 18620 27074 18676 27468
rect 18956 27300 19012 27582
rect 18956 27234 19012 27244
rect 18844 27188 18900 27198
rect 18620 27022 18622 27074
rect 18674 27022 18676 27074
rect 18620 27010 18676 27022
rect 18732 27076 18788 27086
rect 17836 26854 17838 26906
rect 17890 26854 17892 26906
rect 18284 26964 18340 26974
rect 18284 26870 18340 26908
rect 17836 26842 17892 26854
rect 18348 26684 18612 26694
rect 18404 26628 18452 26684
rect 18508 26628 18556 26684
rect 18348 26618 18612 26628
rect 18396 26516 18452 26526
rect 17724 26460 17892 26516
rect 17724 26292 17780 26302
rect 17724 26198 17780 26236
rect 17836 25844 17892 26460
rect 18396 26422 18452 26460
rect 18732 26514 18788 27020
rect 18844 26962 18900 27132
rect 18956 27076 19012 27086
rect 19068 27076 19124 27692
rect 18956 27074 19124 27076
rect 18956 27022 18958 27074
rect 19010 27022 19124 27074
rect 18956 27020 19124 27022
rect 18956 27010 19012 27020
rect 18844 26910 18846 26962
rect 18898 26910 18900 26962
rect 18844 26898 18900 26910
rect 19180 26908 19236 28700
rect 19292 28690 19348 28700
rect 19404 28754 19460 30268
rect 19404 28702 19406 28754
rect 19458 28702 19460 28754
rect 19404 28690 19460 28702
rect 19740 28868 19796 28878
rect 19516 28644 19572 28654
rect 19516 28642 19684 28644
rect 19516 28590 19518 28642
rect 19570 28590 19684 28642
rect 19516 28588 19684 28590
rect 19516 28578 19572 28588
rect 19292 28418 19348 28430
rect 19292 28366 19294 28418
rect 19346 28366 19348 28418
rect 19292 28308 19348 28366
rect 19292 28242 19348 28252
rect 19516 28196 19572 28206
rect 19404 28140 19516 28196
rect 19404 28082 19460 28140
rect 19516 28130 19572 28140
rect 19404 28030 19406 28082
rect 19458 28030 19460 28082
rect 19404 27860 19460 28030
rect 19404 27794 19460 27804
rect 19516 27972 19572 27982
rect 19516 27076 19572 27916
rect 19628 27300 19684 28588
rect 19740 28082 19796 28812
rect 20076 28642 20132 31612
rect 20636 31556 20692 31566
rect 20188 30996 20244 31006
rect 20188 29538 20244 30940
rect 20524 30884 20580 30894
rect 20412 30324 20468 30334
rect 20412 30230 20468 30268
rect 20188 29486 20190 29538
rect 20242 29486 20244 29538
rect 20188 29474 20244 29486
rect 20412 29876 20468 29886
rect 20076 28590 20078 28642
rect 20130 28590 20132 28642
rect 20076 28578 20132 28590
rect 20188 28642 20244 28654
rect 20188 28590 20190 28642
rect 20242 28590 20244 28642
rect 19740 28030 19742 28082
rect 19794 28030 19796 28082
rect 19740 27636 19796 28030
rect 19740 27570 19796 27580
rect 19852 28530 19908 28542
rect 19852 28478 19854 28530
rect 19906 28478 19908 28530
rect 19852 27524 19908 28478
rect 19740 27300 19796 27310
rect 19628 27298 19796 27300
rect 19628 27246 19742 27298
rect 19794 27246 19796 27298
rect 19628 27244 19796 27246
rect 19740 27234 19796 27244
rect 19628 27076 19684 27086
rect 19516 27074 19684 27076
rect 19516 27022 19630 27074
rect 19682 27022 19684 27074
rect 19516 27020 19684 27022
rect 19628 27010 19684 27020
rect 19852 27076 19908 27468
rect 19852 27010 19908 27020
rect 19964 28532 20020 28542
rect 18732 26462 18734 26514
rect 18786 26462 18788 26514
rect 18732 26450 18788 26462
rect 18956 26852 19236 26908
rect 19740 26964 19796 27002
rect 19740 26898 19796 26908
rect 19628 26852 19684 26862
rect 18060 26292 18116 26302
rect 18172 26292 18228 26302
rect 18116 26290 18340 26292
rect 18116 26238 18174 26290
rect 18226 26238 18340 26290
rect 18116 26236 18340 26238
rect 18060 26226 18116 26236
rect 18172 26226 18228 26236
rect 17500 25676 17668 25732
rect 17724 25788 17892 25844
rect 17388 25508 17444 25518
rect 17388 25414 17444 25452
rect 17388 24948 17444 24958
rect 17500 24948 17556 25676
rect 17724 25620 17780 25788
rect 17612 25508 17668 25518
rect 17724 25508 17780 25564
rect 17948 25620 18004 25630
rect 17948 25618 18228 25620
rect 17948 25566 17950 25618
rect 18002 25566 18228 25618
rect 17948 25564 18228 25566
rect 17948 25554 18004 25564
rect 17612 25506 17780 25508
rect 17612 25454 17614 25506
rect 17666 25454 17780 25506
rect 17612 25452 17780 25454
rect 18172 25506 18228 25564
rect 18172 25454 18174 25506
rect 18226 25454 18228 25506
rect 17612 25442 17668 25452
rect 18172 25442 18228 25454
rect 18284 25284 18340 26236
rect 18508 25844 18564 25854
rect 18508 25396 18564 25788
rect 18732 25620 18788 25630
rect 18956 25620 19012 26852
rect 19516 26796 19628 26852
rect 18732 25618 19012 25620
rect 18732 25566 18734 25618
rect 18786 25566 19012 25618
rect 18732 25564 19012 25566
rect 19068 26404 19124 26414
rect 19068 26290 19124 26348
rect 19068 26238 19070 26290
rect 19122 26238 19124 26290
rect 18732 25554 18788 25564
rect 18508 25330 18564 25340
rect 18844 25396 18900 25406
rect 18844 25302 18900 25340
rect 18396 25284 18452 25294
rect 18284 25228 18396 25284
rect 18396 25218 18452 25228
rect 18620 25284 18676 25294
rect 18620 25282 18788 25284
rect 18620 25230 18622 25282
rect 18674 25230 18788 25282
rect 18620 25228 18788 25230
rect 18620 25218 18676 25228
rect 18348 25116 18612 25126
rect 18404 25060 18452 25116
rect 18508 25060 18556 25116
rect 18348 25050 18612 25060
rect 17388 24946 17556 24948
rect 17388 24894 17390 24946
rect 17442 24894 17556 24946
rect 17388 24892 17556 24894
rect 17388 24882 17444 24892
rect 17500 23154 17556 24892
rect 17724 24722 17780 24734
rect 17724 24670 17726 24722
rect 17778 24670 17780 24722
rect 17724 24612 17780 24670
rect 17724 24546 17780 24556
rect 18172 24612 18228 24622
rect 18172 24518 18228 24556
rect 17948 23828 18004 23838
rect 18732 23828 18788 25228
rect 17836 23772 17948 23828
rect 17724 23380 17780 23418
rect 17724 23314 17780 23324
rect 17500 23102 17502 23154
rect 17554 23102 17556 23154
rect 17500 23090 17556 23102
rect 17724 23156 17780 23166
rect 17836 23156 17892 23772
rect 17948 23762 18004 23772
rect 18172 23772 18788 23828
rect 18844 24612 18900 24622
rect 18172 23380 18228 23772
rect 18732 23604 18788 23614
rect 18348 23548 18612 23558
rect 18404 23492 18452 23548
rect 18508 23492 18556 23548
rect 18348 23482 18612 23492
rect 18396 23380 18452 23390
rect 17724 23154 17892 23156
rect 17724 23102 17726 23154
rect 17778 23102 17892 23154
rect 17724 23100 17892 23102
rect 17948 23378 18452 23380
rect 17948 23326 18398 23378
rect 18450 23326 18452 23378
rect 17948 23324 18452 23326
rect 17724 23090 17780 23100
rect 17500 22372 17556 22382
rect 17500 21810 17556 22316
rect 17500 21758 17502 21810
rect 17554 21758 17556 21810
rect 17500 21746 17556 21758
rect 17836 21476 17892 21486
rect 17836 21382 17892 21420
rect 17948 21364 18004 23324
rect 18396 23314 18452 23324
rect 18060 23154 18116 23166
rect 18060 23102 18062 23154
rect 18114 23102 18116 23154
rect 18060 22596 18116 23102
rect 18060 22530 18116 22540
rect 18172 23154 18228 23166
rect 18172 23102 18174 23154
rect 18226 23102 18228 23154
rect 18172 22036 18228 23102
rect 18508 23156 18564 23166
rect 18732 23156 18788 23548
rect 18508 23154 18788 23156
rect 18508 23102 18510 23154
rect 18562 23102 18788 23154
rect 18508 23100 18788 23102
rect 18508 23090 18564 23100
rect 18172 21970 18228 21980
rect 18348 21980 18612 21990
rect 18404 21924 18452 21980
rect 18508 21924 18556 21980
rect 18348 21914 18612 21924
rect 17836 20692 17892 20702
rect 17836 20598 17892 20636
rect 17948 20468 18004 21308
rect 18732 21812 18788 23100
rect 18844 22260 18900 24556
rect 19068 24164 19124 26238
rect 19180 25620 19236 25630
rect 19180 25526 19236 25564
rect 19404 25508 19460 25518
rect 19404 25414 19460 25452
rect 19516 25396 19572 26796
rect 19628 26786 19684 26796
rect 19740 26628 19796 26638
rect 19740 26402 19796 26572
rect 19740 26350 19742 26402
rect 19794 26350 19796 26402
rect 19740 26180 19796 26350
rect 19628 25732 19684 25742
rect 19628 25638 19684 25676
rect 19740 25508 19796 26124
rect 19740 25442 19796 25452
rect 19516 24948 19572 25340
rect 19628 24948 19684 24958
rect 19516 24946 19684 24948
rect 19516 24894 19630 24946
rect 19682 24894 19684 24946
rect 19516 24892 19684 24894
rect 19628 24882 19684 24892
rect 19740 24948 19796 24958
rect 19964 24948 20020 28476
rect 20188 28196 20244 28590
rect 20300 28420 20356 28430
rect 20300 28326 20356 28364
rect 20076 28140 20244 28196
rect 20076 27970 20132 28140
rect 20412 28084 20468 29820
rect 20524 28642 20580 30828
rect 20636 29426 20692 31500
rect 20748 31220 20804 31230
rect 20748 31126 20804 31164
rect 21084 31108 21140 32396
rect 21308 32386 21364 32396
rect 20860 31052 21140 31108
rect 21196 31780 21252 31790
rect 20748 30436 20804 30446
rect 20860 30436 20916 31052
rect 20748 30434 20916 30436
rect 20748 30382 20750 30434
rect 20802 30382 20916 30434
rect 20748 30380 20916 30382
rect 20748 30370 20804 30380
rect 20748 30212 20804 30222
rect 20804 30156 21028 30212
rect 20748 30118 20804 30156
rect 20636 29374 20638 29426
rect 20690 29374 20692 29426
rect 20636 29362 20692 29374
rect 20524 28590 20526 28642
rect 20578 28590 20580 28642
rect 20524 28578 20580 28590
rect 20860 29202 20916 29214
rect 20860 29150 20862 29202
rect 20914 29150 20916 29202
rect 20076 27918 20078 27970
rect 20130 27918 20132 27970
rect 20076 27906 20132 27918
rect 20188 28028 20468 28084
rect 20188 27748 20244 28028
rect 20748 27972 20804 27982
rect 20076 27692 20244 27748
rect 20412 27858 20468 27870
rect 20412 27806 20414 27858
rect 20466 27806 20468 27858
rect 20076 27412 20132 27692
rect 20412 27636 20468 27806
rect 20636 27858 20692 27870
rect 20636 27806 20638 27858
rect 20690 27806 20692 27858
rect 20524 27748 20580 27758
rect 20524 27654 20580 27692
rect 20412 27570 20468 27580
rect 20636 27412 20692 27806
rect 20076 27076 20132 27356
rect 20076 27010 20132 27020
rect 20300 27356 20692 27412
rect 20188 26962 20244 26974
rect 20188 26910 20190 26962
rect 20242 26910 20244 26962
rect 20188 26908 20244 26910
rect 20076 26852 20244 26908
rect 20076 26628 20132 26852
rect 20076 26562 20132 26572
rect 20188 26740 20244 26750
rect 20076 26404 20132 26414
rect 20188 26404 20244 26684
rect 20300 26516 20356 27356
rect 20524 27076 20580 27086
rect 20524 26982 20580 27020
rect 20748 27074 20804 27916
rect 20748 27022 20750 27074
rect 20802 27022 20804 27074
rect 20748 27010 20804 27022
rect 20860 26964 20916 29150
rect 20972 27860 21028 30156
rect 21196 29876 21252 31724
rect 21420 31778 21476 31790
rect 21420 31726 21422 31778
rect 21474 31726 21476 31778
rect 21420 31668 21476 31726
rect 21532 31668 21588 33180
rect 21644 33170 21700 33180
rect 21756 32452 21812 36200
rect 22876 33908 22932 36200
rect 23996 36036 24052 36200
rect 24332 36036 24388 36204
rect 23996 35980 24388 36036
rect 22876 33852 23156 33908
rect 22632 33740 22896 33750
rect 22688 33684 22736 33740
rect 22792 33684 22840 33740
rect 22632 33674 22896 33684
rect 21756 32386 21812 32396
rect 22428 32340 22484 32350
rect 22428 31892 22484 32284
rect 22632 32172 22896 32182
rect 22688 32116 22736 32172
rect 22792 32116 22840 32172
rect 22632 32106 22896 32116
rect 22316 31890 22484 31892
rect 22316 31838 22430 31890
rect 22482 31838 22484 31890
rect 22316 31836 22484 31838
rect 21756 31780 21812 31818
rect 21756 31714 21812 31724
rect 21532 31612 21700 31668
rect 21420 31602 21476 31612
rect 21532 30996 21588 31006
rect 21420 30940 21532 30996
rect 21196 29810 21252 29820
rect 21308 30098 21364 30110
rect 21308 30046 21310 30098
rect 21362 30046 21364 30098
rect 21196 29540 21252 29550
rect 21196 29446 21252 29484
rect 21308 28756 21364 30046
rect 21308 28690 21364 28700
rect 20972 27766 21028 27804
rect 21196 28644 21252 28654
rect 20860 26898 20916 26908
rect 20412 26852 20468 26862
rect 20412 26850 20804 26852
rect 20412 26798 20414 26850
rect 20466 26798 20804 26850
rect 20412 26796 20804 26798
rect 20412 26786 20468 26796
rect 20636 26628 20692 26638
rect 20524 26572 20636 26628
rect 20300 26460 20468 26516
rect 20076 26402 20244 26404
rect 20076 26350 20078 26402
rect 20130 26350 20244 26402
rect 20076 26348 20244 26350
rect 20076 26338 20132 26348
rect 20412 26292 20468 26460
rect 20412 26198 20468 26236
rect 20412 25844 20468 25854
rect 20412 25394 20468 25788
rect 20412 25342 20414 25394
rect 20466 25342 20468 25394
rect 20412 25330 20468 25342
rect 19740 24946 20020 24948
rect 19740 24894 19742 24946
rect 19794 24894 20020 24946
rect 19740 24892 20020 24894
rect 20076 25282 20132 25294
rect 20076 25230 20078 25282
rect 20130 25230 20132 25282
rect 20076 24946 20132 25230
rect 20076 24894 20078 24946
rect 20130 24894 20132 24946
rect 19740 24882 19796 24892
rect 20076 24882 20132 24894
rect 20188 25284 20244 25294
rect 19852 24722 19908 24734
rect 19852 24670 19854 24722
rect 19906 24670 19908 24722
rect 19068 24108 19796 24164
rect 19180 23940 19236 23950
rect 19740 23940 19796 24108
rect 18956 23828 19012 23838
rect 18956 23734 19012 23772
rect 19180 23826 19236 23884
rect 19628 23884 19796 23940
rect 19852 23940 19908 24670
rect 19180 23774 19182 23826
rect 19234 23774 19236 23826
rect 19180 23380 19236 23774
rect 19292 23826 19348 23838
rect 19292 23774 19294 23826
rect 19346 23774 19348 23826
rect 19292 23604 19348 23774
rect 19292 23538 19348 23548
rect 19516 23828 19572 23838
rect 19404 23380 19460 23390
rect 18956 23378 19460 23380
rect 18956 23326 19406 23378
rect 19458 23326 19460 23378
rect 18956 23324 19460 23326
rect 18956 22482 19012 23324
rect 19404 23314 19460 23324
rect 19292 23156 19348 23166
rect 18956 22430 18958 22482
rect 19010 22430 19012 22482
rect 18956 22418 19012 22430
rect 19180 23154 19348 23156
rect 19180 23102 19294 23154
rect 19346 23102 19348 23154
rect 19180 23100 19348 23102
rect 18844 22204 19124 22260
rect 18396 20804 18452 20814
rect 18172 20802 18452 20804
rect 18172 20750 18398 20802
rect 18450 20750 18452 20802
rect 18172 20748 18452 20750
rect 18732 20804 18788 21756
rect 18956 20804 19012 20814
rect 18732 20802 19012 20804
rect 18732 20750 18958 20802
rect 19010 20750 19012 20802
rect 18732 20748 19012 20750
rect 18060 20692 18116 20702
rect 18060 20598 18116 20636
rect 16828 20300 17332 20356
rect 17836 20412 18004 20468
rect 16604 20132 16660 20142
rect 16604 20038 16660 20076
rect 16716 20132 16772 20142
rect 16828 20132 16884 20300
rect 16716 20130 16884 20132
rect 16716 20078 16718 20130
rect 16770 20078 16884 20130
rect 16716 20076 16884 20078
rect 16716 20020 16772 20076
rect 16716 19954 16772 19964
rect 16380 19404 16772 19460
rect 16268 19394 16324 19404
rect 16492 19236 16548 19246
rect 15988 19180 16100 19236
rect 16156 19234 16548 19236
rect 16156 19182 16494 19234
rect 16546 19182 16548 19234
rect 16156 19180 16548 19182
rect 15932 19142 15988 19180
rect 16044 19012 16100 19022
rect 15820 19010 16100 19012
rect 15820 18958 16046 19010
rect 16098 18958 16100 19010
rect 15820 18956 16100 18958
rect 16044 18946 16100 18956
rect 15596 18274 15652 18284
rect 15596 18116 15652 18126
rect 14588 17614 14590 17666
rect 14642 17614 14644 17666
rect 14588 17602 14644 17614
rect 15260 17780 15316 17790
rect 14476 17502 14478 17554
rect 14530 17502 14532 17554
rect 13916 16818 13972 16828
rect 14476 16772 14532 17502
rect 15260 17106 15316 17724
rect 15260 17054 15262 17106
rect 15314 17054 15316 17106
rect 15260 16884 15316 17054
rect 15260 16818 15316 16828
rect 14812 16772 14868 16782
rect 14476 16770 14868 16772
rect 14476 16718 14814 16770
rect 14866 16718 14868 16770
rect 14476 16716 14868 16718
rect 14812 16706 14868 16716
rect 14064 16492 14328 16502
rect 14120 16436 14168 16492
rect 14224 16436 14272 16492
rect 14064 16426 14328 16436
rect 13580 15986 13748 15988
rect 13580 15934 13582 15986
rect 13634 15934 13748 15986
rect 13580 15932 13748 15934
rect 13804 16324 13860 16334
rect 13580 15922 13636 15932
rect 13244 15486 13246 15538
rect 13298 15486 13300 15538
rect 13244 15474 13300 15486
rect 13468 15540 13524 15550
rect 12348 13634 12516 13636
rect 12348 13582 12462 13634
rect 12514 13582 12516 13634
rect 12348 13580 12516 13582
rect 11788 13300 11844 13310
rect 11788 12964 11844 13244
rect 12124 12964 12180 12974
rect 11788 12962 12180 12964
rect 11788 12910 12126 12962
rect 12178 12910 12180 12962
rect 11788 12908 12180 12910
rect 11788 12850 11844 12908
rect 12124 12898 12180 12908
rect 11788 12798 11790 12850
rect 11842 12798 11844 12850
rect 11788 12786 11844 12798
rect 12236 12852 12292 12862
rect 12348 12852 12404 13580
rect 12460 13570 12516 13580
rect 12684 13634 12852 13636
rect 12684 13582 12798 13634
rect 12850 13582 12852 13634
rect 12684 13580 12852 13582
rect 12460 12964 12516 12974
rect 12460 12870 12516 12908
rect 12292 12796 12404 12852
rect 12236 12758 12292 12796
rect 11676 12460 11844 12516
rect 11676 12178 11732 12190
rect 11676 12126 11678 12178
rect 11730 12126 11732 12178
rect 11564 12068 11620 12078
rect 11676 12068 11732 12126
rect 11620 12012 11732 12068
rect 11564 12002 11620 12012
rect 11788 11732 11844 12460
rect 12460 12180 12516 12190
rect 11788 11676 12068 11732
rect 11004 11302 11060 11340
rect 11452 11396 11508 11406
rect 11452 11302 11508 11340
rect 11900 11396 11956 11406
rect 11900 11302 11956 11340
rect 10668 11284 10724 11294
rect 10668 11190 10724 11228
rect 9780 11004 10044 11014
rect 9836 10948 9884 11004
rect 9940 10948 9988 11004
rect 9780 10938 10044 10948
rect 9660 10782 9662 10834
rect 9714 10782 9716 10834
rect 9660 10770 9716 10782
rect 10332 10834 10388 11116
rect 12012 10836 12068 11676
rect 10332 10782 10334 10834
rect 10386 10782 10388 10834
rect 10332 10770 10388 10782
rect 11564 10834 12068 10836
rect 11564 10782 12014 10834
rect 12066 10782 12068 10834
rect 11564 10780 12068 10782
rect 9772 10612 9828 10622
rect 9100 10610 10052 10612
rect 9100 10558 9774 10610
rect 9826 10558 10052 10610
rect 9100 10556 10052 10558
rect 9772 10546 9828 10556
rect 9660 10388 9716 10398
rect 9660 10294 9716 10332
rect 9436 10164 9492 10174
rect 8204 8820 8260 8876
rect 8540 8866 8596 8876
rect 8652 9042 8708 9054
rect 8652 8990 8654 9042
rect 8706 8990 8708 9042
rect 7196 8764 8260 8820
rect 7196 8484 7252 8764
rect 6748 8418 6804 8428
rect 6860 8428 7252 8484
rect 7644 8484 7700 8494
rect 6636 8318 6638 8370
rect 6690 8318 6692 8370
rect 6636 8306 6692 8318
rect 6860 8260 6916 8428
rect 6748 8258 6916 8260
rect 6748 8206 6862 8258
rect 6914 8206 6916 8258
rect 6748 8204 6916 8206
rect 5964 8146 6020 8158
rect 5964 8094 5966 8146
rect 6018 8094 6020 8146
rect 5964 8036 6020 8094
rect 6300 8148 6356 8158
rect 6524 8148 6580 8158
rect 6300 8146 6580 8148
rect 6300 8094 6302 8146
rect 6354 8094 6526 8146
rect 6578 8094 6580 8146
rect 6300 8092 6580 8094
rect 6300 8082 6356 8092
rect 6524 8082 6580 8092
rect 5964 7970 6020 7980
rect 6076 8034 6132 8046
rect 6076 7982 6078 8034
rect 6130 7982 6132 8034
rect 5496 7084 5760 7094
rect 5552 7028 5600 7084
rect 5656 7028 5704 7084
rect 5496 7018 5760 7028
rect 6076 6804 6132 7982
rect 6748 7924 6804 8204
rect 6860 8194 6916 8204
rect 7084 8260 7140 8270
rect 7532 8260 7588 8270
rect 7084 8258 7588 8260
rect 7084 8206 7086 8258
rect 7138 8206 7534 8258
rect 7586 8206 7588 8258
rect 7084 8204 7588 8206
rect 7084 8194 7140 8204
rect 7532 8194 7588 8204
rect 7644 8258 7700 8428
rect 8540 8372 8596 8382
rect 8652 8372 8708 8990
rect 9436 8372 9492 10108
rect 9884 9940 9940 9950
rect 9660 9938 9940 9940
rect 9660 9886 9886 9938
rect 9938 9886 9940 9938
rect 9660 9884 9940 9886
rect 8540 8370 8708 8372
rect 8540 8318 8542 8370
rect 8594 8318 8708 8370
rect 8540 8316 8708 8318
rect 9324 8370 9492 8372
rect 9324 8318 9438 8370
rect 9490 8318 9492 8370
rect 9324 8316 9492 8318
rect 8540 8306 8596 8316
rect 8092 8260 8148 8270
rect 7644 8206 7646 8258
rect 7698 8206 7700 8258
rect 7644 8194 7700 8206
rect 7756 8204 8092 8260
rect 6412 7868 6804 7924
rect 6412 7586 6468 7868
rect 6412 7534 6414 7586
rect 6466 7534 6468 7586
rect 6412 7522 6468 7534
rect 6300 7476 6356 7486
rect 6300 7382 6356 7420
rect 6076 6738 6132 6748
rect 6524 7364 6580 7374
rect 6524 6690 6580 7308
rect 6524 6638 6526 6690
rect 6578 6638 6580 6690
rect 6524 6626 6580 6638
rect 6636 7362 6692 7374
rect 6636 7310 6638 7362
rect 6690 7310 6692 7362
rect 5740 6188 6468 6244
rect 5740 6130 5796 6188
rect 5740 6078 5742 6130
rect 5794 6078 5796 6130
rect 5740 6066 5796 6078
rect 5964 6020 6020 6030
rect 5964 5926 6020 5964
rect 5628 5906 5684 5918
rect 5628 5854 5630 5906
rect 5682 5854 5684 5906
rect 5628 5684 5684 5854
rect 5628 5628 5908 5684
rect 5496 5516 5760 5526
rect 5552 5460 5600 5516
rect 5656 5460 5704 5516
rect 5496 5450 5760 5460
rect 5740 5236 5796 5246
rect 5292 4286 5294 4338
rect 5346 4286 5348 4338
rect 5292 4274 5348 4286
rect 5404 4564 5460 4574
rect 5404 4116 5460 4508
rect 5292 4060 5460 4116
rect 5740 4116 5796 5180
rect 5852 4564 5908 5628
rect 6076 5124 6132 5134
rect 5964 4564 6020 4574
rect 5852 4508 5964 4564
rect 5964 4498 6020 4508
rect 5964 4340 6020 4350
rect 6076 4340 6132 5068
rect 5964 4338 6132 4340
rect 5964 4286 5966 4338
rect 6018 4286 6132 4338
rect 5964 4284 6132 4286
rect 6188 5012 6244 5022
rect 5964 4274 6020 4284
rect 5740 4060 5908 4116
rect 5292 3780 5348 4060
rect 5496 3948 5760 3958
rect 5552 3892 5600 3948
rect 5656 3892 5704 3948
rect 5496 3882 5760 3892
rect 5292 3724 5684 3780
rect 4508 3556 4564 3566
rect 4172 3554 4564 3556
rect 4172 3502 4510 3554
rect 4562 3502 4564 3554
rect 4172 3500 4564 3502
rect 4508 3490 4564 3500
rect 5628 3554 5684 3724
rect 5628 3502 5630 3554
rect 5682 3502 5684 3554
rect 5628 3490 5684 3502
rect 3948 3444 4004 3454
rect 3948 3330 4004 3388
rect 3948 3278 3950 3330
rect 4002 3278 4004 3330
rect 3948 3266 4004 3278
rect 4956 3444 5012 3454
rect 4956 800 5012 3388
rect 5740 3444 5796 3454
rect 5852 3444 5908 4060
rect 5964 3556 6020 3566
rect 6188 3556 6244 4956
rect 6412 4228 6468 6188
rect 6636 5908 6692 7310
rect 6748 6690 6804 7868
rect 7420 8034 7476 8046
rect 7420 7982 7422 8034
rect 7474 7982 7476 8034
rect 7084 7700 7140 7710
rect 7420 7700 7476 7982
rect 7084 7698 7476 7700
rect 7084 7646 7086 7698
rect 7138 7646 7476 7698
rect 7084 7644 7476 7646
rect 7084 7634 7140 7644
rect 7420 7588 7476 7644
rect 7420 7522 7476 7532
rect 6860 7476 6916 7486
rect 7196 7476 7252 7486
rect 6860 7474 7028 7476
rect 6860 7422 6862 7474
rect 6914 7422 7028 7474
rect 6860 7420 7028 7422
rect 6860 7410 6916 7420
rect 6748 6638 6750 6690
rect 6802 6638 6804 6690
rect 6748 6626 6804 6638
rect 6524 5852 6692 5908
rect 6860 6466 6916 6478
rect 6860 6414 6862 6466
rect 6914 6414 6916 6466
rect 6524 4452 6580 5852
rect 6636 5682 6692 5694
rect 6636 5630 6638 5682
rect 6690 5630 6692 5682
rect 6636 4676 6692 5630
rect 6860 5234 6916 6414
rect 6972 5796 7028 7420
rect 7196 7382 7252 7420
rect 7308 7474 7364 7486
rect 7308 7422 7310 7474
rect 7362 7422 7364 7474
rect 7308 6804 7364 7422
rect 7756 7474 7812 8204
rect 8092 8166 8148 8204
rect 9100 8260 9156 8270
rect 9100 8166 9156 8204
rect 8540 8148 8596 8158
rect 8428 8034 8484 8046
rect 8428 7982 8430 8034
rect 8482 7982 8484 8034
rect 7980 7588 8036 7598
rect 7980 7494 8036 7532
rect 8428 7588 8484 7982
rect 8428 7522 8484 7532
rect 7756 7422 7758 7474
rect 7810 7422 7812 7474
rect 7756 7410 7812 7422
rect 8204 7474 8260 7486
rect 8204 7422 8206 7474
rect 8258 7422 8260 7474
rect 8092 7364 8148 7374
rect 8092 7270 8148 7308
rect 7308 6738 7364 6748
rect 6972 5730 7028 5740
rect 7196 6690 7252 6702
rect 7196 6638 7198 6690
rect 7250 6638 7252 6690
rect 6860 5182 6862 5234
rect 6914 5182 6916 5234
rect 6860 5170 6916 5182
rect 6636 4620 6804 4676
rect 6636 4452 6692 4462
rect 6524 4450 6692 4452
rect 6524 4398 6638 4450
rect 6690 4398 6692 4450
rect 6524 4396 6692 4398
rect 6636 4386 6692 4396
rect 6748 4228 6804 4620
rect 6412 4162 6468 4172
rect 6524 4172 6804 4228
rect 5964 3554 6244 3556
rect 5964 3502 5966 3554
rect 6018 3502 6244 3554
rect 5964 3500 6244 3502
rect 5964 3490 6020 3500
rect 5740 3442 5908 3444
rect 5740 3390 5742 3442
rect 5794 3390 5908 3442
rect 5740 3388 5908 3390
rect 5740 3378 5796 3388
rect 6524 800 6580 4172
rect 7196 3780 7252 6638
rect 8204 5572 8260 7422
rect 8540 7474 8596 8092
rect 8540 7422 8542 7474
rect 8594 7422 8596 7474
rect 8540 7410 8596 7422
rect 8652 8034 8708 8046
rect 8652 7982 8654 8034
rect 8706 7982 8708 8034
rect 8652 7028 8708 7982
rect 9100 7700 9156 7710
rect 9100 7606 9156 7644
rect 9324 7364 9380 8316
rect 9436 8306 9492 8316
rect 9548 8372 9604 8382
rect 9548 7812 9604 8316
rect 9324 7298 9380 7308
rect 9436 7756 9604 7812
rect 8652 6962 8708 6972
rect 9436 6916 9492 7756
rect 9548 7588 9604 7598
rect 9548 7494 9604 7532
rect 8540 6804 8596 6814
rect 8204 5506 8260 5516
rect 8316 6578 8372 6590
rect 8316 6526 8318 6578
rect 8370 6526 8372 6578
rect 7196 3714 7252 3724
rect 8316 3444 8372 6526
rect 8540 5908 8596 6748
rect 8764 5908 8820 5918
rect 8540 5906 8820 5908
rect 8540 5854 8766 5906
rect 8818 5854 8820 5906
rect 8540 5852 8820 5854
rect 8764 4226 8820 5852
rect 8988 5572 9044 5582
rect 8988 5236 9044 5516
rect 8764 4174 8766 4226
rect 8818 4174 8820 4226
rect 8764 4162 8820 4174
rect 8876 5234 9044 5236
rect 8876 5182 8990 5234
rect 9042 5182 9044 5234
rect 8876 5180 9044 5182
rect 8764 3556 8820 3566
rect 8876 3556 8932 5180
rect 8988 5170 9044 5180
rect 9324 5010 9380 5022
rect 9324 4958 9326 5010
rect 9378 4958 9380 5010
rect 9324 4564 9380 4958
rect 9436 5010 9492 6860
rect 9660 7028 9716 9884
rect 9884 9874 9940 9884
rect 9996 9604 10052 10556
rect 10892 10500 10948 10510
rect 10668 9828 10724 9838
rect 10892 9828 10948 10444
rect 10668 9826 10948 9828
rect 10668 9774 10670 9826
rect 10722 9774 10948 9826
rect 10668 9772 10948 9774
rect 11116 9826 11172 9838
rect 11116 9774 11118 9826
rect 11170 9774 11172 9826
rect 10668 9762 10724 9772
rect 9996 9548 10164 9604
rect 9780 9436 10044 9446
rect 9836 9380 9884 9436
rect 9940 9380 9988 9436
rect 9780 9370 10044 9380
rect 10108 9268 10164 9548
rect 9996 9212 10164 9268
rect 10332 9602 10388 9614
rect 10332 9550 10334 9602
rect 10386 9550 10388 9602
rect 9772 8372 9828 8382
rect 9772 8278 9828 8316
rect 9996 8036 10052 9212
rect 10332 8260 10388 9550
rect 10332 8194 10388 8204
rect 10052 7980 10500 8036
rect 9996 7970 10052 7980
rect 9780 7868 10044 7878
rect 9836 7812 9884 7868
rect 9940 7812 9988 7868
rect 9780 7802 10044 7812
rect 9996 7474 10052 7486
rect 9996 7422 9998 7474
rect 10050 7422 10052 7474
rect 9996 7364 10052 7422
rect 9996 7298 10052 7308
rect 10220 7476 10276 7486
rect 9660 6690 9716 6972
rect 9660 6638 9662 6690
rect 9714 6638 9716 6690
rect 9548 5908 9604 5918
rect 9548 5814 9604 5852
rect 9660 5684 9716 6638
rect 9780 6300 10044 6310
rect 9836 6244 9884 6300
rect 9940 6244 9988 6300
rect 9780 6234 10044 6244
rect 10220 6132 10276 7420
rect 9996 6076 10276 6132
rect 9436 4958 9438 5010
rect 9490 4958 9492 5010
rect 9436 4946 9492 4958
rect 9548 5628 9716 5684
rect 9772 6018 9828 6030
rect 9772 5966 9774 6018
rect 9826 5966 9828 6018
rect 9548 4788 9604 5628
rect 9772 5236 9828 5966
rect 9884 6020 9940 6030
rect 9996 6020 10052 6076
rect 10332 6020 10388 6030
rect 9884 6018 10052 6020
rect 9884 5966 9886 6018
rect 9938 5966 10052 6018
rect 9884 5964 10052 5966
rect 10220 6018 10388 6020
rect 10220 5966 10334 6018
rect 10386 5966 10388 6018
rect 10220 5964 10388 5966
rect 9884 5954 9940 5964
rect 10108 5906 10164 5918
rect 10108 5854 10110 5906
rect 10162 5854 10164 5906
rect 10108 5796 10164 5854
rect 10108 5730 10164 5740
rect 10108 5572 10164 5582
rect 10220 5572 10276 5964
rect 10332 5954 10388 5964
rect 10164 5516 10276 5572
rect 10444 5906 10500 7980
rect 10780 7700 10836 7710
rect 10780 7606 10836 7644
rect 11116 7698 11172 9774
rect 11564 9826 11620 10780
rect 12012 10770 12068 10780
rect 12460 10612 12516 12124
rect 12684 11396 12740 13580
rect 12796 13570 12852 13580
rect 13356 13746 13412 13758
rect 13356 13694 13358 13746
rect 13410 13694 13412 13746
rect 13356 13636 13412 13694
rect 12908 13524 12964 13534
rect 12796 13076 12852 13086
rect 12908 13076 12964 13468
rect 12852 13020 12964 13076
rect 12796 12982 12852 13020
rect 13244 12292 13300 12302
rect 12908 12290 13300 12292
rect 12908 12238 13246 12290
rect 13298 12238 13300 12290
rect 12908 12236 13300 12238
rect 12796 11396 12852 11406
rect 12684 11340 12796 11396
rect 12796 11330 12852 11340
rect 12460 10610 12628 10612
rect 12460 10558 12462 10610
rect 12514 10558 12628 10610
rect 12460 10556 12628 10558
rect 12460 10546 12516 10556
rect 11564 9774 11566 9826
rect 11618 9774 11620 9826
rect 11564 9762 11620 9774
rect 11788 9828 11844 9838
rect 12348 9828 12404 9838
rect 11788 9826 12404 9828
rect 11788 9774 11790 9826
rect 11842 9774 12350 9826
rect 12402 9774 12404 9826
rect 11788 9772 12404 9774
rect 11788 9762 11844 9772
rect 12348 9762 12404 9772
rect 11452 9602 11508 9614
rect 11452 9550 11454 9602
rect 11506 9550 11508 9602
rect 11452 8820 11508 9550
rect 12236 9604 12292 9614
rect 12124 8932 12180 8942
rect 11452 8764 11732 8820
rect 11676 8372 11732 8764
rect 11900 8372 11956 8382
rect 11676 8370 11956 8372
rect 11676 8318 11902 8370
rect 11954 8318 11956 8370
rect 11676 8316 11956 8318
rect 11900 8306 11956 8316
rect 11116 7646 11118 7698
rect 11170 7646 11172 7698
rect 10780 6020 10836 6030
rect 10780 5926 10836 5964
rect 10444 5854 10446 5906
rect 10498 5854 10500 5906
rect 10108 5506 10164 5516
rect 10444 5348 10500 5854
rect 11004 5908 11060 5918
rect 11004 5814 11060 5852
rect 10892 5794 10948 5806
rect 10892 5742 10894 5794
rect 10946 5742 10948 5794
rect 10892 5348 10948 5742
rect 9772 5170 9828 5180
rect 10108 5292 10500 5348
rect 10668 5292 10948 5348
rect 9884 5124 9940 5134
rect 9884 5030 9940 5068
rect 9660 4900 9716 4910
rect 9660 4806 9716 4844
rect 9324 4498 9380 4508
rect 9436 4732 9604 4788
rect 9780 4732 10044 4742
rect 8764 3554 8932 3556
rect 8764 3502 8766 3554
rect 8818 3502 8932 3554
rect 8764 3500 8932 3502
rect 9212 3780 9268 3790
rect 9212 3554 9268 3724
rect 9212 3502 9214 3554
rect 9266 3502 9268 3554
rect 8764 3490 8820 3500
rect 9212 3490 9268 3502
rect 8316 3378 8372 3388
rect 9436 3442 9492 4732
rect 9836 4676 9884 4732
rect 9940 4676 9988 4732
rect 9780 4666 10044 4676
rect 10108 4564 10164 5292
rect 10668 5234 10724 5292
rect 10668 5182 10670 5234
rect 10722 5182 10724 5234
rect 10668 5170 10724 5182
rect 9996 4508 10164 4564
rect 10444 4788 10500 4798
rect 9548 4228 9604 4238
rect 9548 4134 9604 4172
rect 9548 3556 9604 3566
rect 9996 3556 10052 4508
rect 9548 3554 10052 3556
rect 9548 3502 9550 3554
rect 9602 3502 10052 3554
rect 9548 3500 10052 3502
rect 10444 4228 10500 4732
rect 11116 4564 11172 7646
rect 11564 7588 11620 7598
rect 11564 7586 11732 7588
rect 11564 7534 11566 7586
rect 11618 7534 11732 7586
rect 11564 7532 11732 7534
rect 11564 7522 11620 7532
rect 11452 7476 11508 7486
rect 11452 7382 11508 7420
rect 11564 7250 11620 7262
rect 11564 7198 11566 7250
rect 11618 7198 11620 7250
rect 11116 4498 11172 4508
rect 11228 6578 11284 6590
rect 11228 6526 11230 6578
rect 11282 6526 11284 6578
rect 10444 3554 10500 4172
rect 10444 3502 10446 3554
rect 10498 3502 10500 3554
rect 9548 3490 9604 3500
rect 10444 3490 10500 3502
rect 9436 3390 9438 3442
rect 9490 3390 9492 3442
rect 9436 3378 9492 3390
rect 9660 3388 9716 3398
rect 7756 3332 7812 3342
rect 7756 3330 8148 3332
rect 7756 3278 7758 3330
rect 7810 3278 8148 3330
rect 7756 3276 8148 3278
rect 7756 3266 7812 3276
rect 8092 800 8148 3276
rect 9660 800 9716 3332
rect 9780 3164 10044 3174
rect 9836 3108 9884 3164
rect 9940 3108 9988 3164
rect 9780 3098 10044 3108
rect 11228 800 11284 6526
rect 11340 6020 11396 6030
rect 11340 5926 11396 5964
rect 11564 5684 11620 7198
rect 11564 5618 11620 5628
rect 11676 4788 11732 7532
rect 12124 7474 12180 8876
rect 12236 7700 12292 9548
rect 12236 7634 12292 7644
rect 12460 9602 12516 9614
rect 12460 9550 12462 9602
rect 12514 9550 12516 9602
rect 12124 7422 12126 7474
rect 12178 7422 12180 7474
rect 11788 5908 11844 5918
rect 12124 5908 12180 7422
rect 12460 6916 12516 9550
rect 12460 6690 12516 6860
rect 12460 6638 12462 6690
rect 12514 6638 12516 6690
rect 12460 6626 12516 6638
rect 12572 8258 12628 10556
rect 12908 9828 12964 12236
rect 13244 12226 13300 12236
rect 13132 10498 13188 10510
rect 13132 10446 13134 10498
rect 13186 10446 13188 10498
rect 13132 9940 13188 10446
rect 13244 10500 13300 10510
rect 13356 10500 13412 13580
rect 13300 10444 13412 10500
rect 13244 10434 13300 10444
rect 13132 9874 13188 9884
rect 12908 9734 12964 9772
rect 12572 8206 12574 8258
rect 12626 8206 12628 8258
rect 11788 5906 12180 5908
rect 11788 5854 11790 5906
rect 11842 5854 12180 5906
rect 11788 5852 12180 5854
rect 11788 5124 11844 5852
rect 12460 5796 12516 5806
rect 12460 5702 12516 5740
rect 11788 5058 11844 5068
rect 11676 4722 11732 4732
rect 12460 4340 12516 4350
rect 12572 4340 12628 8206
rect 12908 8036 12964 8046
rect 12908 7586 12964 7980
rect 12908 7534 12910 7586
rect 12962 7534 12964 7586
rect 12908 7522 12964 7534
rect 13244 6132 13300 6142
rect 12796 5908 12852 5918
rect 12796 5236 12852 5852
rect 12796 5142 12852 5180
rect 13020 5684 13076 5694
rect 12516 4284 12628 4340
rect 12684 4900 12740 4910
rect 12684 4338 12740 4844
rect 12684 4286 12686 4338
rect 12738 4286 12740 4338
rect 12460 4246 12516 4284
rect 12684 4274 12740 4286
rect 13020 4338 13076 5628
rect 13020 4286 13022 4338
rect 13074 4286 13076 4338
rect 13020 4274 13076 4286
rect 11676 4228 11732 4238
rect 11676 4134 11732 4172
rect 12908 4228 12964 4238
rect 12908 4134 12964 4172
rect 12348 3666 12404 3678
rect 12348 3614 12350 3666
rect 12402 3614 12404 3666
rect 12348 3388 12404 3614
rect 13244 3554 13300 6076
rect 13468 6020 13524 15484
rect 13804 15538 13860 16268
rect 15260 16324 15316 16334
rect 15316 16268 15428 16324
rect 15260 16258 15316 16268
rect 15372 16212 15428 16268
rect 15372 16118 15428 16156
rect 15260 15986 15316 15998
rect 15260 15934 15262 15986
rect 15314 15934 15316 15986
rect 13916 15876 13972 15886
rect 14924 15876 14980 15886
rect 15260 15876 15316 15934
rect 13916 15874 14420 15876
rect 13916 15822 13918 15874
rect 13970 15822 14420 15874
rect 13916 15820 14420 15822
rect 13916 15810 13972 15820
rect 13804 15486 13806 15538
rect 13858 15486 13860 15538
rect 13804 15474 13860 15486
rect 14140 15428 14196 15438
rect 14140 15334 14196 15372
rect 14364 15314 14420 15820
rect 14924 15874 15316 15876
rect 14924 15822 14926 15874
rect 14978 15822 15316 15874
rect 14924 15820 15316 15822
rect 14924 15810 14980 15820
rect 14812 15540 14868 15550
rect 14812 15426 14868 15484
rect 14812 15374 14814 15426
rect 14866 15374 14868 15426
rect 14812 15362 14868 15374
rect 14364 15262 14366 15314
rect 14418 15262 14420 15314
rect 14364 15092 14420 15262
rect 14924 15202 14980 15214
rect 14924 15150 14926 15202
rect 14978 15150 14980 15202
rect 14924 15148 14980 15150
rect 14364 15026 14420 15036
rect 14476 15092 14980 15148
rect 14064 14924 14328 14934
rect 14120 14868 14168 14924
rect 14224 14868 14272 14924
rect 14064 14858 14328 14868
rect 14476 14642 14532 15092
rect 14812 14980 14868 14990
rect 14868 14924 14980 14980
rect 14812 14914 14868 14924
rect 14476 14590 14478 14642
rect 14530 14590 14532 14642
rect 14476 14578 14532 14590
rect 13804 14532 13860 14542
rect 13804 14530 13972 14532
rect 13804 14478 13806 14530
rect 13858 14478 13972 14530
rect 13804 14476 13972 14478
rect 13804 14466 13860 14476
rect 13804 13636 13860 13646
rect 13804 13542 13860 13580
rect 13580 12404 13636 12414
rect 13580 12310 13636 12348
rect 13916 12180 13972 14476
rect 14924 13970 14980 14924
rect 14924 13918 14926 13970
rect 14978 13918 14980 13970
rect 14364 13748 14420 13758
rect 14700 13748 14756 13758
rect 14364 13746 14756 13748
rect 14364 13694 14366 13746
rect 14418 13694 14702 13746
rect 14754 13694 14756 13746
rect 14364 13692 14756 13694
rect 14364 13682 14420 13692
rect 14700 13636 14756 13692
rect 14700 13570 14756 13580
rect 14064 13356 14328 13366
rect 14120 13300 14168 13356
rect 14224 13300 14272 13356
rect 14064 13290 14328 13300
rect 14924 12740 14980 13918
rect 15036 13636 15092 15820
rect 15596 15540 15652 18060
rect 16156 17780 16212 19180
rect 16492 19170 16548 19180
rect 16268 19010 16324 19022
rect 16268 18958 16270 19010
rect 16322 18958 16324 19010
rect 16268 18452 16324 18958
rect 16268 18386 16324 18396
rect 16380 19012 16436 19022
rect 16156 17686 16212 17724
rect 16380 15986 16436 18956
rect 16716 17108 16772 19404
rect 16828 18338 16884 20076
rect 17388 20132 17444 20142
rect 17388 20038 17444 20076
rect 16940 20018 16996 20030
rect 16940 19966 16942 20018
rect 16994 19966 16996 20018
rect 16940 18452 16996 19966
rect 17724 20018 17780 20030
rect 17724 19966 17726 20018
rect 17778 19966 17780 20018
rect 17276 19124 17332 19134
rect 17276 19122 17556 19124
rect 17276 19070 17278 19122
rect 17330 19070 17556 19122
rect 17276 19068 17556 19070
rect 17276 19058 17332 19068
rect 17500 18674 17556 19068
rect 17500 18622 17502 18674
rect 17554 18622 17556 18674
rect 17500 18610 17556 18622
rect 17276 18452 17332 18462
rect 16940 18450 17332 18452
rect 16940 18398 17278 18450
rect 17330 18398 17332 18450
rect 16940 18396 17332 18398
rect 17276 18386 17332 18396
rect 17612 18452 17668 18462
rect 17612 18358 17668 18396
rect 16828 18286 16830 18338
rect 16882 18286 16884 18338
rect 16828 18274 16884 18286
rect 17724 17892 17780 19966
rect 17836 20020 17892 20412
rect 18172 20356 18228 20748
rect 18396 20738 18452 20748
rect 18956 20738 19012 20748
rect 18620 20692 18676 20702
rect 18284 20580 18340 20618
rect 18620 20598 18676 20636
rect 18284 20514 18340 20524
rect 18844 20578 18900 20590
rect 19068 20580 19124 22204
rect 19180 21700 19236 23100
rect 19292 23090 19348 23100
rect 19404 22932 19460 22942
rect 19404 22838 19460 22876
rect 19404 22596 19460 22606
rect 19404 22502 19460 22540
rect 19180 21634 19236 21644
rect 19292 22258 19348 22270
rect 19292 22206 19294 22258
rect 19346 22206 19348 22258
rect 18844 20526 18846 20578
rect 18898 20526 18900 20578
rect 18844 20468 18900 20526
rect 17948 20300 18228 20356
rect 18348 20412 18612 20422
rect 18404 20356 18452 20412
rect 18508 20356 18556 20412
rect 18844 20402 18900 20412
rect 18956 20524 19124 20580
rect 18348 20346 18612 20356
rect 17948 20242 18004 20300
rect 17948 20190 17950 20242
rect 18002 20190 18004 20242
rect 17948 20178 18004 20190
rect 18172 20130 18228 20142
rect 18172 20078 18174 20130
rect 18226 20078 18228 20130
rect 18172 20020 18228 20078
rect 18284 20132 18340 20142
rect 18284 20038 18340 20076
rect 17836 19964 18228 20020
rect 18732 19012 18788 19022
rect 18348 18844 18612 18854
rect 18404 18788 18452 18844
rect 18508 18788 18556 18844
rect 18348 18778 18612 18788
rect 17836 18450 17892 18462
rect 17836 18398 17838 18450
rect 17890 18398 17892 18450
rect 17836 18340 17892 18398
rect 17836 18274 17892 18284
rect 17724 17826 17780 17836
rect 18060 18116 18116 18126
rect 17052 17780 17108 17790
rect 17052 17686 17108 17724
rect 17612 17612 17892 17668
rect 16828 17108 16884 17118
rect 16716 17052 16828 17108
rect 16380 15934 16382 15986
rect 16434 15934 16436 15986
rect 16380 15922 16436 15934
rect 16492 16098 16548 16110
rect 16492 16046 16494 16098
rect 16546 16046 16548 16098
rect 15148 15538 15652 15540
rect 15148 15486 15598 15538
rect 15650 15486 15652 15538
rect 15148 15484 15652 15486
rect 15148 15314 15204 15484
rect 15596 15474 15652 15484
rect 15148 15262 15150 15314
rect 15202 15262 15204 15314
rect 15148 15250 15204 15262
rect 15596 13858 15652 13870
rect 15596 13806 15598 13858
rect 15650 13806 15652 13858
rect 15036 13570 15092 13580
rect 15372 13746 15428 13758
rect 15372 13694 15374 13746
rect 15426 13694 15428 13746
rect 15372 13636 15428 13694
rect 15596 13748 15652 13806
rect 15596 13682 15652 13692
rect 15372 13570 15428 13580
rect 16156 13636 16212 13646
rect 16492 13636 16548 16046
rect 16716 15316 16772 17052
rect 16828 17014 16884 17052
rect 17612 16994 17668 17612
rect 17836 17556 17892 17612
rect 18060 17666 18116 18060
rect 18060 17614 18062 17666
rect 18114 17614 18116 17666
rect 18060 17602 18116 17614
rect 18284 17668 18340 17678
rect 18284 17574 18340 17612
rect 17836 17462 17892 17500
rect 18620 17556 18676 17566
rect 18620 17462 18676 17500
rect 17612 16942 17614 16994
rect 17666 16942 17668 16994
rect 17612 16930 17668 16942
rect 17724 17444 17780 17454
rect 16716 15250 16772 15260
rect 16828 16210 16884 16222
rect 16828 16158 16830 16210
rect 16882 16158 16884 16210
rect 16828 14756 16884 16158
rect 17724 16100 17780 17388
rect 18348 17276 18612 17286
rect 18404 17220 18452 17276
rect 18508 17220 18556 17276
rect 18348 17210 18612 17220
rect 17836 17108 17892 17118
rect 17836 16994 17892 17052
rect 17836 16942 17838 16994
rect 17890 16942 17892 16994
rect 17836 16930 17892 16942
rect 17948 16996 18004 17006
rect 17948 16994 18116 16996
rect 17948 16942 17950 16994
rect 18002 16942 18116 16994
rect 17948 16940 18116 16942
rect 17948 16930 18004 16940
rect 17948 16770 18004 16782
rect 17948 16718 17950 16770
rect 18002 16718 18004 16770
rect 17836 16100 17892 16110
rect 17724 16098 17892 16100
rect 17724 16046 17838 16098
rect 17890 16046 17892 16098
rect 17724 16044 17892 16046
rect 17836 16034 17892 16044
rect 17500 15314 17556 15326
rect 17500 15262 17502 15314
rect 17554 15262 17556 15314
rect 17052 15204 17108 15214
rect 16828 14690 16884 14700
rect 16940 15092 16996 15102
rect 16604 14642 16660 14654
rect 16604 14590 16606 14642
rect 16658 14590 16660 14642
rect 16604 13972 16660 14590
rect 16940 14644 16996 15036
rect 16940 14550 16996 14588
rect 16604 13906 16660 13916
rect 16212 13580 16324 13636
rect 16156 13542 16212 13580
rect 15148 12740 15204 12750
rect 15484 12740 15540 12750
rect 14924 12738 15204 12740
rect 14924 12686 15150 12738
rect 15202 12686 15204 12738
rect 14924 12684 15204 12686
rect 15148 12404 15204 12684
rect 15148 12338 15204 12348
rect 15260 12738 15540 12740
rect 15260 12686 15486 12738
rect 15538 12686 15540 12738
rect 15260 12684 15540 12686
rect 13916 12086 13972 12124
rect 14700 12068 14756 12078
rect 14700 12066 14980 12068
rect 14700 12014 14702 12066
rect 14754 12014 14980 12066
rect 14700 12012 14980 12014
rect 14700 12002 14756 12012
rect 14064 11788 14328 11798
rect 14120 11732 14168 11788
rect 14224 11732 14272 11788
rect 14064 11722 14328 11732
rect 14924 11506 14980 12012
rect 15148 11844 15204 11854
rect 14924 11454 14926 11506
rect 14978 11454 14980 11506
rect 14924 11442 14980 11454
rect 15036 11788 15148 11844
rect 15036 11394 15092 11788
rect 15148 11778 15204 11788
rect 15036 11342 15038 11394
rect 15090 11342 15092 11394
rect 14812 11282 14868 11294
rect 14812 11230 14814 11282
rect 14866 11230 14868 11282
rect 14588 10500 14644 10510
rect 14064 10220 14328 10230
rect 14120 10164 14168 10220
rect 14224 10164 14272 10220
rect 14064 10154 14328 10164
rect 14476 10052 14532 10062
rect 14140 9940 14196 9950
rect 14140 9846 14196 9884
rect 14028 9716 14084 9726
rect 13916 9714 14084 9716
rect 13916 9662 14030 9714
rect 14082 9662 14084 9714
rect 13916 9660 14084 9662
rect 13580 9604 13636 9614
rect 13580 8932 13636 9548
rect 13580 8866 13636 8876
rect 13916 8484 13972 9660
rect 14028 9650 14084 9660
rect 14364 9716 14420 9726
rect 14476 9716 14532 9996
rect 14588 9826 14644 10444
rect 14588 9774 14590 9826
rect 14642 9774 14644 9826
rect 14588 9762 14644 9774
rect 14364 9714 14532 9716
rect 14364 9662 14366 9714
rect 14418 9662 14532 9714
rect 14364 9660 14532 9662
rect 14364 9650 14420 9660
rect 14064 8652 14328 8662
rect 14120 8596 14168 8652
rect 14224 8596 14272 8652
rect 14064 8586 14328 8596
rect 13916 8418 13972 8428
rect 14140 8484 14196 8494
rect 13692 8204 14084 8260
rect 13580 8146 13636 8158
rect 13580 8094 13582 8146
rect 13634 8094 13636 8146
rect 13580 7476 13636 8094
rect 13692 8146 13748 8204
rect 13692 8094 13694 8146
rect 13746 8094 13748 8146
rect 13692 8082 13748 8094
rect 13916 8036 13972 8046
rect 13580 7410 13636 7420
rect 13804 8034 13972 8036
rect 13804 7982 13918 8034
rect 13970 7982 13972 8034
rect 13804 7980 13972 7982
rect 13468 5348 13524 5964
rect 13356 5292 13468 5348
rect 13356 4450 13412 5292
rect 13468 5282 13524 5292
rect 13580 5796 13636 5806
rect 13580 5234 13636 5740
rect 13580 5182 13582 5234
rect 13634 5182 13636 5234
rect 13580 5170 13636 5182
rect 13468 5124 13524 5134
rect 13468 5030 13524 5068
rect 13804 5122 13860 7980
rect 13916 7970 13972 7980
rect 13916 7476 13972 7486
rect 13916 6690 13972 7420
rect 14028 7364 14084 8204
rect 14140 8258 14196 8428
rect 14140 8206 14142 8258
rect 14194 8206 14196 8258
rect 14140 8194 14196 8206
rect 14476 8258 14532 9660
rect 14476 8206 14478 8258
rect 14530 8206 14532 8258
rect 14476 8194 14532 8206
rect 14700 9604 14756 9614
rect 14700 8258 14756 9548
rect 14812 9492 14868 11230
rect 15036 10052 15092 11342
rect 15260 11172 15316 12684
rect 15484 12674 15540 12684
rect 16156 12738 16212 12750
rect 16156 12686 16158 12738
rect 16210 12686 16212 12738
rect 16156 11844 16212 12686
rect 16268 12180 16324 13580
rect 16492 13570 16548 13580
rect 16716 13748 16772 13758
rect 16492 12738 16548 12750
rect 16492 12686 16494 12738
rect 16546 12686 16548 12738
rect 16492 12404 16548 12686
rect 16492 12338 16548 12348
rect 16268 12124 16548 12180
rect 16156 11778 16212 11788
rect 15932 11508 15988 11518
rect 15372 11396 15428 11406
rect 15820 11396 15876 11406
rect 15372 11394 15876 11396
rect 15372 11342 15374 11394
rect 15426 11342 15822 11394
rect 15874 11342 15876 11394
rect 15372 11340 15876 11342
rect 15372 11330 15428 11340
rect 15820 11330 15876 11340
rect 15932 11394 15988 11452
rect 15932 11342 15934 11394
rect 15986 11342 15988 11394
rect 15932 11330 15988 11342
rect 15708 11172 15764 11182
rect 15260 11106 15316 11116
rect 15596 11170 15764 11172
rect 15596 11118 15710 11170
rect 15762 11118 15764 11170
rect 15596 11116 15764 11118
rect 15596 10612 15652 11116
rect 15708 11106 15764 11116
rect 16156 11172 16212 11182
rect 16156 11078 16212 11116
rect 15596 10518 15652 10556
rect 15820 10610 15876 10622
rect 15820 10558 15822 10610
rect 15874 10558 15876 10610
rect 15260 10498 15316 10510
rect 15260 10446 15262 10498
rect 15314 10446 15316 10498
rect 15260 10276 15316 10446
rect 15708 10500 15764 10510
rect 15708 10406 15764 10444
rect 15820 10276 15876 10558
rect 15260 10220 15876 10276
rect 15036 9986 15092 9996
rect 14924 9828 14980 9838
rect 15820 9828 15876 10220
rect 16156 10610 16212 10622
rect 16156 10558 16158 10610
rect 16210 10558 16212 10610
rect 16044 9828 16100 9838
rect 15820 9826 16100 9828
rect 15820 9774 16046 9826
rect 16098 9774 16100 9826
rect 15820 9772 16100 9774
rect 14924 9734 14980 9772
rect 16044 9762 16100 9772
rect 16156 9828 16212 10558
rect 16492 10388 16548 12124
rect 16492 10322 16548 10332
rect 16604 11282 16660 11294
rect 16604 11230 16606 11282
rect 16658 11230 16660 11282
rect 14812 9426 14868 9436
rect 15260 9602 15316 9614
rect 15260 9550 15262 9602
rect 15314 9550 15316 9602
rect 15260 9156 15316 9550
rect 15372 9604 15428 9614
rect 15372 9510 15428 9548
rect 15484 9602 15540 9614
rect 15484 9550 15486 9602
rect 15538 9550 15540 9602
rect 15484 9268 15540 9550
rect 15484 9202 15540 9212
rect 15820 9602 15876 9614
rect 15820 9550 15822 9602
rect 15874 9550 15876 9602
rect 15820 9156 15876 9550
rect 15932 9604 15988 9614
rect 15932 9510 15988 9548
rect 16156 9266 16212 9772
rect 16156 9214 16158 9266
rect 16210 9214 16212 9266
rect 16156 9202 16212 9214
rect 16268 9602 16324 9614
rect 16268 9550 16270 9602
rect 16322 9550 16324 9602
rect 15260 9100 15428 9156
rect 14812 9044 14868 9054
rect 14812 9042 15316 9044
rect 14812 8990 14814 9042
rect 14866 8990 15316 9042
rect 14812 8988 15316 8990
rect 14812 8978 14868 8988
rect 15260 8930 15316 8988
rect 15260 8878 15262 8930
rect 15314 8878 15316 8930
rect 15036 8820 15092 8830
rect 14700 8206 14702 8258
rect 14754 8206 14756 8258
rect 14700 8194 14756 8206
rect 14924 8764 15036 8820
rect 14252 8036 14308 8046
rect 14252 7942 14308 7980
rect 14028 7308 14644 7364
rect 14064 7084 14328 7094
rect 14120 7028 14168 7084
rect 14224 7028 14272 7084
rect 14064 7018 14328 7028
rect 13916 6638 13918 6690
rect 13970 6638 13972 6690
rect 13916 6626 13972 6638
rect 14476 6578 14532 6590
rect 14476 6526 14478 6578
rect 14530 6526 14532 6578
rect 14028 6466 14084 6478
rect 14028 6414 14030 6466
rect 14082 6414 14084 6466
rect 14028 5684 14084 6414
rect 14252 6466 14308 6478
rect 14252 6414 14254 6466
rect 14306 6414 14308 6466
rect 14252 6020 14308 6414
rect 14476 6132 14532 6526
rect 14476 6066 14532 6076
rect 14588 6466 14644 7308
rect 14924 6804 14980 8764
rect 15036 8754 15092 8764
rect 15260 8260 15316 8878
rect 15260 8194 15316 8204
rect 15372 8036 15428 9100
rect 15260 7980 15428 8036
rect 15596 9100 15820 9156
rect 15260 7700 15316 7980
rect 15036 7644 15260 7700
rect 15036 7362 15092 7644
rect 15260 7606 15316 7644
rect 15596 7698 15652 9100
rect 15820 9062 15876 9100
rect 15708 8932 15764 8942
rect 15708 8838 15764 8876
rect 15596 7646 15598 7698
rect 15650 7646 15652 7698
rect 15596 7634 15652 7646
rect 15708 8148 15764 8158
rect 15708 7698 15764 8092
rect 16268 8148 16324 9550
rect 16604 9268 16660 11230
rect 16716 10388 16772 13692
rect 16828 12066 16884 12078
rect 16828 12014 16830 12066
rect 16882 12014 16884 12066
rect 16828 11508 16884 12014
rect 16828 11442 16884 11452
rect 16716 10322 16772 10332
rect 16940 10052 16996 10062
rect 16940 9826 16996 9996
rect 16940 9774 16942 9826
rect 16994 9774 16996 9826
rect 16940 9762 16996 9774
rect 16604 9202 16660 9212
rect 16716 9714 16772 9726
rect 16716 9662 16718 9714
rect 16770 9662 16772 9714
rect 16380 9042 16436 9054
rect 16380 8990 16382 9042
rect 16434 8990 16436 9042
rect 16380 8820 16436 8990
rect 16492 9044 16548 9054
rect 16716 9044 16772 9662
rect 16492 9042 16772 9044
rect 16492 8990 16494 9042
rect 16546 8990 16772 9042
rect 16492 8988 16772 8990
rect 16492 8978 16548 8988
rect 17052 8932 17108 15148
rect 17500 14420 17556 15262
rect 17948 15314 18004 16718
rect 18060 16324 18116 16940
rect 18172 16882 18228 16894
rect 18732 16884 18788 18956
rect 18844 18338 18900 18350
rect 18844 18286 18846 18338
rect 18898 18286 18900 18338
rect 18844 18116 18900 18286
rect 18844 18050 18900 18060
rect 18844 17108 18900 17118
rect 18844 17014 18900 17052
rect 18172 16830 18174 16882
rect 18226 16830 18228 16882
rect 18172 16436 18228 16830
rect 18172 16370 18228 16380
rect 18284 16828 18788 16884
rect 18060 16258 18116 16268
rect 18284 16100 18340 16828
rect 17948 15262 17950 15314
rect 18002 15262 18004 15314
rect 17948 15250 18004 15262
rect 18060 16044 18340 16100
rect 18732 16212 18788 16222
rect 18732 16098 18788 16156
rect 18732 16046 18734 16098
rect 18786 16046 18788 16098
rect 18060 15148 18116 16044
rect 18732 16034 18788 16046
rect 18956 15876 19012 20524
rect 19292 20356 19348 22206
rect 19404 22260 19460 22270
rect 19516 22260 19572 23772
rect 19404 22258 19572 22260
rect 19404 22206 19406 22258
rect 19458 22206 19572 22258
rect 19404 22204 19572 22206
rect 19404 21476 19460 22204
rect 19628 22148 19684 23884
rect 19852 23874 19908 23884
rect 19740 23716 19796 23726
rect 19740 23622 19796 23660
rect 19964 23156 20020 23166
rect 19964 23062 20020 23100
rect 19404 20468 19460 21420
rect 19404 20402 19460 20412
rect 19516 22092 19684 22148
rect 19740 22820 19796 22830
rect 19068 20300 19348 20356
rect 19068 20132 19124 20300
rect 19516 20132 19572 22092
rect 19740 20356 19796 22764
rect 19964 22258 20020 22270
rect 19964 22206 19966 22258
rect 20018 22206 20020 22258
rect 19964 22148 20020 22206
rect 19964 22082 20020 22092
rect 19964 21474 20020 21486
rect 19964 21422 19966 21474
rect 20018 21422 20020 21474
rect 19964 20580 20020 21422
rect 19964 20514 20020 20524
rect 19068 20066 19124 20076
rect 19180 20076 19572 20132
rect 19628 20300 19796 20356
rect 19068 17556 19124 17566
rect 19180 17556 19236 20076
rect 19404 19460 19460 19470
rect 19404 19346 19460 19404
rect 19404 19294 19406 19346
rect 19458 19294 19460 19346
rect 19404 19282 19460 19294
rect 19404 18116 19460 18126
rect 19124 17500 19236 17556
rect 19292 17668 19348 17678
rect 19068 17490 19124 17500
rect 19292 17108 19348 17612
rect 19404 17554 19460 18060
rect 19628 17668 19684 20300
rect 20188 20244 20244 25228
rect 20524 24948 20580 26572
rect 20636 26562 20692 26572
rect 20300 24892 20580 24948
rect 20636 26290 20692 26302
rect 20636 26238 20638 26290
rect 20690 26238 20692 26290
rect 20300 22258 20356 24892
rect 20300 22206 20302 22258
rect 20354 22206 20356 22258
rect 20300 22194 20356 22206
rect 20412 24724 20468 24734
rect 19852 20188 20244 20244
rect 19740 20132 19796 20142
rect 19852 20132 19908 20188
rect 19740 20130 19908 20132
rect 19740 20078 19742 20130
rect 19794 20078 19908 20130
rect 19740 20076 19908 20078
rect 19740 20066 19796 20076
rect 19628 17574 19684 17612
rect 19964 20018 20020 20030
rect 19964 19966 19966 20018
rect 20018 19966 20020 20018
rect 19404 17502 19406 17554
rect 19458 17502 19460 17554
rect 19404 17490 19460 17502
rect 19516 17444 19572 17454
rect 19964 17444 20020 19966
rect 20076 19234 20132 20188
rect 20076 19182 20078 19234
rect 20130 19182 20132 19234
rect 20076 19170 20132 19182
rect 19572 17388 20020 17444
rect 20076 17668 20132 17678
rect 19516 17350 19572 17388
rect 19292 17042 19348 17052
rect 19404 17106 19460 17118
rect 19404 17054 19406 17106
rect 19458 17054 19460 17106
rect 19404 16996 19460 17054
rect 19852 17108 19908 17118
rect 19404 16930 19460 16940
rect 19740 16994 19796 17006
rect 19740 16942 19742 16994
rect 19794 16942 19796 16994
rect 19628 16436 19684 16446
rect 19068 15876 19124 15886
rect 18956 15874 19236 15876
rect 18956 15822 19070 15874
rect 19122 15822 19236 15874
rect 18956 15820 19236 15822
rect 19068 15810 19124 15820
rect 18348 15708 18612 15718
rect 18404 15652 18452 15708
rect 18508 15652 18556 15708
rect 18348 15642 18612 15652
rect 18060 15092 18228 15148
rect 17948 14420 18004 14430
rect 17500 14364 17948 14420
rect 17388 13972 17444 13982
rect 17388 13878 17444 13916
rect 17948 13858 18004 14364
rect 17948 13806 17950 13858
rect 18002 13806 18004 13858
rect 17948 13794 18004 13806
rect 17164 12404 17220 12414
rect 17164 11394 17220 12348
rect 17948 12180 18004 12190
rect 17948 12086 18004 12124
rect 17164 11342 17166 11394
rect 17218 11342 17220 11394
rect 17164 11330 17220 11342
rect 18172 9940 18228 15092
rect 19068 14644 19124 14654
rect 19068 14550 19124 14588
rect 18348 14140 18612 14150
rect 18404 14084 18452 14140
rect 18508 14084 18556 14140
rect 18348 14074 18612 14084
rect 18620 13636 18676 13646
rect 18620 13542 18676 13580
rect 18956 12740 19012 12750
rect 18732 12684 18956 12740
rect 18348 12572 18612 12582
rect 18404 12516 18452 12572
rect 18508 12516 18556 12572
rect 18348 12506 18612 12516
rect 18732 12290 18788 12684
rect 18956 12674 19012 12684
rect 18732 12238 18734 12290
rect 18786 12238 18788 12290
rect 18732 12226 18788 12238
rect 18348 11004 18612 11014
rect 18404 10948 18452 11004
rect 18508 10948 18556 11004
rect 18348 10938 18612 10948
rect 18284 9940 18340 9950
rect 17948 9938 18340 9940
rect 17948 9886 18286 9938
rect 18338 9886 18340 9938
rect 17948 9884 18340 9886
rect 17276 9716 17332 9726
rect 17500 9716 17556 9726
rect 17276 9714 17556 9716
rect 17276 9662 17278 9714
rect 17330 9662 17502 9714
rect 17554 9662 17556 9714
rect 17276 9660 17556 9662
rect 17276 9650 17332 9660
rect 17500 9650 17556 9660
rect 17836 9714 17892 9726
rect 17836 9662 17838 9714
rect 17890 9662 17892 9714
rect 16380 8754 16436 8764
rect 16828 8876 17052 8932
rect 16716 8260 16772 8270
rect 16716 8166 16772 8204
rect 16268 8082 16324 8092
rect 16828 8036 16884 8876
rect 17052 8866 17108 8876
rect 17164 9602 17220 9614
rect 17164 9550 17166 9602
rect 17218 9550 17220 9602
rect 16716 7980 16884 8036
rect 15708 7646 15710 7698
rect 15762 7646 15764 7698
rect 15708 7634 15764 7646
rect 15820 7700 15876 7710
rect 15820 7606 15876 7644
rect 16492 7586 16548 7598
rect 16492 7534 16494 7586
rect 16546 7534 16548 7586
rect 16268 7476 16324 7486
rect 16268 7382 16324 7420
rect 15036 7310 15038 7362
rect 15090 7310 15092 7362
rect 15036 7298 15092 7310
rect 15036 6804 15092 6814
rect 14924 6802 15092 6804
rect 14924 6750 15038 6802
rect 15090 6750 15092 6802
rect 14924 6748 15092 6750
rect 15036 6738 15092 6748
rect 16492 6580 16548 7534
rect 16716 7474 16772 7980
rect 16716 7422 16718 7474
rect 16770 7422 16772 7474
rect 16716 7410 16772 7422
rect 17164 6690 17220 9550
rect 17724 9602 17780 9614
rect 17724 9550 17726 9602
rect 17778 9550 17780 9602
rect 17388 9156 17444 9166
rect 17388 9062 17444 9100
rect 17612 9042 17668 9054
rect 17612 8990 17614 9042
rect 17666 8990 17668 9042
rect 17500 8930 17556 8942
rect 17500 8878 17502 8930
rect 17554 8878 17556 8930
rect 17500 8484 17556 8878
rect 17612 8820 17668 8990
rect 17612 8754 17668 8764
rect 17500 8418 17556 8428
rect 17724 8484 17780 9550
rect 17836 9156 17892 9662
rect 17836 9090 17892 9100
rect 17948 8596 18004 9884
rect 18284 9874 18340 9884
rect 18348 9436 18612 9446
rect 18404 9380 18452 9436
rect 18508 9380 18556 9436
rect 18348 9370 18612 9380
rect 18284 9156 18340 9166
rect 18284 9062 18340 9100
rect 17724 8418 17780 8428
rect 17836 8540 18004 8596
rect 18060 9042 18116 9054
rect 18060 8990 18062 9042
rect 18114 8990 18116 9042
rect 17388 7812 17444 7822
rect 17388 7698 17444 7756
rect 17388 7646 17390 7698
rect 17442 7646 17444 7698
rect 17388 7634 17444 7646
rect 17724 7700 17780 7710
rect 17836 7700 17892 8540
rect 17724 7698 17892 7700
rect 17724 7646 17726 7698
rect 17778 7646 17892 7698
rect 17724 7644 17892 7646
rect 17724 7634 17780 7644
rect 17164 6638 17166 6690
rect 17218 6638 17220 6690
rect 17164 6626 17220 6638
rect 16492 6514 16548 6524
rect 14588 6414 14590 6466
rect 14642 6414 14644 6466
rect 14252 5954 14308 5964
rect 14588 5796 14644 6414
rect 14812 6468 14868 6478
rect 14812 6374 14868 6412
rect 15820 6468 15876 6478
rect 15484 6018 15540 6030
rect 15484 5966 15486 6018
rect 15538 5966 15540 6018
rect 15148 5908 15204 5918
rect 15372 5908 15428 5918
rect 15148 5906 15428 5908
rect 15148 5854 15150 5906
rect 15202 5854 15374 5906
rect 15426 5854 15428 5906
rect 15148 5852 15428 5854
rect 15148 5842 15204 5852
rect 13804 5070 13806 5122
rect 13858 5070 13860 5122
rect 13804 5058 13860 5070
rect 13916 5628 14084 5684
rect 14476 5794 14644 5796
rect 14476 5742 14590 5794
rect 14642 5742 14644 5794
rect 14476 5740 14644 5742
rect 13356 4398 13358 4450
rect 13410 4398 13412 4450
rect 13356 4386 13412 4398
rect 13916 4226 13972 5628
rect 14064 5516 14328 5526
rect 14120 5460 14168 5516
rect 14224 5460 14272 5516
rect 14064 5450 14328 5460
rect 14028 5348 14084 5358
rect 14028 5122 14084 5292
rect 14028 5070 14030 5122
rect 14082 5070 14084 5122
rect 14028 5058 14084 5070
rect 13916 4174 13918 4226
rect 13970 4174 13972 4226
rect 13244 3502 13246 3554
rect 13298 3502 13300 3554
rect 13244 3490 13300 3502
rect 13580 3556 13636 3566
rect 13356 3444 13412 3482
rect 13580 3462 13636 3500
rect 13916 3556 13972 4174
rect 14064 3948 14328 3958
rect 14120 3892 14168 3948
rect 14224 3892 14272 3948
rect 14064 3882 14328 3892
rect 13916 3490 13972 3500
rect 14252 3556 14308 3566
rect 14476 3556 14532 5740
rect 14588 5730 14644 5740
rect 15372 5684 15428 5852
rect 15372 5618 15428 5628
rect 14588 5236 14644 5246
rect 14588 5142 14644 5180
rect 15484 5236 15540 5966
rect 15484 5170 15540 5180
rect 15708 5906 15764 5918
rect 15708 5854 15710 5906
rect 15762 5854 15764 5906
rect 14252 3554 14532 3556
rect 14252 3502 14254 3554
rect 14306 3502 14532 3554
rect 14252 3500 14532 3502
rect 14588 4900 14644 4910
rect 14252 3490 14308 3500
rect 12348 3332 12852 3388
rect 13356 3378 13412 3388
rect 12796 800 12852 3332
rect 14588 1876 14644 4844
rect 15708 4452 15764 5854
rect 15820 5906 15876 6412
rect 17164 6468 17220 6478
rect 15820 5854 15822 5906
rect 15874 5854 15876 5906
rect 15820 5842 15876 5854
rect 16156 6020 16212 6030
rect 16156 5906 16212 5964
rect 16156 5854 16158 5906
rect 16210 5854 16212 5906
rect 16156 5842 16212 5854
rect 16492 5906 16548 5918
rect 16492 5854 16494 5906
rect 16546 5854 16548 5906
rect 15708 4386 15764 4396
rect 16044 5794 16100 5806
rect 16044 5742 16046 5794
rect 16098 5742 16100 5794
rect 16044 4450 16100 5742
rect 16492 5796 16548 5854
rect 16492 5730 16548 5740
rect 17052 5236 17108 5246
rect 16716 5010 16772 5022
rect 16716 4958 16718 5010
rect 16770 4958 16772 5010
rect 16716 4564 16772 4958
rect 16716 4498 16772 4508
rect 16828 5012 16884 5022
rect 16044 4398 16046 4450
rect 16098 4398 16100 4450
rect 16044 4386 16100 4398
rect 16828 4340 16884 4956
rect 16828 4246 16884 4284
rect 17052 4228 17108 5180
rect 17052 4162 17108 4172
rect 17052 4004 17108 4014
rect 14364 1820 14644 1876
rect 15932 3666 15988 3678
rect 15932 3614 15934 3666
rect 15986 3614 15988 3666
rect 14364 800 14420 1820
rect 15932 800 15988 3614
rect 17052 3554 17108 3948
rect 17052 3502 17054 3554
rect 17106 3502 17108 3554
rect 17052 3490 17108 3502
rect 17164 3442 17220 6412
rect 17388 5908 17444 5918
rect 17388 5814 17444 5852
rect 17836 5684 17892 7644
rect 17388 5124 17444 5134
rect 17276 4338 17332 4350
rect 17276 4286 17278 4338
rect 17330 4286 17332 4338
rect 17276 3780 17332 4286
rect 17276 3714 17332 3724
rect 17388 3554 17444 5068
rect 17500 5122 17556 5134
rect 17500 5070 17502 5122
rect 17554 5070 17556 5122
rect 17500 5012 17556 5070
rect 17500 4946 17556 4956
rect 17500 4564 17556 4574
rect 17500 4470 17556 4508
rect 17836 4564 17892 5628
rect 17948 8372 18004 8382
rect 17948 6690 18004 8316
rect 18060 7364 18116 8990
rect 18620 9044 18676 9054
rect 18620 8950 18676 8988
rect 18348 7868 18612 7878
rect 18404 7812 18452 7868
rect 18508 7812 18556 7868
rect 18348 7802 18612 7812
rect 18396 7700 18452 7710
rect 18396 7606 18452 7644
rect 18508 7588 18564 7598
rect 18508 7494 18564 7532
rect 18844 7586 18900 7598
rect 18844 7534 18846 7586
rect 18898 7534 18900 7586
rect 18172 7476 18228 7486
rect 18172 7382 18228 7420
rect 18060 7298 18116 7308
rect 18844 6804 18900 7534
rect 19180 7586 19236 15820
rect 19404 14308 19460 14318
rect 19404 13858 19460 14252
rect 19516 14084 19572 14094
rect 19516 13970 19572 14028
rect 19516 13918 19518 13970
rect 19570 13918 19572 13970
rect 19516 13906 19572 13918
rect 19628 13972 19684 16380
rect 19740 15876 19796 16942
rect 19852 16882 19908 17052
rect 19852 16830 19854 16882
rect 19906 16830 19908 16882
rect 19852 16818 19908 16830
rect 20076 16660 20132 17612
rect 19852 16604 20132 16660
rect 20300 17666 20356 17678
rect 20300 17614 20302 17666
rect 20354 17614 20356 17666
rect 20300 16660 20356 17614
rect 19852 16210 19908 16604
rect 19852 16158 19854 16210
rect 19906 16158 19908 16210
rect 19852 16146 19908 16158
rect 20300 16210 20356 16604
rect 20412 16548 20468 24668
rect 20636 23828 20692 26238
rect 20748 26292 20804 26796
rect 20860 26516 20916 26554
rect 20860 26450 20916 26460
rect 20860 26292 20916 26302
rect 20748 26290 20916 26292
rect 20748 26238 20862 26290
rect 20914 26238 20916 26290
rect 20748 26236 20916 26238
rect 20860 26226 20916 26236
rect 20972 26290 21028 26302
rect 20972 26238 20974 26290
rect 21026 26238 21028 26290
rect 20748 25282 20804 25294
rect 20748 25230 20750 25282
rect 20802 25230 20804 25282
rect 20748 24724 20804 25230
rect 20972 25284 21028 26238
rect 20972 25218 21028 25228
rect 21084 24724 21140 24734
rect 20748 24722 21140 24724
rect 20748 24670 21086 24722
rect 21138 24670 21140 24722
rect 20748 24668 21140 24670
rect 20636 23762 20692 23772
rect 20860 23716 20916 23726
rect 20636 23044 20692 23054
rect 20636 22950 20692 22988
rect 20748 22260 20804 22270
rect 20748 22166 20804 22204
rect 20748 21586 20804 21598
rect 20748 21534 20750 21586
rect 20802 21534 20804 21586
rect 20748 21476 20804 21534
rect 20748 21410 20804 21420
rect 20748 20356 20804 20366
rect 20636 19908 20692 19918
rect 20636 19814 20692 19852
rect 20524 19236 20580 19246
rect 20524 19142 20580 19180
rect 20636 19012 20692 19022
rect 20412 16482 20468 16492
rect 20524 19010 20692 19012
rect 20524 18958 20638 19010
rect 20690 18958 20692 19010
rect 20524 18956 20692 18958
rect 20300 16158 20302 16210
rect 20354 16158 20356 16210
rect 20300 16146 20356 16158
rect 19740 15148 19796 15820
rect 20412 15202 20468 15214
rect 20412 15150 20414 15202
rect 20466 15150 20468 15202
rect 19740 15092 20356 15148
rect 19852 14530 19908 14542
rect 19852 14478 19854 14530
rect 19906 14478 19908 14530
rect 19852 14420 19908 14478
rect 19852 14354 19908 14364
rect 20076 14196 20132 14206
rect 19740 13972 19796 13982
rect 19628 13970 19796 13972
rect 19628 13918 19742 13970
rect 19794 13918 19796 13970
rect 19628 13916 19796 13918
rect 19740 13906 19796 13916
rect 19404 13806 19406 13858
rect 19458 13806 19460 13858
rect 19404 13794 19460 13806
rect 19964 13860 20020 13870
rect 19964 13766 20020 13804
rect 20076 13858 20132 14140
rect 20300 13972 20356 15092
rect 20412 14530 20468 15150
rect 20412 14478 20414 14530
rect 20466 14478 20468 14530
rect 20412 14308 20468 14478
rect 20412 14242 20468 14252
rect 20412 13972 20468 13982
rect 20300 13970 20468 13972
rect 20300 13918 20414 13970
rect 20466 13918 20468 13970
rect 20300 13916 20468 13918
rect 20412 13906 20468 13916
rect 20076 13806 20078 13858
rect 20130 13806 20132 13858
rect 20076 13794 20132 13806
rect 20524 12962 20580 18956
rect 20636 18946 20692 18956
rect 20748 18116 20804 20300
rect 20860 18340 20916 23660
rect 20860 18274 20916 18284
rect 20748 18050 20804 18060
rect 20636 17892 20692 17902
rect 20972 17892 21028 24668
rect 21084 24658 21140 24668
rect 21084 23716 21140 23726
rect 21196 23716 21252 28588
rect 21308 28532 21364 28542
rect 21308 28438 21364 28476
rect 21420 28420 21476 30940
rect 21532 30930 21588 30940
rect 21532 30100 21588 30110
rect 21532 28642 21588 30044
rect 21532 28590 21534 28642
rect 21586 28590 21588 28642
rect 21532 28578 21588 28590
rect 21420 27858 21476 28364
rect 21644 28082 21700 31612
rect 22092 31666 22148 31678
rect 22092 31614 22094 31666
rect 22146 31614 22148 31666
rect 21756 31554 21812 31566
rect 21756 31502 21758 31554
rect 21810 31502 21812 31554
rect 21756 30434 21812 31502
rect 22092 31444 22148 31614
rect 22148 31388 22260 31444
rect 22092 31378 22148 31388
rect 21756 30382 21758 30434
rect 21810 30382 21812 30434
rect 21756 30370 21812 30382
rect 21868 30324 21924 30334
rect 21756 30212 21812 30222
rect 21756 29986 21812 30156
rect 21868 30210 21924 30268
rect 21868 30158 21870 30210
rect 21922 30158 21924 30210
rect 21868 30146 21924 30158
rect 22092 30100 22148 30110
rect 21980 29988 22036 29998
rect 21756 29934 21758 29986
rect 21810 29934 21812 29986
rect 21756 29922 21812 29934
rect 21868 29932 21980 29988
rect 21868 28866 21924 29932
rect 21980 29922 22036 29932
rect 21868 28814 21870 28866
rect 21922 28814 21924 28866
rect 21868 28802 21924 28814
rect 21980 29204 22036 29214
rect 21980 28642 22036 29148
rect 21980 28590 21982 28642
rect 22034 28590 22036 28642
rect 21980 28578 22036 28590
rect 22092 28418 22148 30044
rect 22204 29540 22260 31388
rect 22204 29474 22260 29484
rect 22092 28366 22094 28418
rect 22146 28366 22148 28418
rect 22092 28354 22148 28366
rect 22316 28308 22372 31836
rect 22428 31826 22484 31836
rect 22540 32004 22596 32014
rect 22540 30772 22596 31948
rect 22652 31778 22708 31790
rect 22652 31726 22654 31778
rect 22706 31726 22708 31778
rect 22652 31332 22708 31726
rect 22988 31556 23044 31566
rect 22988 31462 23044 31500
rect 23100 31332 23156 33852
rect 23772 33458 23828 33470
rect 23772 33406 23774 33458
rect 23826 33406 23828 33458
rect 23324 32564 23380 32574
rect 23324 31778 23380 32508
rect 23436 32450 23492 32462
rect 23436 32398 23438 32450
rect 23490 32398 23492 32450
rect 23436 32340 23492 32398
rect 23436 32274 23492 32284
rect 23772 32004 23828 33406
rect 23884 32564 23940 32574
rect 24108 32564 24164 32574
rect 24556 32564 24612 32574
rect 23940 32562 24612 32564
rect 23940 32510 24110 32562
rect 24162 32510 24558 32562
rect 24610 32510 24612 32562
rect 23940 32508 24612 32510
rect 23884 32498 23940 32508
rect 24108 32498 24164 32508
rect 23772 31938 23828 31948
rect 23324 31726 23326 31778
rect 23378 31726 23380 31778
rect 23324 31714 23380 31726
rect 23548 31668 23604 31678
rect 24108 31668 24164 31678
rect 22652 31266 22708 31276
rect 22988 31276 23156 31332
rect 23212 31332 23268 31342
rect 23268 31276 23380 31332
rect 22764 30996 22820 31006
rect 22764 30902 22820 30940
rect 22652 30882 22708 30894
rect 22652 30830 22654 30882
rect 22706 30830 22708 30882
rect 22652 30772 22708 30830
rect 22428 30716 22708 30772
rect 22428 29428 22484 30716
rect 22632 30604 22896 30614
rect 22688 30548 22736 30604
rect 22792 30548 22840 30604
rect 22632 30538 22896 30548
rect 22652 29988 22708 29998
rect 22652 29986 22932 29988
rect 22652 29934 22654 29986
rect 22706 29934 22932 29986
rect 22652 29932 22932 29934
rect 22652 29922 22708 29932
rect 22764 29428 22820 29438
rect 22428 29372 22764 29428
rect 22764 29334 22820 29372
rect 22876 29204 22932 29932
rect 22876 29138 22932 29148
rect 22632 29036 22896 29046
rect 22688 28980 22736 29036
rect 22792 28980 22840 29036
rect 22632 28970 22896 28980
rect 22204 28196 22260 28206
rect 21644 28030 21646 28082
rect 21698 28030 21700 28082
rect 21644 28018 21700 28030
rect 21756 28084 21812 28094
rect 21420 27806 21422 27858
rect 21474 27806 21476 27858
rect 21420 27794 21476 27806
rect 21756 27970 21812 28028
rect 21756 27918 21758 27970
rect 21810 27918 21812 27970
rect 21308 27748 21364 27758
rect 21308 27654 21364 27692
rect 21756 27300 21812 27918
rect 21756 27234 21812 27244
rect 21868 27860 21924 27870
rect 21868 27076 21924 27804
rect 22204 27300 22260 28140
rect 22316 27858 22372 28252
rect 22988 28084 23044 31276
rect 23212 31266 23268 31276
rect 23324 30436 23380 31276
rect 23548 31106 23604 31612
rect 23548 31054 23550 31106
rect 23602 31054 23604 31106
rect 23548 31042 23604 31054
rect 23884 31666 24164 31668
rect 23884 31614 24110 31666
rect 24162 31614 24164 31666
rect 23884 31612 24164 31614
rect 23436 30996 23492 31006
rect 23436 30902 23492 30940
rect 23548 30884 23604 30894
rect 23548 30790 23604 30828
rect 23324 30380 23492 30436
rect 23324 30210 23380 30222
rect 23324 30158 23326 30210
rect 23378 30158 23380 30210
rect 23100 30098 23156 30110
rect 23100 30046 23102 30098
rect 23154 30046 23156 30098
rect 23100 28308 23156 30046
rect 23212 29988 23268 29998
rect 23212 29894 23268 29932
rect 23324 29876 23380 30158
rect 23324 29810 23380 29820
rect 23212 29314 23268 29326
rect 23212 29262 23214 29314
rect 23266 29262 23268 29314
rect 23212 29204 23268 29262
rect 23212 29138 23268 29148
rect 23100 28252 23268 28308
rect 23100 28084 23156 28094
rect 22988 28082 23156 28084
rect 22988 28030 23102 28082
rect 23154 28030 23156 28082
rect 22988 28028 23156 28030
rect 23100 28018 23156 28028
rect 23212 27972 23268 28252
rect 23212 27906 23268 27916
rect 22316 27806 22318 27858
rect 22370 27806 22372 27858
rect 22316 27794 22372 27806
rect 22428 27860 22484 27870
rect 22204 27244 22372 27300
rect 22204 27076 22260 27086
rect 21756 27074 21924 27076
rect 21756 27022 21870 27074
rect 21922 27022 21924 27074
rect 21756 27020 21924 27022
rect 21308 26962 21364 26974
rect 21308 26910 21310 26962
rect 21362 26910 21364 26962
rect 21308 25844 21364 26910
rect 21420 26852 21476 26862
rect 21420 26758 21476 26796
rect 21644 26850 21700 26862
rect 21644 26798 21646 26850
rect 21698 26798 21700 26850
rect 21308 25778 21364 25788
rect 21420 26068 21476 26078
rect 21420 25730 21476 26012
rect 21420 25678 21422 25730
rect 21474 25678 21476 25730
rect 21420 25666 21476 25678
rect 21532 25732 21588 25742
rect 21644 25732 21700 26798
rect 21756 26628 21812 27020
rect 21868 27010 21924 27020
rect 22092 27074 22260 27076
rect 22092 27022 22206 27074
rect 22258 27022 22260 27074
rect 22092 27020 22260 27022
rect 21756 26562 21812 26572
rect 22092 26516 22148 27020
rect 22204 27010 22260 27020
rect 22316 26908 22372 27244
rect 22428 27076 22484 27804
rect 22632 27468 22896 27478
rect 22688 27412 22736 27468
rect 22792 27412 22840 27468
rect 22632 27402 22896 27412
rect 22428 26982 22484 27020
rect 22652 27300 22708 27310
rect 22652 27074 22708 27244
rect 23100 27300 23156 27310
rect 23436 27300 23492 30380
rect 23884 30212 23940 31612
rect 24108 31602 24164 31612
rect 23884 30146 23940 30156
rect 24220 30884 24276 32508
rect 24556 32498 24612 32508
rect 24220 30210 24276 30828
rect 24220 30158 24222 30210
rect 24274 30158 24276 30210
rect 23660 30098 23716 30110
rect 23660 30046 23662 30098
rect 23714 30046 23716 30098
rect 23660 29652 23716 30046
rect 23660 29586 23716 29596
rect 24108 29652 24164 29662
rect 24108 29558 24164 29596
rect 23772 29316 23828 29326
rect 23772 28644 23828 29260
rect 23772 28550 23828 28588
rect 23156 27244 23268 27300
rect 23100 27234 23156 27244
rect 22652 27022 22654 27074
rect 22706 27022 22708 27074
rect 22652 27010 22708 27022
rect 22092 26450 22148 26460
rect 22204 26852 22372 26908
rect 22540 26964 22596 27002
rect 22540 26898 22596 26908
rect 23212 26908 23268 27244
rect 23436 27234 23492 27244
rect 23324 27076 23380 27086
rect 23772 27076 23828 27086
rect 23324 27074 23828 27076
rect 23324 27022 23326 27074
rect 23378 27022 23774 27074
rect 23826 27022 23828 27074
rect 23324 27020 23828 27022
rect 23324 27010 23380 27020
rect 23772 26908 23828 27020
rect 24220 26908 24276 30158
rect 24556 30994 24612 31006
rect 24556 30942 24558 30994
rect 24610 30942 24612 30994
rect 24556 28308 24612 30942
rect 24668 30660 24724 36204
rect 25088 36200 25200 37000
rect 26208 36200 26320 37000
rect 27328 36200 27440 37000
rect 28448 36200 28560 37000
rect 29568 36200 29680 37000
rect 30688 36200 30800 37000
rect 30940 36204 31668 36260
rect 24780 33346 24836 33358
rect 24780 33294 24782 33346
rect 24834 33294 24836 33346
rect 24780 31892 24836 33294
rect 25116 32004 25172 36200
rect 25564 33572 25620 33582
rect 25564 33478 25620 33516
rect 25228 33460 25284 33470
rect 25228 32562 25284 33404
rect 26236 32676 26292 36200
rect 27356 33348 27412 36200
rect 27356 33282 27412 33292
rect 27580 33124 27636 33134
rect 27356 33122 27636 33124
rect 27356 33070 27582 33122
rect 27634 33070 27636 33122
rect 27356 33068 27636 33070
rect 26916 32956 27180 32966
rect 26972 32900 27020 32956
rect 27076 32900 27124 32956
rect 26916 32890 27180 32900
rect 26236 32620 26516 32676
rect 25228 32510 25230 32562
rect 25282 32510 25284 32562
rect 25228 32498 25284 32510
rect 26236 32452 26292 32462
rect 26236 32358 26292 32396
rect 25116 31948 25284 32004
rect 24780 31826 24836 31836
rect 24668 30594 24724 30604
rect 25228 30548 25284 31948
rect 25340 31556 25396 31566
rect 25340 31218 25396 31500
rect 25340 31166 25342 31218
rect 25394 31166 25396 31218
rect 25340 31154 25396 31166
rect 26348 31554 26404 31566
rect 26348 31502 26350 31554
rect 26402 31502 26404 31554
rect 26348 31444 26404 31502
rect 26460 31556 26516 32620
rect 26460 31490 26516 31500
rect 26684 32228 26740 32238
rect 25452 31108 25508 31118
rect 25452 31014 25508 31052
rect 25900 30884 25956 30894
rect 25340 30772 25396 30782
rect 25340 30678 25396 30716
rect 25228 30492 25508 30548
rect 25340 30324 25396 30334
rect 24892 30100 24948 30110
rect 24892 30006 24948 30044
rect 24556 28242 24612 28252
rect 24668 29652 24724 29662
rect 22652 26852 22708 26862
rect 23212 26852 23380 26908
rect 21868 26292 21924 26302
rect 22204 26292 22260 26852
rect 22540 26740 22596 26750
rect 22540 26514 22596 26684
rect 22540 26462 22542 26514
rect 22594 26462 22596 26514
rect 22540 26450 22596 26462
rect 22652 26514 22708 26796
rect 22652 26462 22654 26514
rect 22706 26462 22708 26514
rect 22652 26450 22708 26462
rect 21756 26180 21812 26190
rect 21756 26086 21812 26124
rect 21868 26066 21924 26236
rect 21868 26014 21870 26066
rect 21922 26014 21924 26066
rect 21868 25844 21924 26014
rect 21868 25778 21924 25788
rect 21980 26236 22260 26292
rect 22428 26404 22484 26414
rect 21532 25730 21700 25732
rect 21532 25678 21534 25730
rect 21586 25678 21700 25730
rect 21532 25676 21700 25678
rect 21756 25732 21812 25742
rect 21532 25666 21588 25676
rect 21756 25394 21812 25676
rect 21756 25342 21758 25394
rect 21810 25342 21812 25394
rect 21756 25330 21812 25342
rect 21756 25172 21812 25182
rect 21532 23940 21588 23950
rect 21532 23846 21588 23884
rect 21140 23660 21252 23716
rect 21308 23826 21364 23838
rect 21308 23774 21310 23826
rect 21362 23774 21364 23826
rect 21084 23650 21140 23660
rect 21308 23604 21364 23774
rect 21756 23826 21812 25116
rect 21980 24610 22036 26236
rect 22092 26066 22148 26078
rect 22092 26014 22094 26066
rect 22146 26014 22148 26066
rect 22092 25844 22148 26014
rect 22204 26068 22260 26078
rect 22204 25974 22260 26012
rect 22428 25844 22484 26348
rect 23212 26404 23268 26414
rect 22764 26292 22820 26302
rect 22764 26198 22820 26236
rect 23212 26290 23268 26348
rect 23212 26238 23214 26290
rect 23266 26238 23268 26290
rect 23212 26226 23268 26238
rect 23324 26290 23380 26852
rect 23324 26238 23326 26290
rect 23378 26238 23380 26290
rect 23324 26226 23380 26238
rect 23660 26852 23716 26862
rect 23660 26290 23716 26796
rect 23660 26238 23662 26290
rect 23714 26238 23716 26290
rect 23548 26068 23604 26078
rect 23324 26066 23604 26068
rect 23324 26014 23550 26066
rect 23602 26014 23604 26066
rect 23324 26012 23604 26014
rect 22092 25788 22484 25844
rect 22632 25900 22896 25910
rect 22688 25844 22736 25900
rect 22792 25844 22840 25900
rect 22632 25834 22896 25844
rect 22428 25620 22484 25630
rect 22428 25618 22932 25620
rect 22428 25566 22430 25618
rect 22482 25566 22932 25618
rect 22428 25564 22932 25566
rect 22428 25554 22484 25564
rect 22092 25396 22148 25406
rect 22092 25302 22148 25340
rect 22316 25394 22372 25406
rect 22316 25342 22318 25394
rect 22370 25342 22372 25394
rect 21980 24558 21982 24610
rect 22034 24558 22036 24610
rect 21980 24546 22036 24558
rect 22316 23940 22372 25342
rect 22876 24834 22932 25564
rect 22988 25396 23044 25406
rect 22988 24946 23044 25340
rect 23100 25284 23156 25294
rect 23100 25190 23156 25228
rect 22988 24894 22990 24946
rect 23042 24894 23044 24946
rect 22988 24882 23044 24894
rect 22876 24782 22878 24834
rect 22930 24782 22932 24834
rect 22876 24770 22932 24782
rect 22652 24722 22708 24734
rect 22652 24670 22654 24722
rect 22706 24670 22708 24722
rect 22652 24500 22708 24670
rect 23324 24722 23380 26012
rect 23548 26002 23604 26012
rect 23324 24670 23326 24722
rect 23378 24670 23380 24722
rect 23324 24658 23380 24670
rect 23436 25506 23492 25518
rect 23436 25454 23438 25506
rect 23490 25454 23492 25506
rect 23436 25284 23492 25454
rect 22316 23874 22372 23884
rect 22428 24444 22708 24500
rect 23436 24500 23492 25228
rect 23660 25172 23716 26238
rect 23660 25106 23716 25116
rect 23772 26852 24276 26908
rect 24444 26964 24500 27002
rect 24444 26898 24500 26908
rect 23772 24724 23828 26852
rect 24668 26516 24724 29596
rect 25228 29428 25284 29438
rect 25228 29334 25284 29372
rect 25228 28308 25284 28318
rect 25228 27858 25284 28252
rect 25228 27806 25230 27858
rect 25282 27806 25284 27858
rect 25228 27794 25284 27806
rect 24668 26422 24724 26460
rect 24892 27636 24948 27646
rect 23884 26404 23940 26414
rect 23884 25620 23940 26348
rect 23884 25554 23940 25564
rect 24220 25396 24276 25406
rect 24220 25302 24276 25340
rect 23772 24610 23828 24668
rect 23772 24558 23774 24610
rect 23826 24558 23828 24610
rect 23772 24500 23828 24558
rect 23436 24444 23828 24500
rect 24220 24948 24276 24958
rect 21756 23774 21758 23826
rect 21810 23774 21812 23826
rect 21756 23762 21812 23774
rect 21308 23538 21364 23548
rect 21868 23714 21924 23726
rect 21868 23662 21870 23714
rect 21922 23662 21924 23714
rect 21644 23044 21700 23054
rect 21532 22932 21588 22942
rect 21532 22370 21588 22876
rect 21532 22318 21534 22370
rect 21586 22318 21588 22370
rect 21532 22306 21588 22318
rect 21308 22260 21364 22270
rect 21308 22166 21364 22204
rect 21644 22146 21700 22988
rect 21868 22370 21924 23662
rect 21868 22318 21870 22370
rect 21922 22318 21924 22370
rect 21868 22306 21924 22318
rect 22316 23716 22372 23726
rect 22428 23716 22484 24444
rect 22632 24332 22896 24342
rect 22688 24276 22736 24332
rect 22792 24276 22840 24332
rect 22632 24266 22896 24276
rect 22316 23714 22484 23716
rect 22316 23662 22318 23714
rect 22370 23662 22484 23714
rect 22316 23660 22484 23662
rect 22764 23940 22820 23950
rect 22316 22260 22372 23660
rect 22764 23042 22820 23884
rect 23212 23156 23268 23166
rect 23436 23156 23492 24444
rect 23996 24276 24052 24286
rect 23996 24162 24052 24220
rect 23996 24110 23998 24162
rect 24050 24110 24052 24162
rect 23996 24098 24052 24110
rect 23884 24052 23940 24062
rect 23548 23940 23604 23950
rect 23884 23940 23940 23996
rect 23548 23938 23940 23940
rect 23548 23886 23550 23938
rect 23602 23886 23886 23938
rect 23938 23886 23940 23938
rect 23548 23884 23940 23886
rect 23548 23874 23604 23884
rect 23884 23874 23940 23884
rect 23268 23100 23492 23156
rect 23548 23492 23604 23502
rect 23212 23062 23268 23100
rect 22764 22990 22766 23042
rect 22818 22990 22820 23042
rect 22764 22978 22820 22990
rect 22632 22764 22896 22774
rect 22688 22708 22736 22764
rect 22792 22708 22840 22764
rect 22632 22698 22896 22708
rect 23548 22596 23604 23436
rect 24220 23380 24276 24892
rect 24332 24610 24388 24622
rect 24332 24558 24334 24610
rect 24386 24558 24388 24610
rect 24332 24052 24388 24558
rect 24332 23986 24388 23996
rect 24780 24610 24836 24622
rect 24780 24558 24782 24610
rect 24834 24558 24836 24610
rect 24780 23940 24836 24558
rect 24556 23884 24836 23940
rect 24332 23826 24388 23838
rect 24332 23774 24334 23826
rect 24386 23774 24388 23826
rect 24332 23604 24388 23774
rect 24332 23538 24388 23548
rect 24444 23716 24500 23726
rect 24556 23716 24612 23884
rect 24444 23714 24612 23716
rect 24444 23662 24446 23714
rect 24498 23662 24612 23714
rect 24444 23660 24612 23662
rect 24668 23714 24724 23726
rect 24668 23662 24670 23714
rect 24722 23662 24724 23714
rect 24332 23380 24388 23390
rect 24220 23378 24388 23380
rect 24220 23326 24334 23378
rect 24386 23326 24388 23378
rect 24220 23324 24388 23326
rect 24332 23314 24388 23324
rect 24444 23268 24500 23660
rect 24668 23380 24724 23662
rect 24668 23314 24724 23324
rect 24444 23202 24500 23212
rect 24556 23266 24612 23278
rect 24556 23214 24558 23266
rect 24610 23214 24612 23266
rect 23660 23044 23716 23054
rect 23660 22950 23716 22988
rect 24108 23044 24164 23054
rect 24556 23044 24612 23214
rect 24108 23042 24612 23044
rect 24108 22990 24110 23042
rect 24162 22990 24612 23042
rect 24108 22988 24612 22990
rect 24668 23154 24724 23166
rect 24668 23102 24670 23154
rect 24722 23102 24724 23154
rect 22316 22194 22372 22204
rect 22876 22370 22932 22382
rect 22876 22318 22878 22370
rect 22930 22318 22932 22370
rect 21644 22094 21646 22146
rect 21698 22094 21700 22146
rect 21644 22082 21700 22094
rect 21084 21812 21140 21822
rect 21084 21718 21140 21756
rect 21420 21586 21476 21598
rect 21420 21534 21422 21586
rect 21474 21534 21476 21586
rect 21420 20244 21476 21534
rect 21868 21476 21924 21486
rect 21868 21382 21924 21420
rect 22540 21474 22596 21486
rect 22540 21422 22542 21474
rect 22594 21422 22596 21474
rect 21644 21362 21700 21374
rect 21644 21310 21646 21362
rect 21698 21310 21700 21362
rect 21420 20178 21476 20188
rect 21532 20580 21588 20590
rect 21644 20580 21700 21310
rect 22540 21364 22596 21422
rect 22876 21476 22932 22318
rect 22876 21410 22932 21420
rect 22988 21474 23044 21486
rect 22988 21422 22990 21474
rect 23042 21422 23044 21474
rect 22540 21298 22596 21308
rect 22988 21362 23044 21422
rect 22988 21310 22990 21362
rect 23042 21310 23044 21362
rect 22988 21298 23044 21310
rect 23324 21474 23380 21486
rect 23324 21422 23326 21474
rect 23378 21422 23380 21474
rect 23324 21362 23380 21422
rect 23324 21310 23326 21362
rect 23378 21310 23380 21362
rect 22632 21196 22896 21206
rect 22688 21140 22736 21196
rect 22792 21140 22840 21196
rect 22632 21130 22896 21140
rect 22764 20916 22820 20926
rect 22764 20822 22820 20860
rect 21532 20578 21700 20580
rect 21532 20526 21534 20578
rect 21586 20526 21700 20578
rect 21532 20524 21700 20526
rect 21868 20690 21924 20702
rect 21868 20638 21870 20690
rect 21922 20638 21924 20690
rect 20636 17890 21028 17892
rect 20636 17838 20638 17890
rect 20690 17838 21028 17890
rect 20636 17836 21028 17838
rect 21084 20018 21140 20030
rect 21084 19966 21086 20018
rect 21138 19966 21140 20018
rect 21084 19124 21140 19966
rect 21420 19124 21476 19134
rect 21532 19124 21588 20524
rect 21084 19122 21588 19124
rect 21084 19070 21422 19122
rect 21474 19070 21588 19122
rect 21084 19068 21588 19070
rect 21644 20018 21700 20030
rect 21644 19966 21646 20018
rect 21698 19966 21700 20018
rect 20636 17826 20692 17836
rect 20748 17554 20804 17566
rect 20748 17502 20750 17554
rect 20802 17502 20804 17554
rect 20748 17220 20804 17502
rect 20860 17220 20916 17230
rect 20748 17164 20860 17220
rect 20860 17106 20916 17164
rect 20860 17054 20862 17106
rect 20914 17054 20916 17106
rect 20860 17042 20916 17054
rect 20636 16884 20692 16894
rect 20636 14642 20692 16828
rect 21084 16772 21140 19068
rect 21420 19058 21476 19068
rect 21644 18564 21700 19966
rect 21756 19906 21812 19918
rect 21756 19854 21758 19906
rect 21810 19854 21812 19906
rect 21756 19236 21812 19854
rect 21756 19170 21812 19180
rect 21644 18498 21700 18508
rect 21644 18340 21700 18350
rect 21420 18116 21476 18126
rect 21420 17778 21476 18060
rect 21420 17726 21422 17778
rect 21474 17726 21476 17778
rect 21420 17714 21476 17726
rect 21644 17556 21700 18284
rect 21308 17500 21700 17556
rect 21868 18228 21924 20638
rect 22876 20580 22932 20590
rect 22092 20018 22148 20030
rect 22092 19966 22094 20018
rect 22146 19966 22148 20018
rect 22092 19908 22148 19966
rect 22876 20018 22932 20524
rect 22876 19966 22878 20018
rect 22930 19966 22932 20018
rect 22876 19954 22932 19966
rect 22092 19124 22148 19852
rect 22988 19908 23044 19918
rect 22988 19814 23044 19852
rect 22632 19628 22896 19638
rect 22688 19572 22736 19628
rect 22792 19572 22840 19628
rect 22632 19562 22896 19572
rect 23212 19234 23268 19246
rect 23212 19182 23214 19234
rect 23266 19182 23268 19234
rect 22428 19124 22484 19134
rect 22092 19122 22484 19124
rect 22092 19070 22430 19122
rect 22482 19070 22484 19122
rect 22092 19068 22484 19070
rect 22428 18788 22484 19068
rect 22764 19122 22820 19134
rect 22764 19070 22766 19122
rect 22818 19070 22820 19122
rect 22652 19012 22708 19022
rect 22652 18918 22708 18956
rect 22428 18722 22484 18732
rect 22764 18228 22820 19070
rect 23212 19012 23268 19182
rect 23212 18946 23268 18956
rect 21868 18172 22820 18228
rect 23212 18452 23268 18462
rect 23324 18452 23380 21310
rect 23436 20916 23492 20926
rect 23548 20916 23604 22540
rect 23660 22258 23716 22270
rect 23660 22206 23662 22258
rect 23714 22206 23716 22258
rect 23660 21812 23716 22206
rect 23660 21746 23716 21756
rect 23772 21474 23828 21486
rect 23772 21422 23774 21474
rect 23826 21422 23828 21474
rect 23772 21362 23828 21422
rect 23772 21310 23774 21362
rect 23826 21310 23828 21362
rect 23772 21298 23828 21310
rect 23436 20914 23604 20916
rect 23436 20862 23438 20914
rect 23490 20862 23604 20914
rect 23436 20860 23604 20862
rect 23996 21252 24052 21262
rect 23996 20916 24052 21196
rect 23436 20850 23492 20860
rect 23548 20244 23604 20254
rect 23548 20150 23604 20188
rect 23996 20130 24052 20860
rect 23996 20078 23998 20130
rect 24050 20078 24052 20130
rect 23996 20066 24052 20078
rect 23660 19908 23716 19918
rect 23660 19010 23716 19852
rect 23660 18958 23662 19010
rect 23714 18958 23716 19010
rect 23268 18396 23380 18452
rect 23436 18450 23492 18462
rect 23436 18398 23438 18450
rect 23490 18398 23492 18450
rect 21196 16772 21252 16782
rect 21084 16716 21196 16772
rect 20748 16100 20804 16110
rect 20748 16006 20804 16044
rect 21196 15538 21252 16716
rect 21196 15486 21198 15538
rect 21250 15486 21252 15538
rect 21196 15474 21252 15486
rect 20748 14756 20804 14766
rect 20748 14662 20804 14700
rect 20636 14590 20638 14642
rect 20690 14590 20692 14642
rect 20636 14578 20692 14590
rect 21308 14308 21364 17500
rect 21868 17442 21924 18172
rect 22632 18060 22896 18070
rect 22688 18004 22736 18060
rect 22792 18004 22840 18060
rect 22632 17994 22896 18004
rect 22988 18004 23044 18014
rect 21868 17390 21870 17442
rect 21922 17390 21924 17442
rect 21420 16884 21476 16894
rect 21756 16884 21812 16894
rect 21420 16882 21812 16884
rect 21420 16830 21422 16882
rect 21474 16830 21758 16882
rect 21810 16830 21812 16882
rect 21420 16828 21812 16830
rect 21420 16818 21476 16828
rect 21420 16548 21476 16558
rect 21420 16322 21476 16492
rect 21420 16270 21422 16322
rect 21474 16270 21476 16322
rect 21420 16258 21476 16270
rect 21756 16324 21812 16828
rect 21868 16772 21924 17390
rect 21980 17668 22036 17678
rect 21980 16996 22036 17612
rect 21980 16902 22036 16940
rect 22316 17666 22372 17678
rect 22316 17614 22318 17666
rect 22370 17614 22372 17666
rect 22316 16996 22372 17614
rect 22988 17668 23044 17948
rect 22988 17574 23044 17612
rect 22428 17556 22484 17566
rect 22428 17462 22484 17500
rect 22652 17556 22708 17566
rect 22652 17462 22708 17500
rect 23212 17444 23268 18396
rect 22988 17388 23268 17444
rect 22372 16940 22484 16996
rect 22316 16930 22372 16940
rect 22204 16884 22260 16894
rect 22204 16790 22260 16828
rect 21868 16716 22036 16772
rect 21756 16268 21924 16324
rect 21756 16100 21812 16110
rect 21756 16006 21812 16044
rect 21868 15988 21924 16268
rect 21980 16212 22036 16716
rect 22092 16212 22148 16222
rect 21980 16156 22092 16212
rect 22092 16146 22148 16156
rect 21980 15988 22036 15998
rect 21868 15986 22148 15988
rect 21868 15934 21982 15986
rect 22034 15934 22148 15986
rect 21868 15932 22148 15934
rect 21980 15922 22036 15932
rect 21756 15316 21812 15326
rect 21756 15222 21812 15260
rect 21980 15314 22036 15326
rect 21980 15262 21982 15314
rect 22034 15262 22036 15314
rect 21420 14308 21476 14318
rect 21308 14252 21420 14308
rect 20748 14084 20804 14094
rect 20748 13970 20804 14028
rect 20748 13918 20750 13970
rect 20802 13918 20804 13970
rect 20748 13906 20804 13918
rect 20524 12910 20526 12962
rect 20578 12910 20580 12962
rect 19404 12850 19460 12862
rect 19404 12798 19406 12850
rect 19458 12798 19460 12850
rect 19404 11506 19460 12798
rect 19740 12850 19796 12862
rect 19740 12798 19742 12850
rect 19794 12798 19796 12850
rect 19516 12740 19572 12750
rect 19516 12646 19572 12684
rect 19740 12740 19796 12798
rect 19740 12674 19796 12684
rect 19964 12850 20020 12862
rect 19964 12798 19966 12850
rect 20018 12798 20020 12850
rect 19404 11454 19406 11506
rect 19458 11454 19460 11506
rect 19404 11442 19460 11454
rect 19516 11508 19572 11518
rect 19516 11394 19572 11452
rect 19964 11508 20020 12798
rect 20300 12740 20356 12750
rect 20300 11620 20356 12684
rect 20524 12404 20580 12910
rect 20524 12338 20580 12348
rect 21196 12404 21252 12414
rect 21196 12310 21252 12348
rect 20300 11554 20356 11564
rect 20860 12066 20916 12078
rect 20860 12014 20862 12066
rect 20914 12014 20916 12066
rect 19964 11442 20020 11452
rect 20636 11508 20692 11518
rect 20636 11414 20692 11452
rect 19516 11342 19518 11394
rect 19570 11342 19572 11394
rect 19516 11330 19572 11342
rect 20188 11394 20244 11406
rect 20188 11342 20190 11394
rect 20242 11342 20244 11394
rect 19292 11170 19348 11182
rect 19292 11118 19294 11170
rect 19346 11118 19348 11170
rect 19292 10836 19348 11118
rect 19292 10770 19348 10780
rect 19740 11170 19796 11182
rect 19740 11118 19742 11170
rect 19794 11118 19796 11170
rect 19740 9156 19796 11118
rect 20188 11172 20244 11342
rect 20188 11106 20244 11116
rect 20524 11170 20580 11182
rect 20524 11118 20526 11170
rect 20578 11118 20580 11170
rect 20524 10948 20580 11118
rect 20748 11172 20804 11182
rect 20748 11078 20804 11116
rect 20748 10948 20804 10958
rect 20860 10948 20916 12014
rect 20524 10892 20748 10948
rect 20804 10892 20916 10948
rect 20972 11620 21028 11630
rect 20748 10882 20804 10892
rect 20636 10724 20692 10734
rect 20860 10724 20916 10734
rect 20972 10724 21028 11564
rect 20692 10668 20804 10724
rect 20636 10658 20692 10668
rect 20524 10612 20580 10622
rect 20524 10518 20580 10556
rect 20636 10498 20692 10510
rect 20636 10446 20638 10498
rect 20690 10446 20692 10498
rect 20636 10276 20692 10446
rect 19740 9090 19796 9100
rect 20076 10220 20692 10276
rect 20076 9154 20132 10220
rect 20748 10164 20804 10668
rect 20860 10722 21028 10724
rect 20860 10670 20862 10722
rect 20914 10670 21028 10722
rect 20860 10668 21028 10670
rect 21084 10724 21140 10734
rect 20860 10658 20916 10668
rect 21084 10630 21140 10668
rect 20524 10108 20804 10164
rect 20300 9828 20356 9838
rect 20356 9772 20468 9828
rect 20300 9734 20356 9772
rect 20076 9102 20078 9154
rect 20130 9102 20132 9154
rect 20076 9090 20132 9102
rect 19292 9042 19348 9054
rect 19292 8990 19294 9042
rect 19346 8990 19348 9042
rect 19292 8372 19348 8990
rect 19292 8278 19348 8316
rect 20188 9044 20244 9054
rect 20188 7698 20244 8988
rect 20188 7646 20190 7698
rect 20242 7646 20244 7698
rect 20188 7634 20244 7646
rect 19180 7534 19182 7586
rect 19234 7534 19236 7586
rect 19180 7140 19236 7534
rect 19516 7588 19572 7598
rect 19516 7494 19572 7532
rect 19852 7588 19908 7598
rect 19852 7494 19908 7532
rect 20412 7588 20468 9772
rect 20524 9714 20580 10108
rect 20524 9662 20526 9714
rect 20578 9662 20580 9714
rect 20524 9650 20580 9662
rect 21308 8372 21364 14252
rect 21420 14214 21476 14252
rect 21980 14084 22036 15262
rect 22092 15204 22148 15932
rect 22316 15204 22372 15214
rect 22092 15202 22372 15204
rect 22092 15150 22318 15202
rect 22370 15150 22372 15202
rect 22092 15148 22372 15150
rect 22316 15138 22372 15148
rect 21980 14018 22036 14028
rect 22316 14196 22372 14206
rect 22316 13858 22372 14140
rect 22316 13806 22318 13858
rect 22370 13806 22372 13858
rect 22316 13794 22372 13806
rect 21868 13636 21924 13646
rect 21868 13542 21924 13580
rect 22428 13074 22484 16940
rect 22540 16884 22596 16894
rect 22540 16790 22596 16828
rect 22632 16492 22896 16502
rect 22688 16436 22736 16492
rect 22792 16436 22840 16492
rect 22632 16426 22896 16436
rect 22876 16212 22932 16222
rect 22988 16212 23044 17388
rect 23436 17220 23492 18398
rect 23660 18340 23716 18958
rect 24108 19012 24164 22988
rect 24668 22484 24724 23102
rect 24668 22418 24724 22428
rect 24780 21700 24836 21710
rect 24780 21606 24836 21644
rect 24220 21476 24276 21486
rect 24220 21382 24276 21420
rect 24444 20692 24500 20702
rect 24444 20130 24500 20636
rect 24444 20078 24446 20130
rect 24498 20078 24500 20130
rect 24444 20066 24500 20078
rect 24556 20020 24612 20030
rect 24556 20018 24724 20020
rect 24556 19966 24558 20018
rect 24610 19966 24724 20018
rect 24556 19964 24724 19966
rect 24556 19954 24612 19964
rect 24108 18918 24164 18956
rect 24668 18788 24724 19964
rect 24892 19460 24948 27580
rect 25340 26908 25396 30268
rect 25228 26852 25396 26908
rect 25228 24948 25284 26852
rect 25340 26292 25396 26302
rect 25340 26198 25396 26236
rect 25228 24882 25284 24892
rect 25452 24948 25508 30492
rect 25900 28754 25956 30828
rect 26236 30660 26292 30670
rect 26236 29650 26292 30604
rect 26236 29598 26238 29650
rect 26290 29598 26292 29650
rect 26236 29586 26292 29598
rect 25900 28702 25902 28754
rect 25954 28702 25956 28754
rect 25900 28690 25956 28702
rect 26236 28420 26292 28430
rect 25564 27972 25620 27982
rect 25564 27746 25620 27916
rect 26236 27860 26292 28364
rect 26236 27766 26292 27804
rect 25564 27694 25566 27746
rect 25618 27694 25620 27746
rect 25564 27682 25620 27694
rect 25788 27746 25844 27758
rect 25788 27694 25790 27746
rect 25842 27694 25844 27746
rect 25788 27300 25844 27694
rect 25564 27244 25844 27300
rect 25564 26740 25620 27244
rect 25900 27188 25956 27198
rect 25564 26674 25620 26684
rect 25676 27132 25900 27188
rect 25564 26516 25620 26526
rect 25564 26422 25620 26460
rect 25676 26402 25732 27132
rect 25900 27122 25956 27132
rect 26348 26908 26404 31388
rect 26572 28756 26628 28766
rect 26572 27188 26628 28700
rect 26572 27094 26628 27132
rect 26348 26852 26628 26908
rect 25676 26350 25678 26402
rect 25730 26350 25732 26402
rect 25676 26338 25732 26350
rect 26572 25732 26628 26852
rect 26684 26292 26740 32172
rect 27356 31892 27412 33068
rect 27580 33058 27636 33068
rect 28476 32900 28532 36200
rect 29596 33572 29652 36200
rect 30044 33572 30100 33582
rect 29596 33570 30100 33572
rect 29596 33518 30046 33570
rect 30098 33518 30100 33570
rect 29596 33516 30100 33518
rect 30044 33506 30100 33516
rect 30156 33460 30212 33470
rect 29036 33346 29092 33358
rect 29036 33294 29038 33346
rect 29090 33294 29092 33346
rect 28476 32834 28532 32844
rect 28700 33124 28756 33134
rect 29036 33124 29092 33294
rect 28700 33122 29092 33124
rect 28700 33070 28702 33122
rect 28754 33070 29092 33122
rect 28700 33068 29092 33070
rect 28588 32788 28644 32798
rect 27804 32564 27860 32574
rect 27356 31890 27748 31892
rect 27356 31838 27358 31890
rect 27410 31838 27748 31890
rect 27356 31836 27748 31838
rect 27356 31826 27412 31836
rect 26908 31780 26964 31790
rect 26908 31686 26964 31724
rect 26796 31554 26852 31566
rect 26796 31502 26798 31554
rect 26850 31502 26852 31554
rect 26796 26852 26852 31502
rect 26916 31388 27180 31398
rect 26972 31332 27020 31388
rect 27076 31332 27124 31388
rect 26916 31322 27180 31332
rect 27468 31108 27524 31118
rect 27468 30994 27524 31052
rect 27468 30942 27470 30994
rect 27522 30942 27524 30994
rect 27468 30930 27524 30942
rect 27692 30884 27748 31836
rect 27692 30322 27748 30828
rect 27692 30270 27694 30322
rect 27746 30270 27748 30322
rect 27692 30258 27748 30270
rect 27804 31778 27860 32508
rect 28476 32562 28532 32574
rect 28476 32510 28478 32562
rect 28530 32510 28532 32562
rect 28028 32452 28084 32462
rect 28028 31890 28084 32396
rect 28252 32340 28308 32350
rect 28028 31838 28030 31890
rect 28082 31838 28084 31890
rect 28028 31826 28084 31838
rect 28140 32284 28252 32340
rect 27804 31726 27806 31778
rect 27858 31726 27860 31778
rect 27804 30324 27860 31726
rect 28140 31666 28196 32284
rect 28252 32274 28308 32284
rect 28476 31892 28532 32510
rect 28140 31614 28142 31666
rect 28194 31614 28196 31666
rect 28140 31602 28196 31614
rect 28252 31668 28308 31678
rect 28252 31574 28308 31612
rect 27804 30258 27860 30268
rect 28028 31554 28084 31566
rect 28028 31502 28030 31554
rect 28082 31502 28084 31554
rect 28028 31220 28084 31502
rect 27132 29988 27188 29998
rect 27132 29986 27300 29988
rect 27132 29934 27134 29986
rect 27186 29934 27300 29986
rect 27132 29932 27300 29934
rect 27132 29922 27188 29932
rect 26916 29820 27180 29830
rect 26972 29764 27020 29820
rect 27076 29764 27124 29820
rect 26916 29754 27180 29764
rect 27132 29540 27188 29550
rect 27244 29540 27300 29932
rect 27188 29484 27300 29540
rect 27132 29474 27188 29484
rect 26916 28252 27180 28262
rect 26972 28196 27020 28252
rect 27076 28196 27124 28252
rect 26916 28186 27180 28196
rect 27356 28196 27412 28206
rect 27132 27746 27188 27758
rect 27132 27694 27134 27746
rect 27186 27694 27188 27746
rect 27132 27636 27188 27694
rect 27132 27570 27188 27580
rect 27020 26962 27076 26974
rect 27020 26910 27022 26962
rect 27074 26910 27076 26962
rect 27020 26908 27076 26910
rect 27020 26852 27300 26908
rect 26796 26786 26852 26796
rect 26916 26684 27180 26694
rect 26972 26628 27020 26684
rect 27076 26628 27124 26684
rect 26916 26618 27180 26628
rect 26684 26226 26740 26236
rect 26572 25676 26740 25732
rect 26460 25620 26516 25630
rect 26460 25526 26516 25564
rect 25452 24882 25508 24892
rect 26012 25284 26068 25294
rect 26012 24834 26068 25228
rect 26012 24782 26014 24834
rect 26066 24782 26068 24834
rect 26012 24770 26068 24782
rect 25228 24724 25284 24734
rect 25228 24630 25284 24668
rect 25564 24164 25620 24174
rect 25564 24050 25620 24108
rect 25564 23998 25566 24050
rect 25618 23998 25620 24050
rect 25564 23986 25620 23998
rect 26012 24052 26068 24062
rect 25452 23938 25508 23950
rect 25452 23886 25454 23938
rect 25506 23886 25508 23938
rect 25116 23826 25172 23838
rect 25116 23774 25118 23826
rect 25170 23774 25172 23826
rect 25116 23604 25172 23774
rect 25452 23716 25508 23886
rect 25452 23650 25508 23660
rect 25788 23716 25844 23726
rect 25788 23714 25956 23716
rect 25788 23662 25790 23714
rect 25842 23662 25956 23714
rect 25788 23660 25956 23662
rect 25788 23650 25844 23660
rect 25116 23538 25172 23548
rect 25452 23268 25508 23278
rect 25340 23266 25508 23268
rect 25340 23214 25454 23266
rect 25506 23214 25508 23266
rect 25340 23212 25508 23214
rect 25228 23044 25284 23054
rect 25340 23044 25396 23212
rect 25452 23202 25508 23212
rect 25284 22988 25396 23044
rect 25564 23154 25620 23166
rect 25564 23102 25566 23154
rect 25618 23102 25620 23154
rect 25228 22978 25284 22988
rect 25452 22930 25508 22942
rect 25452 22878 25454 22930
rect 25506 22878 25508 22930
rect 25228 22148 25284 22158
rect 25228 21810 25284 22092
rect 25228 21758 25230 21810
rect 25282 21758 25284 21810
rect 25228 21746 25284 21758
rect 25340 21812 25396 21822
rect 25340 21718 25396 21756
rect 25452 21810 25508 22878
rect 25564 22484 25620 23102
rect 25788 22484 25844 22494
rect 25564 22482 25844 22484
rect 25564 22430 25790 22482
rect 25842 22430 25844 22482
rect 25564 22428 25844 22430
rect 25788 22036 25844 22428
rect 25788 21970 25844 21980
rect 25452 21758 25454 21810
rect 25506 21758 25508 21810
rect 25452 21746 25508 21758
rect 25900 21586 25956 23660
rect 25900 21534 25902 21586
rect 25954 21534 25956 21586
rect 25900 21522 25956 21534
rect 26012 23714 26068 23996
rect 26012 23662 26014 23714
rect 26066 23662 26068 23714
rect 25788 21476 25844 21486
rect 25564 21474 25844 21476
rect 25564 21422 25790 21474
rect 25842 21422 25844 21474
rect 25564 21420 25844 21422
rect 25228 20916 25284 20926
rect 24892 19394 24948 19404
rect 25004 20132 25060 20142
rect 24780 19124 24836 19134
rect 24780 19030 24836 19068
rect 25004 18900 25060 20076
rect 25228 19572 25284 20860
rect 25564 20914 25620 21420
rect 25788 21410 25844 21420
rect 26012 21252 26068 23662
rect 26124 23826 26180 23838
rect 26124 23774 26126 23826
rect 26178 23774 26180 23826
rect 26124 23492 26180 23774
rect 26460 23716 26516 23754
rect 26460 23650 26516 23660
rect 26124 23426 26180 23436
rect 26460 23492 26516 23502
rect 26348 23380 26404 23390
rect 26348 23286 26404 23324
rect 26124 23154 26180 23166
rect 26124 23102 26126 23154
rect 26178 23102 26180 23154
rect 26124 22594 26180 23102
rect 26124 22542 26126 22594
rect 26178 22542 26180 22594
rect 26124 22530 26180 22542
rect 26236 23154 26292 23166
rect 26236 23102 26238 23154
rect 26290 23102 26292 23154
rect 26236 22372 26292 23102
rect 26124 22316 26292 22372
rect 26348 22594 26404 22606
rect 26348 22542 26350 22594
rect 26402 22542 26404 22594
rect 26124 21586 26180 22316
rect 26124 21534 26126 21586
rect 26178 21534 26180 21586
rect 26124 21522 26180 21534
rect 26236 22146 26292 22158
rect 26236 22094 26238 22146
rect 26290 22094 26292 22146
rect 25564 20862 25566 20914
rect 25618 20862 25620 20914
rect 25564 20850 25620 20862
rect 25900 21196 26068 21252
rect 26236 21476 26292 22094
rect 25900 20132 25956 21196
rect 26236 20804 26292 21420
rect 25900 20066 25956 20076
rect 26012 20802 26292 20804
rect 26012 20750 26238 20802
rect 26290 20750 26292 20802
rect 26012 20748 26292 20750
rect 25340 20020 25396 20030
rect 25340 20018 25508 20020
rect 25340 19966 25342 20018
rect 25394 19966 25508 20018
rect 25340 19964 25508 19966
rect 25340 19954 25396 19964
rect 25228 19236 25284 19516
rect 25340 19460 25396 19470
rect 25340 19366 25396 19404
rect 25228 19180 25396 19236
rect 24668 18722 24724 18732
rect 24780 18844 25060 18900
rect 25228 19012 25284 19022
rect 24556 18676 24612 18686
rect 23660 18274 23716 18284
rect 24220 18340 24276 18350
rect 23548 17892 23604 17902
rect 23548 17798 23604 17836
rect 23996 17666 24052 17678
rect 23996 17614 23998 17666
rect 24050 17614 24052 17666
rect 23996 17444 24052 17614
rect 23996 17378 24052 17388
rect 23100 17164 23604 17220
rect 23100 17106 23156 17164
rect 23100 17054 23102 17106
rect 23154 17054 23156 17106
rect 23100 17042 23156 17054
rect 23436 16884 23492 16894
rect 23436 16790 23492 16828
rect 22876 16210 23044 16212
rect 22876 16158 22878 16210
rect 22930 16158 23044 16210
rect 22876 16156 23044 16158
rect 22876 16146 22932 16156
rect 23436 15988 23492 15998
rect 23436 15894 23492 15932
rect 23100 15874 23156 15886
rect 23100 15822 23102 15874
rect 23154 15822 23156 15874
rect 22632 14924 22896 14934
rect 22688 14868 22736 14924
rect 22792 14868 22840 14924
rect 22632 14858 22896 14868
rect 23100 14084 23156 15822
rect 22764 14028 23156 14084
rect 23212 14530 23268 14542
rect 23212 14478 23214 14530
rect 23266 14478 23268 14530
rect 23212 14308 23268 14478
rect 22764 13746 22820 14028
rect 22764 13694 22766 13746
rect 22818 13694 22820 13746
rect 22764 13682 22820 13694
rect 23100 13858 23156 13870
rect 23100 13806 23102 13858
rect 23154 13806 23156 13858
rect 22632 13356 22896 13366
rect 22688 13300 22736 13356
rect 22792 13300 22840 13356
rect 23100 13300 23156 13806
rect 23212 13412 23268 14252
rect 23212 13346 23268 13356
rect 23324 13972 23380 13982
rect 22632 13290 22896 13300
rect 22988 13244 23100 13300
rect 22988 13188 23044 13244
rect 23100 13234 23156 13244
rect 22428 13022 22430 13074
rect 22482 13022 22484 13074
rect 22428 13010 22484 13022
rect 22764 13132 23044 13188
rect 23212 13188 23268 13198
rect 21868 12964 21924 12974
rect 21868 12962 22148 12964
rect 21868 12910 21870 12962
rect 21922 12910 22148 12962
rect 21868 12908 22148 12910
rect 21868 12898 21924 12908
rect 21756 12404 21812 12414
rect 21644 12348 21756 12404
rect 22092 12404 22148 12908
rect 22540 12962 22596 12974
rect 22540 12910 22542 12962
rect 22594 12910 22596 12962
rect 22316 12628 22372 12638
rect 22204 12404 22260 12414
rect 22092 12402 22260 12404
rect 22092 12350 22206 12402
rect 22258 12350 22260 12402
rect 22092 12348 22260 12350
rect 21644 11396 21700 12348
rect 21756 12338 21812 12348
rect 22204 12338 22260 12348
rect 22316 12290 22372 12572
rect 22540 12516 22596 12910
rect 22764 12850 22820 13132
rect 22988 12964 23044 12974
rect 22988 12870 23044 12908
rect 22764 12798 22766 12850
rect 22818 12798 22820 12850
rect 22764 12786 22820 12798
rect 23212 12850 23268 13132
rect 23324 12962 23380 13916
rect 23324 12910 23326 12962
rect 23378 12910 23380 12962
rect 23324 12898 23380 12910
rect 23212 12798 23214 12850
rect 23266 12798 23268 12850
rect 23212 12628 23268 12798
rect 23212 12562 23268 12572
rect 22540 12450 22596 12460
rect 22316 12238 22318 12290
rect 22370 12238 22372 12290
rect 22316 12226 22372 12238
rect 22652 12292 22708 12302
rect 22652 12290 22932 12292
rect 22652 12238 22654 12290
rect 22706 12238 22932 12290
rect 22652 12236 22932 12238
rect 22652 12226 22708 12236
rect 21756 12066 21812 12078
rect 22764 12068 22820 12078
rect 21756 12014 21758 12066
rect 21810 12014 21812 12066
rect 21756 11508 21812 12014
rect 22428 12066 22820 12068
rect 22428 12014 22766 12066
rect 22818 12014 22820 12066
rect 22428 12012 22820 12014
rect 21756 11452 21924 11508
rect 21644 11394 21812 11396
rect 21644 11342 21646 11394
rect 21698 11342 21812 11394
rect 21644 11340 21812 11342
rect 21644 11330 21700 11340
rect 21644 10948 21700 10958
rect 21420 10836 21476 10846
rect 21420 10052 21476 10780
rect 21644 10834 21700 10892
rect 21644 10782 21646 10834
rect 21698 10782 21700 10834
rect 21644 10770 21700 10782
rect 21532 10612 21588 10622
rect 21532 10518 21588 10556
rect 21420 9986 21476 9996
rect 21532 9156 21588 9166
rect 21588 9100 21700 9156
rect 21532 9090 21588 9100
rect 21532 8372 21588 8382
rect 21308 8370 21588 8372
rect 21308 8318 21534 8370
rect 21586 8318 21588 8370
rect 21308 8316 21588 8318
rect 21308 8260 21364 8316
rect 21532 8306 21588 8316
rect 21308 8194 21364 8204
rect 20748 8148 20804 8158
rect 20524 7700 20580 7710
rect 20580 7644 20692 7700
rect 20524 7634 20580 7644
rect 20412 7474 20468 7532
rect 20412 7422 20414 7474
rect 20466 7422 20468 7474
rect 20412 7410 20468 7422
rect 19180 7074 19236 7084
rect 20188 7364 20244 7374
rect 18844 6748 19348 6804
rect 17948 6638 17950 6690
rect 18002 6638 18004 6690
rect 17948 5122 18004 6638
rect 18732 6690 18788 6702
rect 18732 6638 18734 6690
rect 18786 6638 18788 6690
rect 18172 6580 18228 6590
rect 18284 6580 18340 6590
rect 18228 6578 18340 6580
rect 18228 6526 18286 6578
rect 18338 6526 18340 6578
rect 18228 6524 18340 6526
rect 17948 5070 17950 5122
rect 18002 5070 18004 5122
rect 17948 5012 18004 5070
rect 17948 4946 18004 4956
rect 18060 5796 18116 5806
rect 17612 4452 17668 4462
rect 17612 4338 17668 4396
rect 17612 4286 17614 4338
rect 17666 4286 17668 4338
rect 17612 4274 17668 4286
rect 17836 4004 17892 4508
rect 17948 4452 18004 4462
rect 18060 4452 18116 5740
rect 17948 4450 18116 4452
rect 17948 4398 17950 4450
rect 18002 4398 18116 4450
rect 17948 4396 18116 4398
rect 18172 4452 18228 6524
rect 18284 6514 18340 6524
rect 18620 6580 18676 6590
rect 18396 6468 18452 6506
rect 18620 6486 18676 6524
rect 18396 6402 18452 6412
rect 18348 6300 18612 6310
rect 18404 6244 18452 6300
rect 18508 6244 18556 6300
rect 18348 6234 18612 6244
rect 18732 6020 18788 6638
rect 19292 6692 19348 6748
rect 19180 6578 19236 6590
rect 19180 6526 19182 6578
rect 19234 6526 19236 6578
rect 18508 5964 18788 6020
rect 18956 6466 19012 6478
rect 18956 6414 18958 6466
rect 19010 6414 19012 6466
rect 18508 4900 18564 5964
rect 18956 5796 19012 6414
rect 18620 5740 19012 5796
rect 19068 5794 19124 5806
rect 19068 5742 19070 5794
rect 19122 5742 19124 5794
rect 18620 5234 18676 5740
rect 18620 5182 18622 5234
rect 18674 5182 18676 5234
rect 18620 5170 18676 5182
rect 19068 4900 19124 5742
rect 19180 5124 19236 6526
rect 19292 5796 19348 6636
rect 19628 6690 19684 6702
rect 19628 6638 19630 6690
rect 19682 6638 19684 6690
rect 19516 6580 19572 6590
rect 19628 6580 19684 6638
rect 19572 6524 19684 6580
rect 20076 6578 20132 6590
rect 20076 6526 20078 6578
rect 20130 6526 20132 6578
rect 19516 6514 19572 6524
rect 19292 5730 19348 5740
rect 19964 6466 20020 6478
rect 19964 6414 19966 6466
rect 20018 6414 20020 6466
rect 19180 5058 19236 5068
rect 18508 4844 18788 4900
rect 18348 4732 18612 4742
rect 18404 4676 18452 4732
rect 18508 4676 18556 4732
rect 18348 4666 18612 4676
rect 18620 4564 18676 4574
rect 18732 4564 18788 4844
rect 19068 4834 19124 4844
rect 19292 5012 19348 5022
rect 18620 4562 18788 4564
rect 18620 4510 18622 4562
rect 18674 4510 18788 4562
rect 18620 4508 18788 4510
rect 18956 4564 19012 4574
rect 18620 4498 18676 4508
rect 18956 4470 19012 4508
rect 18284 4452 18340 4462
rect 18172 4450 18340 4452
rect 18172 4398 18286 4450
rect 18338 4398 18340 4450
rect 18172 4396 18340 4398
rect 17948 4386 18004 4396
rect 18284 4386 18340 4396
rect 18396 4450 18452 4462
rect 18396 4398 18398 4450
rect 18450 4398 18452 4450
rect 17836 3938 17892 3948
rect 18396 4228 18452 4398
rect 19292 4338 19348 4956
rect 19964 4452 20020 6414
rect 20076 5012 20132 6526
rect 20188 6130 20244 7308
rect 20300 6692 20356 6702
rect 20300 6598 20356 6636
rect 20188 6078 20190 6130
rect 20242 6078 20244 6130
rect 20188 6066 20244 6078
rect 20412 6020 20468 6030
rect 20412 5926 20468 5964
rect 20524 6020 20580 6030
rect 20636 6020 20692 7644
rect 20748 7698 20804 8092
rect 20748 7646 20750 7698
rect 20802 7646 20804 7698
rect 20748 7634 20804 7646
rect 21084 7700 21140 7710
rect 20972 7588 21028 7598
rect 20972 7494 21028 7532
rect 21084 7588 21140 7644
rect 21420 7588 21476 7598
rect 21084 7586 21476 7588
rect 21084 7534 21086 7586
rect 21138 7534 21422 7586
rect 21474 7534 21476 7586
rect 21084 7532 21476 7534
rect 21084 7522 21140 7532
rect 21420 7522 21476 7532
rect 21532 7588 21588 7598
rect 21532 7494 21588 7532
rect 21532 7252 21588 7262
rect 21644 7252 21700 9100
rect 21532 7250 21700 7252
rect 21532 7198 21534 7250
rect 21586 7198 21700 7250
rect 21532 7196 21700 7198
rect 21532 7186 21588 7196
rect 20860 7140 20916 7150
rect 20860 6690 20916 7084
rect 20860 6638 20862 6690
rect 20914 6638 20916 6690
rect 20860 6626 20916 6638
rect 21308 6692 21364 6702
rect 21308 6598 21364 6636
rect 21756 6692 21812 11340
rect 21868 11172 21924 11452
rect 22428 11506 22484 12012
rect 22764 12002 22820 12012
rect 22876 11956 22932 12236
rect 22988 12180 23044 12190
rect 22988 12178 23156 12180
rect 22988 12126 22990 12178
rect 23042 12126 23156 12178
rect 22988 12124 23156 12126
rect 22988 12114 23044 12124
rect 22876 11900 23044 11956
rect 22632 11788 22896 11798
rect 22688 11732 22736 11788
rect 22792 11732 22840 11788
rect 22632 11722 22896 11732
rect 22428 11454 22430 11506
rect 22482 11454 22484 11506
rect 22428 11442 22484 11454
rect 21868 11060 21924 11116
rect 22764 11284 22820 11294
rect 22316 11060 22372 11070
rect 21868 11004 22316 11060
rect 22316 10834 22372 11004
rect 22316 10782 22318 10834
rect 22370 10782 22372 10834
rect 22316 10770 22372 10782
rect 22764 10836 22820 11228
rect 22764 10742 22820 10780
rect 22428 10724 22484 10734
rect 22428 10630 22484 10668
rect 22092 10610 22148 10622
rect 22092 10558 22094 10610
rect 22146 10558 22148 10610
rect 22092 9714 22148 10558
rect 22540 10610 22596 10622
rect 22540 10558 22542 10610
rect 22594 10558 22596 10610
rect 22540 10388 22596 10558
rect 22428 10332 22596 10388
rect 22428 9828 22484 10332
rect 22632 10220 22896 10230
rect 22688 10164 22736 10220
rect 22792 10164 22840 10220
rect 22632 10154 22896 10164
rect 22092 9662 22094 9714
rect 22146 9662 22148 9714
rect 22092 9650 22148 9662
rect 22204 9772 22484 9828
rect 22204 8930 22260 9772
rect 22316 9602 22372 9614
rect 22316 9550 22318 9602
rect 22370 9550 22372 9602
rect 22316 9268 22372 9550
rect 22428 9604 22484 9772
rect 22540 10052 22596 10062
rect 22988 10052 23044 11900
rect 23100 11620 23156 12124
rect 23100 11554 23156 11564
rect 23212 12178 23268 12190
rect 23212 12126 23214 12178
rect 23266 12126 23268 12178
rect 23212 11284 23268 12126
rect 23212 11218 23268 11228
rect 23324 10836 23380 10846
rect 23324 10742 23380 10780
rect 23548 10836 23604 17164
rect 24220 16994 24276 18284
rect 24556 17778 24612 18620
rect 24780 17890 24836 18844
rect 25116 18338 25172 18350
rect 25116 18286 25118 18338
rect 25170 18286 25172 18338
rect 25116 18228 25172 18286
rect 24780 17838 24782 17890
rect 24834 17838 24836 17890
rect 24780 17826 24836 17838
rect 24892 18172 25172 18228
rect 25228 18228 25284 18956
rect 25340 18564 25396 19180
rect 25452 19012 25508 19964
rect 25564 20018 25620 20030
rect 25564 19966 25566 20018
rect 25618 19966 25620 20018
rect 25564 19796 25620 19966
rect 25788 20018 25844 20030
rect 25788 19966 25790 20018
rect 25842 19966 25844 20018
rect 25564 19730 25620 19740
rect 25676 19906 25732 19918
rect 25676 19854 25678 19906
rect 25730 19854 25732 19906
rect 25564 19234 25620 19246
rect 25564 19182 25566 19234
rect 25618 19182 25620 19234
rect 25564 19124 25620 19182
rect 25676 19236 25732 19854
rect 25788 19908 25844 19966
rect 25788 19842 25844 19852
rect 26012 19796 26068 20748
rect 26236 20738 26292 20748
rect 26348 21364 26404 22542
rect 26460 22148 26516 23436
rect 26460 22054 26516 22092
rect 26572 23266 26628 23278
rect 26572 23214 26574 23266
rect 26626 23214 26628 23266
rect 26460 21364 26516 21374
rect 26348 21362 26516 21364
rect 26348 21310 26462 21362
rect 26514 21310 26516 21362
rect 26348 21308 26516 21310
rect 26348 20580 26404 21308
rect 26460 21298 26516 21308
rect 26124 20524 26404 20580
rect 26124 20130 26180 20524
rect 26124 20078 26126 20130
rect 26178 20078 26180 20130
rect 26124 20066 26180 20078
rect 26236 20132 26292 20142
rect 26236 20038 26292 20076
rect 26460 20132 26516 20142
rect 26572 20132 26628 23214
rect 26684 23044 26740 25676
rect 27132 25508 27188 25518
rect 27132 25414 27188 25452
rect 26916 25116 27180 25126
rect 26972 25060 27020 25116
rect 27076 25060 27124 25116
rect 26916 25050 27180 25060
rect 26796 24388 26852 24398
rect 26796 23826 26852 24332
rect 27132 24276 27188 24286
rect 27132 23938 27188 24220
rect 27132 23886 27134 23938
rect 27186 23886 27188 23938
rect 27132 23874 27188 23886
rect 26796 23774 26798 23826
rect 26850 23774 26852 23826
rect 26796 23762 26852 23774
rect 26916 23548 27180 23558
rect 26972 23492 27020 23548
rect 27076 23492 27124 23548
rect 26916 23482 27180 23492
rect 27132 23268 27188 23278
rect 26684 22978 26740 22988
rect 27020 23154 27076 23166
rect 27020 23102 27022 23154
rect 27074 23102 27076 23154
rect 27020 22932 27076 23102
rect 27020 22260 27076 22876
rect 26684 22204 27076 22260
rect 27132 22370 27188 23212
rect 27132 22318 27134 22370
rect 27186 22318 27188 22370
rect 26684 21700 26740 22204
rect 27132 22148 27188 22318
rect 27244 22372 27300 26852
rect 27356 25394 27412 28140
rect 27804 27636 27860 27646
rect 27468 27186 27524 27198
rect 27468 27134 27470 27186
rect 27522 27134 27524 27186
rect 27468 25732 27524 27134
rect 27580 26516 27636 26526
rect 27580 26422 27636 26460
rect 27804 25732 27860 27580
rect 28028 27186 28084 31164
rect 28476 31108 28532 31836
rect 28476 31042 28532 31052
rect 28028 27134 28030 27186
rect 28082 27134 28084 27186
rect 28028 26908 28084 27134
rect 27916 26852 28084 26908
rect 28140 30882 28196 30894
rect 28140 30830 28142 30882
rect 28194 30830 28196 30882
rect 28140 26908 28196 30830
rect 28588 30436 28644 32732
rect 28476 30380 28644 30436
rect 28476 29988 28532 30380
rect 28588 30212 28644 30222
rect 28588 30118 28644 30156
rect 28476 29932 28644 29988
rect 28476 29652 28532 29662
rect 28476 28756 28532 29596
rect 28476 28662 28532 28700
rect 28364 28420 28420 28430
rect 28364 28326 28420 28364
rect 28364 27074 28420 27086
rect 28364 27022 28366 27074
rect 28418 27022 28420 27074
rect 28140 26852 28308 26908
rect 27916 26068 27972 26852
rect 28140 26292 28196 26302
rect 28140 26198 28196 26236
rect 27916 26002 27972 26012
rect 28028 25732 28084 25742
rect 27804 25676 27972 25732
rect 27468 25666 27524 25676
rect 27356 25342 27358 25394
rect 27410 25342 27412 25394
rect 27356 25330 27412 25342
rect 27692 25508 27748 25518
rect 27468 24612 27524 24622
rect 27468 23826 27524 24556
rect 27468 23774 27470 23826
rect 27522 23774 27524 23826
rect 27468 23762 27524 23774
rect 27580 23716 27636 23726
rect 27356 23380 27412 23390
rect 27356 23286 27412 23324
rect 27244 22306 27300 22316
rect 27468 22370 27524 22382
rect 27468 22318 27470 22370
rect 27522 22318 27524 22370
rect 26684 21634 26740 21644
rect 26796 22092 27188 22148
rect 26796 21588 26852 22092
rect 26916 21980 27180 21990
rect 26972 21924 27020 21980
rect 27076 21924 27124 21980
rect 26916 21914 27180 21924
rect 27468 21812 27524 22318
rect 27244 21756 27468 21812
rect 27020 21588 27076 21598
rect 27244 21588 27300 21756
rect 27468 21746 27524 21756
rect 26796 21586 27076 21588
rect 26796 21534 27022 21586
rect 27074 21534 27076 21586
rect 26796 21532 27076 21534
rect 26684 21476 26740 21486
rect 26684 20580 26740 21420
rect 26796 20804 26852 21532
rect 27020 21476 27076 21532
rect 27020 21410 27076 21420
rect 27132 21586 27300 21588
rect 27132 21534 27246 21586
rect 27298 21534 27300 21586
rect 27132 21532 27300 21534
rect 27132 20916 27188 21532
rect 27244 21522 27300 21532
rect 27468 21588 27524 21598
rect 27468 21494 27524 21532
rect 27580 21028 27636 23660
rect 27692 22596 27748 25452
rect 27804 25506 27860 25518
rect 27804 25454 27806 25506
rect 27858 25454 27860 25506
rect 27804 24388 27860 25454
rect 27804 24322 27860 24332
rect 27804 23828 27860 23838
rect 27804 22932 27860 23772
rect 27916 23604 27972 25676
rect 28028 25638 28084 25676
rect 28252 25618 28308 26852
rect 28252 25566 28254 25618
rect 28306 25566 28308 25618
rect 28252 25554 28308 25566
rect 28364 25394 28420 27022
rect 28588 26908 28644 29932
rect 28700 28532 28756 33068
rect 29148 32452 29204 32462
rect 29148 32358 29204 32396
rect 29260 31892 29316 31902
rect 29260 31778 29316 31836
rect 29260 31726 29262 31778
rect 29314 31726 29316 31778
rect 29260 31714 29316 31726
rect 29708 31892 29764 31902
rect 29260 31220 29316 31230
rect 29148 30996 29204 31006
rect 28924 29316 28980 29326
rect 28700 28466 28756 28476
rect 28812 29204 28868 29214
rect 28812 28084 28868 29148
rect 28924 28644 28980 29260
rect 29148 29204 29204 30940
rect 29260 30212 29316 31164
rect 29708 30212 29764 31836
rect 29932 31666 29988 31678
rect 29932 31614 29934 31666
rect 29986 31614 29988 31666
rect 29932 30884 29988 31614
rect 29932 30818 29988 30828
rect 29260 30118 29316 30156
rect 29372 30210 29876 30212
rect 29372 30158 29710 30210
rect 29762 30158 29876 30210
rect 29372 30156 29876 30158
rect 29260 29428 29316 29438
rect 29372 29428 29428 30156
rect 29708 30146 29764 30156
rect 29260 29426 29428 29428
rect 29260 29374 29262 29426
rect 29314 29374 29428 29426
rect 29260 29372 29428 29374
rect 29260 29362 29316 29372
rect 29148 29148 29428 29204
rect 29148 28644 29204 28654
rect 28924 28642 29204 28644
rect 28924 28590 29150 28642
rect 29202 28590 29204 28642
rect 28924 28588 29204 28590
rect 29148 28578 29204 28588
rect 29260 28084 29316 28094
rect 28812 28028 28980 28084
rect 28588 26852 28868 26908
rect 28812 26516 28868 26852
rect 28812 26450 28868 26460
rect 28364 25342 28366 25394
rect 28418 25342 28420 25394
rect 28364 24836 28420 25342
rect 28140 24610 28196 24622
rect 28140 24558 28142 24610
rect 28194 24558 28196 24610
rect 28140 23826 28196 24558
rect 28364 24276 28420 24780
rect 28364 24210 28420 24220
rect 28476 25396 28532 25406
rect 28476 24050 28532 25340
rect 28588 25396 28644 25406
rect 28588 25394 28756 25396
rect 28588 25342 28590 25394
rect 28642 25342 28756 25394
rect 28588 25340 28756 25342
rect 28588 25330 28644 25340
rect 28476 23998 28478 24050
rect 28530 23998 28532 24050
rect 28476 23986 28532 23998
rect 28588 24164 28644 24174
rect 28588 23938 28644 24108
rect 28588 23886 28590 23938
rect 28642 23886 28644 23938
rect 28588 23874 28644 23886
rect 28140 23774 28142 23826
rect 28194 23774 28196 23826
rect 28028 23604 28084 23614
rect 27916 23548 28028 23604
rect 28028 23538 28084 23548
rect 27804 22866 27860 22876
rect 28028 23266 28084 23278
rect 28028 23214 28030 23266
rect 28082 23214 28084 23266
rect 28028 22820 28084 23214
rect 28028 22754 28084 22764
rect 27692 22540 28084 22596
rect 27692 22372 27748 22382
rect 27916 22372 27972 22382
rect 27692 22370 27916 22372
rect 27692 22318 27694 22370
rect 27746 22318 27916 22370
rect 27692 22316 27916 22318
rect 27692 22306 27748 22316
rect 27580 20962 27636 20972
rect 26796 20738 26852 20748
rect 26908 20860 27188 20916
rect 27244 20916 27300 20926
rect 27244 20914 27524 20916
rect 27244 20862 27246 20914
rect 27298 20862 27524 20914
rect 27244 20860 27524 20862
rect 26908 20802 26964 20860
rect 27244 20850 27300 20860
rect 26908 20750 26910 20802
rect 26962 20750 26964 20802
rect 26908 20738 26964 20750
rect 27468 20804 27524 20860
rect 27804 20804 27860 20814
rect 27468 20802 27860 20804
rect 27468 20750 27806 20802
rect 27858 20750 27860 20802
rect 27468 20748 27860 20750
rect 27804 20738 27860 20748
rect 27020 20690 27076 20702
rect 27020 20638 27022 20690
rect 27074 20638 27076 20690
rect 27020 20580 27076 20638
rect 27356 20692 27412 20702
rect 27356 20598 27412 20636
rect 26684 20524 27076 20580
rect 27580 20580 27636 20590
rect 27580 20486 27636 20524
rect 26916 20412 27180 20422
rect 26972 20356 27020 20412
rect 27076 20356 27124 20412
rect 26916 20346 27180 20356
rect 26460 20130 26628 20132
rect 26460 20078 26462 20130
rect 26514 20078 26628 20130
rect 26460 20076 26628 20078
rect 27132 20244 27188 20254
rect 27804 20244 27860 20254
rect 27132 20130 27188 20188
rect 27468 20188 27804 20244
rect 27132 20078 27134 20130
rect 27186 20078 27188 20130
rect 26460 20066 26516 20076
rect 27132 20066 27188 20078
rect 27356 20130 27412 20142
rect 27356 20078 27358 20130
rect 27410 20078 27412 20130
rect 26796 20018 26852 20030
rect 26796 19966 26798 20018
rect 26850 19966 26852 20018
rect 25900 19740 26068 19796
rect 26572 19908 26628 19918
rect 25788 19684 25844 19694
rect 25788 19458 25844 19628
rect 25788 19406 25790 19458
rect 25842 19406 25844 19458
rect 25788 19394 25844 19406
rect 25676 19180 25844 19236
rect 25564 19068 25732 19124
rect 25452 18956 25620 19012
rect 25452 18564 25508 18574
rect 25340 18562 25508 18564
rect 25340 18510 25454 18562
rect 25506 18510 25508 18562
rect 25340 18508 25508 18510
rect 25340 18452 25396 18508
rect 25452 18498 25508 18508
rect 25340 18386 25396 18396
rect 25564 18452 25620 18956
rect 25564 18386 25620 18396
rect 24556 17726 24558 17778
rect 24610 17726 24612 17778
rect 24556 17714 24612 17726
rect 24332 17668 24388 17678
rect 24332 17574 24388 17612
rect 24220 16942 24222 16994
rect 24274 16942 24276 16994
rect 24220 16930 24276 16942
rect 24444 17108 24500 17118
rect 23884 16100 23940 16110
rect 24220 16100 24276 16110
rect 23884 16006 23940 16044
rect 24108 16044 24220 16100
rect 24108 14756 24164 16044
rect 24220 16006 24276 16044
rect 24444 16098 24500 17052
rect 24444 16046 24446 16098
rect 24498 16046 24500 16098
rect 24444 15428 24500 16046
rect 24444 15362 24500 15372
rect 24556 15988 24612 15998
rect 24108 14690 24164 14700
rect 24220 15314 24276 15326
rect 24220 15262 24222 15314
rect 24274 15262 24276 15314
rect 23996 14420 24052 14430
rect 23996 13300 24052 14364
rect 23996 12852 24052 13244
rect 24220 12962 24276 15262
rect 24556 15202 24612 15932
rect 24668 15986 24724 15998
rect 24668 15934 24670 15986
rect 24722 15934 24724 15986
rect 24668 15876 24724 15934
rect 24668 15810 24724 15820
rect 24556 15150 24558 15202
rect 24610 15150 24612 15202
rect 24556 15148 24612 15150
rect 24892 15148 24948 18172
rect 25228 18162 25284 18172
rect 25340 18004 25396 18014
rect 25116 17890 25172 17902
rect 25116 17838 25118 17890
rect 25170 17838 25172 17890
rect 25004 17556 25060 17566
rect 25004 16324 25060 17500
rect 25116 17442 25172 17838
rect 25116 17390 25118 17442
rect 25170 17390 25172 17442
rect 25116 16548 25172 17390
rect 25228 16996 25284 17006
rect 25340 16996 25396 17948
rect 25452 17666 25508 17678
rect 25452 17614 25454 17666
rect 25506 17614 25508 17666
rect 25452 17444 25508 17614
rect 25676 17668 25732 19068
rect 25452 17378 25508 17388
rect 25564 17442 25620 17454
rect 25564 17390 25566 17442
rect 25618 17390 25620 17442
rect 25452 16996 25508 17006
rect 25340 16994 25508 16996
rect 25340 16942 25454 16994
rect 25506 16942 25508 16994
rect 25340 16940 25508 16942
rect 25228 16882 25284 16940
rect 25452 16930 25508 16940
rect 25228 16830 25230 16882
rect 25282 16830 25284 16882
rect 25228 16818 25284 16830
rect 25116 16492 25284 16548
rect 25116 16324 25172 16334
rect 25004 16322 25172 16324
rect 25004 16270 25118 16322
rect 25170 16270 25172 16322
rect 25004 16268 25172 16270
rect 25116 16258 25172 16268
rect 25228 16100 25284 16492
rect 24556 15092 24724 15148
rect 24668 14644 24724 15092
rect 24556 13748 24612 13758
rect 24332 13746 24612 13748
rect 24332 13694 24558 13746
rect 24610 13694 24612 13746
rect 24332 13692 24612 13694
rect 24332 13076 24388 13692
rect 24556 13682 24612 13692
rect 24668 13524 24724 14588
rect 24332 12982 24388 13020
rect 24556 13468 24724 13524
rect 24780 15092 24948 15148
rect 25116 16044 25284 16100
rect 25340 16436 25396 16446
rect 25116 15092 25172 16044
rect 24220 12910 24222 12962
rect 24274 12910 24276 12962
rect 23996 12850 24164 12852
rect 23996 12798 23998 12850
rect 24050 12798 24164 12850
rect 23996 12796 24164 12798
rect 23996 12786 24052 12796
rect 23660 12404 23716 12414
rect 23660 12310 23716 12348
rect 24108 12290 24164 12796
rect 24220 12516 24276 12910
rect 24220 12450 24276 12460
rect 24108 12238 24110 12290
rect 24162 12238 24164 12290
rect 24108 12226 24164 12238
rect 24556 12178 24612 13468
rect 24668 13188 24724 13198
rect 24668 13074 24724 13132
rect 24668 13022 24670 13074
rect 24722 13022 24724 13074
rect 24668 13010 24724 13022
rect 24556 12126 24558 12178
rect 24610 12126 24612 12178
rect 24556 12114 24612 12126
rect 24668 12180 24724 12190
rect 24668 12066 24724 12124
rect 24668 12014 24670 12066
rect 24722 12014 24724 12066
rect 24668 12002 24724 12014
rect 24556 11508 24612 11518
rect 24332 11506 24612 11508
rect 24332 11454 24558 11506
rect 24610 11454 24612 11506
rect 24332 11452 24612 11454
rect 23548 10770 23604 10780
rect 23660 11284 23716 11294
rect 23660 10834 23716 11228
rect 23660 10782 23662 10834
rect 23714 10782 23716 10834
rect 23660 10770 23716 10782
rect 23772 11060 23828 11070
rect 23772 10834 23828 11004
rect 24332 10836 24388 11452
rect 24556 11442 24612 11452
rect 24780 10836 24836 15092
rect 25116 15026 25172 15036
rect 25228 15204 25284 15214
rect 25228 15090 25284 15148
rect 25228 15038 25230 15090
rect 25282 15038 25284 15090
rect 25228 15026 25284 15038
rect 25340 14642 25396 16380
rect 25452 16100 25508 16110
rect 25452 16006 25508 16044
rect 25340 14590 25342 14642
rect 25394 14590 25396 14642
rect 25228 13972 25284 13982
rect 25228 13878 25284 13916
rect 25340 12404 25396 14590
rect 25452 15204 25508 15214
rect 25452 13748 25508 15148
rect 25564 13972 25620 17390
rect 25676 17106 25732 17612
rect 25676 17054 25678 17106
rect 25730 17054 25732 17106
rect 25676 17042 25732 17054
rect 25788 16996 25844 19180
rect 25788 16930 25844 16940
rect 25788 16772 25844 16782
rect 25676 15986 25732 15998
rect 25676 15934 25678 15986
rect 25730 15934 25732 15986
rect 25676 15876 25732 15934
rect 25676 15810 25732 15820
rect 25788 15426 25844 16716
rect 25900 16436 25956 19740
rect 26012 19572 26068 19582
rect 26012 19234 26068 19516
rect 26012 19182 26014 19234
rect 26066 19182 26068 19234
rect 26012 19170 26068 19182
rect 26348 19124 26404 19134
rect 26124 19122 26404 19124
rect 26124 19070 26350 19122
rect 26402 19070 26404 19122
rect 26124 19068 26404 19070
rect 26012 18900 26068 18910
rect 26012 18564 26068 18844
rect 26012 18470 26068 18508
rect 26124 18452 26180 19068
rect 26348 19058 26404 19068
rect 26572 19124 26628 19852
rect 26684 19796 26740 19806
rect 26684 19702 26740 19740
rect 26796 19684 26852 19966
rect 27356 20020 27412 20078
rect 27356 19954 27412 19964
rect 27468 19906 27524 20188
rect 27804 20178 27860 20188
rect 27468 19854 27470 19906
rect 27522 19854 27524 19906
rect 27468 19842 27524 19854
rect 27916 19906 27972 22316
rect 27916 19854 27918 19906
rect 27970 19854 27972 19906
rect 27916 19842 27972 19854
rect 26796 19618 26852 19628
rect 27580 19460 27636 19470
rect 27020 19348 27076 19358
rect 27020 19254 27076 19292
rect 27580 19234 27636 19404
rect 28028 19460 28084 22540
rect 28140 22370 28196 23774
rect 28252 23826 28308 23838
rect 28252 23774 28254 23826
rect 28306 23774 28308 23826
rect 28252 23716 28308 23774
rect 28252 23650 28308 23660
rect 28364 23714 28420 23726
rect 28364 23662 28366 23714
rect 28418 23662 28420 23714
rect 28364 23492 28420 23662
rect 28364 23426 28420 23436
rect 28588 23604 28644 23614
rect 28700 23604 28756 25340
rect 28812 24498 28868 24510
rect 28812 24446 28814 24498
rect 28866 24446 28868 24498
rect 28812 24276 28868 24446
rect 28812 24210 28868 24220
rect 28924 23716 28980 28028
rect 29260 27970 29316 28028
rect 29260 27918 29262 27970
rect 29314 27918 29316 27970
rect 29260 27906 29316 27918
rect 29148 27074 29204 27086
rect 29148 27022 29150 27074
rect 29202 27022 29204 27074
rect 29148 25620 29204 27022
rect 29372 26908 29428 29148
rect 29820 27860 29876 30156
rect 29932 29316 29988 29326
rect 29932 29314 30100 29316
rect 29932 29262 29934 29314
rect 29986 29262 30100 29314
rect 29932 29260 30100 29262
rect 29932 29250 29988 29260
rect 29932 27860 29988 27870
rect 29820 27858 29988 27860
rect 29820 27806 29934 27858
rect 29986 27806 29988 27858
rect 29820 27804 29988 27806
rect 29932 27794 29988 27804
rect 30044 27636 30100 29260
rect 29148 25554 29204 25564
rect 29260 26852 29428 26908
rect 29820 27580 30100 27636
rect 29036 24724 29092 24734
rect 29036 24630 29092 24668
rect 29260 24388 29316 26852
rect 29596 25732 29652 25742
rect 29596 25638 29652 25676
rect 29484 25508 29540 25518
rect 29484 25414 29540 25452
rect 29372 25282 29428 25294
rect 29820 25284 29876 27580
rect 30044 27412 30100 27422
rect 29932 27188 29988 27198
rect 29932 26402 29988 27132
rect 29932 26350 29934 26402
rect 29986 26350 29988 26402
rect 29932 26338 29988 26350
rect 29372 25230 29374 25282
rect 29426 25230 29428 25282
rect 29372 25060 29428 25230
rect 29372 24994 29428 25004
rect 29484 25228 29876 25284
rect 29932 25508 29988 25518
rect 30044 25508 30100 27356
rect 30156 26908 30212 33404
rect 30380 32900 30436 32910
rect 30436 32844 30548 32900
rect 30380 32834 30436 32844
rect 30268 30882 30324 30894
rect 30268 30830 30270 30882
rect 30322 30830 30324 30882
rect 30268 28420 30324 30830
rect 30380 30772 30436 30782
rect 30492 30772 30548 32844
rect 30604 30996 30660 31006
rect 30604 30902 30660 30940
rect 30492 30716 30660 30772
rect 30380 30210 30436 30716
rect 30380 30158 30382 30210
rect 30434 30158 30436 30210
rect 30380 30146 30436 30158
rect 30268 27524 30324 28364
rect 30380 28084 30436 28094
rect 30380 27990 30436 28028
rect 30492 27860 30548 27870
rect 30492 27766 30548 27804
rect 30268 27458 30324 27468
rect 30604 27298 30660 30716
rect 30716 29764 30772 36200
rect 30828 31220 30884 31230
rect 30828 31126 30884 31164
rect 30828 30884 30884 30894
rect 30828 30790 30884 30828
rect 30716 29708 30884 29764
rect 30604 27246 30606 27298
rect 30658 27246 30660 27298
rect 30604 27234 30660 27246
rect 30716 27972 30772 27982
rect 30716 27634 30772 27916
rect 30716 27582 30718 27634
rect 30770 27582 30772 27634
rect 30156 26852 30324 26908
rect 29932 25506 30100 25508
rect 29932 25454 29934 25506
rect 29986 25454 30100 25506
rect 29932 25452 30100 25454
rect 29372 24836 29428 24846
rect 29372 24742 29428 24780
rect 29372 24612 29428 24622
rect 29484 24612 29540 25228
rect 29932 25172 29988 25452
rect 29372 24610 29540 24612
rect 29372 24558 29374 24610
rect 29426 24558 29540 24610
rect 29372 24556 29540 24558
rect 29708 25116 29988 25172
rect 29372 24546 29428 24556
rect 29596 24500 29652 24510
rect 29596 24406 29652 24444
rect 29260 24332 29540 24388
rect 29372 23938 29428 23950
rect 29372 23886 29374 23938
rect 29426 23886 29428 23938
rect 29260 23716 29316 23726
rect 28924 23660 29204 23716
rect 28700 23548 28980 23604
rect 28252 23268 28308 23278
rect 28252 23174 28308 23212
rect 28476 23268 28532 23278
rect 28588 23268 28644 23548
rect 28924 23378 28980 23548
rect 28924 23326 28926 23378
rect 28978 23326 28980 23378
rect 28924 23314 28980 23326
rect 29036 23492 29092 23502
rect 28476 23266 28644 23268
rect 28476 23214 28478 23266
rect 28530 23214 28644 23266
rect 28476 23212 28644 23214
rect 29036 23266 29092 23436
rect 29036 23214 29038 23266
rect 29090 23214 29092 23266
rect 28476 23202 28532 23212
rect 28812 23154 28868 23166
rect 28812 23102 28814 23154
rect 28866 23102 28868 23154
rect 28364 22932 28420 22942
rect 28140 22318 28142 22370
rect 28194 22318 28196 22370
rect 28140 22306 28196 22318
rect 28252 22930 28420 22932
rect 28252 22878 28366 22930
rect 28418 22878 28420 22930
rect 28252 22876 28420 22878
rect 28252 21812 28308 22876
rect 28364 22866 28420 22876
rect 28812 22932 28868 23102
rect 28812 22866 28868 22876
rect 28924 23156 28980 23166
rect 28364 22148 28420 22158
rect 28364 22146 28532 22148
rect 28364 22094 28366 22146
rect 28418 22094 28532 22146
rect 28364 22092 28532 22094
rect 28364 22082 28420 22092
rect 28252 21756 28420 21812
rect 28252 20804 28308 20814
rect 28252 20710 28308 20748
rect 28364 20802 28420 21756
rect 28364 20750 28366 20802
rect 28418 20750 28420 20802
rect 28364 20738 28420 20750
rect 28476 20580 28532 22092
rect 28588 22146 28644 22158
rect 28588 22094 28590 22146
rect 28642 22094 28644 22146
rect 28588 22036 28644 22094
rect 28588 21970 28644 21980
rect 28700 22146 28756 22158
rect 28700 22094 28702 22146
rect 28754 22094 28756 22146
rect 28588 20916 28644 20926
rect 28700 20916 28756 22094
rect 28588 20914 28756 20916
rect 28588 20862 28590 20914
rect 28642 20862 28756 20914
rect 28588 20860 28756 20862
rect 28812 21698 28868 21710
rect 28812 21646 28814 21698
rect 28866 21646 28868 21698
rect 28812 21252 28868 21646
rect 28588 20850 28644 20860
rect 28588 20692 28644 20702
rect 28812 20692 28868 21196
rect 28644 20636 28756 20692
rect 28588 20626 28644 20636
rect 28364 20524 28532 20580
rect 28364 19796 28420 20524
rect 28588 20244 28644 20254
rect 28364 19730 28420 19740
rect 28476 20188 28588 20244
rect 28028 19394 28084 19404
rect 27580 19182 27582 19234
rect 27634 19182 27636 19234
rect 27580 19170 27636 19182
rect 28364 19348 28420 19358
rect 26572 19030 26628 19068
rect 26460 19010 26516 19022
rect 26460 18958 26462 19010
rect 26514 18958 26516 19010
rect 26348 18900 26404 18910
rect 26012 17556 26068 17566
rect 26012 16994 26068 17500
rect 26012 16942 26014 16994
rect 26066 16942 26068 16994
rect 26012 16884 26068 16942
rect 26012 16818 26068 16828
rect 25900 16370 25956 16380
rect 25788 15374 25790 15426
rect 25842 15374 25844 15426
rect 25788 15362 25844 15374
rect 25900 16212 25956 16222
rect 25900 15426 25956 16156
rect 26124 15652 26180 18396
rect 26236 18844 26348 18900
rect 26236 17556 26292 18844
rect 26348 18834 26404 18844
rect 26348 18450 26404 18462
rect 26348 18398 26350 18450
rect 26402 18398 26404 18450
rect 26348 18116 26404 18398
rect 26348 17780 26404 18060
rect 26348 17714 26404 17724
rect 26236 17554 26404 17556
rect 26236 17502 26238 17554
rect 26290 17502 26404 17554
rect 26236 17500 26404 17502
rect 26236 17490 26292 17500
rect 26124 15586 26180 15596
rect 26236 17108 26292 17118
rect 25900 15374 25902 15426
rect 25954 15374 25956 15426
rect 25900 15362 25956 15374
rect 25676 15316 25732 15326
rect 25676 15148 25732 15260
rect 26236 15148 26292 17052
rect 26348 15876 26404 17500
rect 26460 16098 26516 18958
rect 28028 19012 28084 19022
rect 28364 19012 28420 19292
rect 28476 19234 28532 20188
rect 28588 20178 28644 20188
rect 28700 19684 28756 20636
rect 28812 20626 28868 20636
rect 28476 19182 28478 19234
rect 28530 19182 28532 19234
rect 28476 19170 28532 19182
rect 28588 19628 28756 19684
rect 28588 19122 28644 19628
rect 28588 19070 28590 19122
rect 28642 19070 28644 19122
rect 28588 19012 28644 19070
rect 28364 18956 28532 19012
rect 28028 18918 28084 18956
rect 26916 18844 27180 18854
rect 26972 18788 27020 18844
rect 27076 18788 27124 18844
rect 26916 18778 27180 18788
rect 28028 18788 28084 18798
rect 28028 18676 28084 18732
rect 28028 18674 28308 18676
rect 28028 18622 28030 18674
rect 28082 18622 28308 18674
rect 28028 18620 28308 18622
rect 28028 18610 28084 18620
rect 27804 18562 27860 18574
rect 27804 18510 27806 18562
rect 27858 18510 27860 18562
rect 26796 18450 26852 18462
rect 26796 18398 26798 18450
rect 26850 18398 26852 18450
rect 26796 17892 26852 18398
rect 26796 17826 26852 17836
rect 26908 18450 26964 18462
rect 26908 18398 26910 18450
rect 26962 18398 26964 18450
rect 26572 17668 26628 17678
rect 26796 17668 26852 17678
rect 26572 17666 26852 17668
rect 26572 17614 26574 17666
rect 26626 17614 26798 17666
rect 26850 17614 26852 17666
rect 26572 17612 26852 17614
rect 26572 17602 26628 17612
rect 26796 17602 26852 17612
rect 26684 17444 26740 17454
rect 26908 17444 26964 18398
rect 27020 18452 27076 18462
rect 27020 18358 27076 18396
rect 27356 18452 27412 18462
rect 27580 18452 27636 18462
rect 27412 18396 27524 18452
rect 27356 18386 27412 18396
rect 27468 18338 27524 18396
rect 27468 18286 27470 18338
rect 27522 18286 27524 18338
rect 27468 18274 27524 18286
rect 27132 18228 27188 18238
rect 27020 18172 27132 18228
rect 27020 17666 27076 18172
rect 27132 18162 27188 18172
rect 27356 18228 27412 18238
rect 27020 17614 27022 17666
rect 27074 17614 27076 17666
rect 27020 17602 27076 17614
rect 26460 16046 26462 16098
rect 26514 16046 26516 16098
rect 26460 16034 26516 16046
rect 26572 17388 26684 17444
rect 26348 15820 26516 15876
rect 25676 15092 26292 15148
rect 25788 14532 25844 14542
rect 25564 13916 25732 13972
rect 25564 13748 25620 13758
rect 25452 13746 25620 13748
rect 25452 13694 25566 13746
rect 25618 13694 25620 13746
rect 25452 13692 25620 13694
rect 25564 13682 25620 13692
rect 25340 12338 25396 12348
rect 25452 13076 25508 13086
rect 25452 12740 25508 13020
rect 25452 12178 25508 12684
rect 25452 12126 25454 12178
rect 25506 12126 25508 12178
rect 25452 12114 25508 12126
rect 25676 11732 25732 13916
rect 25788 13860 25844 14476
rect 25788 13766 25844 13804
rect 25900 14084 25956 14094
rect 25900 12404 25956 14028
rect 26236 13748 26292 15092
rect 26348 15202 26404 15214
rect 26348 15150 26350 15202
rect 26402 15150 26404 15202
rect 26348 14196 26404 15150
rect 26348 14130 26404 14140
rect 26460 14084 26516 15820
rect 26460 14018 26516 14028
rect 26236 13692 26516 13748
rect 26348 13524 26404 13534
rect 25676 11666 25732 11676
rect 25788 12348 25956 12404
rect 26012 13522 26404 13524
rect 26012 13470 26350 13522
rect 26402 13470 26404 13522
rect 26012 13468 26404 13470
rect 25564 11620 25620 11630
rect 25452 11394 25508 11406
rect 25452 11342 25454 11394
rect 25506 11342 25508 11394
rect 24892 11170 24948 11182
rect 24892 11118 24894 11170
rect 24946 11118 24948 11170
rect 24892 11060 24948 11118
rect 25004 11172 25060 11182
rect 25004 11078 25060 11116
rect 25116 11170 25172 11182
rect 25116 11118 25118 11170
rect 25170 11118 25172 11170
rect 24892 10994 24948 11004
rect 23772 10782 23774 10834
rect 23826 10782 23828 10834
rect 23772 10770 23828 10782
rect 23884 10834 24388 10836
rect 23884 10782 24334 10834
rect 24386 10782 24388 10834
rect 23884 10780 24388 10782
rect 23548 10610 23604 10622
rect 23548 10558 23550 10610
rect 23602 10558 23604 10610
rect 23548 10388 23604 10558
rect 23884 10388 23940 10780
rect 24332 10770 24388 10780
rect 24556 10780 24836 10836
rect 23548 10332 23940 10388
rect 24108 10610 24164 10622
rect 24108 10558 24110 10610
rect 24162 10558 24164 10610
rect 24108 10164 24164 10558
rect 24220 10612 24276 10622
rect 24220 10518 24276 10556
rect 24108 10098 24164 10108
rect 22540 9826 22596 9996
rect 22652 9996 23044 10052
rect 22652 9938 22708 9996
rect 22652 9886 22654 9938
rect 22706 9886 22708 9938
rect 22652 9874 22708 9886
rect 22540 9774 22542 9826
rect 22594 9774 22596 9826
rect 22540 9762 22596 9774
rect 23212 9828 23268 9838
rect 24108 9828 24164 9838
rect 24556 9828 24612 10780
rect 25116 10724 25172 11118
rect 25116 10658 25172 10668
rect 23212 9826 23828 9828
rect 23212 9774 23214 9826
rect 23266 9774 23828 9826
rect 23212 9772 23828 9774
rect 23212 9762 23268 9772
rect 22764 9604 22820 9614
rect 22428 9602 22820 9604
rect 22428 9550 22766 9602
rect 22818 9550 22820 9602
rect 22428 9548 22820 9550
rect 22764 9538 22820 9548
rect 22428 9268 22484 9278
rect 22316 9266 22484 9268
rect 22316 9214 22430 9266
rect 22482 9214 22484 9266
rect 22316 9212 22484 9214
rect 22428 9202 22484 9212
rect 23772 9266 23828 9772
rect 24108 9826 24276 9828
rect 24108 9774 24110 9826
rect 24162 9774 24276 9826
rect 24108 9772 24276 9774
rect 24108 9762 24164 9772
rect 23772 9214 23774 9266
rect 23826 9214 23828 9266
rect 23772 9202 23828 9214
rect 22204 8878 22206 8930
rect 22258 8878 22260 8930
rect 22204 8866 22260 8878
rect 22652 9154 22708 9166
rect 22652 9102 22654 9154
rect 22706 9102 22708 9154
rect 22652 8820 22708 9102
rect 23996 9154 24052 9166
rect 23996 9102 23998 9154
rect 24050 9102 24052 9154
rect 22764 9044 22820 9054
rect 22764 8950 22820 8988
rect 23996 8820 24052 9102
rect 24108 9156 24164 9166
rect 24108 9062 24164 9100
rect 24220 9044 24276 9772
rect 24556 9762 24612 9772
rect 24668 10610 24724 10622
rect 24668 10558 24670 10610
rect 24722 10558 24724 10610
rect 24668 9268 24724 10558
rect 25228 10612 25284 10622
rect 25228 10518 25284 10556
rect 25340 10498 25396 10510
rect 25340 10446 25342 10498
rect 25394 10446 25396 10498
rect 25340 10276 25396 10446
rect 24780 10220 25396 10276
rect 24780 9938 24836 10220
rect 24780 9886 24782 9938
rect 24834 9886 24836 9938
rect 24780 9874 24836 9886
rect 25228 10052 25284 10062
rect 24780 9268 24836 9278
rect 25228 9268 25284 9996
rect 24668 9266 24836 9268
rect 24668 9214 24782 9266
rect 24834 9214 24836 9266
rect 24668 9212 24836 9214
rect 24780 9202 24836 9212
rect 25004 9212 25228 9268
rect 24332 9156 24388 9166
rect 24556 9156 24612 9166
rect 24388 9100 24500 9156
rect 24332 9090 24388 9100
rect 24220 8978 24276 8988
rect 24444 9042 24500 9100
rect 24556 9062 24612 9100
rect 24444 8990 24446 9042
rect 24498 8990 24500 9042
rect 24444 8978 24500 8990
rect 22652 8764 23044 8820
rect 22632 8652 22896 8662
rect 22688 8596 22736 8652
rect 22792 8596 22840 8652
rect 22632 8586 22896 8596
rect 20524 6018 20692 6020
rect 20524 5966 20526 6018
rect 20578 5966 20692 6018
rect 20524 5964 20692 5966
rect 20748 6468 20804 6478
rect 20524 5954 20580 5964
rect 20748 5908 20804 6412
rect 20860 5908 20916 5918
rect 20748 5906 20916 5908
rect 20748 5854 20862 5906
rect 20914 5854 20916 5906
rect 20748 5852 20916 5854
rect 20076 4946 20132 4956
rect 20636 5684 20692 5694
rect 20076 4452 20132 4462
rect 19964 4450 20132 4452
rect 19964 4398 20078 4450
rect 20130 4398 20132 4450
rect 19964 4396 20132 4398
rect 20076 4386 20132 4396
rect 19292 4286 19294 4338
rect 19346 4286 19348 4338
rect 19292 4274 19348 4286
rect 17388 3502 17390 3554
rect 17442 3502 17444 3554
rect 17388 3490 17444 3502
rect 17500 3668 17556 3678
rect 17164 3390 17166 3442
rect 17218 3390 17220 3442
rect 17164 3378 17220 3390
rect 17500 800 17556 3612
rect 17612 3556 17668 3566
rect 17612 3462 17668 3500
rect 18396 3556 18452 4172
rect 18620 3668 18676 3678
rect 18620 3574 18676 3612
rect 19068 3668 19124 3678
rect 18396 3490 18452 3500
rect 18348 3164 18612 3174
rect 18404 3108 18452 3164
rect 18508 3108 18556 3164
rect 18348 3098 18612 3108
rect 19068 800 19124 3612
rect 20636 800 20692 5628
rect 20748 5234 20804 5852
rect 20860 5842 20916 5852
rect 20748 5182 20750 5234
rect 20802 5182 20804 5234
rect 20748 5170 20804 5182
rect 21756 5122 21812 6636
rect 22092 7364 22148 7374
rect 22092 6690 22148 7308
rect 22632 7084 22896 7094
rect 22688 7028 22736 7084
rect 22792 7028 22840 7084
rect 22632 7018 22896 7028
rect 22092 6638 22094 6690
rect 22146 6638 22148 6690
rect 22092 6626 22148 6638
rect 22988 5796 23044 8764
rect 23996 8754 24052 8764
rect 23772 8484 23828 8494
rect 23660 8428 23772 8484
rect 23436 7476 23492 7486
rect 23436 7382 23492 7420
rect 23548 7364 23604 7374
rect 23548 7270 23604 7308
rect 22988 5730 23044 5740
rect 21868 5684 21924 5694
rect 21868 5590 21924 5628
rect 22632 5516 22896 5526
rect 22688 5460 22736 5516
rect 22792 5460 22840 5516
rect 22632 5450 22896 5460
rect 22540 5236 22596 5246
rect 22540 5142 22596 5180
rect 21756 5070 21758 5122
rect 21810 5070 21812 5122
rect 21756 5058 21812 5070
rect 22876 5012 22932 5022
rect 22764 4564 22820 4574
rect 22652 4452 22708 4462
rect 22204 4396 22652 4452
rect 22204 4226 22260 4396
rect 22652 4358 22708 4396
rect 22764 4450 22820 4508
rect 22764 4398 22766 4450
rect 22818 4398 22820 4450
rect 22764 4386 22820 4398
rect 22204 4174 22206 4226
rect 22258 4174 22260 4226
rect 22204 4162 22260 4174
rect 22652 4116 22708 4126
rect 22876 4116 22932 4956
rect 23660 4788 23716 8428
rect 23772 8418 23828 8428
rect 24444 8484 24500 8494
rect 23884 7812 23940 7822
rect 23772 7474 23828 7486
rect 23772 7422 23774 7474
rect 23826 7422 23828 7474
rect 23772 6804 23828 7422
rect 23772 6738 23828 6748
rect 23884 4900 23940 7756
rect 24444 7698 24500 8428
rect 25004 8370 25060 9212
rect 25228 9174 25284 9212
rect 25452 9268 25508 11342
rect 25564 10722 25620 11564
rect 25564 10670 25566 10722
rect 25618 10670 25620 10722
rect 25564 10658 25620 10670
rect 25676 11172 25732 11182
rect 25676 10610 25732 11116
rect 25676 10558 25678 10610
rect 25730 10558 25732 10610
rect 25676 10546 25732 10558
rect 25564 9268 25620 9278
rect 25452 9266 25620 9268
rect 25452 9214 25566 9266
rect 25618 9214 25620 9266
rect 25452 9212 25620 9214
rect 25004 8318 25006 8370
rect 25058 8318 25060 8370
rect 25004 8306 25060 8318
rect 25452 7812 25508 9212
rect 25564 9202 25620 9212
rect 25788 8260 25844 12348
rect 25900 12180 25956 12218
rect 25900 12114 25956 12124
rect 25900 11956 25956 11966
rect 25900 11862 25956 11900
rect 26012 11394 26068 13468
rect 26348 13458 26404 13468
rect 26348 13076 26404 13086
rect 26012 11342 26014 11394
rect 26066 11342 26068 11394
rect 26012 11330 26068 11342
rect 26236 13020 26348 13076
rect 26236 11282 26292 13020
rect 26348 13010 26404 13020
rect 26236 11230 26238 11282
rect 26290 11230 26292 11282
rect 26236 11218 26292 11230
rect 26460 10836 26516 13692
rect 26572 11788 26628 17388
rect 26684 17378 26740 17388
rect 26796 17388 26964 17444
rect 26796 17108 26852 17388
rect 26916 17276 27180 17286
rect 26972 17220 27020 17276
rect 27076 17220 27124 17276
rect 26916 17210 27180 17220
rect 27356 17108 27412 18172
rect 27580 18116 27636 18396
rect 27468 18060 27636 18116
rect 27468 17554 27524 18060
rect 27468 17502 27470 17554
rect 27522 17502 27524 17554
rect 27468 17444 27524 17502
rect 27468 17378 27524 17388
rect 27580 17556 27636 17566
rect 26796 17052 26964 17108
rect 26684 16996 26740 17006
rect 26684 16902 26740 16940
rect 26908 16882 26964 17052
rect 27356 17042 27412 17052
rect 27580 17106 27636 17500
rect 27580 17054 27582 17106
rect 27634 17054 27636 17106
rect 27580 17042 27636 17054
rect 26908 16830 26910 16882
rect 26962 16830 26964 16882
rect 26796 16660 26852 16670
rect 26796 15986 26852 16604
rect 26908 16436 26964 16830
rect 27804 16884 27860 18510
rect 27916 18564 27972 18574
rect 27916 17554 27972 18508
rect 28140 18228 28196 18238
rect 28140 18134 28196 18172
rect 27916 17502 27918 17554
rect 27970 17502 27972 17554
rect 27916 17490 27972 17502
rect 28028 17892 28084 17902
rect 27916 17108 27972 17118
rect 28028 17108 28084 17836
rect 27916 17106 28084 17108
rect 27916 17054 27918 17106
rect 27970 17054 28084 17106
rect 27916 17052 28084 17054
rect 27916 17042 27972 17052
rect 27804 16828 27972 16884
rect 27244 16660 27300 16670
rect 27244 16566 27300 16604
rect 27468 16660 27524 16670
rect 27468 16658 27636 16660
rect 27468 16606 27470 16658
rect 27522 16606 27636 16658
rect 27468 16604 27636 16606
rect 27468 16594 27524 16604
rect 26908 16380 27188 16436
rect 26796 15934 26798 15986
rect 26850 15934 26852 15986
rect 26796 15876 26852 15934
rect 26908 15988 26964 15998
rect 26908 15894 26964 15932
rect 26796 15810 26852 15820
rect 27020 15876 27076 15914
rect 27020 15810 27076 15820
rect 27132 15876 27188 16380
rect 27468 16324 27524 16334
rect 27468 16098 27524 16268
rect 27468 16046 27470 16098
rect 27522 16046 27524 16098
rect 27468 16034 27524 16046
rect 27132 15874 27300 15876
rect 27132 15822 27134 15874
rect 27186 15822 27300 15874
rect 27132 15820 27300 15822
rect 27132 15810 27188 15820
rect 26916 15708 27180 15718
rect 26972 15652 27020 15708
rect 27076 15652 27124 15708
rect 26916 15642 27180 15652
rect 26908 15314 26964 15326
rect 26908 15262 26910 15314
rect 26962 15262 26964 15314
rect 26908 15092 26964 15262
rect 27132 15316 27188 15326
rect 27132 15222 27188 15260
rect 26908 15026 26964 15036
rect 26916 14140 27180 14150
rect 26972 14084 27020 14140
rect 27076 14084 27124 14140
rect 26916 14074 27180 14084
rect 27244 13972 27300 15820
rect 27580 15652 27636 16604
rect 27916 16098 27972 16828
rect 28028 16772 28084 16782
rect 28028 16678 28084 16716
rect 28028 16548 28084 16558
rect 28028 16210 28084 16492
rect 28028 16158 28030 16210
rect 28082 16158 28084 16210
rect 28028 16146 28084 16158
rect 27916 16046 27918 16098
rect 27970 16046 27972 16098
rect 27692 15876 27748 15886
rect 27692 15782 27748 15820
rect 27580 15596 27748 15652
rect 27468 15540 27524 15550
rect 27356 15202 27412 15214
rect 27356 15150 27358 15202
rect 27410 15150 27412 15202
rect 27356 14980 27412 15150
rect 27356 14914 27412 14924
rect 27468 14530 27524 15484
rect 27468 14478 27470 14530
rect 27522 14478 27524 14530
rect 27468 14466 27524 14478
rect 27580 15314 27636 15326
rect 27580 15262 27582 15314
rect 27634 15262 27636 15314
rect 27580 14980 27636 15262
rect 27692 15148 27748 15596
rect 27804 15316 27860 15326
rect 27804 15222 27860 15260
rect 27692 15092 27860 15148
rect 27580 14532 27636 14924
rect 27580 14466 27636 14476
rect 27692 14868 27748 14878
rect 26908 13916 27300 13972
rect 26684 13522 26740 13534
rect 26684 13470 26686 13522
rect 26738 13470 26740 13522
rect 26684 13188 26740 13470
rect 26684 13122 26740 13132
rect 26796 13076 26852 13086
rect 26796 12982 26852 13020
rect 26908 12740 26964 13916
rect 27356 13860 27412 13870
rect 27580 13860 27636 13870
rect 27356 13858 27580 13860
rect 27356 13806 27358 13858
rect 27410 13806 27580 13858
rect 27356 13804 27580 13806
rect 27356 13794 27412 13804
rect 27580 13794 27636 13804
rect 27132 13746 27188 13758
rect 27132 13694 27134 13746
rect 27186 13694 27188 13746
rect 27132 13524 27188 13694
rect 27132 13458 27188 13468
rect 27580 13636 27636 13646
rect 26796 12684 26964 12740
rect 27244 13412 27300 13422
rect 26796 11956 26852 12684
rect 26916 12572 27180 12582
rect 26972 12516 27020 12572
rect 27076 12516 27124 12572
rect 26916 12506 27180 12516
rect 27244 12178 27300 13356
rect 27244 12126 27246 12178
rect 27298 12126 27300 12178
rect 26908 11956 26964 11966
rect 26796 11900 26908 11956
rect 26908 11890 26964 11900
rect 26572 11732 26852 11788
rect 26796 11506 26852 11732
rect 26796 11454 26798 11506
rect 26850 11454 26852 11506
rect 26796 11442 26852 11454
rect 26916 11004 27180 11014
rect 26972 10948 27020 11004
rect 27076 10948 27124 11004
rect 26916 10938 27180 10948
rect 26572 10836 26628 10846
rect 26460 10834 26628 10836
rect 26460 10782 26574 10834
rect 26626 10782 26628 10834
rect 26460 10780 26628 10782
rect 26572 10770 26628 10780
rect 26908 10724 26964 10734
rect 26908 9938 26964 10668
rect 26908 9886 26910 9938
rect 26962 9886 26964 9938
rect 26908 9874 26964 9886
rect 27244 9940 27300 12126
rect 27468 13412 27524 13422
rect 27468 12628 27524 13356
rect 27580 12962 27636 13580
rect 27580 12910 27582 12962
rect 27634 12910 27636 12962
rect 27580 12898 27636 12910
rect 27356 11396 27412 11406
rect 27468 11396 27524 12572
rect 27356 11394 27524 11396
rect 27356 11342 27358 11394
rect 27410 11342 27524 11394
rect 27356 11340 27524 11342
rect 27580 12180 27636 12190
rect 27580 11394 27636 12124
rect 27580 11342 27582 11394
rect 27634 11342 27636 11394
rect 27356 11330 27412 11340
rect 27580 11330 27636 11342
rect 27692 10948 27748 14812
rect 27804 13188 27860 15092
rect 27916 14756 27972 16046
rect 28140 16100 28196 16110
rect 28252 16100 28308 18620
rect 28364 18450 28420 18462
rect 28364 18398 28366 18450
rect 28418 18398 28420 18450
rect 28364 17220 28420 18398
rect 28476 17890 28532 18956
rect 28588 18946 28644 18956
rect 28700 19236 28756 19246
rect 28700 18450 28756 19180
rect 28924 18788 28980 23100
rect 29036 22372 29092 23214
rect 29148 23156 29204 23660
rect 29148 23090 29204 23100
rect 29260 23154 29316 23660
rect 29260 23102 29262 23154
rect 29314 23102 29316 23154
rect 29036 22306 29092 22316
rect 29148 22484 29204 22494
rect 29148 22370 29204 22428
rect 29148 22318 29150 22370
rect 29202 22318 29204 22370
rect 29148 22306 29204 22318
rect 29260 22372 29316 23102
rect 29260 22306 29316 22316
rect 29260 21700 29316 21710
rect 29260 21586 29316 21644
rect 29260 21534 29262 21586
rect 29314 21534 29316 21586
rect 29260 21522 29316 21534
rect 29372 21028 29428 23886
rect 29484 22932 29540 24332
rect 29596 23156 29652 23166
rect 29708 23156 29764 25116
rect 30044 25060 30100 25070
rect 30100 25004 30212 25060
rect 30044 24994 30100 25004
rect 29596 23154 29764 23156
rect 29596 23102 29598 23154
rect 29650 23102 29764 23154
rect 29596 23100 29764 23102
rect 29820 24276 29876 24286
rect 29596 23090 29652 23100
rect 29820 22932 29876 24220
rect 29932 23156 29988 23166
rect 29932 23062 29988 23100
rect 29484 22876 29764 22932
rect 29484 22260 29540 22270
rect 29484 22258 29652 22260
rect 29484 22206 29486 22258
rect 29538 22206 29652 22258
rect 29484 22204 29652 22206
rect 29484 22194 29540 22204
rect 28700 18398 28702 18450
rect 28754 18398 28756 18450
rect 28700 18386 28756 18398
rect 28812 18732 28980 18788
rect 29036 20972 29428 21028
rect 29596 21698 29652 22204
rect 29708 22146 29764 22876
rect 29820 22866 29876 22876
rect 29708 22094 29710 22146
rect 29762 22094 29764 22146
rect 29708 22082 29764 22094
rect 29820 22484 29876 22494
rect 29820 21812 29876 22428
rect 29932 22258 29988 22270
rect 29932 22206 29934 22258
rect 29986 22206 29988 22258
rect 29932 22148 29988 22206
rect 29932 22082 29988 22092
rect 30044 22260 30100 22270
rect 29596 21646 29598 21698
rect 29650 21646 29652 21698
rect 28476 17838 28478 17890
rect 28530 17838 28532 17890
rect 28476 17826 28532 17838
rect 28700 17892 28756 17902
rect 28588 17668 28644 17678
rect 28588 17574 28644 17612
rect 28476 17444 28532 17454
rect 28476 17350 28532 17388
rect 28700 17332 28756 17836
rect 28588 17276 28756 17332
rect 28364 17164 28532 17220
rect 28364 16996 28420 17006
rect 28364 16902 28420 16940
rect 28476 16436 28532 17164
rect 28476 16370 28532 16380
rect 28588 17106 28644 17276
rect 28588 17054 28590 17106
rect 28642 17054 28644 17106
rect 28140 16098 28308 16100
rect 28140 16046 28142 16098
rect 28194 16046 28308 16098
rect 28140 16044 28308 16046
rect 28140 16034 28196 16044
rect 28252 15316 28308 16044
rect 28252 15250 28308 15260
rect 28364 16324 28420 16334
rect 28140 15092 28196 15102
rect 27916 14690 27972 14700
rect 28028 15090 28196 15092
rect 28028 15038 28142 15090
rect 28194 15038 28196 15090
rect 28028 15036 28196 15038
rect 27916 14420 27972 14430
rect 27916 14326 27972 14364
rect 28028 14196 28084 15036
rect 28140 15026 28196 15036
rect 28252 15092 28308 15102
rect 27916 14140 28084 14196
rect 27916 13412 27972 14140
rect 28140 13860 28196 13870
rect 28140 13766 28196 13804
rect 27916 13346 27972 13356
rect 28028 13746 28084 13758
rect 28028 13694 28030 13746
rect 28082 13694 28084 13746
rect 27916 13188 27972 13198
rect 27804 13186 27972 13188
rect 27804 13134 27918 13186
rect 27970 13134 27972 13186
rect 27804 13132 27972 13134
rect 27916 13122 27972 13132
rect 27804 12852 27860 12862
rect 27804 11282 27860 12796
rect 27916 11620 27972 11630
rect 28028 11620 28084 13694
rect 28252 13186 28308 15036
rect 28364 14756 28420 16268
rect 28588 16212 28644 17054
rect 28588 16098 28644 16156
rect 28588 16046 28590 16098
rect 28642 16046 28644 16098
rect 28588 15988 28644 16046
rect 28812 16882 28868 18732
rect 28924 18564 28980 18574
rect 28924 16994 28980 18508
rect 29036 17892 29092 20972
rect 29148 20802 29204 20814
rect 29148 20750 29150 20802
rect 29202 20750 29204 20802
rect 29148 20692 29204 20750
rect 29148 20626 29204 20636
rect 29372 20802 29428 20814
rect 29372 20750 29374 20802
rect 29426 20750 29428 20802
rect 29372 20244 29428 20750
rect 29372 20178 29428 20188
rect 29260 20130 29316 20142
rect 29260 20078 29262 20130
rect 29314 20078 29316 20130
rect 29260 19796 29316 20078
rect 29484 20020 29540 20030
rect 29484 19926 29540 19964
rect 29260 19730 29316 19740
rect 29036 17826 29092 17836
rect 29148 19684 29204 19694
rect 29148 18450 29204 19628
rect 29148 18398 29150 18450
rect 29202 18398 29204 18450
rect 29148 17332 29204 18398
rect 29260 19460 29316 19470
rect 29260 17778 29316 19404
rect 29484 19236 29540 19246
rect 29596 19236 29652 21646
rect 29708 21756 29876 21812
rect 29708 21026 29764 21756
rect 29932 21700 29988 21710
rect 29708 20974 29710 21026
rect 29762 20974 29764 21026
rect 29708 20962 29764 20974
rect 29820 21644 29932 21700
rect 29708 20018 29764 20030
rect 29708 19966 29710 20018
rect 29762 19966 29764 20018
rect 29708 19460 29764 19966
rect 29708 19394 29764 19404
rect 29540 19180 29652 19236
rect 29484 19170 29540 19180
rect 29260 17726 29262 17778
rect 29314 17726 29316 17778
rect 29260 17714 29316 17726
rect 29372 19124 29428 19134
rect 29372 18676 29428 19068
rect 29820 18900 29876 21644
rect 29932 21634 29988 21644
rect 30044 21588 30100 22204
rect 30044 21474 30100 21532
rect 30044 21422 30046 21474
rect 30098 21422 30100 21474
rect 30044 21410 30100 21422
rect 30156 19684 30212 25004
rect 30268 24610 30324 26852
rect 30716 25620 30772 27582
rect 30268 24558 30270 24610
rect 30322 24558 30324 24610
rect 30268 24546 30324 24558
rect 30604 25564 30772 25620
rect 30604 25172 30660 25564
rect 30492 24164 30548 24174
rect 30604 24164 30660 25116
rect 30548 24108 30660 24164
rect 30716 24500 30772 24510
rect 30492 24098 30548 24108
rect 30268 23156 30324 23166
rect 30268 22708 30324 23100
rect 30268 22642 30324 22652
rect 30604 22932 30660 22942
rect 30604 22370 30660 22876
rect 30716 22482 30772 24444
rect 30828 24162 30884 29708
rect 30940 25730 30996 36204
rect 31612 36036 31668 36204
rect 31808 36200 31920 37000
rect 32928 36200 33040 37000
rect 34048 36200 34160 37000
rect 34412 36204 34916 36260
rect 31836 36036 31892 36200
rect 31612 35980 31892 36036
rect 31200 33740 31464 33750
rect 31256 33684 31304 33740
rect 31360 33684 31408 33740
rect 31200 33674 31464 33684
rect 32956 33460 33012 36200
rect 32956 33394 33012 33404
rect 33740 33684 33796 33694
rect 32172 33346 32228 33358
rect 32172 33294 32174 33346
rect 32226 33294 32228 33346
rect 31724 32676 31780 32686
rect 31612 32674 31780 32676
rect 31612 32622 31726 32674
rect 31778 32622 31780 32674
rect 31612 32620 31780 32622
rect 31276 32452 31332 32462
rect 31612 32452 31668 32620
rect 31724 32610 31780 32620
rect 31836 32564 31892 32574
rect 31836 32470 31892 32508
rect 31052 32450 31668 32452
rect 31052 32398 31278 32450
rect 31330 32398 31668 32450
rect 31052 32396 31668 32398
rect 31052 32228 31108 32396
rect 31276 32386 31332 32396
rect 31724 32340 31780 32350
rect 31724 32246 31780 32284
rect 31052 32162 31108 32172
rect 31200 32172 31464 32182
rect 31256 32116 31304 32172
rect 31360 32116 31408 32172
rect 31200 32106 31464 32116
rect 32060 31892 32116 31902
rect 31948 31890 32116 31892
rect 31948 31838 32062 31890
rect 32114 31838 32116 31890
rect 31948 31836 32116 31838
rect 31388 31668 31444 31678
rect 31052 30996 31108 31006
rect 31052 30902 31108 30940
rect 31388 30994 31444 31612
rect 31724 31108 31780 31118
rect 31724 31014 31780 31052
rect 31836 31108 31892 31118
rect 31948 31108 32004 31836
rect 32060 31826 32116 31836
rect 32172 31892 32228 33294
rect 32956 33236 33012 33246
rect 32956 33234 33572 33236
rect 32956 33182 32958 33234
rect 33010 33182 33572 33234
rect 32956 33180 33572 33182
rect 32956 33170 33012 33180
rect 31836 31106 32004 31108
rect 31836 31054 31838 31106
rect 31890 31054 32004 31106
rect 31836 31052 32004 31054
rect 31388 30942 31390 30994
rect 31442 30942 31444 30994
rect 31388 30884 31444 30942
rect 31388 30818 31444 30828
rect 31200 30604 31464 30614
rect 31256 30548 31304 30604
rect 31360 30548 31408 30604
rect 31200 30538 31464 30548
rect 31200 29036 31464 29046
rect 31256 28980 31304 29036
rect 31360 28980 31408 29036
rect 31200 28970 31464 28980
rect 30940 25678 30942 25730
rect 30994 25678 30996 25730
rect 30940 25666 30996 25678
rect 31052 27858 31108 27870
rect 31052 27806 31054 27858
rect 31106 27806 31108 27858
rect 31052 25620 31108 27806
rect 31612 27858 31668 27870
rect 31612 27806 31614 27858
rect 31666 27806 31668 27858
rect 31276 27748 31332 27758
rect 31276 27654 31332 27692
rect 31612 27636 31668 27806
rect 31612 27570 31668 27580
rect 31200 27468 31464 27478
rect 31256 27412 31304 27468
rect 31360 27412 31408 27468
rect 31200 27402 31464 27412
rect 31836 26908 31892 31052
rect 32060 30996 32116 31006
rect 32060 30902 32116 30940
rect 32060 29316 32116 29326
rect 31500 26852 31892 26908
rect 31948 29314 32116 29316
rect 31948 29262 32062 29314
rect 32114 29262 32116 29314
rect 31948 29260 32116 29262
rect 31948 26908 32004 29260
rect 32060 29250 32116 29260
rect 32172 28756 32228 31836
rect 32284 32676 32340 32686
rect 32284 31780 32340 32620
rect 32732 32004 32788 32014
rect 32284 31714 32340 31724
rect 32396 31778 32452 31790
rect 32396 31726 32398 31778
rect 32450 31726 32452 31778
rect 32396 31332 32452 31726
rect 32284 31276 32452 31332
rect 32284 29652 32340 31276
rect 32396 31106 32452 31118
rect 32396 31054 32398 31106
rect 32450 31054 32452 31106
rect 32396 30996 32452 31054
rect 32396 30930 32452 30940
rect 32508 30996 32564 31006
rect 32508 30994 32676 30996
rect 32508 30942 32510 30994
rect 32562 30942 32676 30994
rect 32508 30940 32676 30942
rect 32508 30930 32564 30940
rect 32396 30772 32452 30782
rect 32396 30678 32452 30716
rect 32508 30324 32564 30334
rect 32508 30230 32564 30268
rect 32620 29988 32676 30940
rect 32620 29922 32676 29932
rect 32284 29586 32340 29596
rect 32508 29540 32564 29550
rect 32508 29314 32564 29484
rect 32508 29262 32510 29314
rect 32562 29262 32564 29314
rect 32172 28754 32340 28756
rect 32172 28702 32174 28754
rect 32226 28702 32340 28754
rect 32172 28700 32340 28702
rect 32172 28690 32228 28700
rect 32060 28196 32116 28206
rect 32060 27970 32116 28140
rect 32060 27918 32062 27970
rect 32114 27918 32116 27970
rect 32060 27906 32116 27918
rect 32172 27972 32228 27982
rect 32172 27878 32228 27916
rect 32060 27748 32116 27758
rect 32060 27654 32116 27692
rect 32172 27636 32228 27646
rect 31948 26852 32116 26908
rect 31500 26290 31556 26852
rect 31500 26238 31502 26290
rect 31554 26238 31556 26290
rect 31500 26226 31556 26238
rect 31948 26178 32004 26190
rect 31948 26126 31950 26178
rect 32002 26126 32004 26178
rect 31200 25900 31464 25910
rect 31256 25844 31304 25900
rect 31360 25844 31408 25900
rect 31200 25834 31464 25844
rect 31052 25564 31220 25620
rect 31052 25060 31108 25070
rect 30828 24110 30830 24162
rect 30882 24110 30884 24162
rect 30828 24098 30884 24110
rect 30940 24948 30996 24958
rect 30940 23378 30996 24892
rect 30940 23326 30942 23378
rect 30994 23326 30996 23378
rect 30940 23314 30996 23326
rect 30716 22430 30718 22482
rect 30770 22430 30772 22482
rect 30716 22418 30772 22430
rect 30828 22932 30884 22942
rect 30604 22318 30606 22370
rect 30658 22318 30660 22370
rect 30604 22306 30660 22318
rect 30828 22260 30884 22876
rect 30828 22166 30884 22204
rect 30940 22372 30996 22382
rect 30940 22258 30996 22316
rect 30940 22206 30942 22258
rect 30994 22206 30996 22258
rect 30492 21588 30548 21598
rect 30940 21588 30996 22206
rect 31052 21700 31108 25004
rect 31164 24612 31220 25564
rect 31164 24546 31220 24556
rect 31612 25508 31668 25518
rect 31612 24388 31668 25452
rect 31200 24332 31464 24342
rect 31256 24276 31304 24332
rect 31360 24276 31408 24332
rect 31612 24322 31668 24332
rect 31200 24266 31464 24276
rect 31948 23604 32004 26126
rect 31836 23548 32004 23604
rect 32060 24722 32116 26852
rect 32172 24948 32228 27580
rect 32284 27074 32340 28700
rect 32396 27860 32452 27870
rect 32396 27766 32452 27804
rect 32284 27022 32286 27074
rect 32338 27022 32340 27074
rect 32284 26908 32340 27022
rect 32284 26852 32452 26908
rect 32172 24882 32228 24892
rect 32284 26178 32340 26190
rect 32284 26126 32286 26178
rect 32338 26126 32340 26178
rect 32060 24670 32062 24722
rect 32114 24670 32116 24722
rect 31836 23156 31892 23548
rect 31724 23044 31780 23054
rect 31200 22764 31464 22774
rect 31256 22708 31304 22764
rect 31360 22708 31408 22764
rect 31200 22698 31464 22708
rect 31612 22596 31668 22606
rect 31388 22372 31444 22382
rect 31388 22278 31444 22316
rect 31612 22370 31668 22540
rect 31612 22318 31614 22370
rect 31666 22318 31668 22370
rect 31612 22306 31668 22318
rect 31052 21634 31108 21644
rect 30380 21476 30436 21486
rect 30268 20692 30324 20702
rect 30268 20130 30324 20636
rect 30268 20078 30270 20130
rect 30322 20078 30324 20130
rect 30268 20066 30324 20078
rect 30156 19618 30212 19628
rect 30156 19460 30212 19470
rect 30044 19346 30100 19358
rect 30044 19294 30046 19346
rect 30098 19294 30100 19346
rect 30044 19236 30100 19294
rect 29932 19124 29988 19134
rect 29932 19030 29988 19068
rect 29820 18844 29988 18900
rect 29596 18676 29652 18686
rect 29372 18674 29652 18676
rect 29372 18622 29598 18674
rect 29650 18622 29652 18674
rect 29372 18620 29652 18622
rect 29148 17266 29204 17276
rect 28924 16942 28926 16994
rect 28978 16942 28980 16994
rect 28924 16930 28980 16942
rect 28812 16830 28814 16882
rect 28866 16830 28868 16882
rect 28812 15988 28868 16830
rect 29148 16770 29204 16782
rect 29148 16718 29150 16770
rect 29202 16718 29204 16770
rect 29148 16324 29204 16718
rect 29148 16258 29204 16268
rect 29260 16212 29316 16222
rect 29260 16118 29316 16156
rect 28812 15932 29316 15988
rect 28588 15922 28644 15932
rect 28476 15874 28532 15886
rect 28476 15822 28478 15874
rect 28530 15822 28532 15874
rect 28476 15316 28532 15822
rect 28700 15876 28756 15886
rect 28476 15260 28644 15316
rect 28476 15092 28532 15102
rect 28476 14998 28532 15036
rect 28588 14868 28644 15260
rect 28588 14802 28644 14812
rect 28700 15314 28756 15820
rect 28700 15262 28702 15314
rect 28754 15262 28756 15314
rect 28476 14756 28532 14766
rect 28364 14754 28532 14756
rect 28364 14702 28478 14754
rect 28530 14702 28532 14754
rect 28364 14700 28532 14702
rect 28476 14690 28532 14700
rect 28588 14418 28644 14430
rect 28588 14366 28590 14418
rect 28642 14366 28644 14418
rect 28476 14308 28532 14318
rect 28252 13134 28254 13186
rect 28306 13134 28308 13186
rect 28252 13122 28308 13134
rect 28364 14306 28532 14308
rect 28364 14254 28478 14306
rect 28530 14254 28532 14306
rect 28364 14252 28532 14254
rect 28364 13076 28420 14252
rect 28476 14242 28532 14252
rect 28588 13300 28644 14366
rect 28588 13234 28644 13244
rect 28364 12852 28420 13020
rect 28476 13076 28532 13086
rect 28700 13076 28756 15262
rect 28924 14980 28980 14990
rect 28476 13074 28756 13076
rect 28476 13022 28478 13074
rect 28530 13022 28756 13074
rect 28476 13020 28756 13022
rect 28812 14756 28868 14766
rect 28812 13746 28868 14700
rect 28812 13694 28814 13746
rect 28866 13694 28868 13746
rect 28476 13010 28532 13020
rect 28364 12786 28420 12796
rect 28812 12628 28868 13694
rect 27916 11618 28084 11620
rect 27916 11566 27918 11618
rect 27970 11566 28084 11618
rect 27916 11564 28084 11566
rect 28140 12572 28868 12628
rect 27916 11554 27972 11564
rect 27804 11230 27806 11282
rect 27858 11230 27860 11282
rect 27804 11218 27860 11230
rect 27356 10892 27748 10948
rect 27356 10834 27412 10892
rect 27356 10782 27358 10834
rect 27410 10782 27412 10834
rect 27356 10770 27412 10782
rect 27580 10500 27636 10510
rect 28140 10500 28196 12572
rect 27580 10498 28196 10500
rect 27580 10446 27582 10498
rect 27634 10446 28196 10498
rect 27580 10444 28196 10446
rect 28252 11732 28308 11742
rect 27580 10434 27636 10444
rect 27356 9940 27412 9950
rect 27244 9938 27412 9940
rect 27244 9886 27358 9938
rect 27410 9886 27412 9938
rect 27244 9884 27412 9886
rect 27356 9874 27412 9884
rect 28252 9826 28308 11676
rect 28476 11620 28532 11630
rect 28476 11526 28532 11564
rect 28364 11282 28420 11294
rect 28364 11230 28366 11282
rect 28418 11230 28420 11282
rect 28364 10724 28420 11230
rect 28364 10658 28420 10668
rect 28252 9774 28254 9826
rect 28306 9774 28308 9826
rect 28028 9604 28084 9614
rect 26916 9436 27180 9446
rect 26972 9380 27020 9436
rect 27076 9380 27124 9436
rect 26916 9370 27180 9380
rect 26012 9268 26068 9278
rect 26348 9268 26404 9278
rect 26068 9266 26404 9268
rect 26068 9214 26350 9266
rect 26402 9214 26404 9266
rect 26068 9212 26404 9214
rect 26012 9174 26068 9212
rect 26348 9202 26404 9212
rect 25788 8194 25844 8204
rect 26684 9154 26740 9166
rect 26684 9102 26686 9154
rect 26738 9102 26740 9154
rect 26684 8148 26740 9102
rect 28028 9154 28084 9548
rect 28028 9102 28030 9154
rect 28082 9102 28084 9154
rect 28028 9090 28084 9102
rect 27356 9044 27412 9054
rect 27356 8950 27412 8988
rect 26684 8082 26740 8092
rect 26796 8260 26852 8270
rect 24444 7646 24446 7698
rect 24498 7646 24500 7698
rect 24444 7634 24500 7646
rect 25228 7756 25508 7812
rect 25900 7812 25956 7822
rect 23996 7476 24052 7486
rect 24220 7476 24276 7486
rect 23996 7474 24164 7476
rect 23996 7422 23998 7474
rect 24050 7422 24164 7474
rect 23996 7420 24164 7422
rect 23996 7410 24052 7420
rect 24108 6132 24164 7420
rect 24220 7382 24276 7420
rect 24556 7474 24612 7486
rect 24556 7422 24558 7474
rect 24610 7422 24612 7474
rect 24220 6802 24276 6814
rect 24220 6750 24222 6802
rect 24274 6750 24276 6802
rect 24220 6356 24276 6750
rect 24556 6580 24612 7422
rect 25116 7474 25172 7486
rect 25116 7422 25118 7474
rect 25170 7422 25172 7474
rect 25116 6690 25172 7422
rect 25116 6638 25118 6690
rect 25170 6638 25172 6690
rect 25116 6626 25172 6638
rect 24556 6486 24612 6524
rect 24332 6468 24388 6478
rect 24332 6356 24388 6412
rect 24668 6466 24724 6478
rect 24668 6414 24670 6466
rect 24722 6414 24724 6466
rect 24220 6300 24388 6356
rect 24220 6132 24276 6142
rect 24108 6130 24276 6132
rect 24108 6078 24222 6130
rect 24274 6078 24276 6130
rect 24108 6076 24276 6078
rect 24220 6066 24276 6076
rect 24332 6130 24388 6300
rect 24332 6078 24334 6130
rect 24386 6078 24388 6130
rect 24332 6066 24388 6078
rect 24556 6356 24612 6366
rect 24556 6130 24612 6300
rect 24556 6078 24558 6130
rect 24610 6078 24612 6130
rect 24444 6020 24500 6030
rect 24108 5906 24164 5918
rect 24108 5854 24110 5906
rect 24162 5854 24164 5906
rect 24108 5124 24164 5854
rect 24108 5058 24164 5068
rect 23884 4844 24164 4900
rect 23660 4732 24052 4788
rect 23212 4564 23268 4574
rect 23212 4470 23268 4508
rect 22652 4114 22932 4116
rect 22652 4062 22654 4114
rect 22706 4062 22932 4114
rect 22652 4060 22932 4062
rect 23772 4226 23828 4238
rect 23772 4174 23774 4226
rect 23826 4174 23828 4226
rect 22652 4050 22708 4060
rect 22632 3948 22896 3958
rect 22688 3892 22736 3948
rect 22792 3892 22840 3948
rect 22632 3882 22896 3892
rect 21868 3668 21924 3678
rect 21868 3574 21924 3612
rect 22204 3668 22260 3678
rect 20748 3556 20804 3566
rect 20748 3462 20804 3500
rect 22204 800 22260 3612
rect 23772 3554 23828 4174
rect 23772 3502 23774 3554
rect 23826 3502 23828 3554
rect 23772 800 23828 3502
rect 23996 3442 24052 4732
rect 24108 4562 24164 4844
rect 24108 4510 24110 4562
rect 24162 4510 24164 4562
rect 24108 4498 24164 4510
rect 24444 4564 24500 5964
rect 24556 5348 24612 6078
rect 24668 6132 24724 6414
rect 24780 6468 24836 6478
rect 24780 6374 24836 6412
rect 25228 6356 25284 7756
rect 25900 7698 25956 7756
rect 25900 7646 25902 7698
rect 25954 7646 25956 7698
rect 25900 7634 25956 7646
rect 25228 6290 25284 6300
rect 25340 7586 25396 7598
rect 25340 7534 25342 7586
rect 25394 7534 25396 7586
rect 24668 6076 25284 6132
rect 25228 6018 25284 6076
rect 25228 5966 25230 6018
rect 25282 5966 25284 6018
rect 25228 5954 25284 5966
rect 25340 6020 25396 7534
rect 26572 7586 26628 7598
rect 26572 7534 26574 7586
rect 26626 7534 26628 7586
rect 25452 7476 25508 7486
rect 25788 7476 25844 7486
rect 25452 7474 25788 7476
rect 25452 7422 25454 7474
rect 25506 7422 25788 7474
rect 25452 7420 25788 7422
rect 25452 7410 25508 7420
rect 25788 7382 25844 7420
rect 26124 7474 26180 7486
rect 26124 7422 26126 7474
rect 26178 7422 26180 7474
rect 25340 5954 25396 5964
rect 25452 6804 25508 6814
rect 25116 5908 25172 5918
rect 25116 5348 25172 5852
rect 25452 5906 25508 6748
rect 25676 6804 25732 6814
rect 25452 5854 25454 5906
rect 25506 5854 25508 5906
rect 24556 5012 24612 5292
rect 24668 5292 25172 5348
rect 24668 5234 24724 5292
rect 24668 5182 24670 5234
rect 24722 5182 24724 5234
rect 24668 5170 24724 5182
rect 25116 5236 25172 5292
rect 25340 5794 25396 5806
rect 25340 5742 25342 5794
rect 25394 5742 25396 5794
rect 25340 5236 25396 5742
rect 25452 5684 25508 5854
rect 25452 5618 25508 5628
rect 25564 6690 25620 6702
rect 25564 6638 25566 6690
rect 25618 6638 25620 6690
rect 25564 5572 25620 6638
rect 25676 6690 25732 6748
rect 25676 6638 25678 6690
rect 25730 6638 25732 6690
rect 25676 6626 25732 6638
rect 26012 6578 26068 6590
rect 26012 6526 26014 6578
rect 26066 6526 26068 6578
rect 25900 6466 25956 6478
rect 25900 6414 25902 6466
rect 25954 6414 25956 6466
rect 25564 5506 25620 5516
rect 25676 5906 25732 5918
rect 25676 5854 25678 5906
rect 25730 5854 25732 5906
rect 25676 5348 25732 5854
rect 25116 5180 25284 5236
rect 24892 5124 24948 5134
rect 24780 5122 24948 5124
rect 24780 5070 24894 5122
rect 24946 5070 24948 5122
rect 24780 5068 24948 5070
rect 24780 5012 24836 5068
rect 24892 5058 24948 5068
rect 24556 4956 24836 5012
rect 25228 5012 25284 5180
rect 25340 5170 25396 5180
rect 25452 5292 25732 5348
rect 25788 5348 25844 5358
rect 25452 5234 25508 5292
rect 25452 5182 25454 5234
rect 25506 5182 25508 5234
rect 25452 5170 25508 5182
rect 25564 5124 25620 5134
rect 25340 5012 25396 5022
rect 25228 5010 25396 5012
rect 25228 4958 25342 5010
rect 25394 4958 25396 5010
rect 25228 4956 25396 4958
rect 25340 4946 25396 4956
rect 25564 5010 25620 5068
rect 25788 5122 25844 5292
rect 25788 5070 25790 5122
rect 25842 5070 25844 5122
rect 25788 5058 25844 5070
rect 25564 4958 25566 5010
rect 25618 4958 25620 5010
rect 25564 4946 25620 4958
rect 24556 4564 24612 4574
rect 24444 4562 24612 4564
rect 24444 4510 24558 4562
rect 24610 4510 24612 4562
rect 24444 4508 24612 4510
rect 24556 4498 24612 4508
rect 24780 4452 24836 4462
rect 25900 4452 25956 6414
rect 26012 5684 26068 6526
rect 26124 5906 26180 7422
rect 26572 7476 26628 7534
rect 26572 7410 26628 7420
rect 26796 7474 26852 8204
rect 27244 8258 27300 8270
rect 27244 8206 27246 8258
rect 27298 8206 27300 8258
rect 27244 8148 27300 8206
rect 27244 8082 27300 8092
rect 28028 8148 28084 8158
rect 28028 8054 28084 8092
rect 27468 8036 27524 8046
rect 27916 8036 27972 8046
rect 27468 8034 27636 8036
rect 27468 7982 27470 8034
rect 27522 7982 27636 8034
rect 27468 7980 27636 7982
rect 27468 7970 27524 7980
rect 26916 7868 27180 7878
rect 26972 7812 27020 7868
rect 27076 7812 27124 7868
rect 26916 7802 27180 7812
rect 26796 7422 26798 7474
rect 26850 7422 26852 7474
rect 26796 7410 26852 7422
rect 27244 7586 27300 7598
rect 27244 7534 27246 7586
rect 27298 7534 27300 7586
rect 26460 6692 26516 6702
rect 26460 6598 26516 6636
rect 26908 6690 26964 6702
rect 26908 6638 26910 6690
rect 26962 6638 26964 6690
rect 26684 6580 26740 6590
rect 26908 6580 26964 6638
rect 27020 6580 27076 6590
rect 26908 6524 27020 6580
rect 26684 6132 26740 6524
rect 27020 6514 27076 6524
rect 26916 6300 27180 6310
rect 26972 6244 27020 6300
rect 27076 6244 27124 6300
rect 26916 6234 27180 6244
rect 27020 6132 27076 6142
rect 27244 6132 27300 7534
rect 27580 7588 27636 7980
rect 27580 7494 27636 7532
rect 27804 7476 27860 7486
rect 27692 7474 27860 7476
rect 27692 7422 27806 7474
rect 27858 7422 27860 7474
rect 27692 7420 27860 7422
rect 27580 6804 27636 6814
rect 27468 6748 27580 6804
rect 27468 6690 27524 6748
rect 27580 6738 27636 6748
rect 27468 6638 27470 6690
rect 27522 6638 27524 6690
rect 27468 6626 27524 6638
rect 26684 6130 27300 6132
rect 26684 6078 26686 6130
rect 26738 6078 27022 6130
rect 27074 6078 27300 6130
rect 26684 6076 27300 6078
rect 27356 6580 27412 6590
rect 26684 6066 26740 6076
rect 27020 6066 27076 6076
rect 27356 6020 27412 6524
rect 26124 5854 26126 5906
rect 26178 5854 26180 5906
rect 26124 5842 26180 5854
rect 26460 5908 26516 5918
rect 26460 5814 26516 5852
rect 27244 5906 27300 5918
rect 27244 5854 27246 5906
rect 27298 5854 27300 5906
rect 26572 5794 26628 5806
rect 26572 5742 26574 5794
rect 26626 5742 26628 5794
rect 26572 5684 26628 5742
rect 26012 5628 26628 5684
rect 27132 5794 27188 5806
rect 27132 5742 27134 5794
rect 27186 5742 27188 5794
rect 26012 5460 26068 5470
rect 26068 5404 26404 5460
rect 26012 5394 26068 5404
rect 26348 5234 26404 5404
rect 26348 5182 26350 5234
rect 26402 5182 26404 5234
rect 26348 5170 26404 5182
rect 26460 5124 26516 5134
rect 26460 5010 26516 5068
rect 27132 5122 27188 5742
rect 27132 5070 27134 5122
rect 27186 5070 27188 5122
rect 27132 5058 27188 5070
rect 26460 4958 26462 5010
rect 26514 4958 26516 5010
rect 26460 4946 26516 4958
rect 26236 4898 26292 4910
rect 26236 4846 26238 4898
rect 26290 4846 26292 4898
rect 26236 4564 26292 4846
rect 26916 4732 27180 4742
rect 26972 4676 27020 4732
rect 27076 4676 27124 4732
rect 26916 4666 27180 4676
rect 26236 4498 26292 4508
rect 27244 4564 27300 5854
rect 27356 5348 27412 5964
rect 27692 5906 27748 7420
rect 27804 7410 27860 7420
rect 27916 7140 27972 7980
rect 28028 7586 28084 7598
rect 28028 7534 28030 7586
rect 28082 7534 28084 7586
rect 28028 7252 28084 7534
rect 28140 7476 28196 7486
rect 28140 7382 28196 7420
rect 28028 7186 28084 7196
rect 27916 7074 27972 7084
rect 28140 6804 28196 6814
rect 28140 6692 28196 6748
rect 28252 6692 28308 9774
rect 28588 9716 28644 9726
rect 28588 9622 28644 9660
rect 28812 9044 28868 9054
rect 28700 8988 28812 9044
rect 28364 8036 28420 8046
rect 28364 7942 28420 7980
rect 28588 7586 28644 7598
rect 28588 7534 28590 7586
rect 28642 7534 28644 7586
rect 28476 7476 28532 7486
rect 28476 7382 28532 7420
rect 28588 7364 28644 7534
rect 28364 7140 28420 7150
rect 28420 7084 28532 7140
rect 28364 7074 28420 7084
rect 28140 6690 28308 6692
rect 28140 6638 28142 6690
rect 28194 6638 28308 6690
rect 28140 6636 28308 6638
rect 28140 6626 28196 6636
rect 27692 5854 27694 5906
rect 27746 5854 27748 5906
rect 27692 5842 27748 5854
rect 27804 6466 27860 6478
rect 27804 6414 27806 6466
rect 27858 6414 27860 6466
rect 27356 5282 27412 5292
rect 27468 5684 27524 5694
rect 27804 5684 27860 6414
rect 28140 6468 28196 6478
rect 28140 6132 28196 6412
rect 28140 6130 28420 6132
rect 28140 6078 28142 6130
rect 28194 6078 28420 6130
rect 28140 6076 28420 6078
rect 28140 6066 28196 6076
rect 27916 6020 27972 6030
rect 27916 5926 27972 5964
rect 28028 5796 28084 5806
rect 27524 5628 27860 5684
rect 27916 5794 28084 5796
rect 27916 5742 28030 5794
rect 28082 5742 28084 5794
rect 27916 5740 28084 5742
rect 27468 5122 27524 5628
rect 27468 5070 27470 5122
rect 27522 5070 27524 5122
rect 27468 5058 27524 5070
rect 27692 5124 27748 5134
rect 27916 5124 27972 5740
rect 28028 5730 28084 5740
rect 28028 5348 28084 5358
rect 28028 5254 28084 5292
rect 27692 5122 27972 5124
rect 27692 5070 27694 5122
rect 27746 5070 27972 5122
rect 27692 5068 27972 5070
rect 27692 5058 27748 5068
rect 28140 5010 28196 5022
rect 28140 4958 28142 5010
rect 28194 4958 28196 5010
rect 27356 4900 27412 4910
rect 27356 4806 27412 4844
rect 27244 4498 27300 4508
rect 28028 4564 28084 4574
rect 26012 4452 26068 4462
rect 25900 4450 26068 4452
rect 25900 4398 26014 4450
rect 26066 4398 26068 4450
rect 25900 4396 26068 4398
rect 24220 4226 24276 4238
rect 24220 4174 24222 4226
rect 24274 4174 24276 4226
rect 24220 3780 24276 4174
rect 24668 4228 24724 4238
rect 24668 4134 24724 4172
rect 24220 3714 24276 3724
rect 24780 3554 24836 4396
rect 26012 4386 26068 4396
rect 25340 4340 25396 4350
rect 25340 4246 25396 4284
rect 27468 4228 27524 4238
rect 28028 4228 28084 4508
rect 28140 4452 28196 4958
rect 28140 4386 28196 4396
rect 28140 4228 28196 4238
rect 28028 4226 28196 4228
rect 28028 4174 28142 4226
rect 28194 4174 28196 4226
rect 28028 4172 28196 4174
rect 28364 4228 28420 6076
rect 28476 5906 28532 7084
rect 28588 6916 28644 7308
rect 28588 6850 28644 6860
rect 28476 5854 28478 5906
rect 28530 5854 28532 5906
rect 28476 5842 28532 5854
rect 28588 6692 28644 6702
rect 28588 5234 28644 6636
rect 28700 5908 28756 8988
rect 28812 8978 28868 8988
rect 28924 7700 28980 14924
rect 29148 14418 29204 14430
rect 29148 14366 29150 14418
rect 29202 14366 29204 14418
rect 29148 13748 29204 14366
rect 29148 13682 29204 13692
rect 29148 13522 29204 13534
rect 29148 13470 29150 13522
rect 29202 13470 29204 13522
rect 29036 13300 29092 13310
rect 29036 12964 29092 13244
rect 29148 13188 29204 13470
rect 29148 13122 29204 13132
rect 29148 12964 29204 12974
rect 29036 12962 29204 12964
rect 29036 12910 29150 12962
rect 29202 12910 29204 12962
rect 29036 12908 29204 12910
rect 29036 12180 29092 12908
rect 29148 12898 29204 12908
rect 29036 12114 29092 12124
rect 29148 11732 29204 11742
rect 29148 11394 29204 11676
rect 29148 11342 29150 11394
rect 29202 11342 29204 11394
rect 29148 11330 29204 11342
rect 29260 10050 29316 15932
rect 29372 15876 29428 18620
rect 29596 18610 29652 18620
rect 29820 18450 29876 18462
rect 29820 18398 29822 18450
rect 29874 18398 29876 18450
rect 29820 18004 29876 18398
rect 29820 17938 29876 17948
rect 29820 17442 29876 17454
rect 29820 17390 29822 17442
rect 29874 17390 29876 17442
rect 29484 16996 29540 17006
rect 29820 16996 29876 17390
rect 29484 16994 29876 16996
rect 29484 16942 29486 16994
rect 29538 16942 29876 16994
rect 29484 16940 29876 16942
rect 29484 16930 29540 16940
rect 29372 15810 29428 15820
rect 29484 16436 29540 16446
rect 29820 16436 29876 16940
rect 29932 16884 29988 18844
rect 30044 18676 30100 19180
rect 30044 18610 30100 18620
rect 30156 19234 30212 19404
rect 30156 19182 30158 19234
rect 30210 19182 30212 19234
rect 30156 18116 30212 19182
rect 30268 19348 30324 19358
rect 30268 18674 30324 19292
rect 30268 18622 30270 18674
rect 30322 18622 30324 18674
rect 30268 18610 30324 18622
rect 30156 18050 30212 18060
rect 30380 17780 30436 21420
rect 30492 20802 30548 21532
rect 30492 20750 30494 20802
rect 30546 20750 30548 20802
rect 30492 20020 30548 20750
rect 30828 21532 30996 21588
rect 31164 21588 31220 21598
rect 31500 21588 31556 21598
rect 31220 21586 31556 21588
rect 31220 21534 31502 21586
rect 31554 21534 31556 21586
rect 31220 21532 31556 21534
rect 30492 19954 30548 19964
rect 30604 20690 30660 20702
rect 30604 20638 30606 20690
rect 30658 20638 30660 20690
rect 30604 19348 30660 20638
rect 30604 19282 30660 19292
rect 30716 19236 30772 19246
rect 30716 19142 30772 19180
rect 30604 18564 30660 18574
rect 30828 18564 30884 21532
rect 31164 21494 31220 21532
rect 31500 21522 31556 21532
rect 30660 18508 30884 18564
rect 30940 21364 30996 21374
rect 30604 18470 30660 18508
rect 30940 18452 30996 21308
rect 31200 21196 31464 21206
rect 31256 21140 31304 21196
rect 31360 21140 31408 21196
rect 31200 21130 31464 21140
rect 31724 20914 31780 22988
rect 31836 21924 31892 23100
rect 31948 23268 32004 23278
rect 31948 22370 32004 23212
rect 31948 22318 31950 22370
rect 32002 22318 32004 22370
rect 31948 22306 32004 22318
rect 32060 23156 32116 24670
rect 32060 22372 32116 23100
rect 32172 23940 32228 23950
rect 32172 22372 32228 23884
rect 32284 23604 32340 26126
rect 32396 23938 32452 26852
rect 32396 23886 32398 23938
rect 32450 23886 32452 23938
rect 32396 23874 32452 23886
rect 32508 23716 32564 29262
rect 32732 27188 32788 31948
rect 33404 31556 33460 31566
rect 33404 31462 33460 31500
rect 33516 31218 33572 33180
rect 33740 32786 33796 33628
rect 33740 32734 33742 32786
rect 33794 32734 33796 32786
rect 33740 32722 33796 32734
rect 33516 31166 33518 31218
rect 33570 31166 33572 31218
rect 33516 31154 33572 31166
rect 33628 32338 33684 32350
rect 33628 32286 33630 32338
rect 33682 32286 33684 32338
rect 33628 31218 33684 32286
rect 34076 32004 34132 36200
rect 34412 32788 34468 36204
rect 34860 36036 34916 36204
rect 35168 36200 35280 37000
rect 35196 36036 35252 36200
rect 34860 35980 35252 36036
rect 35196 34580 35252 34590
rect 35196 33684 35252 34524
rect 35084 33460 35140 33470
rect 34412 32722 34468 32732
rect 34524 33458 35140 33460
rect 34524 33406 35086 33458
rect 35138 33406 35140 33458
rect 34524 33404 35140 33406
rect 34076 31938 34132 31948
rect 34188 32450 34244 32462
rect 34188 32398 34190 32450
rect 34242 32398 34244 32450
rect 33628 31166 33630 31218
rect 33682 31166 33684 31218
rect 33628 31154 33684 31166
rect 33964 31108 34020 31118
rect 33964 31014 34020 31052
rect 32956 30996 33012 31006
rect 32956 30548 33012 30940
rect 33404 30996 33460 31006
rect 33404 30902 33460 30940
rect 32956 30482 33012 30492
rect 33628 30434 33684 30446
rect 33628 30382 33630 30434
rect 33682 30382 33684 30434
rect 33628 30212 33684 30382
rect 33516 30156 33684 30212
rect 34188 30212 34244 32398
rect 34524 32338 34580 33404
rect 35084 33394 35140 33404
rect 34860 32676 34916 32686
rect 34860 32582 34916 32620
rect 35196 32674 35252 33628
rect 35980 33348 36036 33358
rect 35484 32956 35748 32966
rect 35540 32900 35588 32956
rect 35644 32900 35692 32956
rect 35484 32890 35748 32900
rect 35196 32622 35198 32674
rect 35250 32622 35252 32674
rect 35196 32610 35252 32622
rect 34636 32452 34692 32462
rect 34636 32450 35028 32452
rect 34636 32398 34638 32450
rect 34690 32398 35028 32450
rect 34636 32396 35028 32398
rect 34636 32386 34692 32396
rect 34524 32286 34526 32338
rect 34578 32286 34580 32338
rect 34300 30994 34356 31006
rect 34300 30942 34302 30994
rect 34354 30942 34356 30994
rect 34300 30884 34356 30942
rect 34300 30434 34356 30828
rect 34300 30382 34302 30434
rect 34354 30382 34356 30434
rect 34300 30370 34356 30382
rect 34412 30324 34468 30334
rect 34188 30156 34356 30212
rect 33180 29986 33236 29998
rect 33180 29934 33182 29986
rect 33234 29934 33236 29986
rect 33180 29764 33236 29934
rect 33516 29764 33572 30156
rect 33628 30044 34020 30100
rect 33628 29986 33684 30044
rect 33628 29934 33630 29986
rect 33682 29934 33684 29986
rect 33628 29922 33684 29934
rect 33516 29708 33684 29764
rect 33180 29698 33236 29708
rect 33292 29204 33348 29214
rect 33292 29110 33348 29148
rect 33068 28420 33124 28430
rect 33068 27970 33124 28364
rect 33404 28420 33460 28430
rect 33068 27918 33070 27970
rect 33122 27918 33124 27970
rect 33068 27906 33124 27918
rect 33180 28196 33236 28206
rect 32732 27122 32788 27132
rect 33068 26962 33124 26974
rect 33068 26910 33070 26962
rect 33122 26910 33124 26962
rect 32844 26516 32900 26526
rect 32732 26460 32844 26516
rect 32732 23940 32788 26460
rect 32844 26450 32900 26460
rect 33068 26514 33124 26910
rect 33068 26462 33070 26514
rect 33122 26462 33124 26514
rect 33068 26450 33124 26462
rect 33180 26516 33236 28140
rect 33404 27858 33460 28364
rect 33628 28308 33684 29708
rect 33852 29652 33908 29662
rect 33740 29596 33852 29652
rect 33740 29426 33796 29596
rect 33852 29586 33908 29596
rect 33740 29374 33742 29426
rect 33794 29374 33796 29426
rect 33740 29362 33796 29374
rect 33852 29428 33908 29438
rect 33852 29314 33908 29372
rect 33852 29262 33854 29314
rect 33906 29262 33908 29314
rect 33852 29250 33908 29262
rect 33628 28242 33684 28252
rect 33964 28196 34020 30044
rect 34076 29986 34132 29998
rect 34076 29934 34078 29986
rect 34130 29934 34132 29986
rect 34076 28420 34132 29934
rect 34188 29988 34244 29998
rect 34188 29650 34244 29932
rect 34188 29598 34190 29650
rect 34242 29598 34244 29650
rect 34188 29586 34244 29598
rect 34300 29540 34356 30156
rect 34412 29652 34468 30268
rect 34412 29558 34468 29596
rect 34300 29474 34356 29484
rect 34524 29538 34580 32286
rect 34636 30996 34692 31006
rect 34636 30902 34692 30940
rect 34748 30882 34804 30894
rect 34748 30830 34750 30882
rect 34802 30830 34804 30882
rect 34748 30324 34804 30830
rect 34748 30258 34804 30268
rect 34860 30098 34916 30110
rect 34860 30046 34862 30098
rect 34914 30046 34916 30098
rect 34636 29988 34692 29998
rect 34636 29894 34692 29932
rect 34860 29764 34916 30046
rect 34860 29698 34916 29708
rect 34860 29540 34916 29550
rect 34524 29486 34526 29538
rect 34578 29486 34580 29538
rect 34524 29428 34580 29486
rect 34524 29362 34580 29372
rect 34636 29538 34916 29540
rect 34636 29486 34862 29538
rect 34914 29486 34916 29538
rect 34636 29484 34916 29486
rect 34076 28354 34132 28364
rect 34636 28196 34692 29484
rect 34860 29474 34916 29484
rect 34972 28642 35028 32396
rect 35484 31388 35748 31398
rect 35540 31332 35588 31388
rect 35644 31332 35692 31388
rect 35484 31322 35748 31332
rect 35196 30994 35252 31006
rect 35196 30942 35198 30994
rect 35250 30942 35252 30994
rect 35084 30884 35140 30894
rect 35196 30884 35252 30942
rect 35140 30828 35252 30884
rect 35084 30818 35140 30828
rect 35084 30548 35140 30558
rect 35084 29764 35140 30492
rect 35196 29988 35252 29998
rect 35196 29986 35924 29988
rect 35196 29934 35198 29986
rect 35250 29934 35924 29986
rect 35196 29932 35924 29934
rect 35196 29922 35252 29932
rect 35484 29820 35748 29830
rect 35540 29764 35588 29820
rect 35644 29764 35692 29820
rect 35084 29708 35252 29764
rect 35484 29754 35748 29764
rect 35084 29428 35140 29438
rect 35084 29334 35140 29372
rect 34972 28590 34974 28642
rect 35026 28590 35028 28642
rect 34748 28420 34804 28430
rect 34748 28418 34916 28420
rect 34748 28366 34750 28418
rect 34802 28366 34916 28418
rect 34748 28364 34916 28366
rect 34748 28354 34804 28364
rect 33964 28140 34356 28196
rect 33404 27806 33406 27858
rect 33458 27806 33460 27858
rect 33180 26450 33236 26460
rect 33292 27746 33348 27758
rect 33292 27694 33294 27746
rect 33346 27694 33348 27746
rect 33180 26292 33236 26302
rect 33180 26066 33236 26236
rect 33180 26014 33182 26066
rect 33234 26014 33236 26066
rect 33068 25956 33124 25966
rect 32844 25396 32900 25406
rect 32844 25302 32900 25340
rect 33068 25394 33124 25900
rect 33180 25620 33236 26014
rect 33180 25554 33236 25564
rect 33068 25342 33070 25394
rect 33122 25342 33124 25394
rect 33068 25172 33124 25342
rect 33180 25394 33236 25406
rect 33180 25342 33182 25394
rect 33234 25342 33236 25394
rect 33180 25284 33236 25342
rect 33180 25218 33236 25228
rect 32956 25116 33124 25172
rect 32732 23874 32788 23884
rect 32844 24836 32900 24846
rect 32508 23660 32788 23716
rect 32284 23538 32340 23548
rect 32172 22316 32452 22372
rect 32060 22306 32116 22316
rect 32172 22148 32228 22158
rect 31836 21868 32004 21924
rect 31836 21476 31892 21486
rect 31836 21026 31892 21420
rect 31836 20974 31838 21026
rect 31890 20974 31892 21026
rect 31836 20962 31892 20974
rect 31724 20862 31726 20914
rect 31778 20862 31780 20914
rect 31724 20850 31780 20862
rect 31948 20690 32004 21868
rect 32060 21700 32116 21710
rect 32060 21606 32116 21644
rect 32172 21588 32228 22092
rect 32172 21522 32228 21532
rect 32284 22146 32340 22158
rect 32284 22094 32286 22146
rect 32338 22094 32340 22146
rect 32284 20804 32340 22094
rect 32396 21698 32452 22316
rect 32396 21646 32398 21698
rect 32450 21646 32452 21698
rect 32396 21252 32452 21646
rect 32508 21364 32564 21374
rect 32508 21270 32564 21308
rect 32396 21186 32452 21196
rect 32284 20738 32340 20748
rect 32732 20802 32788 23660
rect 32844 21140 32900 24780
rect 32956 24612 33012 25116
rect 32956 24546 33012 24556
rect 33068 24946 33124 24958
rect 33068 24894 33070 24946
rect 33122 24894 33124 24946
rect 33068 24050 33124 24894
rect 33180 24724 33236 24734
rect 33180 24630 33236 24668
rect 33068 23998 33070 24050
rect 33122 23998 33124 24050
rect 33068 23986 33124 23998
rect 33292 23828 33348 27694
rect 33404 26908 33460 27806
rect 34300 27858 34356 28140
rect 34636 28130 34692 28140
rect 34300 27806 34302 27858
rect 34354 27806 34356 27858
rect 33964 27746 34020 27758
rect 33964 27694 33966 27746
rect 34018 27694 34020 27746
rect 33964 26908 34020 27694
rect 33404 26852 33684 26908
rect 33964 26852 34132 26908
rect 33404 26068 33460 26078
rect 33404 26066 33572 26068
rect 33404 26014 33406 26066
rect 33458 26014 33572 26066
rect 33404 26012 33572 26014
rect 33404 26002 33460 26012
rect 33404 25620 33460 25630
rect 33404 25526 33460 25564
rect 33404 24612 33460 24622
rect 33516 24612 33572 26012
rect 33628 25732 33684 26852
rect 34076 26786 34132 26796
rect 34188 26740 34244 26750
rect 34188 26628 34244 26684
rect 34076 26572 34244 26628
rect 33964 26404 34020 26414
rect 33964 26310 34020 26348
rect 33740 26290 33796 26302
rect 33740 26238 33742 26290
rect 33794 26238 33796 26290
rect 33740 25956 33796 26238
rect 33740 25890 33796 25900
rect 33628 25676 33796 25732
rect 33628 25506 33684 25518
rect 33628 25454 33630 25506
rect 33682 25454 33684 25506
rect 33628 25172 33684 25454
rect 33628 25106 33684 25116
rect 33740 24948 33796 25676
rect 33460 24556 33572 24612
rect 33628 24892 33796 24948
rect 33404 24518 33460 24556
rect 32956 23772 33348 23828
rect 32956 21588 33012 23772
rect 33180 23604 33236 23614
rect 33236 23548 33460 23604
rect 33180 23538 33236 23548
rect 33292 23268 33348 23278
rect 33180 23154 33236 23166
rect 33180 23102 33182 23154
rect 33234 23102 33236 23154
rect 33068 22372 33124 22382
rect 33068 22278 33124 22316
rect 33068 21588 33124 21598
rect 32956 21586 33124 21588
rect 32956 21534 33070 21586
rect 33122 21534 33124 21586
rect 32956 21532 33124 21534
rect 33068 21522 33124 21532
rect 32844 21074 32900 21084
rect 32732 20750 32734 20802
rect 32786 20750 32788 20802
rect 32732 20738 32788 20750
rect 31948 20638 31950 20690
rect 32002 20638 32004 20690
rect 31948 20626 32004 20638
rect 32396 20580 32452 20590
rect 31612 20132 31668 20142
rect 31612 20038 31668 20076
rect 31836 20020 31892 20030
rect 31836 19926 31892 19964
rect 31948 20018 32004 20030
rect 31948 19966 31950 20018
rect 32002 19966 32004 20018
rect 31724 19906 31780 19918
rect 31724 19854 31726 19906
rect 31778 19854 31780 19906
rect 31200 19628 31464 19638
rect 31256 19572 31304 19628
rect 31360 19572 31408 19628
rect 31200 19562 31464 19572
rect 31500 19458 31556 19470
rect 31500 19406 31502 19458
rect 31554 19406 31556 19458
rect 30380 17714 30436 17724
rect 30716 18396 30996 18452
rect 31052 19124 31108 19134
rect 30156 17556 30212 17566
rect 30156 17462 30212 17500
rect 30268 17442 30324 17454
rect 30268 17390 30270 17442
rect 30322 17390 30324 17442
rect 30044 16884 30100 16894
rect 29932 16882 30212 16884
rect 29932 16830 30046 16882
rect 30098 16830 30212 16882
rect 29932 16828 30212 16830
rect 30044 16818 30100 16828
rect 29372 14868 29428 14878
rect 29372 12962 29428 14812
rect 29372 12910 29374 12962
rect 29426 12910 29428 12962
rect 29372 12898 29428 12910
rect 29484 12738 29540 16380
rect 29708 16380 29876 16436
rect 29708 15148 29764 16380
rect 30044 16324 30100 16334
rect 29484 12686 29486 12738
rect 29538 12686 29540 12738
rect 29484 12674 29540 12686
rect 29596 15092 29764 15148
rect 29820 15202 29876 15214
rect 29820 15150 29822 15202
rect 29874 15150 29876 15202
rect 29596 11732 29652 15092
rect 29708 13748 29764 13758
rect 29820 13748 29876 15150
rect 29932 14418 29988 14430
rect 29932 14366 29934 14418
rect 29986 14366 29988 14418
rect 29932 14308 29988 14366
rect 29932 14242 29988 14252
rect 29708 13746 29876 13748
rect 29708 13694 29710 13746
rect 29762 13694 29876 13746
rect 29708 13692 29876 13694
rect 29708 13636 29764 13692
rect 29708 13570 29764 13580
rect 29708 13076 29764 13086
rect 29708 12962 29764 13020
rect 29708 12910 29710 12962
rect 29762 12910 29764 12962
rect 29708 12898 29764 12910
rect 30044 12962 30100 16268
rect 30156 14980 30212 16828
rect 30268 16324 30324 17390
rect 30380 17442 30436 17454
rect 30380 17390 30382 17442
rect 30434 17390 30436 17442
rect 30380 16548 30436 17390
rect 30716 17220 30772 18396
rect 30828 18228 30884 18238
rect 30828 17778 30884 18172
rect 30940 17892 30996 17902
rect 30940 17798 30996 17836
rect 30828 17726 30830 17778
rect 30882 17726 30884 17778
rect 30828 17714 30884 17726
rect 30716 17106 30772 17164
rect 30716 17054 30718 17106
rect 30770 17054 30772 17106
rect 30716 17042 30772 17054
rect 31052 16996 31108 19068
rect 31388 19122 31444 19134
rect 31388 19070 31390 19122
rect 31442 19070 31444 19122
rect 31388 18562 31444 19070
rect 31500 18788 31556 19406
rect 31500 18722 31556 18732
rect 31388 18510 31390 18562
rect 31442 18510 31444 18562
rect 31388 18498 31444 18510
rect 31724 18338 31780 19854
rect 31948 18564 32004 19966
rect 32284 19796 32340 19806
rect 32284 19702 32340 19740
rect 32284 19348 32340 19358
rect 32284 19254 32340 19292
rect 32396 19234 32452 20524
rect 33068 20132 33124 20142
rect 33068 20038 33124 20076
rect 33180 20130 33236 23102
rect 33180 20078 33182 20130
rect 33234 20078 33236 20130
rect 33180 20066 33236 20078
rect 33292 21924 33348 23212
rect 32396 19182 32398 19234
rect 32450 19182 32452 19234
rect 32396 19170 32452 19182
rect 32508 19794 32564 19806
rect 32508 19742 32510 19794
rect 32562 19742 32564 19794
rect 31948 18498 32004 18508
rect 31836 18452 31892 18462
rect 31836 18358 31892 18396
rect 32172 18450 32228 18462
rect 32172 18398 32174 18450
rect 32226 18398 32228 18450
rect 31724 18286 31726 18338
rect 31778 18286 31780 18338
rect 31724 18274 31780 18286
rect 31200 18060 31464 18070
rect 31256 18004 31304 18060
rect 31360 18004 31408 18060
rect 31200 17994 31464 18004
rect 32172 17892 32228 18398
rect 32508 18004 32564 19742
rect 33180 18562 33236 18574
rect 33180 18510 33182 18562
rect 33234 18510 33236 18562
rect 33068 18340 33124 18350
rect 32508 17938 32564 17948
rect 32956 18338 33124 18340
rect 32956 18286 33070 18338
rect 33122 18286 33124 18338
rect 32956 18284 33124 18286
rect 32172 17826 32228 17836
rect 31276 17780 31332 17790
rect 31276 17686 31332 17724
rect 32284 17780 32340 17790
rect 32284 17778 32900 17780
rect 32284 17726 32286 17778
rect 32338 17726 32900 17778
rect 32284 17724 32900 17726
rect 32284 17714 32340 17724
rect 31724 17666 31780 17678
rect 31724 17614 31726 17666
rect 31778 17614 31780 17666
rect 31724 17444 31780 17614
rect 31724 17378 31780 17388
rect 32620 17444 32676 17454
rect 30828 16940 31108 16996
rect 32172 16994 32228 17006
rect 32172 16942 32174 16994
rect 32226 16942 32228 16994
rect 30716 16772 30772 16782
rect 30716 16548 30772 16716
rect 30828 16770 30884 16940
rect 31724 16882 31780 16894
rect 31724 16830 31726 16882
rect 31778 16830 31780 16882
rect 30828 16718 30830 16770
rect 30882 16718 30884 16770
rect 30828 16706 30884 16718
rect 30940 16772 30996 16782
rect 30940 16678 30996 16716
rect 31276 16770 31332 16782
rect 31276 16718 31278 16770
rect 31330 16718 31332 16770
rect 31276 16660 31332 16718
rect 31052 16604 31332 16660
rect 31052 16548 31108 16604
rect 30716 16492 31108 16548
rect 31200 16492 31464 16502
rect 30380 16482 30436 16492
rect 31256 16436 31304 16492
rect 31360 16436 31408 16492
rect 31200 16426 31464 16436
rect 30268 16268 30660 16324
rect 30492 15314 30548 15326
rect 30492 15262 30494 15314
rect 30546 15262 30548 15314
rect 30492 15092 30548 15262
rect 30492 15026 30548 15036
rect 30156 14914 30212 14924
rect 30380 13634 30436 13646
rect 30380 13582 30382 13634
rect 30434 13582 30436 13634
rect 30044 12910 30046 12962
rect 30098 12910 30100 12962
rect 30044 12898 30100 12910
rect 30268 12964 30324 12974
rect 30268 12870 30324 12908
rect 29932 12740 29988 12750
rect 29260 9998 29262 10050
rect 29314 9998 29316 10050
rect 29260 9986 29316 9998
rect 29372 11676 29652 11732
rect 29820 12684 29932 12740
rect 29372 9044 29428 11676
rect 29596 11506 29652 11518
rect 29596 11454 29598 11506
rect 29650 11454 29652 11506
rect 29596 10724 29652 11454
rect 29596 10658 29652 10668
rect 29708 10724 29764 10734
rect 29820 10724 29876 12684
rect 29932 12674 29988 12684
rect 30380 12292 30436 13582
rect 30492 13074 30548 13086
rect 30492 13022 30494 13074
rect 30546 13022 30548 13074
rect 30492 12740 30548 13022
rect 30604 12962 30660 16268
rect 31500 15988 31556 15998
rect 30604 12910 30606 12962
rect 30658 12910 30660 12962
rect 30604 12898 30660 12910
rect 30828 15986 31556 15988
rect 30828 15934 31502 15986
rect 31554 15934 31556 15986
rect 30828 15932 31556 15934
rect 30828 12740 30884 15932
rect 31500 15922 31556 15932
rect 31724 15988 31780 16830
rect 32172 16660 32228 16942
rect 32396 16884 32452 16894
rect 32396 16790 32452 16828
rect 32172 16594 32228 16604
rect 32172 16100 32228 16110
rect 31500 15202 31556 15214
rect 31500 15150 31502 15202
rect 31554 15150 31556 15202
rect 31500 15148 31556 15150
rect 31500 15092 31668 15148
rect 31500 15026 31556 15036
rect 31200 14924 31464 14934
rect 31256 14868 31304 14924
rect 31360 14868 31408 14924
rect 31200 14858 31464 14868
rect 30940 14530 30996 14542
rect 30940 14478 30942 14530
rect 30994 14478 30996 14530
rect 30940 13636 30996 14478
rect 30940 13570 30996 13580
rect 31052 14308 31108 14318
rect 30492 12684 30884 12740
rect 30940 12740 30996 12750
rect 30940 12646 30996 12684
rect 30380 12226 30436 12236
rect 29708 10722 29876 10724
rect 29708 10670 29710 10722
rect 29762 10670 29876 10722
rect 29708 10668 29876 10670
rect 30044 12066 30100 12078
rect 30044 12014 30046 12066
rect 30098 12014 30100 12066
rect 30044 11394 30100 12014
rect 31052 11732 31108 14252
rect 31612 13860 31668 15092
rect 31724 14754 31780 15932
rect 32060 16098 32228 16100
rect 32060 16046 32174 16098
rect 32226 16046 32228 16098
rect 32060 16044 32228 16046
rect 31724 14702 31726 14754
rect 31778 14702 31780 14754
rect 31724 14690 31780 14702
rect 31836 15316 31892 15326
rect 32060 15316 32116 16044
rect 32172 16034 32228 16044
rect 32620 15540 32676 17388
rect 32844 16436 32900 17724
rect 32956 16548 33012 18284
rect 33068 18274 33124 18284
rect 33180 17892 33236 18510
rect 33180 17826 33236 17836
rect 33292 17668 33348 21868
rect 33068 17612 33348 17668
rect 33404 18450 33460 23548
rect 33628 23268 33684 24892
rect 33740 24722 33796 24734
rect 33740 24670 33742 24722
rect 33794 24670 33796 24722
rect 33740 24500 33796 24670
rect 33740 24434 33796 24444
rect 33964 24500 34020 24510
rect 33964 24406 34020 24444
rect 33852 24388 33908 24398
rect 33628 23212 33796 23268
rect 33628 23044 33684 23054
rect 33628 22950 33684 22988
rect 33628 21588 33684 21598
rect 33628 21494 33684 21532
rect 33740 20018 33796 23212
rect 33852 23044 33908 24332
rect 33964 23044 34020 23054
rect 33852 23042 34020 23044
rect 33852 22990 33966 23042
rect 34018 22990 34020 23042
rect 33852 22988 34020 22990
rect 33964 22978 34020 22988
rect 34076 21700 34132 26572
rect 34300 26516 34356 27806
rect 34412 28084 34468 28094
rect 34412 27860 34468 28028
rect 34748 28084 34804 28094
rect 34748 27990 34804 28028
rect 34412 26908 34468 27804
rect 34412 26852 34804 26908
rect 34188 26460 34356 26516
rect 34188 25844 34244 26460
rect 34412 26404 34468 26414
rect 34412 26310 34468 26348
rect 34524 26404 34580 26414
rect 34524 26402 34692 26404
rect 34524 26350 34526 26402
rect 34578 26350 34692 26402
rect 34524 26348 34692 26350
rect 34524 26338 34580 26348
rect 34300 26292 34356 26302
rect 34300 26198 34356 26236
rect 34188 25778 34244 25788
rect 34188 25284 34244 25322
rect 34524 25284 34580 25294
rect 34188 25218 34244 25228
rect 34300 25282 34580 25284
rect 34300 25230 34526 25282
rect 34578 25230 34580 25282
rect 34300 25228 34580 25230
rect 34188 24948 34244 24958
rect 34188 23380 34244 24892
rect 34188 23314 34244 23324
rect 34300 24946 34356 25228
rect 34524 25218 34580 25228
rect 34300 24894 34302 24946
rect 34354 24894 34356 24946
rect 34188 23154 34244 23166
rect 34188 23102 34190 23154
rect 34242 23102 34244 23154
rect 34188 22148 34244 23102
rect 34300 22932 34356 24894
rect 34524 24836 34580 24846
rect 34636 24836 34692 26348
rect 34300 22866 34356 22876
rect 34412 24834 34692 24836
rect 34412 24782 34526 24834
rect 34578 24782 34692 24834
rect 34412 24780 34692 24782
rect 34748 26290 34804 26852
rect 34860 26740 34916 28364
rect 34860 26674 34916 26684
rect 34972 26516 35028 28590
rect 35084 28084 35140 28094
rect 35196 28084 35252 29708
rect 35484 28252 35748 28262
rect 35540 28196 35588 28252
rect 35644 28196 35692 28252
rect 35484 28186 35748 28196
rect 35140 28028 35252 28084
rect 35084 28018 35140 28028
rect 35084 27860 35140 27870
rect 35084 27766 35140 27804
rect 35196 27186 35252 27198
rect 35196 27134 35198 27186
rect 35250 27134 35252 27186
rect 34972 26450 35028 26460
rect 35084 26852 35140 26862
rect 34748 26238 34750 26290
rect 34802 26238 34804 26290
rect 34412 24612 34468 24780
rect 34524 24770 34580 24780
rect 34748 24722 34804 26238
rect 34860 26404 34916 26414
rect 34860 25732 34916 26348
rect 34860 25666 34916 25676
rect 34972 25618 35028 25630
rect 34972 25566 34974 25618
rect 35026 25566 35028 25618
rect 34972 25396 35028 25566
rect 34748 24670 34750 24722
rect 34802 24670 34804 24722
rect 34748 24658 34804 24670
rect 34860 25340 35028 25396
rect 34860 24724 34916 25340
rect 35084 24948 35140 26796
rect 35196 26404 35252 27134
rect 35484 26684 35748 26694
rect 35540 26628 35588 26684
rect 35644 26628 35692 26684
rect 35484 26618 35748 26628
rect 35196 26338 35252 26348
rect 35484 25116 35748 25126
rect 35540 25060 35588 25116
rect 35644 25060 35692 25116
rect 35484 25050 35748 25060
rect 35084 24892 35252 24948
rect 34860 24658 34916 24668
rect 35084 24722 35140 24734
rect 35084 24670 35086 24722
rect 35138 24670 35140 24722
rect 34412 22484 34468 24556
rect 34636 24610 34692 24622
rect 34636 24558 34638 24610
rect 34690 24558 34692 24610
rect 34636 24500 34692 24558
rect 34636 24434 34692 24444
rect 35084 24052 35140 24670
rect 35196 24276 35252 24892
rect 35196 24220 35364 24276
rect 35196 24052 35252 24062
rect 35084 24050 35252 24052
rect 35084 23998 35198 24050
rect 35250 23998 35252 24050
rect 35084 23996 35252 23998
rect 35196 23268 35252 23996
rect 34412 22418 34468 22428
rect 34524 23212 35252 23268
rect 34300 22148 34356 22158
rect 34188 22092 34300 22148
rect 34300 22082 34356 22092
rect 34076 21588 34132 21644
rect 34412 21924 34468 21934
rect 34412 21698 34468 21868
rect 34412 21646 34414 21698
rect 34466 21646 34468 21698
rect 34412 21634 34468 21646
rect 34076 21532 34356 21588
rect 33964 21476 34020 21486
rect 33964 21382 34020 21420
rect 33740 19966 33742 20018
rect 33794 19966 33796 20018
rect 33628 19794 33684 19806
rect 33628 19742 33630 19794
rect 33682 19742 33684 19794
rect 33628 18676 33684 19742
rect 33404 18398 33406 18450
rect 33458 18398 33460 18450
rect 33404 18116 33460 18398
rect 33516 18620 33684 18676
rect 33516 18340 33572 18620
rect 33516 18274 33572 18284
rect 33404 17668 33460 18060
rect 33068 16882 33124 17612
rect 33404 17602 33460 17612
rect 33628 17556 33684 17566
rect 33068 16830 33070 16882
rect 33122 16830 33124 16882
rect 33068 16818 33124 16830
rect 33516 17332 33572 17342
rect 33516 16882 33572 17276
rect 33516 16830 33518 16882
rect 33570 16830 33572 16882
rect 33516 16818 33572 16830
rect 32956 16492 33236 16548
rect 32844 16380 33124 16436
rect 33068 16322 33124 16380
rect 33068 16270 33070 16322
rect 33122 16270 33124 16322
rect 33068 16258 33124 16270
rect 32732 16100 32788 16110
rect 33180 16100 33236 16492
rect 32732 16006 32788 16044
rect 32956 16044 33236 16100
rect 31836 15314 32116 15316
rect 31836 15262 31838 15314
rect 31890 15262 32116 15314
rect 31836 15260 32116 15262
rect 32172 15260 32564 15316
rect 31836 14308 31892 15260
rect 32172 15148 32228 15260
rect 32508 15202 32564 15260
rect 32508 15150 32510 15202
rect 32562 15150 32564 15202
rect 32508 15138 32564 15150
rect 32172 15082 32228 15092
rect 32396 15090 32452 15102
rect 32396 15038 32398 15090
rect 32450 15038 32452 15090
rect 31836 14242 31892 14252
rect 31948 14868 32004 14878
rect 31612 13794 31668 13804
rect 31724 13524 31780 13534
rect 31200 13356 31464 13366
rect 31256 13300 31304 13356
rect 31360 13300 31408 13356
rect 31200 13290 31464 13300
rect 31164 13188 31220 13198
rect 31164 12962 31220 13132
rect 31724 13186 31780 13468
rect 31724 13134 31726 13186
rect 31778 13134 31780 13186
rect 31724 13122 31780 13134
rect 31948 13076 32004 14812
rect 32396 14868 32452 15038
rect 32396 14802 32452 14812
rect 32620 14868 32676 15484
rect 32620 14802 32676 14812
rect 32732 15092 32788 15102
rect 32172 14756 32228 14766
rect 31948 13010 32004 13020
rect 32060 14532 32116 14542
rect 31164 12910 31166 12962
rect 31218 12910 31220 12962
rect 31164 12898 31220 12910
rect 31836 12850 31892 12862
rect 31836 12798 31838 12850
rect 31890 12798 31892 12850
rect 31724 12738 31780 12750
rect 31724 12686 31726 12738
rect 31778 12686 31780 12738
rect 31724 11956 31780 12686
rect 31836 12628 31892 12798
rect 31836 12562 31892 12572
rect 32060 12402 32116 14476
rect 32060 12350 32062 12402
rect 32114 12350 32116 12402
rect 32060 12338 32116 12350
rect 32172 12404 32228 14700
rect 32284 14644 32340 14654
rect 32732 14644 32788 15036
rect 32284 14642 32788 14644
rect 32284 14590 32286 14642
rect 32338 14590 32788 14642
rect 32284 14588 32788 14590
rect 32284 14578 32340 14588
rect 32508 13634 32564 13646
rect 32508 13582 32510 13634
rect 32562 13582 32564 13634
rect 32396 13524 32452 13534
rect 32284 13468 32396 13524
rect 32284 13074 32340 13468
rect 32396 13458 32452 13468
rect 32284 13022 32286 13074
rect 32338 13022 32340 13074
rect 32284 13010 32340 13022
rect 32284 12404 32340 12414
rect 32172 12402 32340 12404
rect 32172 12350 32286 12402
rect 32338 12350 32340 12402
rect 32172 12348 32340 12350
rect 32284 12338 32340 12348
rect 31724 11890 31780 11900
rect 32396 12178 32452 12190
rect 32396 12126 32398 12178
rect 32450 12126 32452 12178
rect 30044 11342 30046 11394
rect 30098 11342 30100 11394
rect 29708 10658 29764 10668
rect 29820 10500 29876 10510
rect 29484 10050 29540 10062
rect 29484 9998 29486 10050
rect 29538 9998 29540 10050
rect 29484 9938 29540 9998
rect 29484 9886 29486 9938
rect 29538 9886 29540 9938
rect 29484 9874 29540 9886
rect 29820 9826 29876 10444
rect 29820 9774 29822 9826
rect 29874 9774 29876 9826
rect 29820 9762 29876 9774
rect 29932 9716 29988 9754
rect 29932 9650 29988 9660
rect 29932 9492 29988 9502
rect 29372 8988 29540 9044
rect 28924 7634 28980 7644
rect 29372 8820 29428 8830
rect 29372 7700 29428 8764
rect 29484 8484 29540 8988
rect 29484 8418 29540 8428
rect 29932 8370 29988 9436
rect 29932 8318 29934 8370
rect 29986 8318 29988 8370
rect 29932 8306 29988 8318
rect 30044 9044 30100 11342
rect 30940 11676 31108 11732
rect 31200 11788 31464 11798
rect 31256 11732 31304 11788
rect 31360 11732 31408 11788
rect 31200 11722 31464 11732
rect 30828 11284 30884 11294
rect 30156 11282 30884 11284
rect 30156 11230 30830 11282
rect 30882 11230 30884 11282
rect 30156 11228 30884 11230
rect 30156 9938 30212 11228
rect 30828 11218 30884 11228
rect 30940 11060 30996 11676
rect 32396 11620 32452 12126
rect 32508 11956 32564 13582
rect 32508 11890 32564 11900
rect 32396 11554 32452 11564
rect 32732 11620 32788 11630
rect 30492 11004 30996 11060
rect 31052 11508 31108 11518
rect 30492 10610 30548 11004
rect 31052 10834 31108 11452
rect 31052 10782 31054 10834
rect 31106 10782 31108 10834
rect 31052 10770 31108 10782
rect 31276 11396 31332 11406
rect 31276 10834 31332 11340
rect 31276 10782 31278 10834
rect 31330 10782 31332 10834
rect 31276 10770 31332 10782
rect 32284 11396 32340 11406
rect 32284 10834 32340 11340
rect 32284 10782 32286 10834
rect 32338 10782 32340 10834
rect 32284 10770 32340 10782
rect 32620 10836 32676 10846
rect 30492 10558 30494 10610
rect 30546 10558 30548 10610
rect 30492 10546 30548 10558
rect 30828 10724 30884 10734
rect 30828 10052 30884 10668
rect 31836 10724 31892 10734
rect 31836 10630 31892 10668
rect 30940 10500 30996 10510
rect 30940 10406 30996 10444
rect 31200 10220 31464 10230
rect 31256 10164 31304 10220
rect 31360 10164 31408 10220
rect 31200 10154 31464 10164
rect 30828 9996 31108 10052
rect 30156 9886 30158 9938
rect 30210 9886 30212 9938
rect 30156 9874 30212 9886
rect 30380 9828 30436 9838
rect 30380 9826 30548 9828
rect 30380 9774 30382 9826
rect 30434 9774 30548 9826
rect 30380 9772 30548 9774
rect 30380 9762 30436 9772
rect 30492 9268 30548 9772
rect 30828 9826 30884 9838
rect 30828 9774 30830 9826
rect 30882 9774 30884 9826
rect 30604 9714 30660 9726
rect 30604 9662 30606 9714
rect 30658 9662 30660 9714
rect 30604 9492 30660 9662
rect 30828 9716 30884 9774
rect 30716 9604 30772 9614
rect 30716 9510 30772 9548
rect 30604 9426 30660 9436
rect 30604 9268 30660 9278
rect 30492 9266 30660 9268
rect 30492 9214 30606 9266
rect 30658 9214 30660 9266
rect 30492 9212 30660 9214
rect 30604 9202 30660 9212
rect 30380 9044 30436 9054
rect 30044 8372 30100 8988
rect 30156 8988 30380 9044
rect 30156 8930 30212 8988
rect 30380 8978 30436 8988
rect 30492 9042 30548 9054
rect 30492 8990 30494 9042
rect 30546 8990 30548 9042
rect 30156 8878 30158 8930
rect 30210 8878 30212 8930
rect 30156 8866 30212 8878
rect 30492 8372 30548 8990
rect 30716 9044 30772 9054
rect 30716 8950 30772 8988
rect 30828 8708 30884 9660
rect 31052 9380 31108 9996
rect 31164 9716 31220 9726
rect 31164 9714 31556 9716
rect 31164 9662 31166 9714
rect 31218 9662 31556 9714
rect 31164 9660 31556 9662
rect 31164 9650 31220 9660
rect 31052 9324 31444 9380
rect 31388 9266 31444 9324
rect 31388 9214 31390 9266
rect 31442 9214 31444 9266
rect 31164 9042 31220 9054
rect 31164 8990 31166 9042
rect 31218 8990 31220 9042
rect 31164 8820 31220 8990
rect 31388 8820 31444 9214
rect 31500 9266 31556 9660
rect 31500 9214 31502 9266
rect 31554 9214 31556 9266
rect 31500 9202 31556 9214
rect 32396 9156 32452 9166
rect 32396 9062 32452 9100
rect 31612 9044 31668 9054
rect 31612 8950 31668 8988
rect 31948 9042 32004 9054
rect 31948 8990 31950 9042
rect 32002 8990 32004 9042
rect 31388 8764 31668 8820
rect 31164 8754 31220 8764
rect 30828 8652 31108 8708
rect 30044 8306 30100 8316
rect 30156 8316 30548 8372
rect 29820 8260 29876 8270
rect 29820 8166 29876 8204
rect 30044 8148 30100 8158
rect 30156 8148 30212 8316
rect 30716 8260 30772 8270
rect 30716 8166 30772 8204
rect 29932 8146 30212 8148
rect 29932 8094 30046 8146
rect 30098 8094 30212 8146
rect 29932 8092 30212 8094
rect 29372 7606 29428 7644
rect 29596 8034 29652 8046
rect 29596 7982 29598 8034
rect 29650 7982 29652 8034
rect 29596 7698 29652 7982
rect 29932 8036 29988 8092
rect 30044 8082 30100 8092
rect 29596 7646 29598 7698
rect 29650 7646 29652 7698
rect 29596 7634 29652 7646
rect 29820 7700 29876 7710
rect 29932 7700 29988 7980
rect 30492 8034 30548 8046
rect 30492 7982 30494 8034
rect 30546 7982 30548 8034
rect 30492 7924 30548 7982
rect 30492 7858 30548 7868
rect 30828 8034 30884 8046
rect 30828 7982 30830 8034
rect 30882 7982 30884 8034
rect 29820 7698 29988 7700
rect 29820 7646 29822 7698
rect 29874 7646 29988 7698
rect 29820 7644 29988 7646
rect 29260 7588 29316 7598
rect 28812 7474 28868 7486
rect 28812 7422 28814 7474
rect 28866 7422 28868 7474
rect 28812 6692 28868 7422
rect 29260 7474 29316 7532
rect 29260 7422 29262 7474
rect 29314 7422 29316 7474
rect 29260 7364 29316 7422
rect 29260 7308 29540 7364
rect 29260 6916 29316 6926
rect 29036 6692 29092 6702
rect 28812 6690 29092 6692
rect 28812 6638 29038 6690
rect 29090 6638 29092 6690
rect 28812 6636 29092 6638
rect 29036 6626 29092 6636
rect 29036 5908 29092 5918
rect 28700 5906 29092 5908
rect 28700 5854 29038 5906
rect 29090 5854 29092 5906
rect 28700 5852 29092 5854
rect 28588 5182 28590 5234
rect 28642 5182 28644 5234
rect 28588 5170 28644 5182
rect 29036 5012 29092 5852
rect 29260 5346 29316 6860
rect 29484 6804 29540 7308
rect 29820 6916 29876 7644
rect 30044 7588 30100 7598
rect 30044 7494 30100 7532
rect 30268 7586 30324 7598
rect 30268 7534 30270 7586
rect 30322 7534 30324 7586
rect 29932 7476 29988 7486
rect 29932 7382 29988 7420
rect 29820 6860 30100 6916
rect 29484 6738 29540 6748
rect 29596 6692 29652 6702
rect 29932 6692 29988 6702
rect 29596 6690 29988 6692
rect 29596 6638 29598 6690
rect 29650 6638 29934 6690
rect 29986 6638 29988 6690
rect 29596 6636 29988 6638
rect 29596 6626 29652 6636
rect 29932 6626 29988 6636
rect 29484 6468 29540 6478
rect 29484 6374 29540 6412
rect 29708 6468 29764 6478
rect 30044 6468 30100 6860
rect 29708 6466 30100 6468
rect 29708 6414 29710 6466
rect 29762 6414 30100 6466
rect 29708 6412 30100 6414
rect 30156 6466 30212 6478
rect 30156 6414 30158 6466
rect 30210 6414 30212 6466
rect 29708 6402 29764 6412
rect 30156 6132 30212 6414
rect 30268 6468 30324 7534
rect 30828 7474 30884 7982
rect 30940 8036 30996 8046
rect 30940 7942 30996 7980
rect 30828 7422 30830 7474
rect 30882 7422 30884 7474
rect 30828 7410 30884 7422
rect 31052 7474 31108 8652
rect 31200 8652 31464 8662
rect 31256 8596 31304 8652
rect 31360 8596 31408 8652
rect 31200 8586 31464 8596
rect 31276 8372 31332 8382
rect 31276 8258 31332 8316
rect 31276 8206 31278 8258
rect 31330 8206 31332 8258
rect 31276 8194 31332 8206
rect 31164 8148 31220 8158
rect 31164 7698 31220 8092
rect 31164 7646 31166 7698
rect 31218 7646 31220 7698
rect 31164 7634 31220 7646
rect 31612 8036 31668 8764
rect 31612 7698 31668 7980
rect 31948 7924 32004 8990
rect 32284 9042 32340 9054
rect 32284 8990 32286 9042
rect 32338 8990 32340 9042
rect 32060 8148 32116 8158
rect 32060 8054 32116 8092
rect 32060 7924 32116 7934
rect 31948 7868 32060 7924
rect 31612 7646 31614 7698
rect 31666 7646 31668 7698
rect 31612 7634 31668 7646
rect 32060 7698 32116 7868
rect 32060 7646 32062 7698
rect 32114 7646 32116 7698
rect 32060 7634 32116 7646
rect 32172 7700 32228 7710
rect 31836 7588 31892 7598
rect 31892 7532 32004 7588
rect 31836 7494 31892 7532
rect 31052 7422 31054 7474
rect 31106 7422 31108 7474
rect 31052 7028 31108 7422
rect 31276 7476 31332 7486
rect 31276 7382 31332 7420
rect 31724 7362 31780 7374
rect 31724 7310 31726 7362
rect 31778 7310 31780 7362
rect 30380 6972 31108 7028
rect 31200 7084 31464 7094
rect 31256 7028 31304 7084
rect 31360 7028 31408 7084
rect 31200 7018 31464 7028
rect 30380 6690 30436 6972
rect 31724 6916 31780 7310
rect 30380 6638 30382 6690
rect 30434 6638 30436 6690
rect 30380 6626 30436 6638
rect 30604 6860 31780 6916
rect 30604 6690 30660 6860
rect 30604 6638 30606 6690
rect 30658 6638 30660 6690
rect 30604 6626 30660 6638
rect 31164 6692 31220 6702
rect 31164 6598 31220 6636
rect 30828 6468 30884 6478
rect 30268 6466 30884 6468
rect 30268 6414 30830 6466
rect 30882 6414 30884 6466
rect 30268 6412 30884 6414
rect 30828 6402 30884 6412
rect 31052 6466 31108 6478
rect 31052 6414 31054 6466
rect 31106 6414 31108 6466
rect 29820 6076 30212 6132
rect 29820 6018 29876 6076
rect 29820 5966 29822 6018
rect 29874 5966 29876 6018
rect 29820 5954 29876 5966
rect 31052 5796 31108 6414
rect 31052 5730 31108 5740
rect 31724 5796 31780 5806
rect 31200 5516 31464 5526
rect 31256 5460 31304 5516
rect 31360 5460 31408 5516
rect 31200 5450 31464 5460
rect 29260 5294 29262 5346
rect 29314 5294 29316 5346
rect 29260 5282 29316 5294
rect 28924 4452 28980 4462
rect 28476 4228 28532 4238
rect 28364 4226 28532 4228
rect 28364 4174 28478 4226
rect 28530 4174 28532 4226
rect 28364 4172 28532 4174
rect 27244 3892 27300 3902
rect 25564 3668 25620 3678
rect 25564 3574 25620 3612
rect 24780 3502 24782 3554
rect 24834 3502 24836 3554
rect 24780 3490 24836 3502
rect 23996 3390 23998 3442
rect 24050 3390 24052 3442
rect 23996 3378 24052 3390
rect 25340 3444 25396 3454
rect 25340 800 25396 3388
rect 26916 3164 27180 3174
rect 26972 3108 27020 3164
rect 27076 3108 27124 3164
rect 26916 3098 27180 3108
rect 27244 2772 27300 3836
rect 27468 3442 27524 4172
rect 28140 4162 28196 4172
rect 28476 4162 28532 4172
rect 28700 3892 28756 3902
rect 28364 3780 28420 3790
rect 27468 3390 27470 3442
rect 27522 3390 27524 3442
rect 27468 3378 27524 3390
rect 27804 3444 27860 3482
rect 27804 3378 27860 3388
rect 28364 3442 28420 3724
rect 28364 3390 28366 3442
rect 28418 3390 28420 3442
rect 28364 3378 28420 3390
rect 28476 3556 28532 3566
rect 26908 2716 27300 2772
rect 26908 800 26964 2716
rect 28476 800 28532 3500
rect 28700 3554 28756 3836
rect 28700 3502 28702 3554
rect 28754 3502 28756 3554
rect 28700 3490 28756 3502
rect 28924 3444 28980 4396
rect 29036 4340 29092 4956
rect 29036 4274 29092 4284
rect 29372 5010 29428 5022
rect 29372 4958 29374 5010
rect 29426 4958 29428 5010
rect 29372 4228 29428 4958
rect 31276 5012 31332 5022
rect 29372 4162 29428 4172
rect 29820 4898 29876 4910
rect 29820 4846 29822 4898
rect 29874 4846 29876 4898
rect 29820 3892 29876 4846
rect 30604 4900 30660 4910
rect 30604 4450 30660 4844
rect 30604 4398 30606 4450
rect 30658 4398 30660 4450
rect 30604 4386 30660 4398
rect 31276 4338 31332 4956
rect 31724 4562 31780 5740
rect 31948 5794 32004 7532
rect 31948 5742 31950 5794
rect 32002 5742 32004 5794
rect 31948 5730 32004 5742
rect 31724 4510 31726 4562
rect 31778 4510 31780 4562
rect 31724 4498 31780 4510
rect 32172 4562 32228 7644
rect 32284 6804 32340 8990
rect 32396 8820 32452 8830
rect 32396 8726 32452 8764
rect 32284 6738 32340 6748
rect 32172 4510 32174 4562
rect 32226 4510 32228 4562
rect 32172 4498 32228 4510
rect 31276 4286 31278 4338
rect 31330 4286 31332 4338
rect 31276 4274 31332 4286
rect 29820 3826 29876 3836
rect 30268 4228 30324 4238
rect 29372 3556 29428 3566
rect 29372 3462 29428 3500
rect 29036 3444 29092 3454
rect 28924 3442 29092 3444
rect 28924 3390 29038 3442
rect 29090 3390 29092 3442
rect 28924 3388 29092 3390
rect 29036 3378 29092 3388
rect 29820 3444 29876 3482
rect 29820 3378 29876 3388
rect 30044 3444 30100 3454
rect 30044 800 30100 3388
rect 30268 3442 30324 4172
rect 31836 4228 31892 4238
rect 31836 4226 32116 4228
rect 31836 4174 31838 4226
rect 31890 4174 32116 4226
rect 31836 4172 32116 4174
rect 31836 4162 31892 4172
rect 31200 3948 31464 3958
rect 31256 3892 31304 3948
rect 31360 3892 31408 3948
rect 31200 3882 31464 3892
rect 31052 3556 31108 3566
rect 30268 3390 30270 3442
rect 30322 3390 30324 3442
rect 30268 3378 30324 3390
rect 30604 3444 30660 3482
rect 31052 3462 31108 3500
rect 31612 3556 31668 3566
rect 30604 3378 30660 3388
rect 31500 3444 31556 3482
rect 31500 3378 31556 3388
rect 31612 800 31668 3500
rect 32060 3444 32116 4172
rect 32284 4226 32340 4238
rect 32284 4174 32286 4226
rect 32338 4174 32340 4226
rect 32172 3444 32228 3454
rect 32060 3442 32228 3444
rect 32060 3390 32174 3442
rect 32226 3390 32228 3442
rect 32060 3388 32228 3390
rect 32172 3378 32228 3388
rect 32284 3332 32340 4174
rect 32396 3556 32452 3566
rect 32396 3462 32452 3500
rect 32284 3266 32340 3276
rect 32620 2324 32676 10780
rect 32732 9938 32788 11564
rect 32956 11508 33012 16044
rect 33292 15988 33348 15998
rect 33292 15894 33348 15932
rect 33628 15986 33684 17500
rect 33740 16884 33796 19966
rect 34076 21364 34132 21374
rect 34076 20018 34132 21308
rect 34076 19966 34078 20018
rect 34130 19966 34132 20018
rect 33852 19796 33908 19806
rect 33908 19740 34020 19796
rect 33852 19730 33908 19740
rect 33852 19012 33908 19022
rect 33852 18450 33908 18956
rect 33964 18676 34020 19740
rect 34076 19012 34132 19966
rect 34300 19908 34356 21532
rect 34412 20132 34468 20142
rect 34524 20132 34580 23212
rect 35196 23044 35252 23054
rect 35196 22950 35252 22988
rect 35084 22932 35140 22942
rect 34636 22930 35140 22932
rect 34636 22878 35086 22930
rect 35138 22878 35140 22930
rect 34636 22876 35140 22878
rect 34636 21586 34692 22876
rect 35084 22866 35140 22876
rect 35308 22820 35364 24220
rect 35484 23548 35748 23558
rect 35540 23492 35588 23548
rect 35644 23492 35692 23548
rect 35484 23482 35748 23492
rect 35196 22764 35364 22820
rect 34636 21534 34638 21586
rect 34690 21534 34692 21586
rect 34636 21522 34692 21534
rect 34748 22596 34804 22606
rect 34748 21252 34804 22540
rect 34972 22596 35028 22606
rect 34972 22502 35028 22540
rect 34860 22484 34916 22494
rect 34860 21810 34916 22428
rect 34860 21758 34862 21810
rect 34914 21758 34916 21810
rect 34860 21746 34916 21758
rect 35196 21812 35252 22764
rect 35484 21980 35748 21990
rect 35540 21924 35588 21980
rect 35644 21924 35692 21980
rect 35484 21914 35748 21924
rect 35084 21698 35140 21710
rect 35084 21646 35086 21698
rect 35138 21646 35140 21698
rect 35084 21588 35140 21646
rect 35196 21698 35252 21756
rect 35196 21646 35198 21698
rect 35250 21646 35252 21698
rect 35196 21634 35252 21646
rect 35084 21252 35140 21532
rect 34748 21196 35028 21252
rect 35084 21196 35252 21252
rect 34748 21028 34804 21038
rect 34748 20934 34804 20972
rect 34468 20076 34580 20132
rect 34412 20066 34468 20076
rect 34636 20018 34692 20030
rect 34636 19966 34638 20018
rect 34690 19966 34692 20018
rect 34300 19852 34580 19908
rect 34300 19460 34356 19470
rect 34300 19366 34356 19404
rect 34524 19236 34580 19852
rect 34636 19460 34692 19966
rect 34636 19394 34692 19404
rect 34524 19234 34916 19236
rect 34524 19182 34526 19234
rect 34578 19182 34916 19234
rect 34524 19180 34916 19182
rect 34524 19170 34580 19180
rect 34076 18956 34580 19012
rect 34300 18676 34356 18686
rect 33964 18674 34356 18676
rect 33964 18622 34302 18674
rect 34354 18622 34356 18674
rect 33964 18620 34356 18622
rect 34300 18610 34356 18620
rect 33852 18398 33854 18450
rect 33906 18398 33908 18450
rect 33852 18386 33908 18398
rect 34076 18452 34132 18462
rect 34076 18358 34132 18396
rect 34076 18116 34132 18126
rect 33964 17332 34020 17342
rect 33964 17106 34020 17276
rect 33964 17054 33966 17106
rect 34018 17054 34020 17106
rect 33964 17042 34020 17054
rect 33740 16828 34020 16884
rect 33628 15934 33630 15986
rect 33682 15934 33684 15986
rect 33180 15428 33236 15438
rect 33180 15334 33236 15372
rect 33516 15092 33572 15102
rect 33516 14998 33572 15036
rect 33180 14420 33236 14430
rect 33180 13970 33236 14364
rect 33180 13918 33182 13970
rect 33234 13918 33236 13970
rect 33180 13906 33236 13918
rect 33516 13524 33572 13534
rect 33516 13430 33572 13468
rect 33180 12404 33236 12414
rect 33180 12310 33236 12348
rect 33628 12180 33684 15934
rect 33852 16660 33908 16670
rect 33852 15876 33908 16604
rect 33852 15810 33908 15820
rect 33964 15988 34020 16828
rect 34076 15988 34132 18060
rect 34412 17556 34468 17566
rect 34412 17462 34468 17500
rect 34524 17108 34580 18956
rect 34860 18562 34916 19180
rect 34860 18510 34862 18562
rect 34914 18510 34916 18562
rect 34636 18226 34692 18238
rect 34636 18174 34638 18226
rect 34690 18174 34692 18226
rect 34636 18116 34692 18174
rect 34860 18228 34916 18510
rect 34860 18162 34916 18172
rect 34972 19234 35028 21196
rect 34972 19182 34974 19234
rect 35026 19182 35028 19234
rect 34636 18050 34692 18060
rect 34972 17780 35028 19182
rect 35084 19906 35140 19918
rect 35084 19854 35086 19906
rect 35138 19854 35140 19906
rect 35084 19012 35140 19854
rect 35084 18946 35140 18956
rect 34860 17724 35028 17780
rect 34636 17108 34692 17118
rect 34524 17106 34692 17108
rect 34524 17054 34638 17106
rect 34690 17054 34692 17106
rect 34524 17052 34692 17054
rect 34636 17042 34692 17052
rect 34188 16882 34244 16894
rect 34188 16830 34190 16882
rect 34242 16830 34244 16882
rect 34188 16772 34244 16830
rect 34188 16706 34244 16716
rect 34524 16156 34692 16212
rect 34300 15988 34356 15998
rect 34076 15986 34356 15988
rect 34076 15934 34302 15986
rect 34354 15934 34356 15986
rect 34076 15932 34356 15934
rect 33740 15764 33796 15774
rect 33740 15426 33796 15708
rect 33740 15374 33742 15426
rect 33794 15374 33796 15426
rect 33740 13858 33796 15374
rect 33964 15148 34020 15932
rect 34300 15922 34356 15932
rect 34300 15426 34356 15438
rect 34300 15374 34302 15426
rect 34354 15374 34356 15426
rect 33964 15092 34132 15148
rect 33740 13806 33742 13858
rect 33794 13806 33796 13858
rect 33740 13794 33796 13806
rect 33740 13524 33796 13534
rect 33740 12290 33796 13468
rect 33964 13076 34020 13086
rect 33740 12238 33742 12290
rect 33794 12238 33796 12290
rect 33740 12226 33796 12238
rect 33852 13020 33964 13076
rect 33628 12114 33684 12124
rect 33516 11956 33572 11994
rect 33516 11890 33572 11900
rect 33516 11732 33572 11742
rect 32956 11414 33012 11452
rect 33404 11676 33516 11732
rect 33404 10836 33460 11676
rect 33516 11666 33572 11676
rect 33516 11508 33572 11518
rect 33516 11414 33572 11452
rect 33852 11394 33908 13020
rect 33964 13010 34020 13020
rect 34076 12516 34132 15092
rect 34300 14420 34356 15374
rect 34412 14420 34468 14430
rect 34300 14418 34468 14420
rect 34300 14366 34414 14418
rect 34466 14366 34468 14418
rect 34300 14364 34468 14366
rect 34188 13858 34244 13870
rect 34188 13806 34190 13858
rect 34242 13806 34244 13858
rect 34188 12852 34244 13806
rect 34188 12786 34244 12796
rect 34076 12460 34244 12516
rect 34076 12292 34132 12302
rect 34076 11956 34132 12236
rect 33852 11342 33854 11394
rect 33906 11342 33908 11394
rect 33852 11284 33908 11342
rect 33628 11228 33908 11284
rect 33964 11900 34132 11956
rect 33516 10836 33572 10846
rect 33404 10834 33572 10836
rect 33404 10782 33518 10834
rect 33570 10782 33572 10834
rect 33404 10780 33572 10782
rect 33516 10770 33572 10780
rect 32732 9886 32734 9938
rect 32786 9886 32788 9938
rect 32732 9874 32788 9886
rect 33180 10388 33236 10398
rect 33180 9938 33236 10332
rect 33180 9886 33182 9938
rect 33234 9886 33236 9938
rect 33180 9874 33236 9886
rect 33628 9938 33684 11228
rect 33852 10836 33908 10846
rect 33964 10836 34020 11900
rect 33852 10834 34020 10836
rect 33852 10782 33854 10834
rect 33906 10782 34020 10834
rect 33852 10780 34020 10782
rect 34076 11732 34132 11742
rect 33852 10770 33908 10780
rect 33628 9886 33630 9938
rect 33682 9886 33684 9938
rect 33628 9874 33684 9886
rect 34076 9938 34132 11676
rect 34188 11508 34244 12460
rect 34188 11442 34244 11452
rect 34188 11284 34244 11294
rect 34300 11284 34356 14364
rect 34412 14354 34468 14364
rect 34524 12964 34580 16156
rect 34636 16100 34692 16156
rect 34860 16100 34916 17724
rect 35084 17668 35140 17678
rect 34636 16098 34916 16100
rect 34636 16046 34638 16098
rect 34690 16046 34916 16098
rect 34636 16044 34916 16046
rect 34972 17666 35140 17668
rect 34972 17614 35086 17666
rect 35138 17614 35140 17666
rect 34972 17612 35140 17614
rect 34636 16034 34692 16044
rect 34636 15876 34692 15886
rect 34636 15148 34692 15820
rect 34748 15540 34804 15550
rect 34748 15446 34804 15484
rect 34636 15092 34916 15148
rect 34748 13860 34804 13870
rect 34748 13766 34804 13804
rect 34524 12908 34692 12964
rect 34412 12852 34468 12862
rect 34468 12796 34580 12852
rect 34412 12758 34468 12796
rect 34188 11282 34356 11284
rect 34188 11230 34190 11282
rect 34242 11230 34356 11282
rect 34188 11228 34356 11230
rect 34412 11508 34468 11518
rect 34188 11218 34244 11228
rect 34188 10610 34244 10622
rect 34188 10558 34190 10610
rect 34242 10558 34244 10610
rect 34188 10388 34244 10558
rect 34188 10322 34244 10332
rect 34412 10612 34468 11452
rect 34076 9886 34078 9938
rect 34130 9886 34132 9938
rect 34076 9874 34132 9886
rect 34412 9940 34468 10556
rect 34524 10388 34580 12796
rect 34636 11732 34692 12908
rect 34860 12404 34916 15092
rect 34972 14532 35028 17612
rect 35084 17602 35140 17612
rect 35084 17332 35140 17342
rect 35084 16322 35140 17276
rect 35196 16882 35252 21196
rect 35484 20412 35748 20422
rect 35540 20356 35588 20412
rect 35644 20356 35692 20412
rect 35484 20346 35748 20356
rect 35484 18844 35748 18854
rect 35540 18788 35588 18844
rect 35644 18788 35692 18844
rect 35484 18778 35748 18788
rect 35196 16830 35198 16882
rect 35250 16830 35252 16882
rect 35196 16818 35252 16830
rect 35308 18452 35364 18462
rect 35084 16270 35086 16322
rect 35138 16270 35140 16322
rect 35084 16258 35140 16270
rect 35196 16100 35252 16110
rect 35196 16006 35252 16044
rect 35084 15988 35140 15998
rect 35084 15894 35140 15932
rect 35308 15876 35364 18396
rect 35484 17276 35748 17286
rect 35540 17220 35588 17276
rect 35644 17220 35692 17276
rect 35484 17210 35748 17220
rect 35868 16100 35924 29932
rect 35980 21028 36036 33292
rect 36204 31668 36260 31678
rect 36204 22596 36260 31612
rect 36204 22530 36260 22540
rect 35980 20962 36036 20972
rect 35868 16034 35924 16044
rect 35196 15820 35364 15876
rect 35084 15540 35140 15550
rect 35084 15446 35140 15484
rect 35084 14532 35140 14542
rect 34972 14530 35140 14532
rect 34972 14478 35086 14530
rect 35138 14478 35140 14530
rect 34972 14476 35140 14478
rect 35084 13970 35140 14476
rect 35084 13918 35086 13970
rect 35138 13918 35140 13970
rect 35084 13906 35140 13918
rect 35084 13524 35140 13534
rect 35084 12962 35140 13468
rect 35084 12910 35086 12962
rect 35138 12910 35140 12962
rect 35084 12898 35140 12910
rect 34636 11666 34692 11676
rect 34748 12402 34916 12404
rect 34748 12350 34862 12402
rect 34914 12350 34916 12402
rect 34748 12348 34916 12350
rect 34636 11508 34692 11518
rect 34636 11414 34692 11452
rect 34636 10612 34692 10622
rect 34748 10612 34804 12348
rect 34860 12338 34916 12348
rect 34636 10610 34804 10612
rect 34636 10558 34638 10610
rect 34690 10558 34804 10610
rect 34636 10556 34804 10558
rect 34860 12180 34916 12190
rect 35084 12180 35140 12190
rect 35196 12180 35252 15820
rect 35484 15708 35748 15718
rect 35540 15652 35588 15708
rect 35644 15652 35692 15708
rect 35484 15642 35748 15652
rect 34636 10546 34692 10556
rect 34524 10332 34804 10388
rect 34412 9884 34580 9940
rect 33964 9828 34020 9838
rect 34524 9828 34580 9884
rect 34636 9828 34692 9838
rect 34524 9826 34692 9828
rect 34524 9774 34638 9826
rect 34690 9774 34692 9826
rect 34524 9772 34692 9774
rect 33964 9266 34020 9772
rect 34636 9762 34692 9772
rect 33964 9214 33966 9266
rect 34018 9214 34020 9266
rect 33964 9202 34020 9214
rect 34412 9492 34468 9502
rect 34412 9266 34468 9436
rect 34412 9214 34414 9266
rect 34466 9214 34468 9266
rect 34412 9202 34468 9214
rect 33852 9156 33908 9166
rect 33852 7700 33908 9100
rect 34188 8370 34244 8382
rect 34188 8318 34190 8370
rect 34242 8318 34244 8370
rect 34188 8260 34244 8318
rect 34188 8194 34244 8204
rect 34748 8148 34804 10332
rect 34860 9714 34916 12124
rect 34860 9662 34862 9714
rect 34914 9662 34916 9714
rect 34860 9650 34916 9662
rect 34972 12178 35252 12180
rect 34972 12126 35086 12178
rect 35138 12126 35252 12178
rect 34972 12124 35252 12126
rect 35308 15540 35364 15550
rect 34860 9492 34916 9502
rect 34972 9492 35028 12124
rect 35084 12114 35140 12124
rect 35084 11396 35140 11406
rect 35140 11340 35252 11396
rect 35084 11302 35140 11340
rect 35196 10724 35252 11340
rect 35084 10612 35140 10622
rect 35084 10518 35140 10556
rect 35196 10052 35252 10668
rect 34916 9436 35028 9492
rect 35084 9996 35252 10052
rect 34860 9426 34916 9436
rect 34860 9268 34916 9278
rect 35084 9268 35140 9996
rect 35196 9828 35252 9838
rect 35308 9828 35364 15484
rect 35484 14140 35748 14150
rect 35540 14084 35588 14140
rect 35644 14084 35692 14140
rect 35484 14074 35748 14084
rect 35484 12572 35748 12582
rect 35540 12516 35588 12572
rect 35644 12516 35692 12572
rect 35484 12506 35748 12516
rect 35484 11004 35748 11014
rect 35540 10948 35588 11004
rect 35644 10948 35692 11004
rect 35484 10938 35748 10948
rect 35252 9772 35364 9828
rect 35196 9734 35252 9772
rect 35484 9436 35748 9446
rect 35540 9380 35588 9436
rect 35644 9380 35692 9436
rect 35484 9370 35748 9380
rect 35196 9268 35252 9278
rect 34860 9266 35252 9268
rect 34860 9214 34862 9266
rect 34914 9214 35198 9266
rect 35250 9214 35252 9266
rect 34860 9212 35252 9214
rect 34860 9202 34916 9212
rect 35196 9202 35252 9212
rect 34972 8484 35028 8494
rect 34860 8148 34916 8158
rect 34748 8146 34916 8148
rect 34748 8094 34862 8146
rect 34914 8094 34916 8146
rect 34748 8092 34916 8094
rect 34860 8082 34916 8092
rect 34972 7924 35028 8428
rect 35196 8148 35252 8158
rect 35196 8146 35364 8148
rect 35196 8094 35198 8146
rect 35250 8094 35364 8146
rect 35196 8092 35364 8094
rect 35196 8082 35252 8092
rect 34860 7868 35028 7924
rect 33964 7700 34020 7710
rect 33852 7698 34020 7700
rect 33852 7646 33966 7698
rect 34018 7646 34020 7698
rect 33852 7644 34020 7646
rect 33964 7634 34020 7644
rect 34076 7364 34132 7374
rect 34076 7362 34804 7364
rect 34076 7310 34078 7362
rect 34130 7310 34804 7362
rect 34076 7308 34804 7310
rect 34076 7298 34132 7308
rect 34636 5124 34692 5134
rect 34636 5030 34692 5068
rect 34748 4676 34804 7308
rect 34860 5010 34916 7868
rect 35308 7700 35364 8092
rect 35484 7868 35748 7878
rect 35540 7812 35588 7868
rect 35644 7812 35692 7868
rect 35484 7802 35748 7812
rect 35308 7606 35364 7644
rect 35484 6300 35748 6310
rect 35540 6244 35588 6300
rect 35644 6244 35692 6300
rect 35484 6234 35748 6244
rect 35196 5124 35252 5134
rect 35196 5030 35252 5068
rect 34860 4958 34862 5010
rect 34914 4958 34916 5010
rect 34860 4946 34916 4958
rect 35484 4732 35748 4742
rect 35540 4676 35588 4732
rect 35644 4676 35692 4732
rect 34748 4620 34916 4676
rect 35484 4666 35748 4676
rect 33292 4228 33348 4238
rect 33180 4226 33348 4228
rect 33180 4174 33294 4226
rect 33346 4174 33348 4226
rect 33180 4172 33348 4174
rect 32956 3556 33012 3566
rect 32956 3462 33012 3500
rect 33180 3556 33236 4172
rect 33292 4162 33348 4172
rect 33628 3556 33684 3566
rect 33180 3554 33684 3556
rect 33180 3502 33630 3554
rect 33682 3502 33684 3554
rect 33180 3500 33684 3502
rect 32620 2258 32676 2268
rect 33180 800 33236 3500
rect 33628 3490 33684 3500
rect 34636 3442 34692 3454
rect 34636 3390 34638 3442
rect 34690 3390 34692 3442
rect 34636 3388 34692 3390
rect 33404 3332 33460 3342
rect 34636 3332 34804 3388
rect 33404 3238 33460 3276
rect 34748 3108 34804 3332
rect 34860 3330 34916 4620
rect 34860 3278 34862 3330
rect 34914 3278 34916 3330
rect 34860 3266 34916 3278
rect 35084 3554 35140 3566
rect 35084 3502 35086 3554
rect 35138 3502 35140 3554
rect 35084 3108 35140 3502
rect 34748 3052 35140 3108
rect 35484 3164 35748 3174
rect 35540 3108 35588 3164
rect 35644 3108 35692 3164
rect 35484 3098 35748 3108
rect 34748 800 34804 3052
rect 1792 0 1904 800
rect 3360 0 3472 800
rect 4928 0 5040 800
rect 6496 0 6608 800
rect 8064 0 8176 800
rect 9632 0 9744 800
rect 11200 0 11312 800
rect 12768 0 12880 800
rect 14336 0 14448 800
rect 15904 0 16016 800
rect 17472 0 17584 800
rect 19040 0 19152 800
rect 20608 0 20720 800
rect 22176 0 22288 800
rect 23744 0 23856 800
rect 25312 0 25424 800
rect 26880 0 26992 800
rect 28448 0 28560 800
rect 30016 0 30128 800
rect 31584 0 31696 800
rect 33152 0 33264 800
rect 34720 0 34832 800
<< via2 >>
rect 5496 33738 5552 33740
rect 5496 33686 5498 33738
rect 5498 33686 5550 33738
rect 5550 33686 5552 33738
rect 5496 33684 5552 33686
rect 5600 33738 5656 33740
rect 5600 33686 5602 33738
rect 5602 33686 5654 33738
rect 5654 33686 5656 33738
rect 5600 33684 5656 33686
rect 5704 33738 5760 33740
rect 5704 33686 5706 33738
rect 5706 33686 5758 33738
rect 5758 33686 5760 33738
rect 5704 33684 5760 33686
rect 5496 32170 5552 32172
rect 5496 32118 5498 32170
rect 5498 32118 5550 32170
rect 5550 32118 5552 32170
rect 5496 32116 5552 32118
rect 5600 32170 5656 32172
rect 5600 32118 5602 32170
rect 5602 32118 5654 32170
rect 5654 32118 5656 32170
rect 5600 32116 5656 32118
rect 5704 32170 5760 32172
rect 5704 32118 5706 32170
rect 5706 32118 5758 32170
rect 5758 32118 5760 32170
rect 5704 32116 5760 32118
rect 6300 31836 6356 31892
rect 4620 29932 4676 29988
rect 5496 30602 5552 30604
rect 5496 30550 5498 30602
rect 5498 30550 5550 30602
rect 5550 30550 5552 30602
rect 5496 30548 5552 30550
rect 5600 30602 5656 30604
rect 5600 30550 5602 30602
rect 5602 30550 5654 30602
rect 5654 30550 5656 30602
rect 5600 30548 5656 30550
rect 5704 30602 5760 30604
rect 5704 30550 5706 30602
rect 5706 30550 5758 30602
rect 5758 30550 5760 30602
rect 5704 30548 5760 30550
rect 6860 32450 6916 32452
rect 6860 32398 6862 32450
rect 6862 32398 6914 32450
rect 6914 32398 6916 32450
rect 6860 32396 6916 32398
rect 6524 31836 6580 31892
rect 6412 30210 6468 30212
rect 6412 30158 6414 30210
rect 6414 30158 6466 30210
rect 6466 30158 6468 30210
rect 6412 30156 6468 30158
rect 5628 29986 5684 29988
rect 5628 29934 5630 29986
rect 5630 29934 5682 29986
rect 5682 29934 5684 29986
rect 5628 29932 5684 29934
rect 5740 29484 5796 29540
rect 5496 29034 5552 29036
rect 5496 28982 5498 29034
rect 5498 28982 5550 29034
rect 5550 28982 5552 29034
rect 5496 28980 5552 28982
rect 5600 29034 5656 29036
rect 5600 28982 5602 29034
rect 5602 28982 5654 29034
rect 5654 28982 5656 29034
rect 5600 28980 5656 28982
rect 5704 29034 5760 29036
rect 5704 28982 5706 29034
rect 5706 28982 5758 29034
rect 5758 28982 5760 29034
rect 5704 28980 5760 28982
rect 5180 28812 5236 28868
rect 5964 27692 6020 27748
rect 5496 27466 5552 27468
rect 5496 27414 5498 27466
rect 5498 27414 5550 27466
rect 5550 27414 5552 27466
rect 5496 27412 5552 27414
rect 5600 27466 5656 27468
rect 5600 27414 5602 27466
rect 5602 27414 5654 27466
rect 5654 27414 5656 27466
rect 5600 27412 5656 27414
rect 5704 27466 5760 27468
rect 5704 27414 5706 27466
rect 5706 27414 5758 27466
rect 5758 27414 5760 27466
rect 5704 27412 5760 27414
rect 4284 27244 4340 27300
rect 5628 27298 5684 27300
rect 5628 27246 5630 27298
rect 5630 27246 5682 27298
rect 5682 27246 5684 27298
rect 5628 27244 5684 27246
rect 6524 29372 6580 29428
rect 8204 33516 8260 33572
rect 8316 32732 8372 32788
rect 8988 33292 9044 33348
rect 7868 32396 7924 32452
rect 10556 33516 10612 33572
rect 9996 33346 10052 33348
rect 9996 33294 9998 33346
rect 9998 33294 10050 33346
rect 10050 33294 10052 33346
rect 9996 33292 10052 33294
rect 9780 32954 9836 32956
rect 9780 32902 9782 32954
rect 9782 32902 9834 32954
rect 9834 32902 9836 32954
rect 9780 32900 9836 32902
rect 9884 32954 9940 32956
rect 9884 32902 9886 32954
rect 9886 32902 9938 32954
rect 9938 32902 9940 32954
rect 9884 32900 9940 32902
rect 9988 32954 10044 32956
rect 9988 32902 9990 32954
rect 9990 32902 10042 32954
rect 10042 32902 10044 32954
rect 9988 32900 10044 32902
rect 9548 32786 9604 32788
rect 9548 32734 9550 32786
rect 9550 32734 9602 32786
rect 9602 32734 9604 32786
rect 9548 32732 9604 32734
rect 8652 31836 8708 31892
rect 8092 31724 8148 31780
rect 7308 30940 7364 30996
rect 7084 30210 7140 30212
rect 7084 30158 7086 30210
rect 7086 30158 7138 30210
rect 7138 30158 7140 30210
rect 7084 30156 7140 30158
rect 6748 29708 6804 29764
rect 7308 29986 7364 29988
rect 7308 29934 7310 29986
rect 7310 29934 7362 29986
rect 7362 29934 7364 29986
rect 7308 29932 7364 29934
rect 7980 30994 8036 30996
rect 7980 30942 7982 30994
rect 7982 30942 8034 30994
rect 8034 30942 8036 30994
rect 7980 30940 8036 30942
rect 7532 29372 7588 29428
rect 7868 29596 7924 29652
rect 8204 31666 8260 31668
rect 8204 31614 8206 31666
rect 8206 31614 8258 31666
rect 8258 31614 8260 31666
rect 8204 31612 8260 31614
rect 9212 31612 9268 31668
rect 9780 31386 9836 31388
rect 9780 31334 9782 31386
rect 9782 31334 9834 31386
rect 9834 31334 9836 31386
rect 9780 31332 9836 31334
rect 9884 31386 9940 31388
rect 9884 31334 9886 31386
rect 9886 31334 9938 31386
rect 9938 31334 9940 31386
rect 9884 31332 9940 31334
rect 9988 31386 10044 31388
rect 9988 31334 9990 31386
rect 9990 31334 10042 31386
rect 10042 31334 10044 31386
rect 9988 31332 10044 31334
rect 10220 31836 10276 31892
rect 9548 30268 9604 30324
rect 8204 30098 8260 30100
rect 8204 30046 8206 30098
rect 8206 30046 8258 30098
rect 8258 30046 8260 30098
rect 8204 30044 8260 30046
rect 8204 29708 8260 29764
rect 8316 29932 8372 29988
rect 9212 29708 9268 29764
rect 9548 29708 9604 29764
rect 8876 29650 8932 29652
rect 8876 29598 8878 29650
rect 8878 29598 8930 29650
rect 8930 29598 8932 29650
rect 8876 29596 8932 29598
rect 7756 29372 7812 29428
rect 6860 28866 6916 28868
rect 6860 28814 6862 28866
rect 6862 28814 6914 28866
rect 6914 28814 6916 28866
rect 6860 28812 6916 28814
rect 6636 28700 6692 28756
rect 6860 28642 6916 28644
rect 6860 28590 6862 28642
rect 6862 28590 6914 28642
rect 6914 28590 6916 28642
rect 6860 28588 6916 28590
rect 7308 28700 7364 28756
rect 6524 27580 6580 27636
rect 6300 27356 6356 27412
rect 6972 27746 7028 27748
rect 6972 27694 6974 27746
rect 6974 27694 7026 27746
rect 7026 27694 7028 27746
rect 6972 27692 7028 27694
rect 7196 27356 7252 27412
rect 6972 27132 7028 27188
rect 6860 27020 6916 27076
rect 5740 26460 5796 26516
rect 4396 26178 4452 26180
rect 4396 26126 4398 26178
rect 4398 26126 4450 26178
rect 4450 26126 4452 26178
rect 4396 26124 4452 26126
rect 6188 26124 6244 26180
rect 5496 25898 5552 25900
rect 5496 25846 5498 25898
rect 5498 25846 5550 25898
rect 5550 25846 5552 25898
rect 5496 25844 5552 25846
rect 5600 25898 5656 25900
rect 5600 25846 5602 25898
rect 5602 25846 5654 25898
rect 5654 25846 5656 25898
rect 5600 25844 5656 25846
rect 5704 25898 5760 25900
rect 5704 25846 5706 25898
rect 5706 25846 5758 25898
rect 5758 25846 5760 25898
rect 5704 25844 5760 25846
rect 6860 26572 6916 26628
rect 6300 25394 6356 25396
rect 6300 25342 6302 25394
rect 6302 25342 6354 25394
rect 6354 25342 6356 25394
rect 6300 25340 6356 25342
rect 3612 25228 3668 25284
rect 7420 28028 7476 28084
rect 7420 27132 7476 27188
rect 7644 28754 7700 28756
rect 7644 28702 7646 28754
rect 7646 28702 7698 28754
rect 7698 28702 7700 28754
rect 7644 28700 7700 28702
rect 7308 26572 7364 26628
rect 7420 26402 7476 26404
rect 7420 26350 7422 26402
rect 7422 26350 7474 26402
rect 7474 26350 7476 26402
rect 7420 26348 7476 26350
rect 8092 27580 8148 27636
rect 8652 29426 8708 29428
rect 8652 29374 8654 29426
rect 8654 29374 8706 29426
rect 8706 29374 8708 29426
rect 8652 29372 8708 29374
rect 9324 29372 9380 29428
rect 8988 29202 9044 29204
rect 8988 29150 8990 29202
rect 8990 29150 9042 29202
rect 9042 29150 9044 29202
rect 8988 29148 9044 29150
rect 8764 28924 8820 28980
rect 8540 28252 8596 28308
rect 8540 28082 8596 28084
rect 8540 28030 8542 28082
rect 8542 28030 8594 28082
rect 8594 28030 8596 28082
rect 8540 28028 8596 28030
rect 7868 27020 7924 27076
rect 8540 27074 8596 27076
rect 8540 27022 8542 27074
rect 8542 27022 8594 27074
rect 8594 27022 8596 27074
rect 8540 27020 8596 27022
rect 7644 26572 7700 26628
rect 7868 26684 7924 26740
rect 6860 25228 6916 25284
rect 6636 24722 6692 24724
rect 6636 24670 6638 24722
rect 6638 24670 6690 24722
rect 6690 24670 6692 24722
rect 6636 24668 6692 24670
rect 5496 24330 5552 24332
rect 5496 24278 5498 24330
rect 5498 24278 5550 24330
rect 5550 24278 5552 24330
rect 5496 24276 5552 24278
rect 5600 24330 5656 24332
rect 5600 24278 5602 24330
rect 5602 24278 5654 24330
rect 5654 24278 5656 24330
rect 5600 24276 5656 24278
rect 5704 24330 5760 24332
rect 5704 24278 5706 24330
rect 5706 24278 5758 24330
rect 5758 24278 5760 24330
rect 5704 24276 5760 24278
rect 8204 26572 8260 26628
rect 8540 26572 8596 26628
rect 8428 26514 8484 26516
rect 8428 26462 8430 26514
rect 8430 26462 8482 26514
rect 8482 26462 8484 26514
rect 8428 26460 8484 26462
rect 8204 26348 8260 26404
rect 8092 25228 8148 25284
rect 8540 25900 8596 25956
rect 9548 29260 9604 29316
rect 9996 29986 10052 29988
rect 9996 29934 9998 29986
rect 9998 29934 10050 29986
rect 10050 29934 10052 29986
rect 9996 29932 10052 29934
rect 9780 29818 9836 29820
rect 9780 29766 9782 29818
rect 9782 29766 9834 29818
rect 9834 29766 9836 29818
rect 9780 29764 9836 29766
rect 9884 29818 9940 29820
rect 9884 29766 9886 29818
rect 9886 29766 9938 29818
rect 9938 29766 9940 29818
rect 9884 29764 9940 29766
rect 9988 29818 10044 29820
rect 9988 29766 9990 29818
rect 9990 29766 10042 29818
rect 10042 29766 10044 29818
rect 9988 29764 10044 29766
rect 10444 30994 10500 30996
rect 10444 30942 10446 30994
rect 10446 30942 10498 30994
rect 10498 30942 10500 30994
rect 10444 30940 10500 30942
rect 10668 30156 10724 30212
rect 10892 29932 10948 29988
rect 10108 29650 10164 29652
rect 10108 29598 10110 29650
rect 10110 29598 10162 29650
rect 10162 29598 10164 29650
rect 10108 29596 10164 29598
rect 10332 29820 10388 29876
rect 9996 29484 10052 29540
rect 9884 29426 9940 29428
rect 9884 29374 9886 29426
rect 9886 29374 9938 29426
rect 9938 29374 9940 29426
rect 9884 29372 9940 29374
rect 9324 28924 9380 28980
rect 10780 29148 10836 29204
rect 8764 28028 8820 28084
rect 9996 28530 10052 28532
rect 9996 28478 9998 28530
rect 9998 28478 10050 28530
rect 10050 28478 10052 28530
rect 9996 28476 10052 28478
rect 9324 28252 9380 28308
rect 9100 27916 9156 27972
rect 8988 27804 9044 27860
rect 9780 28250 9836 28252
rect 9780 28198 9782 28250
rect 9782 28198 9834 28250
rect 9834 28198 9836 28250
rect 9780 28196 9836 28198
rect 9884 28250 9940 28252
rect 9884 28198 9886 28250
rect 9886 28198 9938 28250
rect 9938 28198 9940 28250
rect 9884 28196 9940 28198
rect 9988 28250 10044 28252
rect 9988 28198 9990 28250
rect 9990 28198 10042 28250
rect 10042 28198 10044 28250
rect 9988 28196 10044 28198
rect 9884 27746 9940 27748
rect 9884 27694 9886 27746
rect 9886 27694 9938 27746
rect 9938 27694 9940 27746
rect 9884 27692 9940 27694
rect 9884 27186 9940 27188
rect 9884 27134 9886 27186
rect 9886 27134 9938 27186
rect 9938 27134 9940 27186
rect 9884 27132 9940 27134
rect 10108 27074 10164 27076
rect 10108 27022 10110 27074
rect 10110 27022 10162 27074
rect 10162 27022 10164 27074
rect 10108 27020 10164 27022
rect 10332 27916 10388 27972
rect 10332 27244 10388 27300
rect 9884 26796 9940 26852
rect 9780 26682 9836 26684
rect 9780 26630 9782 26682
rect 9782 26630 9834 26682
rect 9834 26630 9836 26682
rect 9780 26628 9836 26630
rect 9884 26682 9940 26684
rect 9884 26630 9886 26682
rect 9886 26630 9938 26682
rect 9938 26630 9940 26682
rect 9884 26628 9940 26630
rect 9988 26682 10044 26684
rect 9988 26630 9990 26682
rect 9990 26630 10042 26682
rect 10042 26630 10044 26682
rect 9988 26628 10044 26630
rect 9772 26514 9828 26516
rect 9772 26462 9774 26514
rect 9774 26462 9826 26514
rect 9826 26462 9828 26514
rect 9772 26460 9828 26462
rect 9884 26402 9940 26404
rect 9884 26350 9886 26402
rect 9886 26350 9938 26402
rect 9938 26350 9940 26402
rect 9884 26348 9940 26350
rect 9436 26236 9492 26292
rect 10892 28924 10948 28980
rect 11116 29596 11172 29652
rect 11228 30716 11284 30772
rect 10892 27858 10948 27860
rect 10892 27806 10894 27858
rect 10894 27806 10946 27858
rect 10946 27806 10948 27858
rect 10892 27804 10948 27806
rect 12348 33570 12404 33572
rect 12348 33518 12350 33570
rect 12350 33518 12402 33570
rect 12402 33518 12404 33570
rect 12348 33516 12404 33518
rect 14064 33738 14120 33740
rect 14064 33686 14066 33738
rect 14066 33686 14118 33738
rect 14118 33686 14120 33738
rect 14064 33684 14120 33686
rect 14168 33738 14224 33740
rect 14168 33686 14170 33738
rect 14170 33686 14222 33738
rect 14222 33686 14224 33738
rect 14168 33684 14224 33686
rect 14272 33738 14328 33740
rect 14272 33686 14274 33738
rect 14274 33686 14326 33738
rect 14326 33686 14328 33738
rect 14272 33684 14328 33686
rect 13916 33516 13972 33572
rect 11900 31890 11956 31892
rect 11900 31838 11902 31890
rect 11902 31838 11954 31890
rect 11954 31838 11956 31890
rect 11900 31836 11956 31838
rect 11564 30994 11620 30996
rect 11564 30942 11566 30994
rect 11566 30942 11618 30994
rect 11618 30942 11620 30994
rect 11564 30940 11620 30942
rect 12124 31500 12180 31556
rect 12460 31500 12516 31556
rect 12572 30380 12628 30436
rect 12572 30156 12628 30212
rect 11452 29596 11508 29652
rect 12572 29650 12628 29652
rect 12572 29598 12574 29650
rect 12574 29598 12626 29650
rect 12626 29598 12628 29650
rect 12572 29596 12628 29598
rect 11228 28812 11284 28868
rect 11564 29148 11620 29204
rect 11788 28700 11844 28756
rect 11340 28476 11396 28532
rect 10892 27580 10948 27636
rect 13244 31500 13300 31556
rect 12236 28700 12292 28756
rect 12460 28588 12516 28644
rect 11452 27132 11508 27188
rect 11004 27074 11060 27076
rect 11004 27022 11006 27074
rect 11006 27022 11058 27074
rect 11058 27022 11060 27074
rect 11004 27020 11060 27022
rect 12012 27804 12068 27860
rect 14064 32170 14120 32172
rect 14064 32118 14066 32170
rect 14066 32118 14118 32170
rect 14118 32118 14120 32170
rect 14064 32116 14120 32118
rect 14168 32170 14224 32172
rect 14168 32118 14170 32170
rect 14170 32118 14222 32170
rect 14222 32118 14224 32170
rect 14168 32116 14224 32118
rect 14272 32170 14328 32172
rect 14272 32118 14274 32170
rect 14274 32118 14326 32170
rect 14326 32118 14328 32170
rect 14272 32116 14328 32118
rect 14588 31778 14644 31780
rect 14588 31726 14590 31778
rect 14590 31726 14642 31778
rect 14642 31726 14644 31778
rect 14588 31724 14644 31726
rect 13804 31554 13860 31556
rect 13804 31502 13806 31554
rect 13806 31502 13858 31554
rect 13858 31502 13860 31554
rect 13804 31500 13860 31502
rect 14064 30602 14120 30604
rect 14064 30550 14066 30602
rect 14066 30550 14118 30602
rect 14118 30550 14120 30602
rect 14064 30548 14120 30550
rect 14168 30602 14224 30604
rect 14168 30550 14170 30602
rect 14170 30550 14222 30602
rect 14222 30550 14224 30602
rect 14168 30548 14224 30550
rect 14272 30602 14328 30604
rect 14272 30550 14274 30602
rect 14274 30550 14326 30602
rect 14326 30550 14328 30602
rect 14272 30548 14328 30550
rect 14028 30380 14084 30436
rect 13020 30044 13076 30100
rect 14588 30940 14644 30996
rect 14924 30882 14980 30884
rect 14924 30830 14926 30882
rect 14926 30830 14978 30882
rect 14978 30830 14980 30882
rect 14924 30828 14980 30830
rect 14064 29034 14120 29036
rect 14064 28982 14066 29034
rect 14066 28982 14118 29034
rect 14118 28982 14120 29034
rect 14064 28980 14120 28982
rect 14168 29034 14224 29036
rect 14168 28982 14170 29034
rect 14170 28982 14222 29034
rect 14222 28982 14224 29034
rect 14168 28980 14224 28982
rect 14272 29034 14328 29036
rect 14272 28982 14274 29034
rect 14274 28982 14326 29034
rect 14326 28982 14328 29034
rect 14272 28980 14328 28982
rect 12684 28588 12740 28644
rect 11900 27244 11956 27300
rect 12796 27634 12852 27636
rect 12796 27582 12798 27634
rect 12798 27582 12850 27634
rect 12850 27582 12852 27634
rect 12796 27580 12852 27582
rect 12908 27356 12964 27412
rect 12572 27074 12628 27076
rect 12572 27022 12574 27074
rect 12574 27022 12626 27074
rect 12626 27022 12628 27074
rect 12572 27020 12628 27022
rect 12348 26908 12404 26964
rect 10780 26572 10836 26628
rect 10444 26012 10500 26068
rect 9884 25900 9940 25956
rect 11564 26348 11620 26404
rect 12124 26124 12180 26180
rect 9780 25114 9836 25116
rect 9780 25062 9782 25114
rect 9782 25062 9834 25114
rect 9834 25062 9836 25114
rect 9780 25060 9836 25062
rect 9884 25114 9940 25116
rect 9884 25062 9886 25114
rect 9886 25062 9938 25114
rect 9938 25062 9940 25114
rect 9884 25060 9940 25062
rect 9988 25114 10044 25116
rect 9988 25062 9990 25114
rect 9990 25062 10042 25114
rect 10042 25062 10044 25114
rect 9988 25060 10044 25062
rect 7196 24722 7252 24724
rect 7196 24670 7198 24722
rect 7198 24670 7250 24722
rect 7250 24670 7252 24722
rect 7196 24668 7252 24670
rect 7756 24722 7812 24724
rect 7756 24670 7758 24722
rect 7758 24670 7810 24722
rect 7810 24670 7812 24722
rect 7756 24668 7812 24670
rect 6748 23714 6804 23716
rect 6748 23662 6750 23714
rect 6750 23662 6802 23714
rect 6802 23662 6804 23714
rect 6748 23660 6804 23662
rect 4732 23042 4788 23044
rect 4732 22990 4734 23042
rect 4734 22990 4786 23042
rect 4786 22990 4788 23042
rect 4732 22988 4788 22990
rect 5496 22762 5552 22764
rect 5496 22710 5498 22762
rect 5498 22710 5550 22762
rect 5550 22710 5552 22762
rect 5496 22708 5552 22710
rect 5600 22762 5656 22764
rect 5600 22710 5602 22762
rect 5602 22710 5654 22762
rect 5654 22710 5656 22762
rect 5600 22708 5656 22710
rect 5704 22762 5760 22764
rect 5704 22710 5706 22762
rect 5706 22710 5758 22762
rect 5758 22710 5760 22762
rect 5704 22708 5760 22710
rect 4396 22092 4452 22148
rect 6636 22146 6692 22148
rect 6636 22094 6638 22146
rect 6638 22094 6690 22146
rect 6690 22094 6692 22146
rect 6636 22092 6692 22094
rect 6972 23436 7028 23492
rect 7084 22540 7140 22596
rect 7308 23826 7364 23828
rect 7308 23774 7310 23826
rect 7310 23774 7362 23826
rect 7362 23774 7364 23826
rect 7308 23772 7364 23774
rect 7756 23772 7812 23828
rect 7420 23660 7476 23716
rect 7308 23042 7364 23044
rect 7308 22990 7310 23042
rect 7310 22990 7362 23042
rect 7362 22990 7364 23042
rect 7308 22988 7364 22990
rect 7868 23660 7924 23716
rect 10220 25340 10276 25396
rect 11900 26066 11956 26068
rect 11900 26014 11902 26066
rect 11902 26014 11954 26066
rect 11954 26014 11956 26066
rect 11900 26012 11956 26014
rect 13804 28530 13860 28532
rect 13804 28478 13806 28530
rect 13806 28478 13858 28530
rect 13858 28478 13860 28530
rect 13804 28476 13860 28478
rect 12460 26402 12516 26404
rect 12460 26350 12462 26402
rect 12462 26350 12514 26402
rect 12514 26350 12516 26402
rect 12460 26348 12516 26350
rect 12908 25452 12964 25508
rect 12236 25282 12292 25284
rect 12236 25230 12238 25282
rect 12238 25230 12290 25282
rect 12290 25230 12292 25282
rect 12236 25228 12292 25230
rect 8316 24722 8372 24724
rect 8316 24670 8318 24722
rect 8318 24670 8370 24722
rect 8370 24670 8372 24722
rect 8316 24668 8372 24670
rect 7980 23436 8036 23492
rect 6524 21474 6580 21476
rect 6524 21422 6526 21474
rect 6526 21422 6578 21474
rect 6578 21422 6580 21474
rect 6524 21420 6580 21422
rect 5496 21194 5552 21196
rect 5496 21142 5498 21194
rect 5498 21142 5550 21194
rect 5550 21142 5552 21194
rect 5496 21140 5552 21142
rect 5600 21194 5656 21196
rect 5600 21142 5602 21194
rect 5602 21142 5654 21194
rect 5654 21142 5656 21194
rect 5600 21140 5656 21142
rect 5704 21194 5760 21196
rect 5704 21142 5706 21194
rect 5706 21142 5758 21194
rect 5758 21142 5760 21194
rect 5704 21140 5760 21142
rect 7196 21420 7252 21476
rect 7756 22540 7812 22596
rect 8204 22652 8260 22708
rect 7532 21420 7588 21476
rect 3724 20188 3780 20244
rect 5068 20188 5124 20244
rect 6524 20524 6580 20580
rect 6300 20188 6356 20244
rect 5740 19906 5796 19908
rect 5740 19854 5742 19906
rect 5742 19854 5794 19906
rect 5794 19854 5796 19906
rect 5740 19852 5796 19854
rect 5496 19626 5552 19628
rect 5496 19574 5498 19626
rect 5498 19574 5550 19626
rect 5550 19574 5552 19626
rect 5496 19572 5552 19574
rect 5600 19626 5656 19628
rect 5600 19574 5602 19626
rect 5602 19574 5654 19626
rect 5654 19574 5656 19626
rect 5600 19572 5656 19574
rect 5704 19626 5760 19628
rect 5704 19574 5706 19626
rect 5706 19574 5758 19626
rect 5758 19574 5760 19626
rect 5704 19572 5760 19574
rect 6860 19740 6916 19796
rect 6972 18732 7028 18788
rect 7420 20578 7476 20580
rect 7420 20526 7422 20578
rect 7422 20526 7474 20578
rect 7474 20526 7476 20578
rect 7420 20524 7476 20526
rect 7308 18620 7364 18676
rect 7532 19292 7588 19348
rect 6076 18508 6132 18564
rect 7420 18562 7476 18564
rect 7420 18510 7422 18562
rect 7422 18510 7474 18562
rect 7474 18510 7476 18562
rect 7420 18508 7476 18510
rect 7308 18396 7364 18452
rect 5496 18058 5552 18060
rect 5496 18006 5498 18058
rect 5498 18006 5550 18058
rect 5550 18006 5552 18058
rect 5496 18004 5552 18006
rect 5600 18058 5656 18060
rect 5600 18006 5602 18058
rect 5602 18006 5654 18058
rect 5654 18006 5656 18058
rect 5600 18004 5656 18006
rect 5704 18058 5760 18060
rect 5704 18006 5706 18058
rect 5706 18006 5758 18058
rect 5758 18006 5760 18058
rect 5704 18004 5760 18006
rect 7868 20188 7924 20244
rect 7980 20076 8036 20132
rect 7868 19740 7924 19796
rect 7868 18620 7924 18676
rect 8204 20188 8260 20244
rect 8428 23154 8484 23156
rect 8428 23102 8430 23154
rect 8430 23102 8482 23154
rect 8482 23102 8484 23154
rect 8428 23100 8484 23102
rect 8428 21586 8484 21588
rect 8428 21534 8430 21586
rect 8430 21534 8482 21586
rect 8482 21534 8484 21586
rect 8428 21532 8484 21534
rect 12236 24892 12292 24948
rect 9548 24668 9604 24724
rect 9100 24444 9156 24500
rect 9884 24444 9940 24500
rect 10220 23772 10276 23828
rect 9780 23546 9836 23548
rect 9780 23494 9782 23546
rect 9782 23494 9834 23546
rect 9834 23494 9836 23546
rect 9780 23492 9836 23494
rect 9884 23546 9940 23548
rect 9884 23494 9886 23546
rect 9886 23494 9938 23546
rect 9938 23494 9940 23546
rect 9884 23492 9940 23494
rect 9988 23546 10044 23548
rect 9988 23494 9990 23546
rect 9990 23494 10042 23546
rect 10042 23494 10044 23546
rect 9988 23492 10044 23494
rect 7980 18508 8036 18564
rect 8540 20802 8596 20804
rect 8540 20750 8542 20802
rect 8542 20750 8594 20802
rect 8594 20750 8596 20802
rect 8540 20748 8596 20750
rect 9436 23154 9492 23156
rect 9436 23102 9438 23154
rect 9438 23102 9490 23154
rect 9490 23102 9492 23154
rect 9436 23100 9492 23102
rect 9660 22652 9716 22708
rect 10108 22540 10164 22596
rect 8876 22428 8932 22484
rect 11564 24834 11620 24836
rect 11564 24782 11566 24834
rect 11566 24782 11618 24834
rect 11618 24782 11620 24834
rect 11564 24780 11620 24782
rect 12012 24780 12068 24836
rect 10332 22482 10388 22484
rect 10332 22430 10334 22482
rect 10334 22430 10386 22482
rect 10386 22430 10388 22482
rect 10332 22428 10388 22430
rect 10556 23154 10612 23156
rect 10556 23102 10558 23154
rect 10558 23102 10610 23154
rect 10610 23102 10612 23154
rect 10556 23100 10612 23102
rect 10108 22092 10164 22148
rect 9780 21978 9836 21980
rect 9780 21926 9782 21978
rect 9782 21926 9834 21978
rect 9834 21926 9836 21978
rect 9780 21924 9836 21926
rect 9884 21978 9940 21980
rect 9884 21926 9886 21978
rect 9886 21926 9938 21978
rect 9938 21926 9940 21978
rect 9884 21924 9940 21926
rect 9988 21978 10044 21980
rect 9988 21926 9990 21978
rect 9990 21926 10042 21978
rect 10042 21926 10044 21978
rect 9988 21924 10044 21926
rect 11116 24444 11172 24500
rect 11564 22540 11620 22596
rect 11564 22258 11620 22260
rect 11564 22206 11566 22258
rect 11566 22206 11618 22258
rect 11618 22206 11620 22258
rect 11564 22204 11620 22206
rect 10444 21756 10500 21812
rect 12796 24946 12852 24948
rect 12796 24894 12798 24946
rect 12798 24894 12850 24946
rect 12850 24894 12852 24946
rect 12796 24892 12852 24894
rect 12348 24834 12404 24836
rect 12348 24782 12350 24834
rect 12350 24782 12402 24834
rect 12402 24782 12404 24834
rect 12348 24780 12404 24782
rect 13692 28418 13748 28420
rect 13692 28366 13694 28418
rect 13694 28366 13746 28418
rect 13746 28366 13748 28418
rect 13692 28364 13748 28366
rect 13692 27858 13748 27860
rect 13692 27806 13694 27858
rect 13694 27806 13746 27858
rect 13746 27806 13748 27858
rect 13692 27804 13748 27806
rect 13468 27356 13524 27412
rect 13804 27580 13860 27636
rect 14252 27970 14308 27972
rect 14252 27918 14254 27970
rect 14254 27918 14306 27970
rect 14306 27918 14308 27970
rect 14252 27916 14308 27918
rect 14064 27466 14120 27468
rect 14064 27414 14066 27466
rect 14066 27414 14118 27466
rect 14118 27414 14120 27466
rect 14064 27412 14120 27414
rect 14168 27466 14224 27468
rect 14168 27414 14170 27466
rect 14170 27414 14222 27466
rect 14222 27414 14224 27466
rect 14168 27412 14224 27414
rect 14272 27466 14328 27468
rect 14272 27414 14274 27466
rect 14274 27414 14326 27466
rect 14326 27414 14328 27466
rect 14272 27412 14328 27414
rect 13132 26178 13188 26180
rect 13132 26126 13134 26178
rect 13134 26126 13186 26178
rect 13186 26126 13188 26178
rect 13132 26124 13188 26126
rect 13356 26460 13412 26516
rect 13916 26850 13972 26852
rect 13916 26798 13918 26850
rect 13918 26798 13970 26850
rect 13970 26798 13972 26850
rect 13916 26796 13972 26798
rect 14064 25898 14120 25900
rect 14064 25846 14066 25898
rect 14066 25846 14118 25898
rect 14118 25846 14120 25898
rect 14064 25844 14120 25846
rect 14168 25898 14224 25900
rect 14168 25846 14170 25898
rect 14170 25846 14222 25898
rect 14222 25846 14224 25898
rect 14168 25844 14224 25846
rect 14272 25898 14328 25900
rect 14272 25846 14274 25898
rect 14274 25846 14326 25898
rect 14326 25846 14328 25898
rect 14272 25844 14328 25846
rect 13692 25564 13748 25620
rect 14028 25564 14084 25620
rect 13244 25004 13300 25060
rect 13692 25116 13748 25172
rect 13132 24444 13188 24500
rect 12012 23548 12068 23604
rect 11900 22092 11956 22148
rect 11900 21868 11956 21924
rect 10332 21532 10388 21588
rect 8764 20636 8820 20692
rect 8876 21474 8932 21476
rect 8876 21422 8878 21474
rect 8878 21422 8930 21474
rect 8930 21422 8932 21474
rect 8876 21420 8932 21422
rect 8540 20018 8596 20020
rect 8540 19966 8542 20018
rect 8542 19966 8594 20018
rect 8594 19966 8596 20018
rect 8540 19964 8596 19966
rect 8652 19906 8708 19908
rect 8652 19854 8654 19906
rect 8654 19854 8706 19906
rect 8706 19854 8708 19906
rect 8652 19852 8708 19854
rect 8428 19740 8484 19796
rect 8540 19346 8596 19348
rect 8540 19294 8542 19346
rect 8542 19294 8594 19346
rect 8594 19294 8596 19346
rect 8540 19292 8596 19294
rect 8204 18732 8260 18788
rect 8092 18284 8148 18340
rect 9324 21308 9380 21364
rect 9324 20802 9380 20804
rect 9324 20750 9326 20802
rect 9326 20750 9378 20802
rect 9378 20750 9380 20802
rect 9324 20748 9380 20750
rect 9548 20690 9604 20692
rect 9548 20638 9550 20690
rect 9550 20638 9602 20690
rect 9602 20638 9604 20690
rect 9548 20636 9604 20638
rect 9780 20410 9836 20412
rect 9780 20358 9782 20410
rect 9782 20358 9834 20410
rect 9834 20358 9836 20410
rect 9780 20356 9836 20358
rect 9884 20410 9940 20412
rect 9884 20358 9886 20410
rect 9886 20358 9938 20410
rect 9938 20358 9940 20410
rect 9884 20356 9940 20358
rect 9988 20410 10044 20412
rect 9988 20358 9990 20410
rect 9990 20358 10042 20410
rect 10042 20358 10044 20410
rect 9988 20356 10044 20358
rect 10332 20188 10388 20244
rect 9436 20018 9492 20020
rect 9436 19966 9438 20018
rect 9438 19966 9490 20018
rect 9490 19966 9492 20018
rect 9436 19964 9492 19966
rect 9772 20130 9828 20132
rect 9772 20078 9774 20130
rect 9774 20078 9826 20130
rect 9826 20078 9828 20130
rect 9772 20076 9828 20078
rect 10780 21532 10836 21588
rect 9660 19740 9716 19796
rect 10220 19852 10276 19908
rect 8988 19292 9044 19348
rect 9100 18732 9156 18788
rect 8876 18396 8932 18452
rect 9780 18842 9836 18844
rect 9780 18790 9782 18842
rect 9782 18790 9834 18842
rect 9834 18790 9836 18842
rect 9780 18788 9836 18790
rect 9884 18842 9940 18844
rect 9884 18790 9886 18842
rect 9886 18790 9938 18842
rect 9938 18790 9940 18842
rect 9884 18788 9940 18790
rect 9988 18842 10044 18844
rect 9988 18790 9990 18842
rect 9990 18790 10042 18842
rect 10042 18790 10044 18842
rect 9988 18788 10044 18790
rect 10892 21474 10948 21476
rect 10892 21422 10894 21474
rect 10894 21422 10946 21474
rect 10946 21422 10948 21474
rect 10892 21420 10948 21422
rect 11564 20860 11620 20916
rect 10892 20412 10948 20468
rect 11452 20412 11508 20468
rect 11228 20018 11284 20020
rect 11228 19966 11230 20018
rect 11230 19966 11282 20018
rect 11282 19966 11284 20018
rect 11228 19964 11284 19966
rect 12908 23938 12964 23940
rect 12908 23886 12910 23938
rect 12910 23886 12962 23938
rect 12962 23886 12964 23938
rect 12908 23884 12964 23886
rect 13356 23548 13412 23604
rect 12460 22258 12516 22260
rect 12460 22206 12462 22258
rect 12462 22206 12514 22258
rect 12514 22206 12516 22258
rect 12460 22204 12516 22206
rect 12908 22204 12964 22260
rect 12908 21810 12964 21812
rect 12908 21758 12910 21810
rect 12910 21758 12962 21810
rect 12962 21758 12964 21810
rect 12908 21756 12964 21758
rect 13580 24444 13636 24500
rect 13580 23938 13636 23940
rect 13580 23886 13582 23938
rect 13582 23886 13634 23938
rect 13634 23886 13636 23938
rect 13580 23884 13636 23886
rect 13356 21868 13412 21924
rect 13580 22092 13636 22148
rect 13244 20748 13300 20804
rect 14252 25004 14308 25060
rect 14588 28476 14644 28532
rect 14700 28418 14756 28420
rect 14700 28366 14702 28418
rect 14702 28366 14754 28418
rect 14754 28366 14756 28418
rect 14700 28364 14756 28366
rect 14588 27244 14644 27300
rect 16044 33458 16100 33460
rect 16044 33406 16046 33458
rect 16046 33406 16098 33458
rect 16098 33406 16100 33458
rect 16044 33404 16100 33406
rect 15820 32786 15876 32788
rect 15820 32734 15822 32786
rect 15822 32734 15874 32786
rect 15874 32734 15876 32786
rect 15820 32732 15876 32734
rect 15372 32450 15428 32452
rect 15372 32398 15374 32450
rect 15374 32398 15426 32450
rect 15426 32398 15428 32450
rect 15372 32396 15428 32398
rect 15372 31218 15428 31220
rect 15372 31166 15374 31218
rect 15374 31166 15426 31218
rect 15426 31166 15428 31218
rect 15372 31164 15428 31166
rect 15708 31164 15764 31220
rect 15596 30994 15652 30996
rect 15596 30942 15598 30994
rect 15598 30942 15650 30994
rect 15650 30942 15652 30994
rect 15596 30940 15652 30942
rect 16828 32674 16884 32676
rect 16828 32622 16830 32674
rect 16830 32622 16882 32674
rect 16882 32622 16884 32674
rect 16828 32620 16884 32622
rect 16268 32396 16324 32452
rect 16156 31276 16212 31332
rect 16044 30994 16100 30996
rect 16044 30942 16046 30994
rect 16046 30942 16098 30994
rect 16098 30942 16100 30994
rect 16044 30940 16100 30942
rect 16268 30940 16324 30996
rect 16380 29820 16436 29876
rect 15372 28754 15428 28756
rect 15372 28702 15374 28754
rect 15374 28702 15426 28754
rect 15426 28702 15428 28754
rect 15372 28700 15428 28702
rect 15036 28642 15092 28644
rect 15036 28590 15038 28642
rect 15038 28590 15090 28642
rect 15090 28590 15092 28642
rect 15036 28588 15092 28590
rect 16268 29426 16324 29428
rect 16268 29374 16270 29426
rect 16270 29374 16322 29426
rect 16322 29374 16324 29426
rect 16268 29372 16324 29374
rect 15932 28754 15988 28756
rect 15932 28702 15934 28754
rect 15934 28702 15986 28754
rect 15986 28702 15988 28754
rect 15932 28700 15988 28702
rect 16268 29148 16324 29204
rect 15820 28588 15876 28644
rect 15596 28140 15652 28196
rect 14812 27804 14868 27860
rect 14700 27132 14756 27188
rect 14700 26962 14756 26964
rect 14700 26910 14702 26962
rect 14702 26910 14754 26962
rect 14754 26910 14756 26962
rect 14700 26908 14756 26910
rect 15148 27970 15204 27972
rect 15148 27918 15150 27970
rect 15150 27918 15202 27970
rect 15202 27918 15204 27970
rect 15148 27916 15204 27918
rect 15036 27692 15092 27748
rect 15260 27132 15316 27188
rect 14812 26796 14868 26852
rect 14700 26012 14756 26068
rect 14924 26348 14980 26404
rect 14924 26012 14980 26068
rect 15036 25900 15092 25956
rect 15036 25452 15092 25508
rect 14476 24444 14532 24500
rect 14064 24330 14120 24332
rect 14064 24278 14066 24330
rect 14066 24278 14118 24330
rect 14118 24278 14120 24330
rect 14064 24276 14120 24278
rect 14168 24330 14224 24332
rect 14168 24278 14170 24330
rect 14170 24278 14222 24330
rect 14222 24278 14224 24330
rect 14168 24276 14224 24278
rect 14272 24330 14328 24332
rect 14272 24278 14274 24330
rect 14274 24278 14326 24330
rect 14326 24278 14328 24330
rect 14272 24276 14328 24278
rect 14252 23884 14308 23940
rect 13804 23100 13860 23156
rect 14064 22762 14120 22764
rect 14064 22710 14066 22762
rect 14066 22710 14118 22762
rect 14118 22710 14120 22762
rect 14064 22708 14120 22710
rect 14168 22762 14224 22764
rect 14168 22710 14170 22762
rect 14170 22710 14222 22762
rect 14222 22710 14224 22762
rect 14168 22708 14224 22710
rect 14272 22762 14328 22764
rect 14272 22710 14274 22762
rect 14274 22710 14326 22762
rect 14326 22710 14328 22762
rect 14272 22708 14328 22710
rect 13804 22428 13860 22484
rect 14476 21756 14532 21812
rect 12236 20412 12292 20468
rect 12908 20188 12964 20244
rect 11004 19740 11060 19796
rect 9548 18396 9604 18452
rect 8988 17836 9044 17892
rect 9884 17836 9940 17892
rect 10220 18284 10276 18340
rect 9780 17274 9836 17276
rect 9780 17222 9782 17274
rect 9782 17222 9834 17274
rect 9834 17222 9836 17274
rect 9780 17220 9836 17222
rect 9884 17274 9940 17276
rect 9884 17222 9886 17274
rect 9886 17222 9938 17274
rect 9938 17222 9940 17274
rect 9884 17220 9940 17222
rect 9988 17274 10044 17276
rect 9988 17222 9990 17274
rect 9990 17222 10042 17274
rect 10042 17222 10044 17274
rect 9988 17220 10044 17222
rect 11004 19292 11060 19348
rect 10556 18450 10612 18452
rect 10556 18398 10558 18450
rect 10558 18398 10610 18450
rect 10610 18398 10612 18450
rect 10556 18396 10612 18398
rect 10444 18284 10500 18340
rect 10332 17052 10388 17108
rect 8316 16604 8372 16660
rect 5496 16490 5552 16492
rect 5496 16438 5498 16490
rect 5498 16438 5550 16490
rect 5550 16438 5552 16490
rect 5496 16436 5552 16438
rect 5600 16490 5656 16492
rect 5600 16438 5602 16490
rect 5602 16438 5654 16490
rect 5654 16438 5656 16490
rect 5600 16436 5656 16438
rect 5704 16490 5760 16492
rect 5704 16438 5706 16490
rect 5706 16438 5758 16490
rect 5758 16438 5760 16490
rect 5704 16436 5760 16438
rect 5496 14922 5552 14924
rect 5496 14870 5498 14922
rect 5498 14870 5550 14922
rect 5550 14870 5552 14922
rect 5496 14868 5552 14870
rect 5600 14922 5656 14924
rect 5600 14870 5602 14922
rect 5602 14870 5654 14922
rect 5654 14870 5656 14922
rect 5600 14868 5656 14870
rect 5704 14922 5760 14924
rect 5704 14870 5706 14922
rect 5706 14870 5758 14922
rect 5758 14870 5760 14922
rect 5704 14868 5760 14870
rect 9772 16882 9828 16884
rect 9772 16830 9774 16882
rect 9774 16830 9826 16882
rect 9826 16830 9828 16882
rect 9772 16828 9828 16830
rect 10892 17388 10948 17444
rect 10780 17106 10836 17108
rect 10780 17054 10782 17106
rect 10782 17054 10834 17106
rect 10834 17054 10836 17106
rect 10780 17052 10836 17054
rect 10444 16828 10500 16884
rect 10108 16716 10164 16772
rect 9212 16210 9268 16212
rect 9212 16158 9214 16210
rect 9214 16158 9266 16210
rect 9266 16158 9268 16210
rect 9212 16156 9268 16158
rect 12348 19740 12404 19796
rect 12572 20018 12628 20020
rect 12572 19966 12574 20018
rect 12574 19966 12626 20018
rect 12626 19966 12628 20018
rect 12572 19964 12628 19966
rect 12796 19906 12852 19908
rect 12796 19854 12798 19906
rect 12798 19854 12850 19906
rect 12850 19854 12852 19906
rect 12796 19852 12852 19854
rect 13468 20188 13524 20244
rect 12684 19234 12740 19236
rect 12684 19182 12686 19234
rect 12686 19182 12738 19234
rect 12738 19182 12740 19234
rect 12684 19180 12740 19182
rect 12796 19122 12852 19124
rect 12796 19070 12798 19122
rect 12798 19070 12850 19122
rect 12850 19070 12852 19122
rect 12796 19068 12852 19070
rect 12684 18508 12740 18564
rect 13468 19180 13524 19236
rect 12908 17666 12964 17668
rect 12908 17614 12910 17666
rect 12910 17614 12962 17666
rect 12962 17614 12964 17666
rect 12908 17612 12964 17614
rect 13020 18732 13076 18788
rect 12460 17442 12516 17444
rect 12460 17390 12462 17442
rect 12462 17390 12514 17442
rect 12514 17390 12516 17442
rect 12460 17388 12516 17390
rect 12796 17052 12852 17108
rect 12684 16994 12740 16996
rect 12684 16942 12686 16994
rect 12686 16942 12738 16994
rect 12738 16942 12740 16994
rect 12684 16940 12740 16942
rect 12012 16882 12068 16884
rect 12012 16830 12014 16882
rect 12014 16830 12066 16882
rect 12066 16830 12068 16882
rect 12012 16828 12068 16830
rect 11004 16604 11060 16660
rect 11676 16156 11732 16212
rect 9780 15706 9836 15708
rect 9780 15654 9782 15706
rect 9782 15654 9834 15706
rect 9834 15654 9836 15706
rect 9780 15652 9836 15654
rect 9884 15706 9940 15708
rect 9884 15654 9886 15706
rect 9886 15654 9938 15706
rect 9938 15654 9940 15706
rect 9884 15652 9940 15654
rect 9988 15706 10044 15708
rect 9988 15654 9990 15706
rect 9990 15654 10042 15706
rect 10042 15654 10044 15706
rect 9988 15652 10044 15654
rect 9212 14700 9268 14756
rect 6860 13746 6916 13748
rect 6860 13694 6862 13746
rect 6862 13694 6914 13746
rect 6914 13694 6916 13746
rect 6860 13692 6916 13694
rect 5496 13354 5552 13356
rect 5496 13302 5498 13354
rect 5498 13302 5550 13354
rect 5550 13302 5552 13354
rect 5496 13300 5552 13302
rect 5600 13354 5656 13356
rect 5600 13302 5602 13354
rect 5602 13302 5654 13354
rect 5654 13302 5656 13354
rect 5600 13300 5656 13302
rect 5704 13354 5760 13356
rect 5704 13302 5706 13354
rect 5706 13302 5758 13354
rect 5758 13302 5760 13354
rect 5704 13300 5760 13302
rect 6972 12850 7028 12852
rect 6972 12798 6974 12850
rect 6974 12798 7026 12850
rect 7026 12798 7028 12850
rect 6972 12796 7028 12798
rect 6300 12572 6356 12628
rect 6188 12460 6244 12516
rect 4844 12348 4900 12404
rect 4172 8428 4228 8484
rect 5496 11786 5552 11788
rect 5496 11734 5498 11786
rect 5498 11734 5550 11786
rect 5550 11734 5552 11786
rect 5496 11732 5552 11734
rect 5600 11786 5656 11788
rect 5600 11734 5602 11786
rect 5602 11734 5654 11786
rect 5654 11734 5656 11786
rect 5600 11732 5656 11734
rect 5704 11786 5760 11788
rect 5704 11734 5706 11786
rect 5706 11734 5758 11786
rect 5758 11734 5760 11786
rect 5704 11732 5760 11734
rect 7196 13132 7252 13188
rect 7420 13132 7476 13188
rect 7868 13692 7924 13748
rect 7532 12738 7588 12740
rect 7532 12686 7534 12738
rect 7534 12686 7586 12738
rect 7586 12686 7588 12738
rect 7532 12684 7588 12686
rect 7756 12348 7812 12404
rect 9780 14138 9836 14140
rect 9780 14086 9782 14138
rect 9782 14086 9834 14138
rect 9834 14086 9836 14138
rect 9780 14084 9836 14086
rect 9884 14138 9940 14140
rect 9884 14086 9886 14138
rect 9886 14086 9938 14138
rect 9938 14086 9940 14138
rect 9884 14084 9940 14086
rect 9988 14138 10044 14140
rect 9988 14086 9990 14138
rect 9990 14086 10042 14138
rect 10042 14086 10044 14138
rect 9988 14084 10044 14086
rect 8092 12962 8148 12964
rect 8092 12910 8094 12962
rect 8094 12910 8146 12962
rect 8146 12910 8148 12962
rect 8092 12908 8148 12910
rect 8316 13244 8372 13300
rect 8540 13132 8596 13188
rect 8876 12908 8932 12964
rect 8764 12796 8820 12852
rect 8428 12738 8484 12740
rect 8428 12686 8430 12738
rect 8430 12686 8482 12738
rect 8482 12686 8484 12738
rect 8428 12684 8484 12686
rect 8316 12572 8372 12628
rect 7644 12178 7700 12180
rect 7644 12126 7646 12178
rect 7646 12126 7698 12178
rect 7698 12126 7700 12178
rect 7644 12124 7700 12126
rect 7980 11564 8036 11620
rect 5496 10218 5552 10220
rect 5496 10166 5498 10218
rect 5498 10166 5550 10218
rect 5550 10166 5552 10218
rect 5496 10164 5552 10166
rect 5600 10218 5656 10220
rect 5600 10166 5602 10218
rect 5602 10166 5654 10218
rect 5654 10166 5656 10218
rect 5600 10164 5656 10166
rect 5704 10218 5760 10220
rect 5704 10166 5706 10218
rect 5706 10166 5758 10218
rect 5758 10166 5760 10218
rect 5704 10164 5760 10166
rect 7644 10108 7700 10164
rect 6748 9884 6804 9940
rect 5496 8650 5552 8652
rect 5496 8598 5498 8650
rect 5498 8598 5550 8650
rect 5550 8598 5552 8650
rect 5496 8596 5552 8598
rect 5600 8650 5656 8652
rect 5600 8598 5602 8650
rect 5602 8598 5654 8650
rect 5654 8598 5656 8650
rect 5600 8596 5656 8598
rect 5704 8650 5760 8652
rect 5704 8598 5706 8650
rect 5706 8598 5758 8650
rect 5758 8598 5760 8650
rect 5704 8596 5760 8598
rect 7084 8876 7140 8932
rect 8428 12460 8484 12516
rect 8540 12124 8596 12180
rect 11228 14588 11284 14644
rect 11340 13244 11396 13300
rect 11564 13020 11620 13076
rect 9100 12124 9156 12180
rect 10332 12962 10388 12964
rect 10332 12910 10334 12962
rect 10334 12910 10386 12962
rect 10386 12910 10388 12962
rect 10332 12908 10388 12910
rect 9996 12796 10052 12852
rect 10780 12850 10836 12852
rect 10780 12798 10782 12850
rect 10782 12798 10834 12850
rect 10834 12798 10836 12850
rect 10780 12796 10836 12798
rect 9780 12570 9836 12572
rect 9780 12518 9782 12570
rect 9782 12518 9834 12570
rect 9834 12518 9836 12570
rect 9780 12516 9836 12518
rect 9884 12570 9940 12572
rect 9884 12518 9886 12570
rect 9886 12518 9938 12570
rect 9938 12518 9940 12570
rect 9884 12516 9940 12518
rect 9988 12570 10044 12572
rect 9988 12518 9990 12570
rect 9990 12518 10042 12570
rect 10042 12518 10044 12570
rect 9988 12516 10044 12518
rect 8988 11564 9044 11620
rect 8204 9884 8260 9940
rect 8428 10332 8484 10388
rect 10444 12684 10500 12740
rect 10108 12012 10164 12068
rect 10332 12124 10388 12180
rect 9772 11452 9828 11508
rect 9884 11564 9940 11620
rect 9660 11228 9716 11284
rect 9436 11170 9492 11172
rect 9436 11118 9438 11170
rect 9438 11118 9490 11170
rect 9490 11118 9492 11170
rect 9436 11116 9492 11118
rect 10556 11506 10612 11508
rect 10556 11454 10558 11506
rect 10558 11454 10610 11506
rect 10610 11454 10612 11506
rect 10556 11452 10612 11454
rect 11564 12572 11620 12628
rect 11788 14642 11844 14644
rect 11788 14590 11790 14642
rect 11790 14590 11842 14642
rect 11842 14590 11844 14642
rect 11788 14588 11844 14590
rect 13132 18284 13188 18340
rect 14064 21194 14120 21196
rect 14064 21142 14066 21194
rect 14066 21142 14118 21194
rect 14118 21142 14120 21194
rect 14064 21140 14120 21142
rect 14168 21194 14224 21196
rect 14168 21142 14170 21194
rect 14170 21142 14222 21194
rect 14222 21142 14224 21194
rect 14168 21140 14224 21142
rect 14272 21194 14328 21196
rect 14272 21142 14274 21194
rect 14274 21142 14326 21194
rect 14326 21142 14328 21194
rect 14272 21140 14328 21142
rect 13804 20802 13860 20804
rect 13804 20750 13806 20802
rect 13806 20750 13858 20802
rect 13858 20750 13860 20802
rect 13804 20748 13860 20750
rect 13692 19404 13748 19460
rect 13692 19122 13748 19124
rect 13692 19070 13694 19122
rect 13694 19070 13746 19122
rect 13746 19070 13748 19122
rect 13692 19068 13748 19070
rect 13804 18844 13860 18900
rect 13468 18508 13524 18564
rect 13580 18450 13636 18452
rect 13580 18398 13582 18450
rect 13582 18398 13634 18450
rect 13634 18398 13636 18450
rect 13580 18396 13636 18398
rect 13580 16940 13636 16996
rect 13244 16828 13300 16884
rect 14064 19626 14120 19628
rect 14064 19574 14066 19626
rect 14066 19574 14118 19626
rect 14118 19574 14120 19626
rect 14064 19572 14120 19574
rect 14168 19626 14224 19628
rect 14168 19574 14170 19626
rect 14170 19574 14222 19626
rect 14222 19574 14224 19626
rect 14168 19572 14224 19574
rect 14272 19626 14328 19628
rect 14272 19574 14274 19626
rect 14274 19574 14326 19626
rect 14326 19574 14328 19626
rect 14272 19572 14328 19574
rect 14812 24892 14868 24948
rect 15484 27692 15540 27748
rect 16380 28924 16436 28980
rect 17500 32508 17556 32564
rect 17388 31836 17444 31892
rect 16716 31106 16772 31108
rect 16716 31054 16718 31106
rect 16718 31054 16770 31106
rect 16770 31054 16772 31106
rect 16716 31052 16772 31054
rect 17612 32396 17668 32452
rect 17724 31724 17780 31780
rect 17500 31276 17556 31332
rect 17388 31052 17444 31108
rect 17612 31106 17668 31108
rect 17612 31054 17614 31106
rect 17614 31054 17666 31106
rect 17666 31054 17668 31106
rect 17612 31052 17668 31054
rect 17500 30940 17556 30996
rect 17724 30380 17780 30436
rect 16828 29596 16884 29652
rect 18348 32954 18404 32956
rect 18348 32902 18350 32954
rect 18350 32902 18402 32954
rect 18402 32902 18404 32954
rect 18348 32900 18404 32902
rect 18452 32954 18508 32956
rect 18452 32902 18454 32954
rect 18454 32902 18506 32954
rect 18506 32902 18508 32954
rect 18452 32900 18508 32902
rect 18556 32954 18612 32956
rect 18556 32902 18558 32954
rect 18558 32902 18610 32954
rect 18610 32902 18612 32954
rect 18556 32900 18612 32902
rect 18284 32620 18340 32676
rect 18844 31724 18900 31780
rect 18348 31386 18404 31388
rect 18348 31334 18350 31386
rect 18350 31334 18402 31386
rect 18402 31334 18404 31386
rect 18348 31332 18404 31334
rect 18452 31386 18508 31388
rect 18452 31334 18454 31386
rect 18454 31334 18506 31386
rect 18506 31334 18508 31386
rect 18452 31332 18508 31334
rect 18556 31386 18612 31388
rect 18556 31334 18558 31386
rect 18558 31334 18610 31386
rect 18610 31334 18612 31386
rect 18556 31332 18612 31334
rect 17948 31164 18004 31220
rect 18732 31106 18788 31108
rect 18732 31054 18734 31106
rect 18734 31054 18786 31106
rect 18786 31054 18788 31106
rect 18732 31052 18788 31054
rect 18396 30994 18452 30996
rect 18396 30942 18398 30994
rect 18398 30942 18450 30994
rect 18450 30942 18452 30994
rect 18396 30940 18452 30942
rect 20636 33516 20692 33572
rect 19516 31164 19572 31220
rect 19852 32732 19908 32788
rect 16940 29484 16996 29540
rect 19068 31106 19124 31108
rect 19068 31054 19070 31106
rect 19070 31054 19122 31106
rect 19122 31054 19124 31106
rect 19068 31052 19124 31054
rect 18348 29818 18404 29820
rect 18348 29766 18350 29818
rect 18350 29766 18402 29818
rect 18402 29766 18404 29818
rect 18348 29764 18404 29766
rect 18452 29818 18508 29820
rect 18452 29766 18454 29818
rect 18454 29766 18506 29818
rect 18506 29766 18508 29818
rect 18452 29764 18508 29766
rect 18556 29818 18612 29820
rect 18556 29766 18558 29818
rect 18558 29766 18610 29818
rect 18610 29766 18612 29818
rect 18556 29764 18612 29766
rect 18844 29538 18900 29540
rect 18844 29486 18846 29538
rect 18846 29486 18898 29538
rect 18898 29486 18900 29538
rect 18844 29484 18900 29486
rect 17276 29426 17332 29428
rect 17276 29374 17278 29426
rect 17278 29374 17330 29426
rect 17330 29374 17332 29426
rect 17276 29372 17332 29374
rect 16604 29314 16660 29316
rect 16604 29262 16606 29314
rect 16606 29262 16658 29314
rect 16658 29262 16660 29314
rect 16604 29260 16660 29262
rect 16604 29036 16660 29092
rect 15708 27244 15764 27300
rect 15260 26290 15316 26292
rect 15260 26238 15262 26290
rect 15262 26238 15314 26290
rect 15314 26238 15316 26290
rect 15260 26236 15316 26238
rect 15708 26460 15764 26516
rect 16044 27692 16100 27748
rect 15820 26348 15876 26404
rect 15484 25788 15540 25844
rect 14700 21474 14756 21476
rect 14700 21422 14702 21474
rect 14702 21422 14754 21474
rect 14754 21422 14756 21474
rect 14700 21420 14756 21422
rect 14588 20802 14644 20804
rect 14588 20750 14590 20802
rect 14590 20750 14642 20802
rect 14642 20750 14644 20802
rect 14588 20748 14644 20750
rect 15596 24722 15652 24724
rect 15596 24670 15598 24722
rect 15598 24670 15650 24722
rect 15650 24670 15652 24722
rect 15596 24668 15652 24670
rect 16156 26290 16212 26292
rect 16156 26238 16158 26290
rect 16158 26238 16210 26290
rect 16210 26238 16212 26290
rect 16156 26236 16212 26238
rect 17164 29148 17220 29204
rect 17052 29036 17108 29092
rect 17388 29148 17444 29204
rect 16940 28530 16996 28532
rect 16940 28478 16942 28530
rect 16942 28478 16994 28530
rect 16994 28478 16996 28530
rect 16940 28476 16996 28478
rect 17500 28700 17556 28756
rect 16380 27356 16436 27412
rect 16828 26962 16884 26964
rect 16828 26910 16830 26962
rect 16830 26910 16882 26962
rect 16882 26910 16884 26962
rect 16828 26908 16884 26910
rect 16940 26684 16996 26740
rect 16492 26124 16548 26180
rect 16716 26290 16772 26292
rect 16716 26238 16718 26290
rect 16718 26238 16770 26290
rect 16770 26238 16772 26290
rect 16716 26236 16772 26238
rect 16268 25788 16324 25844
rect 16716 25676 16772 25732
rect 17500 28252 17556 28308
rect 17388 27970 17444 27972
rect 17388 27918 17390 27970
rect 17390 27918 17442 27970
rect 17442 27918 17444 27970
rect 17388 27916 17444 27918
rect 17836 29372 17892 29428
rect 18620 29426 18676 29428
rect 18620 29374 18622 29426
rect 18622 29374 18674 29426
rect 18674 29374 18676 29426
rect 18620 29372 18676 29374
rect 17724 29260 17780 29316
rect 18060 29314 18116 29316
rect 18060 29262 18062 29314
rect 18062 29262 18114 29314
rect 18114 29262 18116 29314
rect 18060 29260 18116 29262
rect 17836 29202 17892 29204
rect 17836 29150 17838 29202
rect 17838 29150 17890 29202
rect 17890 29150 17892 29202
rect 17836 29148 17892 29150
rect 17836 28924 17892 28980
rect 17612 28140 17668 28196
rect 17724 28252 17780 28308
rect 17724 27804 17780 27860
rect 17500 27020 17556 27076
rect 17164 26348 17220 26404
rect 17276 26908 17332 26964
rect 16716 24722 16772 24724
rect 16716 24670 16718 24722
rect 16718 24670 16770 24722
rect 16770 24670 16772 24722
rect 16716 24668 16772 24670
rect 17052 24668 17108 24724
rect 17164 24556 17220 24612
rect 17164 23324 17220 23380
rect 16044 22370 16100 22372
rect 16044 22318 16046 22370
rect 16046 22318 16098 22370
rect 16098 22318 16100 22370
rect 16044 22316 16100 22318
rect 15484 21756 15540 21812
rect 14700 19740 14756 19796
rect 15260 21308 15316 21364
rect 14924 20690 14980 20692
rect 14924 20638 14926 20690
rect 14926 20638 14978 20690
rect 14978 20638 14980 20690
rect 14924 20636 14980 20638
rect 15708 20636 15764 20692
rect 15260 20188 15316 20244
rect 14812 19404 14868 19460
rect 14140 19234 14196 19236
rect 14140 19182 14142 19234
rect 14142 19182 14194 19234
rect 14194 19182 14196 19234
rect 14140 19180 14196 19182
rect 15036 19180 15092 19236
rect 14700 18956 14756 19012
rect 14588 18844 14644 18900
rect 13804 17554 13860 17556
rect 13804 17502 13806 17554
rect 13806 17502 13858 17554
rect 13858 17502 13860 17554
rect 13804 17500 13860 17502
rect 14064 18058 14120 18060
rect 14064 18006 14066 18058
rect 14066 18006 14118 18058
rect 14118 18006 14120 18058
rect 14064 18004 14120 18006
rect 14168 18058 14224 18060
rect 14168 18006 14170 18058
rect 14170 18006 14222 18058
rect 14222 18006 14224 18058
rect 14168 18004 14224 18006
rect 14272 18058 14328 18060
rect 14272 18006 14274 18058
rect 14274 18006 14326 18058
rect 14326 18006 14328 18058
rect 14272 18004 14328 18006
rect 14028 17666 14084 17668
rect 14028 17614 14030 17666
rect 14030 17614 14082 17666
rect 14082 17614 14084 17666
rect 14028 17612 14084 17614
rect 14252 17554 14308 17556
rect 14252 17502 14254 17554
rect 14254 17502 14306 17554
rect 14306 17502 14308 17554
rect 14252 17500 14308 17502
rect 16828 21980 16884 22036
rect 16604 21420 16660 21476
rect 17052 21308 17108 21364
rect 16940 20636 16996 20692
rect 16156 20076 16212 20132
rect 15932 19964 15988 20020
rect 15148 19010 15204 19012
rect 15148 18958 15150 19010
rect 15150 18958 15202 19010
rect 15202 18958 15204 19010
rect 15148 18956 15204 18958
rect 14924 18844 14980 18900
rect 15932 19404 15988 19460
rect 16268 19404 16324 19460
rect 17388 26684 17444 26740
rect 19404 30994 19460 30996
rect 19404 30942 19406 30994
rect 19406 30942 19458 30994
rect 19458 30942 19460 30994
rect 19404 30940 19460 30942
rect 20524 32562 20580 32564
rect 20524 32510 20526 32562
rect 20526 32510 20578 32562
rect 20578 32510 20580 32562
rect 20524 32508 20580 32510
rect 20972 32508 21028 32564
rect 20412 31890 20468 31892
rect 20412 31838 20414 31890
rect 20414 31838 20466 31890
rect 20466 31838 20468 31890
rect 20412 31836 20468 31838
rect 20076 31612 20132 31668
rect 19404 30268 19460 30324
rect 19068 29650 19124 29652
rect 19068 29598 19070 29650
rect 19070 29598 19122 29650
rect 19122 29598 19124 29650
rect 19068 29596 19124 29598
rect 18956 28924 19012 28980
rect 19292 28700 19348 28756
rect 18732 28588 18788 28644
rect 18956 28364 19012 28420
rect 18172 28252 18228 28308
rect 18348 28250 18404 28252
rect 18348 28198 18350 28250
rect 18350 28198 18402 28250
rect 18402 28198 18404 28250
rect 18348 28196 18404 28198
rect 18452 28250 18508 28252
rect 18452 28198 18454 28250
rect 18454 28198 18506 28250
rect 18506 28198 18508 28250
rect 18452 28196 18508 28198
rect 18556 28250 18612 28252
rect 18556 28198 18558 28250
rect 18558 28198 18610 28250
rect 18610 28198 18612 28250
rect 18556 28196 18612 28198
rect 18844 28252 18900 28308
rect 17836 27020 17892 27076
rect 19068 27692 19124 27748
rect 18284 27244 18340 27300
rect 18508 27244 18564 27300
rect 18956 27244 19012 27300
rect 18844 27132 18900 27188
rect 18732 27020 18788 27076
rect 18284 26962 18340 26964
rect 18284 26910 18286 26962
rect 18286 26910 18338 26962
rect 18338 26910 18340 26962
rect 18284 26908 18340 26910
rect 18348 26682 18404 26684
rect 18348 26630 18350 26682
rect 18350 26630 18402 26682
rect 18402 26630 18404 26682
rect 18348 26628 18404 26630
rect 18452 26682 18508 26684
rect 18452 26630 18454 26682
rect 18454 26630 18506 26682
rect 18506 26630 18508 26682
rect 18452 26628 18508 26630
rect 18556 26682 18612 26684
rect 18556 26630 18558 26682
rect 18558 26630 18610 26682
rect 18610 26630 18612 26682
rect 18556 26628 18612 26630
rect 17724 26290 17780 26292
rect 17724 26238 17726 26290
rect 17726 26238 17778 26290
rect 17778 26238 17780 26290
rect 17724 26236 17780 26238
rect 18396 26514 18452 26516
rect 18396 26462 18398 26514
rect 18398 26462 18450 26514
rect 18450 26462 18452 26514
rect 18396 26460 18452 26462
rect 19740 28812 19796 28868
rect 19292 28252 19348 28308
rect 19516 28140 19572 28196
rect 19404 27804 19460 27860
rect 19516 27916 19572 27972
rect 20636 31500 20692 31556
rect 20188 30940 20244 30996
rect 20524 30828 20580 30884
rect 20412 30322 20468 30324
rect 20412 30270 20414 30322
rect 20414 30270 20466 30322
rect 20466 30270 20468 30322
rect 20412 30268 20468 30270
rect 20412 29820 20468 29876
rect 19740 27580 19796 27636
rect 19852 27468 19908 27524
rect 19852 27020 19908 27076
rect 19964 28476 20020 28532
rect 19740 26962 19796 26964
rect 19740 26910 19742 26962
rect 19742 26910 19794 26962
rect 19794 26910 19796 26962
rect 19740 26908 19796 26910
rect 18060 26236 18116 26292
rect 17388 25506 17444 25508
rect 17388 25454 17390 25506
rect 17390 25454 17442 25506
rect 17442 25454 17444 25506
rect 17388 25452 17444 25454
rect 17724 25564 17780 25620
rect 18508 25788 18564 25844
rect 19628 26796 19684 26852
rect 19068 26348 19124 26404
rect 18508 25340 18564 25396
rect 18844 25394 18900 25396
rect 18844 25342 18846 25394
rect 18846 25342 18898 25394
rect 18898 25342 18900 25394
rect 18844 25340 18900 25342
rect 18396 25228 18452 25284
rect 18348 25114 18404 25116
rect 18348 25062 18350 25114
rect 18350 25062 18402 25114
rect 18402 25062 18404 25114
rect 18348 25060 18404 25062
rect 18452 25114 18508 25116
rect 18452 25062 18454 25114
rect 18454 25062 18506 25114
rect 18506 25062 18508 25114
rect 18452 25060 18508 25062
rect 18556 25114 18612 25116
rect 18556 25062 18558 25114
rect 18558 25062 18610 25114
rect 18610 25062 18612 25114
rect 18556 25060 18612 25062
rect 17724 24556 17780 24612
rect 18172 24610 18228 24612
rect 18172 24558 18174 24610
rect 18174 24558 18226 24610
rect 18226 24558 18228 24610
rect 18172 24556 18228 24558
rect 17948 23772 18004 23828
rect 17724 23378 17780 23380
rect 17724 23326 17726 23378
rect 17726 23326 17778 23378
rect 17778 23326 17780 23378
rect 17724 23324 17780 23326
rect 18844 24556 18900 24612
rect 18348 23546 18404 23548
rect 18348 23494 18350 23546
rect 18350 23494 18402 23546
rect 18402 23494 18404 23546
rect 18348 23492 18404 23494
rect 18452 23546 18508 23548
rect 18452 23494 18454 23546
rect 18454 23494 18506 23546
rect 18506 23494 18508 23546
rect 18452 23492 18508 23494
rect 18556 23546 18612 23548
rect 18556 23494 18558 23546
rect 18558 23494 18610 23546
rect 18610 23494 18612 23546
rect 18556 23492 18612 23494
rect 18732 23548 18788 23604
rect 17500 22316 17556 22372
rect 17836 21474 17892 21476
rect 17836 21422 17838 21474
rect 17838 21422 17890 21474
rect 17890 21422 17892 21474
rect 17836 21420 17892 21422
rect 18060 22540 18116 22596
rect 18172 21980 18228 22036
rect 18348 21978 18404 21980
rect 18348 21926 18350 21978
rect 18350 21926 18402 21978
rect 18402 21926 18404 21978
rect 18348 21924 18404 21926
rect 18452 21978 18508 21980
rect 18452 21926 18454 21978
rect 18454 21926 18506 21978
rect 18506 21926 18508 21978
rect 18452 21924 18508 21926
rect 18556 21978 18612 21980
rect 18556 21926 18558 21978
rect 18558 21926 18610 21978
rect 18610 21926 18612 21978
rect 18556 21924 18612 21926
rect 17948 21308 18004 21364
rect 17836 20690 17892 20692
rect 17836 20638 17838 20690
rect 17838 20638 17890 20690
rect 17890 20638 17892 20690
rect 17836 20636 17892 20638
rect 19180 25618 19236 25620
rect 19180 25566 19182 25618
rect 19182 25566 19234 25618
rect 19234 25566 19236 25618
rect 19180 25564 19236 25566
rect 19404 25506 19460 25508
rect 19404 25454 19406 25506
rect 19406 25454 19458 25506
rect 19458 25454 19460 25506
rect 19404 25452 19460 25454
rect 19740 26572 19796 26628
rect 19740 26124 19796 26180
rect 19628 25730 19684 25732
rect 19628 25678 19630 25730
rect 19630 25678 19682 25730
rect 19682 25678 19684 25730
rect 19628 25676 19684 25678
rect 19740 25452 19796 25508
rect 19516 25340 19572 25396
rect 20300 28418 20356 28420
rect 20300 28366 20302 28418
rect 20302 28366 20354 28418
rect 20354 28366 20356 28418
rect 20300 28364 20356 28366
rect 20748 31218 20804 31220
rect 20748 31166 20750 31218
rect 20750 31166 20802 31218
rect 20802 31166 20804 31218
rect 20748 31164 20804 31166
rect 21196 31724 21252 31780
rect 20748 30210 20804 30212
rect 20748 30158 20750 30210
rect 20750 30158 20802 30210
rect 20802 30158 20804 30210
rect 20748 30156 20804 30158
rect 20748 27916 20804 27972
rect 20524 27746 20580 27748
rect 20524 27694 20526 27746
rect 20526 27694 20578 27746
rect 20578 27694 20580 27746
rect 20524 27692 20580 27694
rect 20412 27580 20468 27636
rect 20076 27356 20132 27412
rect 20076 27020 20132 27076
rect 20076 26572 20132 26628
rect 20188 26684 20244 26740
rect 20524 27074 20580 27076
rect 20524 27022 20526 27074
rect 20526 27022 20578 27074
rect 20578 27022 20580 27074
rect 20524 27020 20580 27022
rect 21420 31612 21476 31668
rect 22632 33738 22688 33740
rect 22632 33686 22634 33738
rect 22634 33686 22686 33738
rect 22686 33686 22688 33738
rect 22632 33684 22688 33686
rect 22736 33738 22792 33740
rect 22736 33686 22738 33738
rect 22738 33686 22790 33738
rect 22790 33686 22792 33738
rect 22736 33684 22792 33686
rect 22840 33738 22896 33740
rect 22840 33686 22842 33738
rect 22842 33686 22894 33738
rect 22894 33686 22896 33738
rect 22840 33684 22896 33686
rect 21756 32396 21812 32452
rect 22428 32284 22484 32340
rect 22632 32170 22688 32172
rect 22632 32118 22634 32170
rect 22634 32118 22686 32170
rect 22686 32118 22688 32170
rect 22632 32116 22688 32118
rect 22736 32170 22792 32172
rect 22736 32118 22738 32170
rect 22738 32118 22790 32170
rect 22790 32118 22792 32170
rect 22736 32116 22792 32118
rect 22840 32170 22896 32172
rect 22840 32118 22842 32170
rect 22842 32118 22894 32170
rect 22894 32118 22896 32170
rect 22840 32116 22896 32118
rect 21756 31778 21812 31780
rect 21756 31726 21758 31778
rect 21758 31726 21810 31778
rect 21810 31726 21812 31778
rect 21756 31724 21812 31726
rect 21532 30940 21588 30996
rect 21196 29820 21252 29876
rect 21196 29538 21252 29540
rect 21196 29486 21198 29538
rect 21198 29486 21250 29538
rect 21250 29486 21252 29538
rect 21196 29484 21252 29486
rect 21308 28700 21364 28756
rect 20972 27858 21028 27860
rect 20972 27806 20974 27858
rect 20974 27806 21026 27858
rect 21026 27806 21028 27858
rect 20972 27804 21028 27806
rect 21196 28588 21252 28644
rect 20860 26908 20916 26964
rect 20636 26572 20692 26628
rect 20412 26290 20468 26292
rect 20412 26238 20414 26290
rect 20414 26238 20466 26290
rect 20466 26238 20468 26290
rect 20412 26236 20468 26238
rect 20412 25788 20468 25844
rect 20188 25228 20244 25284
rect 19180 23884 19236 23940
rect 18956 23826 19012 23828
rect 18956 23774 18958 23826
rect 18958 23774 19010 23826
rect 19010 23774 19012 23826
rect 18956 23772 19012 23774
rect 19852 23884 19908 23940
rect 19292 23548 19348 23604
rect 19516 23772 19572 23828
rect 18732 21756 18788 21812
rect 18060 20690 18116 20692
rect 18060 20638 18062 20690
rect 18062 20638 18114 20690
rect 18114 20638 18116 20690
rect 18060 20636 18116 20638
rect 16604 20130 16660 20132
rect 16604 20078 16606 20130
rect 16606 20078 16658 20130
rect 16658 20078 16660 20130
rect 16604 20076 16660 20078
rect 16716 19964 16772 20020
rect 15932 19234 15988 19236
rect 15932 19182 15934 19234
rect 15934 19182 15986 19234
rect 15986 19182 15988 19234
rect 15932 19180 15988 19182
rect 15596 18284 15652 18340
rect 15596 18060 15652 18116
rect 15260 17724 15316 17780
rect 13916 16828 13972 16884
rect 15260 16828 15316 16884
rect 14064 16490 14120 16492
rect 14064 16438 14066 16490
rect 14066 16438 14118 16490
rect 14118 16438 14120 16490
rect 14064 16436 14120 16438
rect 14168 16490 14224 16492
rect 14168 16438 14170 16490
rect 14170 16438 14222 16490
rect 14222 16438 14224 16490
rect 14168 16436 14224 16438
rect 14272 16490 14328 16492
rect 14272 16438 14274 16490
rect 14274 16438 14326 16490
rect 14326 16438 14328 16490
rect 14272 16436 14328 16438
rect 13804 16268 13860 16324
rect 13468 15538 13524 15540
rect 13468 15486 13470 15538
rect 13470 15486 13522 15538
rect 13522 15486 13524 15538
rect 13468 15484 13524 15486
rect 11788 13244 11844 13300
rect 12460 12962 12516 12964
rect 12460 12910 12462 12962
rect 12462 12910 12514 12962
rect 12514 12910 12516 12962
rect 12460 12908 12516 12910
rect 12236 12850 12292 12852
rect 12236 12798 12238 12850
rect 12238 12798 12290 12850
rect 12290 12798 12292 12850
rect 12236 12796 12292 12798
rect 11564 12012 11620 12068
rect 12460 12178 12516 12180
rect 12460 12126 12462 12178
rect 12462 12126 12514 12178
rect 12514 12126 12516 12178
rect 12460 12124 12516 12126
rect 11004 11394 11060 11396
rect 11004 11342 11006 11394
rect 11006 11342 11058 11394
rect 11058 11342 11060 11394
rect 11004 11340 11060 11342
rect 11452 11394 11508 11396
rect 11452 11342 11454 11394
rect 11454 11342 11506 11394
rect 11506 11342 11508 11394
rect 11452 11340 11508 11342
rect 11900 11394 11956 11396
rect 11900 11342 11902 11394
rect 11902 11342 11954 11394
rect 11954 11342 11956 11394
rect 11900 11340 11956 11342
rect 10668 11282 10724 11284
rect 10668 11230 10670 11282
rect 10670 11230 10722 11282
rect 10722 11230 10724 11282
rect 10668 11228 10724 11230
rect 10332 11116 10388 11172
rect 9780 11002 9836 11004
rect 9780 10950 9782 11002
rect 9782 10950 9834 11002
rect 9834 10950 9836 11002
rect 9780 10948 9836 10950
rect 9884 11002 9940 11004
rect 9884 10950 9886 11002
rect 9886 10950 9938 11002
rect 9938 10950 9940 11002
rect 9884 10948 9940 10950
rect 9988 11002 10044 11004
rect 9988 10950 9990 11002
rect 9990 10950 10042 11002
rect 10042 10950 10044 11002
rect 9988 10948 10044 10950
rect 9660 10386 9716 10388
rect 9660 10334 9662 10386
rect 9662 10334 9714 10386
rect 9714 10334 9716 10386
rect 9660 10332 9716 10334
rect 9436 10108 9492 10164
rect 8540 8876 8596 8932
rect 6748 8428 6804 8484
rect 7644 8428 7700 8484
rect 5964 7980 6020 8036
rect 5496 7082 5552 7084
rect 5496 7030 5498 7082
rect 5498 7030 5550 7082
rect 5550 7030 5552 7082
rect 5496 7028 5552 7030
rect 5600 7082 5656 7084
rect 5600 7030 5602 7082
rect 5602 7030 5654 7082
rect 5654 7030 5656 7082
rect 5600 7028 5656 7030
rect 5704 7082 5760 7084
rect 5704 7030 5706 7082
rect 5706 7030 5758 7082
rect 5758 7030 5760 7082
rect 5704 7028 5760 7030
rect 8092 8258 8148 8260
rect 8092 8206 8094 8258
rect 8094 8206 8146 8258
rect 8146 8206 8148 8258
rect 8092 8204 8148 8206
rect 6300 7474 6356 7476
rect 6300 7422 6302 7474
rect 6302 7422 6354 7474
rect 6354 7422 6356 7474
rect 6300 7420 6356 7422
rect 6076 6748 6132 6804
rect 6524 7308 6580 7364
rect 5964 6018 6020 6020
rect 5964 5966 5966 6018
rect 5966 5966 6018 6018
rect 6018 5966 6020 6018
rect 5964 5964 6020 5966
rect 5496 5514 5552 5516
rect 5496 5462 5498 5514
rect 5498 5462 5550 5514
rect 5550 5462 5552 5514
rect 5496 5460 5552 5462
rect 5600 5514 5656 5516
rect 5600 5462 5602 5514
rect 5602 5462 5654 5514
rect 5654 5462 5656 5514
rect 5600 5460 5656 5462
rect 5704 5514 5760 5516
rect 5704 5462 5706 5514
rect 5706 5462 5758 5514
rect 5758 5462 5760 5514
rect 5704 5460 5760 5462
rect 5740 5180 5796 5236
rect 5404 4508 5460 4564
rect 6076 5122 6132 5124
rect 6076 5070 6078 5122
rect 6078 5070 6130 5122
rect 6130 5070 6132 5122
rect 6076 5068 6132 5070
rect 5964 4508 6020 4564
rect 6188 4956 6244 5012
rect 5496 3946 5552 3948
rect 5496 3894 5498 3946
rect 5498 3894 5550 3946
rect 5550 3894 5552 3946
rect 5496 3892 5552 3894
rect 5600 3946 5656 3948
rect 5600 3894 5602 3946
rect 5602 3894 5654 3946
rect 5654 3894 5656 3946
rect 5600 3892 5656 3894
rect 5704 3946 5760 3948
rect 5704 3894 5706 3946
rect 5706 3894 5758 3946
rect 5758 3894 5760 3946
rect 5704 3892 5760 3894
rect 3948 3388 4004 3444
rect 4956 3388 5012 3444
rect 7420 7532 7476 7588
rect 7196 7474 7252 7476
rect 7196 7422 7198 7474
rect 7198 7422 7250 7474
rect 7250 7422 7252 7474
rect 7196 7420 7252 7422
rect 9100 8258 9156 8260
rect 9100 8206 9102 8258
rect 9102 8206 9154 8258
rect 9154 8206 9156 8258
rect 9100 8204 9156 8206
rect 8540 8092 8596 8148
rect 7980 7586 8036 7588
rect 7980 7534 7982 7586
rect 7982 7534 8034 7586
rect 8034 7534 8036 7586
rect 7980 7532 8036 7534
rect 8428 7532 8484 7588
rect 8092 7362 8148 7364
rect 8092 7310 8094 7362
rect 8094 7310 8146 7362
rect 8146 7310 8148 7362
rect 8092 7308 8148 7310
rect 7308 6748 7364 6804
rect 6972 5740 7028 5796
rect 6412 4172 6468 4228
rect 9100 7698 9156 7700
rect 9100 7646 9102 7698
rect 9102 7646 9154 7698
rect 9154 7646 9156 7698
rect 9100 7644 9156 7646
rect 9548 8316 9604 8372
rect 9324 7308 9380 7364
rect 8652 6972 8708 7028
rect 9548 7586 9604 7588
rect 9548 7534 9550 7586
rect 9550 7534 9602 7586
rect 9602 7534 9604 7586
rect 9548 7532 9604 7534
rect 9436 6860 9492 6916
rect 8540 6748 8596 6804
rect 8204 5516 8260 5572
rect 7196 3724 7252 3780
rect 8988 5516 9044 5572
rect 10892 10498 10948 10500
rect 10892 10446 10894 10498
rect 10894 10446 10946 10498
rect 10946 10446 10948 10498
rect 10892 10444 10948 10446
rect 9780 9434 9836 9436
rect 9780 9382 9782 9434
rect 9782 9382 9834 9434
rect 9834 9382 9836 9434
rect 9780 9380 9836 9382
rect 9884 9434 9940 9436
rect 9884 9382 9886 9434
rect 9886 9382 9938 9434
rect 9938 9382 9940 9434
rect 9884 9380 9940 9382
rect 9988 9434 10044 9436
rect 9988 9382 9990 9434
rect 9990 9382 10042 9434
rect 10042 9382 10044 9434
rect 9988 9380 10044 9382
rect 9772 8370 9828 8372
rect 9772 8318 9774 8370
rect 9774 8318 9826 8370
rect 9826 8318 9828 8370
rect 9772 8316 9828 8318
rect 10332 8204 10388 8260
rect 9996 7980 10052 8036
rect 9780 7866 9836 7868
rect 9780 7814 9782 7866
rect 9782 7814 9834 7866
rect 9834 7814 9836 7866
rect 9780 7812 9836 7814
rect 9884 7866 9940 7868
rect 9884 7814 9886 7866
rect 9886 7814 9938 7866
rect 9938 7814 9940 7866
rect 9884 7812 9940 7814
rect 9988 7866 10044 7868
rect 9988 7814 9990 7866
rect 9990 7814 10042 7866
rect 10042 7814 10044 7866
rect 9988 7812 10044 7814
rect 9996 7308 10052 7364
rect 10220 7420 10276 7476
rect 9660 6972 9716 7028
rect 9548 5906 9604 5908
rect 9548 5854 9550 5906
rect 9550 5854 9602 5906
rect 9602 5854 9604 5906
rect 9548 5852 9604 5854
rect 9780 6298 9836 6300
rect 9780 6246 9782 6298
rect 9782 6246 9834 6298
rect 9834 6246 9836 6298
rect 9780 6244 9836 6246
rect 9884 6298 9940 6300
rect 9884 6246 9886 6298
rect 9886 6246 9938 6298
rect 9938 6246 9940 6298
rect 9884 6244 9940 6246
rect 9988 6298 10044 6300
rect 9988 6246 9990 6298
rect 9990 6246 10042 6298
rect 10042 6246 10044 6298
rect 9988 6244 10044 6246
rect 10108 5740 10164 5796
rect 10108 5516 10164 5572
rect 10780 7698 10836 7700
rect 10780 7646 10782 7698
rect 10782 7646 10834 7698
rect 10834 7646 10836 7698
rect 10780 7644 10836 7646
rect 13356 13580 13412 13636
rect 12908 13468 12964 13524
rect 12796 13074 12852 13076
rect 12796 13022 12798 13074
rect 12798 13022 12850 13074
rect 12850 13022 12852 13074
rect 12796 13020 12852 13022
rect 12796 11340 12852 11396
rect 12236 9602 12292 9604
rect 12236 9550 12238 9602
rect 12238 9550 12290 9602
rect 12290 9550 12292 9602
rect 12236 9548 12292 9550
rect 12124 8930 12180 8932
rect 12124 8878 12126 8930
rect 12126 8878 12178 8930
rect 12178 8878 12180 8930
rect 12124 8876 12180 8878
rect 10780 6018 10836 6020
rect 10780 5966 10782 6018
rect 10782 5966 10834 6018
rect 10834 5966 10836 6018
rect 10780 5964 10836 5966
rect 11004 5906 11060 5908
rect 11004 5854 11006 5906
rect 11006 5854 11058 5906
rect 11058 5854 11060 5906
rect 11004 5852 11060 5854
rect 9772 5180 9828 5236
rect 9884 5122 9940 5124
rect 9884 5070 9886 5122
rect 9886 5070 9938 5122
rect 9938 5070 9940 5122
rect 9884 5068 9940 5070
rect 9660 4898 9716 4900
rect 9660 4846 9662 4898
rect 9662 4846 9714 4898
rect 9714 4846 9716 4898
rect 9660 4844 9716 4846
rect 9324 4508 9380 4564
rect 9212 3724 9268 3780
rect 8316 3388 8372 3444
rect 9780 4730 9836 4732
rect 9780 4678 9782 4730
rect 9782 4678 9834 4730
rect 9834 4678 9836 4730
rect 9780 4676 9836 4678
rect 9884 4730 9940 4732
rect 9884 4678 9886 4730
rect 9886 4678 9938 4730
rect 9938 4678 9940 4730
rect 9884 4676 9940 4678
rect 9988 4730 10044 4732
rect 9988 4678 9990 4730
rect 9990 4678 10042 4730
rect 10042 4678 10044 4730
rect 9988 4676 10044 4678
rect 10444 4732 10500 4788
rect 9548 4226 9604 4228
rect 9548 4174 9550 4226
rect 9550 4174 9602 4226
rect 9602 4174 9604 4226
rect 9548 4172 9604 4174
rect 11452 7474 11508 7476
rect 11452 7422 11454 7474
rect 11454 7422 11506 7474
rect 11506 7422 11508 7474
rect 11452 7420 11508 7422
rect 11116 4508 11172 4564
rect 10444 4172 10500 4228
rect 9660 3332 9716 3388
rect 9780 3162 9836 3164
rect 9780 3110 9782 3162
rect 9782 3110 9834 3162
rect 9834 3110 9836 3162
rect 9780 3108 9836 3110
rect 9884 3162 9940 3164
rect 9884 3110 9886 3162
rect 9886 3110 9938 3162
rect 9938 3110 9940 3162
rect 9884 3108 9940 3110
rect 9988 3162 10044 3164
rect 9988 3110 9990 3162
rect 9990 3110 10042 3162
rect 10042 3110 10044 3162
rect 9988 3108 10044 3110
rect 11340 6018 11396 6020
rect 11340 5966 11342 6018
rect 11342 5966 11394 6018
rect 11394 5966 11396 6018
rect 11340 5964 11396 5966
rect 11564 5628 11620 5684
rect 12236 7644 12292 7700
rect 12460 6860 12516 6916
rect 13244 10444 13300 10500
rect 13132 9884 13188 9940
rect 12908 9826 12964 9828
rect 12908 9774 12910 9826
rect 12910 9774 12962 9826
rect 12962 9774 12964 9826
rect 12908 9772 12964 9774
rect 12460 5794 12516 5796
rect 12460 5742 12462 5794
rect 12462 5742 12514 5794
rect 12514 5742 12516 5794
rect 12460 5740 12516 5742
rect 11788 5068 11844 5124
rect 11676 4732 11732 4788
rect 12908 7980 12964 8036
rect 13244 6076 13300 6132
rect 12796 5852 12852 5908
rect 12796 5234 12852 5236
rect 12796 5182 12798 5234
rect 12798 5182 12850 5234
rect 12850 5182 12852 5234
rect 12796 5180 12852 5182
rect 13020 5628 13076 5684
rect 12460 4338 12516 4340
rect 12460 4286 12462 4338
rect 12462 4286 12514 4338
rect 12514 4286 12516 4338
rect 12460 4284 12516 4286
rect 12684 4844 12740 4900
rect 11676 4226 11732 4228
rect 11676 4174 11678 4226
rect 11678 4174 11730 4226
rect 11730 4174 11732 4226
rect 11676 4172 11732 4174
rect 12908 4226 12964 4228
rect 12908 4174 12910 4226
rect 12910 4174 12962 4226
rect 12962 4174 12964 4226
rect 12908 4172 12964 4174
rect 15260 16268 15316 16324
rect 15372 16210 15428 16212
rect 15372 16158 15374 16210
rect 15374 16158 15426 16210
rect 15426 16158 15428 16210
rect 15372 16156 15428 16158
rect 14140 15426 14196 15428
rect 14140 15374 14142 15426
rect 14142 15374 14194 15426
rect 14194 15374 14196 15426
rect 14140 15372 14196 15374
rect 14812 15484 14868 15540
rect 14364 15036 14420 15092
rect 14064 14922 14120 14924
rect 14064 14870 14066 14922
rect 14066 14870 14118 14922
rect 14118 14870 14120 14922
rect 14064 14868 14120 14870
rect 14168 14922 14224 14924
rect 14168 14870 14170 14922
rect 14170 14870 14222 14922
rect 14222 14870 14224 14922
rect 14168 14868 14224 14870
rect 14272 14922 14328 14924
rect 14272 14870 14274 14922
rect 14274 14870 14326 14922
rect 14326 14870 14328 14922
rect 14272 14868 14328 14870
rect 14812 14924 14868 14980
rect 13804 13634 13860 13636
rect 13804 13582 13806 13634
rect 13806 13582 13858 13634
rect 13858 13582 13860 13634
rect 13804 13580 13860 13582
rect 13580 12402 13636 12404
rect 13580 12350 13582 12402
rect 13582 12350 13634 12402
rect 13634 12350 13636 12402
rect 13580 12348 13636 12350
rect 14700 13580 14756 13636
rect 14064 13354 14120 13356
rect 14064 13302 14066 13354
rect 14066 13302 14118 13354
rect 14118 13302 14120 13354
rect 14064 13300 14120 13302
rect 14168 13354 14224 13356
rect 14168 13302 14170 13354
rect 14170 13302 14222 13354
rect 14222 13302 14224 13354
rect 14168 13300 14224 13302
rect 14272 13354 14328 13356
rect 14272 13302 14274 13354
rect 14274 13302 14326 13354
rect 14326 13302 14328 13354
rect 14272 13300 14328 13302
rect 16268 18396 16324 18452
rect 16380 18956 16436 19012
rect 16156 17778 16212 17780
rect 16156 17726 16158 17778
rect 16158 17726 16210 17778
rect 16210 17726 16212 17778
rect 16156 17724 16212 17726
rect 17388 20130 17444 20132
rect 17388 20078 17390 20130
rect 17390 20078 17442 20130
rect 17442 20078 17444 20130
rect 17388 20076 17444 20078
rect 17612 18450 17668 18452
rect 17612 18398 17614 18450
rect 17614 18398 17666 18450
rect 17666 18398 17668 18450
rect 17612 18396 17668 18398
rect 18620 20690 18676 20692
rect 18620 20638 18622 20690
rect 18622 20638 18674 20690
rect 18674 20638 18676 20690
rect 18620 20636 18676 20638
rect 18284 20578 18340 20580
rect 18284 20526 18286 20578
rect 18286 20526 18338 20578
rect 18338 20526 18340 20578
rect 18284 20524 18340 20526
rect 19404 22930 19460 22932
rect 19404 22878 19406 22930
rect 19406 22878 19458 22930
rect 19458 22878 19460 22930
rect 19404 22876 19460 22878
rect 19404 22594 19460 22596
rect 19404 22542 19406 22594
rect 19406 22542 19458 22594
rect 19458 22542 19460 22594
rect 19404 22540 19460 22542
rect 19180 21644 19236 21700
rect 18348 20410 18404 20412
rect 18348 20358 18350 20410
rect 18350 20358 18402 20410
rect 18402 20358 18404 20410
rect 18348 20356 18404 20358
rect 18452 20410 18508 20412
rect 18452 20358 18454 20410
rect 18454 20358 18506 20410
rect 18506 20358 18508 20410
rect 18452 20356 18508 20358
rect 18556 20410 18612 20412
rect 18556 20358 18558 20410
rect 18558 20358 18610 20410
rect 18610 20358 18612 20410
rect 18844 20412 18900 20468
rect 18556 20356 18612 20358
rect 18284 20130 18340 20132
rect 18284 20078 18286 20130
rect 18286 20078 18338 20130
rect 18338 20078 18340 20130
rect 18284 20076 18340 20078
rect 18732 18956 18788 19012
rect 18348 18842 18404 18844
rect 18348 18790 18350 18842
rect 18350 18790 18402 18842
rect 18402 18790 18404 18842
rect 18348 18788 18404 18790
rect 18452 18842 18508 18844
rect 18452 18790 18454 18842
rect 18454 18790 18506 18842
rect 18506 18790 18508 18842
rect 18452 18788 18508 18790
rect 18556 18842 18612 18844
rect 18556 18790 18558 18842
rect 18558 18790 18610 18842
rect 18610 18790 18612 18842
rect 18556 18788 18612 18790
rect 17836 18284 17892 18340
rect 17724 17836 17780 17892
rect 18060 18060 18116 18116
rect 17052 17778 17108 17780
rect 17052 17726 17054 17778
rect 17054 17726 17106 17778
rect 17106 17726 17108 17778
rect 17052 17724 17108 17726
rect 16828 17106 16884 17108
rect 16828 17054 16830 17106
rect 16830 17054 16882 17106
rect 16882 17054 16884 17106
rect 16828 17052 16884 17054
rect 15036 13580 15092 13636
rect 15596 13692 15652 13748
rect 15372 13580 15428 13636
rect 18284 17666 18340 17668
rect 18284 17614 18286 17666
rect 18286 17614 18338 17666
rect 18338 17614 18340 17666
rect 18284 17612 18340 17614
rect 17836 17554 17892 17556
rect 17836 17502 17838 17554
rect 17838 17502 17890 17554
rect 17890 17502 17892 17554
rect 17836 17500 17892 17502
rect 18620 17554 18676 17556
rect 18620 17502 18622 17554
rect 18622 17502 18674 17554
rect 18674 17502 18676 17554
rect 18620 17500 18676 17502
rect 17724 17388 17780 17444
rect 16716 15260 16772 15316
rect 18348 17274 18404 17276
rect 18348 17222 18350 17274
rect 18350 17222 18402 17274
rect 18402 17222 18404 17274
rect 18348 17220 18404 17222
rect 18452 17274 18508 17276
rect 18452 17222 18454 17274
rect 18454 17222 18506 17274
rect 18506 17222 18508 17274
rect 18452 17220 18508 17222
rect 18556 17274 18612 17276
rect 18556 17222 18558 17274
rect 18558 17222 18610 17274
rect 18610 17222 18612 17274
rect 18556 17220 18612 17222
rect 17836 17052 17892 17108
rect 17052 15148 17108 15204
rect 16828 14700 16884 14756
rect 16940 15036 16996 15092
rect 16940 14642 16996 14644
rect 16940 14590 16942 14642
rect 16942 14590 16994 14642
rect 16994 14590 16996 14642
rect 16940 14588 16996 14590
rect 16604 13916 16660 13972
rect 16156 13634 16212 13636
rect 16156 13582 16158 13634
rect 16158 13582 16210 13634
rect 16210 13582 16212 13634
rect 16156 13580 16212 13582
rect 15148 12348 15204 12404
rect 13916 12178 13972 12180
rect 13916 12126 13918 12178
rect 13918 12126 13970 12178
rect 13970 12126 13972 12178
rect 13916 12124 13972 12126
rect 14064 11786 14120 11788
rect 14064 11734 14066 11786
rect 14066 11734 14118 11786
rect 14118 11734 14120 11786
rect 14064 11732 14120 11734
rect 14168 11786 14224 11788
rect 14168 11734 14170 11786
rect 14170 11734 14222 11786
rect 14222 11734 14224 11786
rect 14168 11732 14224 11734
rect 14272 11786 14328 11788
rect 14272 11734 14274 11786
rect 14274 11734 14326 11786
rect 14326 11734 14328 11786
rect 14272 11732 14328 11734
rect 15148 11788 15204 11844
rect 14588 10444 14644 10500
rect 14064 10218 14120 10220
rect 14064 10166 14066 10218
rect 14066 10166 14118 10218
rect 14118 10166 14120 10218
rect 14064 10164 14120 10166
rect 14168 10218 14224 10220
rect 14168 10166 14170 10218
rect 14170 10166 14222 10218
rect 14222 10166 14224 10218
rect 14168 10164 14224 10166
rect 14272 10218 14328 10220
rect 14272 10166 14274 10218
rect 14274 10166 14326 10218
rect 14326 10166 14328 10218
rect 14272 10164 14328 10166
rect 14476 9996 14532 10052
rect 14140 9938 14196 9940
rect 14140 9886 14142 9938
rect 14142 9886 14194 9938
rect 14194 9886 14196 9938
rect 14140 9884 14196 9886
rect 13580 9602 13636 9604
rect 13580 9550 13582 9602
rect 13582 9550 13634 9602
rect 13634 9550 13636 9602
rect 13580 9548 13636 9550
rect 13580 8876 13636 8932
rect 14064 8650 14120 8652
rect 14064 8598 14066 8650
rect 14066 8598 14118 8650
rect 14118 8598 14120 8650
rect 14064 8596 14120 8598
rect 14168 8650 14224 8652
rect 14168 8598 14170 8650
rect 14170 8598 14222 8650
rect 14222 8598 14224 8650
rect 14168 8596 14224 8598
rect 14272 8650 14328 8652
rect 14272 8598 14274 8650
rect 14274 8598 14326 8650
rect 14326 8598 14328 8650
rect 14272 8596 14328 8598
rect 13916 8428 13972 8484
rect 14140 8428 14196 8484
rect 13580 7420 13636 7476
rect 13468 5964 13524 6020
rect 13468 5292 13524 5348
rect 13580 5740 13636 5796
rect 13468 5122 13524 5124
rect 13468 5070 13470 5122
rect 13470 5070 13522 5122
rect 13522 5070 13524 5122
rect 13468 5068 13524 5070
rect 13916 7420 13972 7476
rect 14700 9548 14756 9604
rect 16492 13580 16548 13636
rect 16716 13692 16772 13748
rect 16492 12348 16548 12404
rect 16156 11788 16212 11844
rect 15932 11452 15988 11508
rect 15260 11116 15316 11172
rect 16156 11170 16212 11172
rect 16156 11118 16158 11170
rect 16158 11118 16210 11170
rect 16210 11118 16212 11170
rect 16156 11116 16212 11118
rect 15596 10610 15652 10612
rect 15596 10558 15598 10610
rect 15598 10558 15650 10610
rect 15650 10558 15652 10610
rect 15596 10556 15652 10558
rect 15708 10498 15764 10500
rect 15708 10446 15710 10498
rect 15710 10446 15762 10498
rect 15762 10446 15764 10498
rect 15708 10444 15764 10446
rect 15036 9996 15092 10052
rect 14924 9826 14980 9828
rect 14924 9774 14926 9826
rect 14926 9774 14978 9826
rect 14978 9774 14980 9826
rect 14924 9772 14980 9774
rect 16492 10332 16548 10388
rect 16156 9772 16212 9828
rect 14812 9436 14868 9492
rect 15372 9602 15428 9604
rect 15372 9550 15374 9602
rect 15374 9550 15426 9602
rect 15426 9550 15428 9602
rect 15372 9548 15428 9550
rect 15484 9212 15540 9268
rect 15932 9602 15988 9604
rect 15932 9550 15934 9602
rect 15934 9550 15986 9602
rect 15986 9550 15988 9602
rect 15932 9548 15988 9550
rect 15036 8764 15092 8820
rect 14252 8034 14308 8036
rect 14252 7982 14254 8034
rect 14254 7982 14306 8034
rect 14306 7982 14308 8034
rect 14252 7980 14308 7982
rect 14064 7082 14120 7084
rect 14064 7030 14066 7082
rect 14066 7030 14118 7082
rect 14118 7030 14120 7082
rect 14064 7028 14120 7030
rect 14168 7082 14224 7084
rect 14168 7030 14170 7082
rect 14170 7030 14222 7082
rect 14222 7030 14224 7082
rect 14168 7028 14224 7030
rect 14272 7082 14328 7084
rect 14272 7030 14274 7082
rect 14274 7030 14326 7082
rect 14326 7030 14328 7082
rect 14272 7028 14328 7030
rect 14476 6076 14532 6132
rect 15260 8204 15316 8260
rect 15820 9100 15876 9156
rect 15260 7644 15316 7700
rect 15708 8930 15764 8932
rect 15708 8878 15710 8930
rect 15710 8878 15762 8930
rect 15762 8878 15764 8930
rect 15708 8876 15764 8878
rect 15708 8092 15764 8148
rect 16828 11452 16884 11508
rect 16716 10332 16772 10388
rect 16940 9996 16996 10052
rect 16604 9266 16660 9268
rect 16604 9214 16606 9266
rect 16606 9214 16658 9266
rect 16658 9214 16660 9266
rect 16604 9212 16660 9214
rect 18844 18060 18900 18116
rect 18844 17106 18900 17108
rect 18844 17054 18846 17106
rect 18846 17054 18898 17106
rect 18898 17054 18900 17106
rect 18844 17052 18900 17054
rect 18172 16380 18228 16436
rect 18060 16268 18116 16324
rect 18732 16156 18788 16212
rect 19740 23714 19796 23716
rect 19740 23662 19742 23714
rect 19742 23662 19794 23714
rect 19794 23662 19796 23714
rect 19740 23660 19796 23662
rect 19964 23154 20020 23156
rect 19964 23102 19966 23154
rect 19966 23102 20018 23154
rect 20018 23102 20020 23154
rect 19964 23100 20020 23102
rect 19404 21420 19460 21476
rect 19404 20412 19460 20468
rect 19740 22764 19796 22820
rect 19964 22092 20020 22148
rect 19964 20524 20020 20580
rect 19068 20076 19124 20132
rect 19404 19404 19460 19460
rect 19404 18060 19460 18116
rect 19068 17500 19124 17556
rect 19292 17612 19348 17668
rect 20412 24668 20468 24724
rect 19628 17666 19684 17668
rect 19628 17614 19630 17666
rect 19630 17614 19682 17666
rect 19682 17614 19684 17666
rect 19628 17612 19684 17614
rect 19516 17442 19572 17444
rect 19516 17390 19518 17442
rect 19518 17390 19570 17442
rect 19570 17390 19572 17442
rect 19516 17388 19572 17390
rect 20076 17612 20132 17668
rect 19292 17052 19348 17108
rect 19852 17052 19908 17108
rect 19404 16940 19460 16996
rect 19628 16380 19684 16436
rect 18348 15706 18404 15708
rect 18348 15654 18350 15706
rect 18350 15654 18402 15706
rect 18402 15654 18404 15706
rect 18348 15652 18404 15654
rect 18452 15706 18508 15708
rect 18452 15654 18454 15706
rect 18454 15654 18506 15706
rect 18506 15654 18508 15706
rect 18452 15652 18508 15654
rect 18556 15706 18612 15708
rect 18556 15654 18558 15706
rect 18558 15654 18610 15706
rect 18610 15654 18612 15706
rect 18556 15652 18612 15654
rect 17948 14364 18004 14420
rect 17388 13970 17444 13972
rect 17388 13918 17390 13970
rect 17390 13918 17442 13970
rect 17442 13918 17444 13970
rect 17388 13916 17444 13918
rect 17164 12348 17220 12404
rect 17948 12178 18004 12180
rect 17948 12126 17950 12178
rect 17950 12126 18002 12178
rect 18002 12126 18004 12178
rect 17948 12124 18004 12126
rect 19068 14642 19124 14644
rect 19068 14590 19070 14642
rect 19070 14590 19122 14642
rect 19122 14590 19124 14642
rect 19068 14588 19124 14590
rect 18348 14138 18404 14140
rect 18348 14086 18350 14138
rect 18350 14086 18402 14138
rect 18402 14086 18404 14138
rect 18348 14084 18404 14086
rect 18452 14138 18508 14140
rect 18452 14086 18454 14138
rect 18454 14086 18506 14138
rect 18506 14086 18508 14138
rect 18452 14084 18508 14086
rect 18556 14138 18612 14140
rect 18556 14086 18558 14138
rect 18558 14086 18610 14138
rect 18610 14086 18612 14138
rect 18556 14084 18612 14086
rect 18620 13634 18676 13636
rect 18620 13582 18622 13634
rect 18622 13582 18674 13634
rect 18674 13582 18676 13634
rect 18620 13580 18676 13582
rect 18956 12684 19012 12740
rect 18348 12570 18404 12572
rect 18348 12518 18350 12570
rect 18350 12518 18402 12570
rect 18402 12518 18404 12570
rect 18348 12516 18404 12518
rect 18452 12570 18508 12572
rect 18452 12518 18454 12570
rect 18454 12518 18506 12570
rect 18506 12518 18508 12570
rect 18452 12516 18508 12518
rect 18556 12570 18612 12572
rect 18556 12518 18558 12570
rect 18558 12518 18610 12570
rect 18610 12518 18612 12570
rect 18556 12516 18612 12518
rect 18348 11002 18404 11004
rect 18348 10950 18350 11002
rect 18350 10950 18402 11002
rect 18402 10950 18404 11002
rect 18348 10948 18404 10950
rect 18452 11002 18508 11004
rect 18452 10950 18454 11002
rect 18454 10950 18506 11002
rect 18506 10950 18508 11002
rect 18452 10948 18508 10950
rect 18556 11002 18612 11004
rect 18556 10950 18558 11002
rect 18558 10950 18610 11002
rect 18610 10950 18612 11002
rect 18556 10948 18612 10950
rect 16380 8764 16436 8820
rect 17052 8876 17108 8932
rect 16716 8258 16772 8260
rect 16716 8206 16718 8258
rect 16718 8206 16770 8258
rect 16770 8206 16772 8258
rect 16716 8204 16772 8206
rect 16268 8092 16324 8148
rect 15820 7698 15876 7700
rect 15820 7646 15822 7698
rect 15822 7646 15874 7698
rect 15874 7646 15876 7698
rect 15820 7644 15876 7646
rect 16268 7474 16324 7476
rect 16268 7422 16270 7474
rect 16270 7422 16322 7474
rect 16322 7422 16324 7474
rect 16268 7420 16324 7422
rect 17388 9154 17444 9156
rect 17388 9102 17390 9154
rect 17390 9102 17442 9154
rect 17442 9102 17444 9154
rect 17388 9100 17444 9102
rect 17612 8764 17668 8820
rect 17500 8428 17556 8484
rect 17836 9100 17892 9156
rect 18348 9434 18404 9436
rect 18348 9382 18350 9434
rect 18350 9382 18402 9434
rect 18402 9382 18404 9434
rect 18348 9380 18404 9382
rect 18452 9434 18508 9436
rect 18452 9382 18454 9434
rect 18454 9382 18506 9434
rect 18506 9382 18508 9434
rect 18452 9380 18508 9382
rect 18556 9434 18612 9436
rect 18556 9382 18558 9434
rect 18558 9382 18610 9434
rect 18610 9382 18612 9434
rect 18556 9380 18612 9382
rect 18284 9154 18340 9156
rect 18284 9102 18286 9154
rect 18286 9102 18338 9154
rect 18338 9102 18340 9154
rect 18284 9100 18340 9102
rect 17724 8428 17780 8484
rect 17388 7756 17444 7812
rect 16492 6524 16548 6580
rect 14252 5964 14308 6020
rect 14812 6466 14868 6468
rect 14812 6414 14814 6466
rect 14814 6414 14866 6466
rect 14866 6414 14868 6466
rect 14812 6412 14868 6414
rect 15820 6412 15876 6468
rect 14064 5514 14120 5516
rect 14064 5462 14066 5514
rect 14066 5462 14118 5514
rect 14118 5462 14120 5514
rect 14064 5460 14120 5462
rect 14168 5514 14224 5516
rect 14168 5462 14170 5514
rect 14170 5462 14222 5514
rect 14222 5462 14224 5514
rect 14168 5460 14224 5462
rect 14272 5514 14328 5516
rect 14272 5462 14274 5514
rect 14274 5462 14326 5514
rect 14326 5462 14328 5514
rect 14272 5460 14328 5462
rect 14028 5292 14084 5348
rect 13580 3554 13636 3556
rect 13580 3502 13582 3554
rect 13582 3502 13634 3554
rect 13634 3502 13636 3554
rect 13580 3500 13636 3502
rect 14064 3946 14120 3948
rect 14064 3894 14066 3946
rect 14066 3894 14118 3946
rect 14118 3894 14120 3946
rect 14064 3892 14120 3894
rect 14168 3946 14224 3948
rect 14168 3894 14170 3946
rect 14170 3894 14222 3946
rect 14222 3894 14224 3946
rect 14168 3892 14224 3894
rect 14272 3946 14328 3948
rect 14272 3894 14274 3946
rect 14274 3894 14326 3946
rect 14326 3894 14328 3946
rect 14272 3892 14328 3894
rect 13916 3500 13972 3556
rect 15372 5628 15428 5684
rect 14588 5234 14644 5236
rect 14588 5182 14590 5234
rect 14590 5182 14642 5234
rect 14642 5182 14644 5234
rect 14588 5180 14644 5182
rect 15484 5180 15540 5236
rect 14588 4844 14644 4900
rect 13356 3442 13412 3444
rect 13356 3390 13358 3442
rect 13358 3390 13410 3442
rect 13410 3390 13412 3442
rect 13356 3388 13412 3390
rect 17164 6412 17220 6468
rect 16156 5964 16212 6020
rect 15708 4396 15764 4452
rect 16492 5740 16548 5796
rect 17052 5180 17108 5236
rect 16716 4508 16772 4564
rect 16828 4956 16884 5012
rect 16828 4338 16884 4340
rect 16828 4286 16830 4338
rect 16830 4286 16882 4338
rect 16882 4286 16884 4338
rect 16828 4284 16884 4286
rect 17052 4172 17108 4228
rect 17052 3948 17108 4004
rect 17388 5906 17444 5908
rect 17388 5854 17390 5906
rect 17390 5854 17442 5906
rect 17442 5854 17444 5906
rect 17388 5852 17444 5854
rect 17836 5628 17892 5684
rect 17388 5068 17444 5124
rect 17276 3724 17332 3780
rect 17500 4956 17556 5012
rect 17500 4562 17556 4564
rect 17500 4510 17502 4562
rect 17502 4510 17554 4562
rect 17554 4510 17556 4562
rect 17500 4508 17556 4510
rect 17948 8316 18004 8372
rect 18620 9042 18676 9044
rect 18620 8990 18622 9042
rect 18622 8990 18674 9042
rect 18674 8990 18676 9042
rect 18620 8988 18676 8990
rect 18348 7866 18404 7868
rect 18348 7814 18350 7866
rect 18350 7814 18402 7866
rect 18402 7814 18404 7866
rect 18348 7812 18404 7814
rect 18452 7866 18508 7868
rect 18452 7814 18454 7866
rect 18454 7814 18506 7866
rect 18506 7814 18508 7866
rect 18452 7812 18508 7814
rect 18556 7866 18612 7868
rect 18556 7814 18558 7866
rect 18558 7814 18610 7866
rect 18610 7814 18612 7866
rect 18556 7812 18612 7814
rect 18396 7698 18452 7700
rect 18396 7646 18398 7698
rect 18398 7646 18450 7698
rect 18450 7646 18452 7698
rect 18396 7644 18452 7646
rect 18508 7586 18564 7588
rect 18508 7534 18510 7586
rect 18510 7534 18562 7586
rect 18562 7534 18564 7586
rect 18508 7532 18564 7534
rect 18172 7474 18228 7476
rect 18172 7422 18174 7474
rect 18174 7422 18226 7474
rect 18226 7422 18228 7474
rect 18172 7420 18228 7422
rect 18060 7308 18116 7364
rect 19404 14252 19460 14308
rect 19516 14028 19572 14084
rect 20300 16604 20356 16660
rect 20860 26514 20916 26516
rect 20860 26462 20862 26514
rect 20862 26462 20914 26514
rect 20914 26462 20916 26514
rect 20860 26460 20916 26462
rect 20972 25228 21028 25284
rect 20636 23772 20692 23828
rect 20860 23660 20916 23716
rect 20636 23042 20692 23044
rect 20636 22990 20638 23042
rect 20638 22990 20690 23042
rect 20690 22990 20692 23042
rect 20636 22988 20692 22990
rect 20748 22258 20804 22260
rect 20748 22206 20750 22258
rect 20750 22206 20802 22258
rect 20802 22206 20804 22258
rect 20748 22204 20804 22206
rect 20748 21420 20804 21476
rect 20748 20300 20804 20356
rect 20636 19906 20692 19908
rect 20636 19854 20638 19906
rect 20638 19854 20690 19906
rect 20690 19854 20692 19906
rect 20636 19852 20692 19854
rect 20524 19234 20580 19236
rect 20524 19182 20526 19234
rect 20526 19182 20578 19234
rect 20578 19182 20580 19234
rect 20524 19180 20580 19182
rect 20412 16492 20468 16548
rect 19740 15820 19796 15876
rect 19852 14364 19908 14420
rect 20076 14140 20132 14196
rect 19964 13858 20020 13860
rect 19964 13806 19966 13858
rect 19966 13806 20018 13858
rect 20018 13806 20020 13858
rect 19964 13804 20020 13806
rect 20412 14252 20468 14308
rect 20860 18284 20916 18340
rect 20748 18060 20804 18116
rect 21308 28530 21364 28532
rect 21308 28478 21310 28530
rect 21310 28478 21362 28530
rect 21362 28478 21364 28530
rect 21308 28476 21364 28478
rect 21532 30098 21588 30100
rect 21532 30046 21534 30098
rect 21534 30046 21586 30098
rect 21586 30046 21588 30098
rect 21532 30044 21588 30046
rect 21420 28364 21476 28420
rect 22092 31388 22148 31444
rect 21868 30268 21924 30324
rect 21756 30156 21812 30212
rect 22092 30044 22148 30100
rect 21980 29932 22036 29988
rect 21980 29148 22036 29204
rect 22204 29484 22260 29540
rect 22540 31948 22596 32004
rect 22988 31554 23044 31556
rect 22988 31502 22990 31554
rect 22990 31502 23042 31554
rect 23042 31502 23044 31554
rect 22988 31500 23044 31502
rect 23324 32508 23380 32564
rect 23436 32284 23492 32340
rect 23884 32508 23940 32564
rect 23772 31948 23828 32004
rect 23548 31612 23604 31668
rect 22652 31276 22708 31332
rect 23212 31276 23268 31332
rect 22764 30994 22820 30996
rect 22764 30942 22766 30994
rect 22766 30942 22818 30994
rect 22818 30942 22820 30994
rect 22764 30940 22820 30942
rect 22632 30602 22688 30604
rect 22632 30550 22634 30602
rect 22634 30550 22686 30602
rect 22686 30550 22688 30602
rect 22632 30548 22688 30550
rect 22736 30602 22792 30604
rect 22736 30550 22738 30602
rect 22738 30550 22790 30602
rect 22790 30550 22792 30602
rect 22736 30548 22792 30550
rect 22840 30602 22896 30604
rect 22840 30550 22842 30602
rect 22842 30550 22894 30602
rect 22894 30550 22896 30602
rect 22840 30548 22896 30550
rect 22764 29426 22820 29428
rect 22764 29374 22766 29426
rect 22766 29374 22818 29426
rect 22818 29374 22820 29426
rect 22764 29372 22820 29374
rect 22876 29148 22932 29204
rect 22632 29034 22688 29036
rect 22632 28982 22634 29034
rect 22634 28982 22686 29034
rect 22686 28982 22688 29034
rect 22632 28980 22688 28982
rect 22736 29034 22792 29036
rect 22736 28982 22738 29034
rect 22738 28982 22790 29034
rect 22790 28982 22792 29034
rect 22736 28980 22792 28982
rect 22840 29034 22896 29036
rect 22840 28982 22842 29034
rect 22842 28982 22894 29034
rect 22894 28982 22896 29034
rect 22840 28980 22896 28982
rect 22316 28252 22372 28308
rect 22204 28140 22260 28196
rect 21756 28028 21812 28084
rect 21308 27746 21364 27748
rect 21308 27694 21310 27746
rect 21310 27694 21362 27746
rect 21362 27694 21364 27746
rect 21308 27692 21364 27694
rect 21756 27244 21812 27300
rect 21868 27804 21924 27860
rect 23436 30994 23492 30996
rect 23436 30942 23438 30994
rect 23438 30942 23490 30994
rect 23490 30942 23492 30994
rect 23436 30940 23492 30942
rect 23548 30882 23604 30884
rect 23548 30830 23550 30882
rect 23550 30830 23602 30882
rect 23602 30830 23604 30882
rect 23548 30828 23604 30830
rect 23212 29986 23268 29988
rect 23212 29934 23214 29986
rect 23214 29934 23266 29986
rect 23266 29934 23268 29986
rect 23212 29932 23268 29934
rect 23324 29820 23380 29876
rect 23212 29148 23268 29204
rect 23212 27916 23268 27972
rect 22428 27804 22484 27860
rect 21420 26850 21476 26852
rect 21420 26798 21422 26850
rect 21422 26798 21474 26850
rect 21474 26798 21476 26850
rect 21420 26796 21476 26798
rect 21308 25788 21364 25844
rect 21420 26012 21476 26068
rect 21756 26572 21812 26628
rect 22632 27466 22688 27468
rect 22632 27414 22634 27466
rect 22634 27414 22686 27466
rect 22686 27414 22688 27466
rect 22632 27412 22688 27414
rect 22736 27466 22792 27468
rect 22736 27414 22738 27466
rect 22738 27414 22790 27466
rect 22790 27414 22792 27466
rect 22736 27412 22792 27414
rect 22840 27466 22896 27468
rect 22840 27414 22842 27466
rect 22842 27414 22894 27466
rect 22894 27414 22896 27466
rect 22840 27412 22896 27414
rect 22428 27074 22484 27076
rect 22428 27022 22430 27074
rect 22430 27022 22482 27074
rect 22482 27022 22484 27074
rect 22428 27020 22484 27022
rect 22652 27244 22708 27300
rect 23884 30156 23940 30212
rect 24220 30828 24276 30884
rect 23660 29596 23716 29652
rect 24108 29650 24164 29652
rect 24108 29598 24110 29650
rect 24110 29598 24162 29650
rect 24162 29598 24164 29650
rect 24108 29596 24164 29598
rect 23772 29314 23828 29316
rect 23772 29262 23774 29314
rect 23774 29262 23826 29314
rect 23826 29262 23828 29314
rect 23772 29260 23828 29262
rect 23772 28642 23828 28644
rect 23772 28590 23774 28642
rect 23774 28590 23826 28642
rect 23826 28590 23828 28642
rect 23772 28588 23828 28590
rect 23100 27244 23156 27300
rect 22092 26460 22148 26516
rect 22540 26962 22596 26964
rect 22540 26910 22542 26962
rect 22542 26910 22594 26962
rect 22594 26910 22596 26962
rect 22540 26908 22596 26910
rect 23436 27244 23492 27300
rect 25564 33570 25620 33572
rect 25564 33518 25566 33570
rect 25566 33518 25618 33570
rect 25618 33518 25620 33570
rect 25564 33516 25620 33518
rect 25228 33404 25284 33460
rect 27356 33292 27412 33348
rect 26916 32954 26972 32956
rect 26916 32902 26918 32954
rect 26918 32902 26970 32954
rect 26970 32902 26972 32954
rect 26916 32900 26972 32902
rect 27020 32954 27076 32956
rect 27020 32902 27022 32954
rect 27022 32902 27074 32954
rect 27074 32902 27076 32954
rect 27020 32900 27076 32902
rect 27124 32954 27180 32956
rect 27124 32902 27126 32954
rect 27126 32902 27178 32954
rect 27178 32902 27180 32954
rect 27124 32900 27180 32902
rect 26236 32450 26292 32452
rect 26236 32398 26238 32450
rect 26238 32398 26290 32450
rect 26290 32398 26292 32450
rect 26236 32396 26292 32398
rect 24780 31836 24836 31892
rect 24668 30604 24724 30660
rect 25340 31500 25396 31556
rect 26460 31500 26516 31556
rect 26684 32172 26740 32228
rect 26348 31388 26404 31444
rect 25452 31106 25508 31108
rect 25452 31054 25454 31106
rect 25454 31054 25506 31106
rect 25506 31054 25508 31106
rect 25452 31052 25508 31054
rect 25900 30882 25956 30884
rect 25900 30830 25902 30882
rect 25902 30830 25954 30882
rect 25954 30830 25956 30882
rect 25900 30828 25956 30830
rect 25340 30770 25396 30772
rect 25340 30718 25342 30770
rect 25342 30718 25394 30770
rect 25394 30718 25396 30770
rect 25340 30716 25396 30718
rect 25340 30268 25396 30324
rect 24892 30098 24948 30100
rect 24892 30046 24894 30098
rect 24894 30046 24946 30098
rect 24946 30046 24948 30098
rect 24892 30044 24948 30046
rect 24556 28252 24612 28308
rect 24668 29596 24724 29652
rect 22652 26796 22708 26852
rect 22540 26684 22596 26740
rect 21868 26236 21924 26292
rect 21756 26178 21812 26180
rect 21756 26126 21758 26178
rect 21758 26126 21810 26178
rect 21810 26126 21812 26178
rect 21756 26124 21812 26126
rect 21868 25788 21924 25844
rect 22428 26348 22484 26404
rect 21756 25676 21812 25732
rect 21756 25116 21812 25172
rect 21532 23938 21588 23940
rect 21532 23886 21534 23938
rect 21534 23886 21586 23938
rect 21586 23886 21588 23938
rect 21532 23884 21588 23886
rect 21084 23660 21140 23716
rect 22204 26066 22260 26068
rect 22204 26014 22206 26066
rect 22206 26014 22258 26066
rect 22258 26014 22260 26066
rect 22204 26012 22260 26014
rect 23212 26348 23268 26404
rect 22764 26290 22820 26292
rect 22764 26238 22766 26290
rect 22766 26238 22818 26290
rect 22818 26238 22820 26290
rect 22764 26236 22820 26238
rect 23660 26796 23716 26852
rect 22632 25898 22688 25900
rect 22632 25846 22634 25898
rect 22634 25846 22686 25898
rect 22686 25846 22688 25898
rect 22632 25844 22688 25846
rect 22736 25898 22792 25900
rect 22736 25846 22738 25898
rect 22738 25846 22790 25898
rect 22790 25846 22792 25898
rect 22736 25844 22792 25846
rect 22840 25898 22896 25900
rect 22840 25846 22842 25898
rect 22842 25846 22894 25898
rect 22894 25846 22896 25898
rect 22840 25844 22896 25846
rect 22092 25394 22148 25396
rect 22092 25342 22094 25394
rect 22094 25342 22146 25394
rect 22146 25342 22148 25394
rect 22092 25340 22148 25342
rect 22988 25340 23044 25396
rect 23100 25282 23156 25284
rect 23100 25230 23102 25282
rect 23102 25230 23154 25282
rect 23154 25230 23156 25282
rect 23100 25228 23156 25230
rect 23436 25228 23492 25284
rect 22316 23884 22372 23940
rect 23660 25116 23716 25172
rect 24444 26962 24500 26964
rect 24444 26910 24446 26962
rect 24446 26910 24498 26962
rect 24498 26910 24500 26962
rect 24444 26908 24500 26910
rect 25228 29426 25284 29428
rect 25228 29374 25230 29426
rect 25230 29374 25282 29426
rect 25282 29374 25284 29426
rect 25228 29372 25284 29374
rect 25228 28252 25284 28308
rect 24668 26514 24724 26516
rect 24668 26462 24670 26514
rect 24670 26462 24722 26514
rect 24722 26462 24724 26514
rect 24668 26460 24724 26462
rect 24892 27580 24948 27636
rect 23884 26402 23940 26404
rect 23884 26350 23886 26402
rect 23886 26350 23938 26402
rect 23938 26350 23940 26402
rect 23884 26348 23940 26350
rect 23884 25564 23940 25620
rect 24220 25394 24276 25396
rect 24220 25342 24222 25394
rect 24222 25342 24274 25394
rect 24274 25342 24276 25394
rect 24220 25340 24276 25342
rect 23772 24668 23828 24724
rect 24220 24892 24276 24948
rect 21308 23548 21364 23604
rect 21644 22988 21700 23044
rect 21532 22876 21588 22932
rect 21308 22258 21364 22260
rect 21308 22206 21310 22258
rect 21310 22206 21362 22258
rect 21362 22206 21364 22258
rect 21308 22204 21364 22206
rect 22632 24330 22688 24332
rect 22632 24278 22634 24330
rect 22634 24278 22686 24330
rect 22686 24278 22688 24330
rect 22632 24276 22688 24278
rect 22736 24330 22792 24332
rect 22736 24278 22738 24330
rect 22738 24278 22790 24330
rect 22790 24278 22792 24330
rect 22736 24276 22792 24278
rect 22840 24330 22896 24332
rect 22840 24278 22842 24330
rect 22842 24278 22894 24330
rect 22894 24278 22896 24330
rect 22840 24276 22896 24278
rect 22764 23884 22820 23940
rect 23996 24220 24052 24276
rect 23884 23996 23940 24052
rect 23212 23154 23268 23156
rect 23212 23102 23214 23154
rect 23214 23102 23266 23154
rect 23266 23102 23268 23154
rect 23212 23100 23268 23102
rect 23548 23436 23604 23492
rect 22632 22762 22688 22764
rect 22632 22710 22634 22762
rect 22634 22710 22686 22762
rect 22686 22710 22688 22762
rect 22632 22708 22688 22710
rect 22736 22762 22792 22764
rect 22736 22710 22738 22762
rect 22738 22710 22790 22762
rect 22790 22710 22792 22762
rect 22736 22708 22792 22710
rect 22840 22762 22896 22764
rect 22840 22710 22842 22762
rect 22842 22710 22894 22762
rect 22894 22710 22896 22762
rect 22840 22708 22896 22710
rect 24332 23996 24388 24052
rect 24332 23548 24388 23604
rect 24668 23324 24724 23380
rect 24444 23212 24500 23268
rect 23660 23042 23716 23044
rect 23660 22990 23662 23042
rect 23662 22990 23714 23042
rect 23714 22990 23716 23042
rect 23660 22988 23716 22990
rect 23548 22540 23604 22596
rect 22316 22204 22372 22260
rect 21084 21810 21140 21812
rect 21084 21758 21086 21810
rect 21086 21758 21138 21810
rect 21138 21758 21140 21810
rect 21084 21756 21140 21758
rect 21868 21474 21924 21476
rect 21868 21422 21870 21474
rect 21870 21422 21922 21474
rect 21922 21422 21924 21474
rect 21868 21420 21924 21422
rect 21420 20188 21476 20244
rect 22876 21420 22932 21476
rect 22540 21308 22596 21364
rect 22632 21194 22688 21196
rect 22632 21142 22634 21194
rect 22634 21142 22686 21194
rect 22686 21142 22688 21194
rect 22632 21140 22688 21142
rect 22736 21194 22792 21196
rect 22736 21142 22738 21194
rect 22738 21142 22790 21194
rect 22790 21142 22792 21194
rect 22736 21140 22792 21142
rect 22840 21194 22896 21196
rect 22840 21142 22842 21194
rect 22842 21142 22894 21194
rect 22894 21142 22896 21194
rect 22840 21140 22896 21142
rect 22764 20914 22820 20916
rect 22764 20862 22766 20914
rect 22766 20862 22818 20914
rect 22818 20862 22820 20914
rect 22764 20860 22820 20862
rect 20860 17164 20916 17220
rect 20636 16828 20692 16884
rect 21756 19180 21812 19236
rect 21644 18508 21700 18564
rect 21644 18338 21700 18340
rect 21644 18286 21646 18338
rect 21646 18286 21698 18338
rect 21698 18286 21700 18338
rect 21644 18284 21700 18286
rect 21420 18060 21476 18116
rect 22876 20524 22932 20580
rect 22092 19852 22148 19908
rect 22988 19906 23044 19908
rect 22988 19854 22990 19906
rect 22990 19854 23042 19906
rect 23042 19854 23044 19906
rect 22988 19852 23044 19854
rect 22632 19626 22688 19628
rect 22632 19574 22634 19626
rect 22634 19574 22686 19626
rect 22686 19574 22688 19626
rect 22632 19572 22688 19574
rect 22736 19626 22792 19628
rect 22736 19574 22738 19626
rect 22738 19574 22790 19626
rect 22790 19574 22792 19626
rect 22736 19572 22792 19574
rect 22840 19626 22896 19628
rect 22840 19574 22842 19626
rect 22842 19574 22894 19626
rect 22894 19574 22896 19626
rect 22840 19572 22896 19574
rect 22652 19010 22708 19012
rect 22652 18958 22654 19010
rect 22654 18958 22706 19010
rect 22706 18958 22708 19010
rect 22652 18956 22708 18958
rect 22428 18732 22484 18788
rect 23212 18956 23268 19012
rect 23660 21756 23716 21812
rect 23996 21196 24052 21252
rect 23996 20860 24052 20916
rect 23548 20242 23604 20244
rect 23548 20190 23550 20242
rect 23550 20190 23602 20242
rect 23602 20190 23604 20242
rect 23548 20188 23604 20190
rect 23660 19852 23716 19908
rect 23212 18396 23268 18452
rect 21196 16716 21252 16772
rect 20748 16098 20804 16100
rect 20748 16046 20750 16098
rect 20750 16046 20802 16098
rect 20802 16046 20804 16098
rect 20748 16044 20804 16046
rect 20748 14754 20804 14756
rect 20748 14702 20750 14754
rect 20750 14702 20802 14754
rect 20802 14702 20804 14754
rect 20748 14700 20804 14702
rect 22632 18058 22688 18060
rect 22632 18006 22634 18058
rect 22634 18006 22686 18058
rect 22686 18006 22688 18058
rect 22632 18004 22688 18006
rect 22736 18058 22792 18060
rect 22736 18006 22738 18058
rect 22738 18006 22790 18058
rect 22790 18006 22792 18058
rect 22736 18004 22792 18006
rect 22840 18058 22896 18060
rect 22840 18006 22842 18058
rect 22842 18006 22894 18058
rect 22894 18006 22896 18058
rect 22840 18004 22896 18006
rect 22988 17948 23044 18004
rect 21420 16492 21476 16548
rect 21980 17612 22036 17668
rect 21980 16994 22036 16996
rect 21980 16942 21982 16994
rect 21982 16942 22034 16994
rect 22034 16942 22036 16994
rect 21980 16940 22036 16942
rect 22988 17666 23044 17668
rect 22988 17614 22990 17666
rect 22990 17614 23042 17666
rect 23042 17614 23044 17666
rect 22988 17612 23044 17614
rect 22428 17554 22484 17556
rect 22428 17502 22430 17554
rect 22430 17502 22482 17554
rect 22482 17502 22484 17554
rect 22428 17500 22484 17502
rect 22652 17554 22708 17556
rect 22652 17502 22654 17554
rect 22654 17502 22706 17554
rect 22706 17502 22708 17554
rect 22652 17500 22708 17502
rect 22316 16940 22372 16996
rect 22204 16882 22260 16884
rect 22204 16830 22206 16882
rect 22206 16830 22258 16882
rect 22258 16830 22260 16882
rect 22204 16828 22260 16830
rect 21756 16098 21812 16100
rect 21756 16046 21758 16098
rect 21758 16046 21810 16098
rect 21810 16046 21812 16098
rect 21756 16044 21812 16046
rect 22092 16156 22148 16212
rect 21756 15314 21812 15316
rect 21756 15262 21758 15314
rect 21758 15262 21810 15314
rect 21810 15262 21812 15314
rect 21756 15260 21812 15262
rect 21420 14306 21476 14308
rect 21420 14254 21422 14306
rect 21422 14254 21474 14306
rect 21474 14254 21476 14306
rect 21420 14252 21476 14254
rect 20748 14028 20804 14084
rect 19516 12738 19572 12740
rect 19516 12686 19518 12738
rect 19518 12686 19570 12738
rect 19570 12686 19572 12738
rect 19516 12684 19572 12686
rect 19740 12684 19796 12740
rect 19516 11452 19572 11508
rect 20300 12738 20356 12740
rect 20300 12686 20302 12738
rect 20302 12686 20354 12738
rect 20354 12686 20356 12738
rect 20300 12684 20356 12686
rect 20524 12348 20580 12404
rect 21196 12402 21252 12404
rect 21196 12350 21198 12402
rect 21198 12350 21250 12402
rect 21250 12350 21252 12402
rect 21196 12348 21252 12350
rect 20300 11564 20356 11620
rect 19964 11452 20020 11508
rect 20636 11506 20692 11508
rect 20636 11454 20638 11506
rect 20638 11454 20690 11506
rect 20690 11454 20692 11506
rect 20636 11452 20692 11454
rect 19292 10780 19348 10836
rect 20188 11116 20244 11172
rect 20748 11170 20804 11172
rect 20748 11118 20750 11170
rect 20750 11118 20802 11170
rect 20802 11118 20804 11170
rect 20748 11116 20804 11118
rect 20748 10892 20804 10948
rect 20972 11564 21028 11620
rect 20636 10668 20692 10724
rect 20524 10610 20580 10612
rect 20524 10558 20526 10610
rect 20526 10558 20578 10610
rect 20578 10558 20580 10610
rect 20524 10556 20580 10558
rect 19740 9100 19796 9156
rect 21084 10722 21140 10724
rect 21084 10670 21086 10722
rect 21086 10670 21138 10722
rect 21138 10670 21140 10722
rect 21084 10668 21140 10670
rect 20300 9826 20356 9828
rect 20300 9774 20302 9826
rect 20302 9774 20354 9826
rect 20354 9774 20356 9826
rect 20300 9772 20356 9774
rect 19292 8370 19348 8372
rect 19292 8318 19294 8370
rect 19294 8318 19346 8370
rect 19346 8318 19348 8370
rect 19292 8316 19348 8318
rect 20188 8988 20244 9044
rect 19516 7586 19572 7588
rect 19516 7534 19518 7586
rect 19518 7534 19570 7586
rect 19570 7534 19572 7586
rect 19516 7532 19572 7534
rect 19852 7586 19908 7588
rect 19852 7534 19854 7586
rect 19854 7534 19906 7586
rect 19906 7534 19908 7586
rect 19852 7532 19908 7534
rect 21980 14028 22036 14084
rect 22316 14140 22372 14196
rect 21868 13634 21924 13636
rect 21868 13582 21870 13634
rect 21870 13582 21922 13634
rect 21922 13582 21924 13634
rect 21868 13580 21924 13582
rect 22540 16882 22596 16884
rect 22540 16830 22542 16882
rect 22542 16830 22594 16882
rect 22594 16830 22596 16882
rect 22540 16828 22596 16830
rect 22632 16490 22688 16492
rect 22632 16438 22634 16490
rect 22634 16438 22686 16490
rect 22686 16438 22688 16490
rect 22632 16436 22688 16438
rect 22736 16490 22792 16492
rect 22736 16438 22738 16490
rect 22738 16438 22790 16490
rect 22790 16438 22792 16490
rect 22736 16436 22792 16438
rect 22840 16490 22896 16492
rect 22840 16438 22842 16490
rect 22842 16438 22894 16490
rect 22894 16438 22896 16490
rect 22840 16436 22896 16438
rect 24668 22428 24724 22484
rect 24780 21698 24836 21700
rect 24780 21646 24782 21698
rect 24782 21646 24834 21698
rect 24834 21646 24836 21698
rect 24780 21644 24836 21646
rect 24220 21474 24276 21476
rect 24220 21422 24222 21474
rect 24222 21422 24274 21474
rect 24274 21422 24276 21474
rect 24220 21420 24276 21422
rect 24444 20636 24500 20692
rect 24108 19010 24164 19012
rect 24108 18958 24110 19010
rect 24110 18958 24162 19010
rect 24162 18958 24164 19010
rect 24108 18956 24164 18958
rect 25340 26290 25396 26292
rect 25340 26238 25342 26290
rect 25342 26238 25394 26290
rect 25394 26238 25396 26290
rect 25340 26236 25396 26238
rect 25228 24892 25284 24948
rect 26236 30604 26292 30660
rect 26236 28364 26292 28420
rect 25564 27916 25620 27972
rect 26236 27858 26292 27860
rect 26236 27806 26238 27858
rect 26238 27806 26290 27858
rect 26290 27806 26292 27858
rect 26236 27804 26292 27806
rect 25564 26684 25620 26740
rect 25900 27132 25956 27188
rect 25564 26514 25620 26516
rect 25564 26462 25566 26514
rect 25566 26462 25618 26514
rect 25618 26462 25620 26514
rect 25564 26460 25620 26462
rect 26572 28700 26628 28756
rect 26572 27186 26628 27188
rect 26572 27134 26574 27186
rect 26574 27134 26626 27186
rect 26626 27134 26628 27186
rect 26572 27132 26628 27134
rect 30156 33404 30212 33460
rect 28476 32844 28532 32900
rect 28588 32732 28644 32788
rect 27804 32508 27860 32564
rect 26908 31778 26964 31780
rect 26908 31726 26910 31778
rect 26910 31726 26962 31778
rect 26962 31726 26964 31778
rect 26908 31724 26964 31726
rect 26916 31386 26972 31388
rect 26916 31334 26918 31386
rect 26918 31334 26970 31386
rect 26970 31334 26972 31386
rect 26916 31332 26972 31334
rect 27020 31386 27076 31388
rect 27020 31334 27022 31386
rect 27022 31334 27074 31386
rect 27074 31334 27076 31386
rect 27020 31332 27076 31334
rect 27124 31386 27180 31388
rect 27124 31334 27126 31386
rect 27126 31334 27178 31386
rect 27178 31334 27180 31386
rect 27124 31332 27180 31334
rect 27468 31052 27524 31108
rect 27692 30828 27748 30884
rect 28028 32396 28084 32452
rect 28252 32284 28308 32340
rect 28476 31836 28532 31892
rect 28252 31666 28308 31668
rect 28252 31614 28254 31666
rect 28254 31614 28306 31666
rect 28306 31614 28308 31666
rect 28252 31612 28308 31614
rect 27804 30268 27860 30324
rect 28028 31164 28084 31220
rect 26916 29818 26972 29820
rect 26916 29766 26918 29818
rect 26918 29766 26970 29818
rect 26970 29766 26972 29818
rect 26916 29764 26972 29766
rect 27020 29818 27076 29820
rect 27020 29766 27022 29818
rect 27022 29766 27074 29818
rect 27074 29766 27076 29818
rect 27020 29764 27076 29766
rect 27124 29818 27180 29820
rect 27124 29766 27126 29818
rect 27126 29766 27178 29818
rect 27178 29766 27180 29818
rect 27124 29764 27180 29766
rect 27132 29484 27188 29540
rect 26916 28250 26972 28252
rect 26916 28198 26918 28250
rect 26918 28198 26970 28250
rect 26970 28198 26972 28250
rect 26916 28196 26972 28198
rect 27020 28250 27076 28252
rect 27020 28198 27022 28250
rect 27022 28198 27074 28250
rect 27074 28198 27076 28250
rect 27020 28196 27076 28198
rect 27124 28250 27180 28252
rect 27124 28198 27126 28250
rect 27126 28198 27178 28250
rect 27178 28198 27180 28250
rect 27124 28196 27180 28198
rect 27356 28140 27412 28196
rect 27132 27580 27188 27636
rect 26796 26796 26852 26852
rect 26916 26682 26972 26684
rect 26916 26630 26918 26682
rect 26918 26630 26970 26682
rect 26970 26630 26972 26682
rect 26916 26628 26972 26630
rect 27020 26682 27076 26684
rect 27020 26630 27022 26682
rect 27022 26630 27074 26682
rect 27074 26630 27076 26682
rect 27020 26628 27076 26630
rect 27124 26682 27180 26684
rect 27124 26630 27126 26682
rect 27126 26630 27178 26682
rect 27178 26630 27180 26682
rect 27124 26628 27180 26630
rect 26684 26236 26740 26292
rect 26460 25618 26516 25620
rect 26460 25566 26462 25618
rect 26462 25566 26514 25618
rect 26514 25566 26516 25618
rect 26460 25564 26516 25566
rect 25452 24892 25508 24948
rect 26012 25228 26068 25284
rect 25228 24722 25284 24724
rect 25228 24670 25230 24722
rect 25230 24670 25282 24722
rect 25282 24670 25284 24722
rect 25228 24668 25284 24670
rect 25564 24108 25620 24164
rect 26012 23996 26068 24052
rect 25452 23660 25508 23716
rect 25116 23548 25172 23604
rect 25228 22988 25284 23044
rect 25228 22092 25284 22148
rect 25340 21810 25396 21812
rect 25340 21758 25342 21810
rect 25342 21758 25394 21810
rect 25394 21758 25396 21810
rect 25340 21756 25396 21758
rect 25788 21980 25844 22036
rect 25228 20860 25284 20916
rect 24892 19404 24948 19460
rect 25004 20076 25060 20132
rect 24780 19122 24836 19124
rect 24780 19070 24782 19122
rect 24782 19070 24834 19122
rect 24834 19070 24836 19122
rect 24780 19068 24836 19070
rect 26460 23714 26516 23716
rect 26460 23662 26462 23714
rect 26462 23662 26514 23714
rect 26514 23662 26516 23714
rect 26460 23660 26516 23662
rect 26124 23436 26180 23492
rect 26460 23436 26516 23492
rect 26348 23378 26404 23380
rect 26348 23326 26350 23378
rect 26350 23326 26402 23378
rect 26402 23326 26404 23378
rect 26348 23324 26404 23326
rect 26236 21420 26292 21476
rect 25900 20076 25956 20132
rect 25228 19516 25284 19572
rect 25340 19458 25396 19460
rect 25340 19406 25342 19458
rect 25342 19406 25394 19458
rect 25394 19406 25396 19458
rect 25340 19404 25396 19406
rect 24668 18732 24724 18788
rect 25228 18956 25284 19012
rect 24556 18620 24612 18676
rect 23660 18284 23716 18340
rect 24220 18284 24276 18340
rect 23548 17890 23604 17892
rect 23548 17838 23550 17890
rect 23550 17838 23602 17890
rect 23602 17838 23604 17890
rect 23548 17836 23604 17838
rect 23996 17388 24052 17444
rect 23436 16882 23492 16884
rect 23436 16830 23438 16882
rect 23438 16830 23490 16882
rect 23490 16830 23492 16882
rect 23436 16828 23492 16830
rect 23436 15986 23492 15988
rect 23436 15934 23438 15986
rect 23438 15934 23490 15986
rect 23490 15934 23492 15986
rect 23436 15932 23492 15934
rect 22632 14922 22688 14924
rect 22632 14870 22634 14922
rect 22634 14870 22686 14922
rect 22686 14870 22688 14922
rect 22632 14868 22688 14870
rect 22736 14922 22792 14924
rect 22736 14870 22738 14922
rect 22738 14870 22790 14922
rect 22790 14870 22792 14922
rect 22736 14868 22792 14870
rect 22840 14922 22896 14924
rect 22840 14870 22842 14922
rect 22842 14870 22894 14922
rect 22894 14870 22896 14922
rect 22840 14868 22896 14870
rect 23212 14252 23268 14308
rect 22632 13354 22688 13356
rect 22632 13302 22634 13354
rect 22634 13302 22686 13354
rect 22686 13302 22688 13354
rect 22632 13300 22688 13302
rect 22736 13354 22792 13356
rect 22736 13302 22738 13354
rect 22738 13302 22790 13354
rect 22790 13302 22792 13354
rect 22736 13300 22792 13302
rect 22840 13354 22896 13356
rect 22840 13302 22842 13354
rect 22842 13302 22894 13354
rect 22894 13302 22896 13354
rect 22840 13300 22896 13302
rect 23212 13356 23268 13412
rect 23324 13916 23380 13972
rect 23100 13244 23156 13300
rect 23212 13132 23268 13188
rect 21756 12348 21812 12404
rect 22316 12572 22372 12628
rect 22988 12962 23044 12964
rect 22988 12910 22990 12962
rect 22990 12910 23042 12962
rect 23042 12910 23044 12962
rect 22988 12908 23044 12910
rect 23212 12572 23268 12628
rect 22540 12460 22596 12516
rect 21644 10892 21700 10948
rect 21420 10834 21476 10836
rect 21420 10782 21422 10834
rect 21422 10782 21474 10834
rect 21474 10782 21476 10834
rect 21420 10780 21476 10782
rect 21532 10610 21588 10612
rect 21532 10558 21534 10610
rect 21534 10558 21586 10610
rect 21586 10558 21588 10610
rect 21532 10556 21588 10558
rect 21420 9996 21476 10052
rect 21532 9100 21588 9156
rect 21308 8204 21364 8260
rect 20748 8092 20804 8148
rect 20524 7644 20580 7700
rect 20412 7532 20468 7588
rect 19180 7084 19236 7140
rect 20188 7308 20244 7364
rect 18172 6524 18228 6580
rect 17948 4956 18004 5012
rect 18060 5740 18116 5796
rect 17836 4508 17892 4564
rect 17612 4396 17668 4452
rect 18620 6578 18676 6580
rect 18620 6526 18622 6578
rect 18622 6526 18674 6578
rect 18674 6526 18676 6578
rect 18620 6524 18676 6526
rect 18396 6466 18452 6468
rect 18396 6414 18398 6466
rect 18398 6414 18450 6466
rect 18450 6414 18452 6466
rect 18396 6412 18452 6414
rect 18348 6298 18404 6300
rect 18348 6246 18350 6298
rect 18350 6246 18402 6298
rect 18402 6246 18404 6298
rect 18348 6244 18404 6246
rect 18452 6298 18508 6300
rect 18452 6246 18454 6298
rect 18454 6246 18506 6298
rect 18506 6246 18508 6298
rect 18452 6244 18508 6246
rect 18556 6298 18612 6300
rect 18556 6246 18558 6298
rect 18558 6246 18610 6298
rect 18610 6246 18612 6298
rect 18556 6244 18612 6246
rect 19292 6690 19348 6692
rect 19292 6638 19294 6690
rect 19294 6638 19346 6690
rect 19346 6638 19348 6690
rect 19292 6636 19348 6638
rect 19516 6524 19572 6580
rect 19292 5740 19348 5796
rect 19180 5068 19236 5124
rect 18348 4730 18404 4732
rect 18348 4678 18350 4730
rect 18350 4678 18402 4730
rect 18402 4678 18404 4730
rect 18348 4676 18404 4678
rect 18452 4730 18508 4732
rect 18452 4678 18454 4730
rect 18454 4678 18506 4730
rect 18506 4678 18508 4730
rect 18452 4676 18508 4678
rect 18556 4730 18612 4732
rect 18556 4678 18558 4730
rect 18558 4678 18610 4730
rect 18610 4678 18612 4730
rect 18556 4676 18612 4678
rect 19068 4844 19124 4900
rect 19292 4956 19348 5012
rect 18956 4562 19012 4564
rect 18956 4510 18958 4562
rect 18958 4510 19010 4562
rect 19010 4510 19012 4562
rect 18956 4508 19012 4510
rect 17836 3948 17892 4004
rect 20300 6690 20356 6692
rect 20300 6638 20302 6690
rect 20302 6638 20354 6690
rect 20354 6638 20356 6690
rect 20300 6636 20356 6638
rect 20412 6018 20468 6020
rect 20412 5966 20414 6018
rect 20414 5966 20466 6018
rect 20466 5966 20468 6018
rect 20412 5964 20468 5966
rect 21084 7644 21140 7700
rect 20972 7586 21028 7588
rect 20972 7534 20974 7586
rect 20974 7534 21026 7586
rect 21026 7534 21028 7586
rect 20972 7532 21028 7534
rect 21532 7586 21588 7588
rect 21532 7534 21534 7586
rect 21534 7534 21586 7586
rect 21586 7534 21588 7586
rect 21532 7532 21588 7534
rect 20860 7084 20916 7140
rect 21308 6690 21364 6692
rect 21308 6638 21310 6690
rect 21310 6638 21362 6690
rect 21362 6638 21364 6690
rect 21308 6636 21364 6638
rect 22632 11786 22688 11788
rect 22632 11734 22634 11786
rect 22634 11734 22686 11786
rect 22686 11734 22688 11786
rect 22632 11732 22688 11734
rect 22736 11786 22792 11788
rect 22736 11734 22738 11786
rect 22738 11734 22790 11786
rect 22790 11734 22792 11786
rect 22736 11732 22792 11734
rect 22840 11786 22896 11788
rect 22840 11734 22842 11786
rect 22842 11734 22894 11786
rect 22894 11734 22896 11786
rect 22840 11732 22896 11734
rect 21868 11116 21924 11172
rect 22764 11228 22820 11284
rect 22316 11004 22372 11060
rect 22764 10834 22820 10836
rect 22764 10782 22766 10834
rect 22766 10782 22818 10834
rect 22818 10782 22820 10834
rect 22764 10780 22820 10782
rect 22428 10722 22484 10724
rect 22428 10670 22430 10722
rect 22430 10670 22482 10722
rect 22482 10670 22484 10722
rect 22428 10668 22484 10670
rect 22632 10218 22688 10220
rect 22632 10166 22634 10218
rect 22634 10166 22686 10218
rect 22686 10166 22688 10218
rect 22632 10164 22688 10166
rect 22736 10218 22792 10220
rect 22736 10166 22738 10218
rect 22738 10166 22790 10218
rect 22790 10166 22792 10218
rect 22736 10164 22792 10166
rect 22840 10218 22896 10220
rect 22840 10166 22842 10218
rect 22842 10166 22894 10218
rect 22894 10166 22896 10218
rect 22840 10164 22896 10166
rect 23100 11564 23156 11620
rect 23212 11228 23268 11284
rect 23324 10834 23380 10836
rect 23324 10782 23326 10834
rect 23326 10782 23378 10834
rect 23378 10782 23380 10834
rect 23324 10780 23380 10782
rect 25564 19740 25620 19796
rect 25788 19852 25844 19908
rect 26460 22146 26516 22148
rect 26460 22094 26462 22146
rect 26462 22094 26514 22146
rect 26514 22094 26516 22146
rect 26460 22092 26516 22094
rect 26236 20130 26292 20132
rect 26236 20078 26238 20130
rect 26238 20078 26290 20130
rect 26290 20078 26292 20130
rect 26236 20076 26292 20078
rect 27132 25506 27188 25508
rect 27132 25454 27134 25506
rect 27134 25454 27186 25506
rect 27186 25454 27188 25506
rect 27132 25452 27188 25454
rect 26916 25114 26972 25116
rect 26916 25062 26918 25114
rect 26918 25062 26970 25114
rect 26970 25062 26972 25114
rect 26916 25060 26972 25062
rect 27020 25114 27076 25116
rect 27020 25062 27022 25114
rect 27022 25062 27074 25114
rect 27074 25062 27076 25114
rect 27020 25060 27076 25062
rect 27124 25114 27180 25116
rect 27124 25062 27126 25114
rect 27126 25062 27178 25114
rect 27178 25062 27180 25114
rect 27124 25060 27180 25062
rect 26796 24332 26852 24388
rect 27132 24220 27188 24276
rect 26916 23546 26972 23548
rect 26916 23494 26918 23546
rect 26918 23494 26970 23546
rect 26970 23494 26972 23546
rect 26916 23492 26972 23494
rect 27020 23546 27076 23548
rect 27020 23494 27022 23546
rect 27022 23494 27074 23546
rect 27074 23494 27076 23546
rect 27020 23492 27076 23494
rect 27124 23546 27180 23548
rect 27124 23494 27126 23546
rect 27126 23494 27178 23546
rect 27178 23494 27180 23546
rect 27124 23492 27180 23494
rect 27132 23212 27188 23268
rect 26684 22988 26740 23044
rect 27020 22876 27076 22932
rect 27804 27580 27860 27636
rect 27580 26514 27636 26516
rect 27580 26462 27582 26514
rect 27582 26462 27634 26514
rect 27634 26462 27636 26514
rect 27580 26460 27636 26462
rect 27468 25676 27524 25732
rect 28476 31052 28532 31108
rect 28588 30210 28644 30212
rect 28588 30158 28590 30210
rect 28590 30158 28642 30210
rect 28642 30158 28644 30210
rect 28588 30156 28644 30158
rect 28476 29596 28532 29652
rect 28476 28754 28532 28756
rect 28476 28702 28478 28754
rect 28478 28702 28530 28754
rect 28530 28702 28532 28754
rect 28476 28700 28532 28702
rect 28364 28418 28420 28420
rect 28364 28366 28366 28418
rect 28366 28366 28418 28418
rect 28418 28366 28420 28418
rect 28364 28364 28420 28366
rect 28140 26290 28196 26292
rect 28140 26238 28142 26290
rect 28142 26238 28194 26290
rect 28194 26238 28196 26290
rect 28140 26236 28196 26238
rect 27916 26012 27972 26068
rect 27692 25452 27748 25508
rect 27468 24556 27524 24612
rect 27580 23660 27636 23716
rect 27356 23378 27412 23380
rect 27356 23326 27358 23378
rect 27358 23326 27410 23378
rect 27410 23326 27412 23378
rect 27356 23324 27412 23326
rect 27244 22316 27300 22372
rect 26684 21644 26740 21700
rect 26916 21978 26972 21980
rect 26916 21926 26918 21978
rect 26918 21926 26970 21978
rect 26970 21926 26972 21978
rect 26916 21924 26972 21926
rect 27020 21978 27076 21980
rect 27020 21926 27022 21978
rect 27022 21926 27074 21978
rect 27074 21926 27076 21978
rect 27020 21924 27076 21926
rect 27124 21978 27180 21980
rect 27124 21926 27126 21978
rect 27126 21926 27178 21978
rect 27178 21926 27180 21978
rect 27124 21924 27180 21926
rect 27468 21756 27524 21812
rect 26684 21420 26740 21476
rect 27020 21420 27076 21476
rect 27468 21586 27524 21588
rect 27468 21534 27470 21586
rect 27470 21534 27522 21586
rect 27522 21534 27524 21586
rect 27468 21532 27524 21534
rect 27804 24332 27860 24388
rect 27804 23772 27860 23828
rect 28028 25730 28084 25732
rect 28028 25678 28030 25730
rect 28030 25678 28082 25730
rect 28082 25678 28084 25730
rect 28028 25676 28084 25678
rect 29148 32450 29204 32452
rect 29148 32398 29150 32450
rect 29150 32398 29202 32450
rect 29202 32398 29204 32450
rect 29148 32396 29204 32398
rect 29260 31836 29316 31892
rect 29708 31836 29764 31892
rect 29260 31164 29316 31220
rect 29148 30940 29204 30996
rect 28924 29314 28980 29316
rect 28924 29262 28926 29314
rect 28926 29262 28978 29314
rect 28978 29262 28980 29314
rect 28924 29260 28980 29262
rect 28700 28476 28756 28532
rect 28812 29148 28868 29204
rect 29932 30828 29988 30884
rect 29260 30210 29316 30212
rect 29260 30158 29262 30210
rect 29262 30158 29314 30210
rect 29314 30158 29316 30210
rect 29260 30156 29316 30158
rect 28812 26460 28868 26516
rect 28364 24780 28420 24836
rect 28364 24220 28420 24276
rect 28476 25340 28532 25396
rect 28588 24108 28644 24164
rect 28028 23548 28084 23604
rect 27804 22876 27860 22932
rect 28028 22764 28084 22820
rect 27916 22316 27972 22372
rect 27580 20972 27636 21028
rect 26796 20748 26852 20804
rect 27356 20690 27412 20692
rect 27356 20638 27358 20690
rect 27358 20638 27410 20690
rect 27410 20638 27412 20690
rect 27356 20636 27412 20638
rect 27580 20578 27636 20580
rect 27580 20526 27582 20578
rect 27582 20526 27634 20578
rect 27634 20526 27636 20578
rect 27580 20524 27636 20526
rect 26916 20410 26972 20412
rect 26916 20358 26918 20410
rect 26918 20358 26970 20410
rect 26970 20358 26972 20410
rect 26916 20356 26972 20358
rect 27020 20410 27076 20412
rect 27020 20358 27022 20410
rect 27022 20358 27074 20410
rect 27074 20358 27076 20410
rect 27020 20356 27076 20358
rect 27124 20410 27180 20412
rect 27124 20358 27126 20410
rect 27126 20358 27178 20410
rect 27178 20358 27180 20410
rect 27124 20356 27180 20358
rect 27132 20188 27188 20244
rect 27804 20188 27860 20244
rect 26572 19852 26628 19908
rect 25788 19628 25844 19684
rect 25340 18396 25396 18452
rect 25564 18396 25620 18452
rect 25228 18172 25284 18228
rect 24332 17666 24388 17668
rect 24332 17614 24334 17666
rect 24334 17614 24386 17666
rect 24386 17614 24388 17666
rect 24332 17612 24388 17614
rect 24444 17052 24500 17108
rect 23884 16098 23940 16100
rect 23884 16046 23886 16098
rect 23886 16046 23938 16098
rect 23938 16046 23940 16098
rect 23884 16044 23940 16046
rect 24220 16098 24276 16100
rect 24220 16046 24222 16098
rect 24222 16046 24274 16098
rect 24274 16046 24276 16098
rect 24220 16044 24276 16046
rect 24444 15372 24500 15428
rect 24556 15932 24612 15988
rect 24108 14700 24164 14756
rect 23996 14364 24052 14420
rect 23996 13244 24052 13300
rect 24668 15820 24724 15876
rect 25340 17948 25396 18004
rect 25004 17500 25060 17556
rect 25228 16940 25284 16996
rect 25676 17612 25732 17668
rect 25452 17388 25508 17444
rect 24668 14588 24724 14644
rect 24332 13074 24388 13076
rect 24332 13022 24334 13074
rect 24334 13022 24386 13074
rect 24386 13022 24388 13074
rect 24332 13020 24388 13022
rect 25340 16380 25396 16436
rect 23660 12402 23716 12404
rect 23660 12350 23662 12402
rect 23662 12350 23714 12402
rect 23714 12350 23716 12402
rect 23660 12348 23716 12350
rect 24220 12460 24276 12516
rect 24668 13132 24724 13188
rect 24668 12124 24724 12180
rect 23548 10780 23604 10836
rect 23660 11228 23716 11284
rect 23772 11004 23828 11060
rect 25116 15036 25172 15092
rect 25228 15148 25284 15204
rect 25452 16098 25508 16100
rect 25452 16046 25454 16098
rect 25454 16046 25506 16098
rect 25506 16046 25508 16098
rect 25452 16044 25508 16046
rect 25228 13970 25284 13972
rect 25228 13918 25230 13970
rect 25230 13918 25282 13970
rect 25282 13918 25284 13970
rect 25228 13916 25284 13918
rect 25452 15148 25508 15204
rect 25788 16940 25844 16996
rect 25788 16716 25844 16772
rect 25676 15820 25732 15876
rect 26012 19516 26068 19572
rect 26012 18844 26068 18900
rect 26012 18562 26068 18564
rect 26012 18510 26014 18562
rect 26014 18510 26066 18562
rect 26066 18510 26068 18562
rect 26012 18508 26068 18510
rect 26684 19794 26740 19796
rect 26684 19742 26686 19794
rect 26686 19742 26738 19794
rect 26738 19742 26740 19794
rect 26684 19740 26740 19742
rect 27356 19964 27412 20020
rect 26796 19628 26852 19684
rect 27580 19404 27636 19460
rect 27020 19346 27076 19348
rect 27020 19294 27022 19346
rect 27022 19294 27074 19346
rect 27074 19294 27076 19346
rect 27020 19292 27076 19294
rect 28252 23660 28308 23716
rect 28364 23436 28420 23492
rect 28588 23548 28644 23604
rect 28812 24220 28868 24276
rect 29260 28028 29316 28084
rect 29148 25564 29204 25620
rect 29036 24722 29092 24724
rect 29036 24670 29038 24722
rect 29038 24670 29090 24722
rect 29090 24670 29092 24722
rect 29036 24668 29092 24670
rect 29596 25730 29652 25732
rect 29596 25678 29598 25730
rect 29598 25678 29650 25730
rect 29650 25678 29652 25730
rect 29596 25676 29652 25678
rect 29484 25506 29540 25508
rect 29484 25454 29486 25506
rect 29486 25454 29538 25506
rect 29538 25454 29540 25506
rect 29484 25452 29540 25454
rect 30044 27356 30100 27412
rect 29932 27132 29988 27188
rect 29372 25004 29428 25060
rect 30380 32844 30436 32900
rect 30380 30716 30436 30772
rect 30604 30994 30660 30996
rect 30604 30942 30606 30994
rect 30606 30942 30658 30994
rect 30658 30942 30660 30994
rect 30604 30940 30660 30942
rect 30268 28364 30324 28420
rect 30380 28082 30436 28084
rect 30380 28030 30382 28082
rect 30382 28030 30434 28082
rect 30434 28030 30436 28082
rect 30380 28028 30436 28030
rect 30492 27858 30548 27860
rect 30492 27806 30494 27858
rect 30494 27806 30546 27858
rect 30546 27806 30548 27858
rect 30492 27804 30548 27806
rect 30268 27468 30324 27524
rect 30828 31218 30884 31220
rect 30828 31166 30830 31218
rect 30830 31166 30882 31218
rect 30882 31166 30884 31218
rect 30828 31164 30884 31166
rect 30828 30882 30884 30884
rect 30828 30830 30830 30882
rect 30830 30830 30882 30882
rect 30882 30830 30884 30882
rect 30828 30828 30884 30830
rect 30716 27916 30772 27972
rect 29372 24834 29428 24836
rect 29372 24782 29374 24834
rect 29374 24782 29426 24834
rect 29426 24782 29428 24834
rect 29372 24780 29428 24782
rect 29596 24498 29652 24500
rect 29596 24446 29598 24498
rect 29598 24446 29650 24498
rect 29650 24446 29652 24498
rect 29596 24444 29652 24446
rect 28252 23266 28308 23268
rect 28252 23214 28254 23266
rect 28254 23214 28306 23266
rect 28306 23214 28308 23266
rect 28252 23212 28308 23214
rect 29036 23436 29092 23492
rect 28812 22876 28868 22932
rect 28924 23100 28980 23156
rect 28252 20802 28308 20804
rect 28252 20750 28254 20802
rect 28254 20750 28306 20802
rect 28306 20750 28308 20802
rect 28252 20748 28308 20750
rect 28588 21980 28644 22036
rect 28812 21196 28868 21252
rect 28588 20636 28644 20692
rect 28364 19740 28420 19796
rect 28588 20188 28644 20244
rect 28028 19404 28084 19460
rect 28364 19292 28420 19348
rect 26572 19122 26628 19124
rect 26572 19070 26574 19122
rect 26574 19070 26626 19122
rect 26626 19070 26628 19122
rect 26572 19068 26628 19070
rect 26124 18396 26180 18452
rect 26012 17500 26068 17556
rect 26012 16828 26068 16884
rect 25900 16380 25956 16436
rect 25900 16156 25956 16212
rect 26348 18844 26404 18900
rect 26348 18060 26404 18116
rect 26348 17724 26404 17780
rect 26124 15596 26180 15652
rect 26236 17052 26292 17108
rect 25676 15314 25732 15316
rect 25676 15262 25678 15314
rect 25678 15262 25730 15314
rect 25730 15262 25732 15314
rect 25676 15260 25732 15262
rect 28028 19010 28084 19012
rect 28028 18958 28030 19010
rect 28030 18958 28082 19010
rect 28082 18958 28084 19010
rect 28028 18956 28084 18958
rect 28812 20636 28868 20692
rect 26916 18842 26972 18844
rect 26916 18790 26918 18842
rect 26918 18790 26970 18842
rect 26970 18790 26972 18842
rect 26916 18788 26972 18790
rect 27020 18842 27076 18844
rect 27020 18790 27022 18842
rect 27022 18790 27074 18842
rect 27074 18790 27076 18842
rect 27020 18788 27076 18790
rect 27124 18842 27180 18844
rect 27124 18790 27126 18842
rect 27126 18790 27178 18842
rect 27178 18790 27180 18842
rect 27124 18788 27180 18790
rect 28028 18732 28084 18788
rect 26796 17836 26852 17892
rect 27020 18450 27076 18452
rect 27020 18398 27022 18450
rect 27022 18398 27074 18450
rect 27074 18398 27076 18450
rect 27020 18396 27076 18398
rect 27356 18396 27412 18452
rect 27580 18396 27636 18452
rect 27132 18172 27188 18228
rect 27356 18172 27412 18228
rect 26684 17388 26740 17444
rect 25788 14476 25844 14532
rect 25340 12348 25396 12404
rect 25452 13020 25508 13076
rect 25452 12684 25508 12740
rect 25788 13858 25844 13860
rect 25788 13806 25790 13858
rect 25790 13806 25842 13858
rect 25842 13806 25844 13858
rect 25788 13804 25844 13806
rect 25900 14028 25956 14084
rect 26348 14140 26404 14196
rect 26460 14028 26516 14084
rect 25676 11676 25732 11732
rect 25564 11564 25620 11620
rect 25004 11170 25060 11172
rect 25004 11118 25006 11170
rect 25006 11118 25058 11170
rect 25058 11118 25060 11170
rect 25004 11116 25060 11118
rect 24892 11004 24948 11060
rect 24220 10610 24276 10612
rect 24220 10558 24222 10610
rect 24222 10558 24274 10610
rect 24274 10558 24276 10610
rect 24220 10556 24276 10558
rect 24108 10108 24164 10164
rect 22540 9996 22596 10052
rect 25116 10668 25172 10724
rect 22764 9042 22820 9044
rect 22764 8990 22766 9042
rect 22766 8990 22818 9042
rect 22818 8990 22820 9042
rect 22764 8988 22820 8990
rect 24108 9154 24164 9156
rect 24108 9102 24110 9154
rect 24110 9102 24162 9154
rect 24162 9102 24164 9154
rect 24108 9100 24164 9102
rect 24556 9772 24612 9828
rect 25228 10610 25284 10612
rect 25228 10558 25230 10610
rect 25230 10558 25282 10610
rect 25282 10558 25284 10610
rect 25228 10556 25284 10558
rect 25228 9996 25284 10052
rect 25228 9266 25284 9268
rect 25228 9214 25230 9266
rect 25230 9214 25282 9266
rect 25282 9214 25284 9266
rect 25228 9212 25284 9214
rect 24332 9100 24388 9156
rect 24220 8988 24276 9044
rect 24556 9154 24612 9156
rect 24556 9102 24558 9154
rect 24558 9102 24610 9154
rect 24610 9102 24612 9154
rect 24556 9100 24612 9102
rect 22632 8650 22688 8652
rect 22632 8598 22634 8650
rect 22634 8598 22686 8650
rect 22686 8598 22688 8650
rect 22632 8596 22688 8598
rect 22736 8650 22792 8652
rect 22736 8598 22738 8650
rect 22738 8598 22790 8650
rect 22790 8598 22792 8650
rect 22736 8596 22792 8598
rect 22840 8650 22896 8652
rect 22840 8598 22842 8650
rect 22842 8598 22894 8650
rect 22894 8598 22896 8650
rect 22840 8596 22896 8598
rect 21756 6636 21812 6692
rect 20748 6412 20804 6468
rect 20076 4956 20132 5012
rect 20636 5628 20692 5684
rect 18396 4172 18452 4228
rect 17500 3612 17556 3668
rect 17612 3554 17668 3556
rect 17612 3502 17614 3554
rect 17614 3502 17666 3554
rect 17666 3502 17668 3554
rect 17612 3500 17668 3502
rect 18620 3666 18676 3668
rect 18620 3614 18622 3666
rect 18622 3614 18674 3666
rect 18674 3614 18676 3666
rect 18620 3612 18676 3614
rect 19068 3612 19124 3668
rect 18396 3500 18452 3556
rect 18348 3162 18404 3164
rect 18348 3110 18350 3162
rect 18350 3110 18402 3162
rect 18402 3110 18404 3162
rect 18348 3108 18404 3110
rect 18452 3162 18508 3164
rect 18452 3110 18454 3162
rect 18454 3110 18506 3162
rect 18506 3110 18508 3162
rect 18452 3108 18508 3110
rect 18556 3162 18612 3164
rect 18556 3110 18558 3162
rect 18558 3110 18610 3162
rect 18610 3110 18612 3162
rect 18556 3108 18612 3110
rect 22092 7308 22148 7364
rect 22632 7082 22688 7084
rect 22632 7030 22634 7082
rect 22634 7030 22686 7082
rect 22686 7030 22688 7082
rect 22632 7028 22688 7030
rect 22736 7082 22792 7084
rect 22736 7030 22738 7082
rect 22738 7030 22790 7082
rect 22790 7030 22792 7082
rect 22736 7028 22792 7030
rect 22840 7082 22896 7084
rect 22840 7030 22842 7082
rect 22842 7030 22894 7082
rect 22894 7030 22896 7082
rect 22840 7028 22896 7030
rect 23996 8764 24052 8820
rect 23772 8428 23828 8484
rect 23436 7474 23492 7476
rect 23436 7422 23438 7474
rect 23438 7422 23490 7474
rect 23490 7422 23492 7474
rect 23436 7420 23492 7422
rect 23548 7362 23604 7364
rect 23548 7310 23550 7362
rect 23550 7310 23602 7362
rect 23602 7310 23604 7362
rect 23548 7308 23604 7310
rect 22988 5740 23044 5796
rect 21868 5682 21924 5684
rect 21868 5630 21870 5682
rect 21870 5630 21922 5682
rect 21922 5630 21924 5682
rect 21868 5628 21924 5630
rect 22632 5514 22688 5516
rect 22632 5462 22634 5514
rect 22634 5462 22686 5514
rect 22686 5462 22688 5514
rect 22632 5460 22688 5462
rect 22736 5514 22792 5516
rect 22736 5462 22738 5514
rect 22738 5462 22790 5514
rect 22790 5462 22792 5514
rect 22736 5460 22792 5462
rect 22840 5514 22896 5516
rect 22840 5462 22842 5514
rect 22842 5462 22894 5514
rect 22894 5462 22896 5514
rect 22840 5460 22896 5462
rect 22540 5234 22596 5236
rect 22540 5182 22542 5234
rect 22542 5182 22594 5234
rect 22594 5182 22596 5234
rect 22540 5180 22596 5182
rect 22876 4956 22932 5012
rect 22764 4508 22820 4564
rect 22652 4450 22708 4452
rect 22652 4398 22654 4450
rect 22654 4398 22706 4450
rect 22706 4398 22708 4450
rect 22652 4396 22708 4398
rect 24444 8428 24500 8484
rect 23884 7756 23940 7812
rect 23772 6748 23828 6804
rect 25676 11116 25732 11172
rect 25900 12178 25956 12180
rect 25900 12126 25902 12178
rect 25902 12126 25954 12178
rect 25954 12126 25956 12178
rect 25900 12124 25956 12126
rect 25900 11954 25956 11956
rect 25900 11902 25902 11954
rect 25902 11902 25954 11954
rect 25954 11902 25956 11954
rect 25900 11900 25956 11902
rect 26348 13020 26404 13076
rect 26916 17274 26972 17276
rect 26916 17222 26918 17274
rect 26918 17222 26970 17274
rect 26970 17222 26972 17274
rect 26916 17220 26972 17222
rect 27020 17274 27076 17276
rect 27020 17222 27022 17274
rect 27022 17222 27074 17274
rect 27074 17222 27076 17274
rect 27020 17220 27076 17222
rect 27124 17274 27180 17276
rect 27124 17222 27126 17274
rect 27126 17222 27178 17274
rect 27178 17222 27180 17274
rect 27124 17220 27180 17222
rect 27468 17388 27524 17444
rect 27580 17500 27636 17556
rect 26684 16994 26740 16996
rect 26684 16942 26686 16994
rect 26686 16942 26738 16994
rect 26738 16942 26740 16994
rect 26684 16940 26740 16942
rect 27356 17052 27412 17108
rect 26796 16604 26852 16660
rect 27916 18508 27972 18564
rect 28140 18226 28196 18228
rect 28140 18174 28142 18226
rect 28142 18174 28194 18226
rect 28194 18174 28196 18226
rect 28140 18172 28196 18174
rect 28028 17836 28084 17892
rect 27244 16658 27300 16660
rect 27244 16606 27246 16658
rect 27246 16606 27298 16658
rect 27298 16606 27300 16658
rect 27244 16604 27300 16606
rect 26908 15986 26964 15988
rect 26908 15934 26910 15986
rect 26910 15934 26962 15986
rect 26962 15934 26964 15986
rect 26908 15932 26964 15934
rect 26796 15820 26852 15876
rect 27020 15874 27076 15876
rect 27020 15822 27022 15874
rect 27022 15822 27074 15874
rect 27074 15822 27076 15874
rect 27020 15820 27076 15822
rect 27468 16268 27524 16324
rect 26916 15706 26972 15708
rect 26916 15654 26918 15706
rect 26918 15654 26970 15706
rect 26970 15654 26972 15706
rect 26916 15652 26972 15654
rect 27020 15706 27076 15708
rect 27020 15654 27022 15706
rect 27022 15654 27074 15706
rect 27074 15654 27076 15706
rect 27020 15652 27076 15654
rect 27124 15706 27180 15708
rect 27124 15654 27126 15706
rect 27126 15654 27178 15706
rect 27178 15654 27180 15706
rect 27124 15652 27180 15654
rect 27132 15314 27188 15316
rect 27132 15262 27134 15314
rect 27134 15262 27186 15314
rect 27186 15262 27188 15314
rect 27132 15260 27188 15262
rect 26908 15036 26964 15092
rect 26916 14138 26972 14140
rect 26916 14086 26918 14138
rect 26918 14086 26970 14138
rect 26970 14086 26972 14138
rect 26916 14084 26972 14086
rect 27020 14138 27076 14140
rect 27020 14086 27022 14138
rect 27022 14086 27074 14138
rect 27074 14086 27076 14138
rect 27020 14084 27076 14086
rect 27124 14138 27180 14140
rect 27124 14086 27126 14138
rect 27126 14086 27178 14138
rect 27178 14086 27180 14138
rect 27124 14084 27180 14086
rect 28028 16770 28084 16772
rect 28028 16718 28030 16770
rect 28030 16718 28082 16770
rect 28082 16718 28084 16770
rect 28028 16716 28084 16718
rect 28028 16492 28084 16548
rect 27692 15874 27748 15876
rect 27692 15822 27694 15874
rect 27694 15822 27746 15874
rect 27746 15822 27748 15874
rect 27692 15820 27748 15822
rect 27468 15484 27524 15540
rect 27356 14924 27412 14980
rect 27804 15314 27860 15316
rect 27804 15262 27806 15314
rect 27806 15262 27858 15314
rect 27858 15262 27860 15314
rect 27804 15260 27860 15262
rect 27580 14924 27636 14980
rect 27580 14476 27636 14532
rect 27692 14812 27748 14868
rect 26684 13132 26740 13188
rect 26796 13074 26852 13076
rect 26796 13022 26798 13074
rect 26798 13022 26850 13074
rect 26850 13022 26852 13074
rect 26796 13020 26852 13022
rect 27580 13804 27636 13860
rect 27132 13468 27188 13524
rect 27580 13580 27636 13636
rect 27244 13356 27300 13412
rect 26916 12570 26972 12572
rect 26916 12518 26918 12570
rect 26918 12518 26970 12570
rect 26970 12518 26972 12570
rect 26916 12516 26972 12518
rect 27020 12570 27076 12572
rect 27020 12518 27022 12570
rect 27022 12518 27074 12570
rect 27074 12518 27076 12570
rect 27020 12516 27076 12518
rect 27124 12570 27180 12572
rect 27124 12518 27126 12570
rect 27126 12518 27178 12570
rect 27178 12518 27180 12570
rect 27124 12516 27180 12518
rect 26908 11900 26964 11956
rect 26916 11002 26972 11004
rect 26916 10950 26918 11002
rect 26918 10950 26970 11002
rect 26970 10950 26972 11002
rect 26916 10948 26972 10950
rect 27020 11002 27076 11004
rect 27020 10950 27022 11002
rect 27022 10950 27074 11002
rect 27074 10950 27076 11002
rect 27020 10948 27076 10950
rect 27124 11002 27180 11004
rect 27124 10950 27126 11002
rect 27126 10950 27178 11002
rect 27178 10950 27180 11002
rect 27124 10948 27180 10950
rect 26908 10668 26964 10724
rect 27468 13356 27524 13412
rect 27468 12572 27524 12628
rect 27580 12124 27636 12180
rect 28588 18956 28644 19012
rect 28700 19180 28756 19236
rect 29148 23100 29204 23156
rect 29260 23660 29316 23716
rect 29036 22316 29092 22372
rect 29148 22428 29204 22484
rect 29260 22316 29316 22372
rect 29260 21644 29316 21700
rect 30044 25004 30100 25060
rect 29820 24220 29876 24276
rect 29932 23154 29988 23156
rect 29932 23102 29934 23154
rect 29934 23102 29986 23154
rect 29986 23102 29988 23154
rect 29932 23100 29988 23102
rect 29820 22876 29876 22932
rect 29820 22428 29876 22484
rect 29932 22092 29988 22148
rect 30044 22204 30100 22260
rect 28700 17836 28756 17892
rect 28588 17666 28644 17668
rect 28588 17614 28590 17666
rect 28590 17614 28642 17666
rect 28642 17614 28644 17666
rect 28588 17612 28644 17614
rect 28476 17442 28532 17444
rect 28476 17390 28478 17442
rect 28478 17390 28530 17442
rect 28530 17390 28532 17442
rect 28476 17388 28532 17390
rect 28364 16994 28420 16996
rect 28364 16942 28366 16994
rect 28366 16942 28418 16994
rect 28418 16942 28420 16994
rect 28364 16940 28420 16942
rect 28476 16380 28532 16436
rect 28252 15260 28308 15316
rect 28364 16268 28420 16324
rect 27916 14700 27972 14756
rect 27916 14418 27972 14420
rect 27916 14366 27918 14418
rect 27918 14366 27970 14418
rect 27970 14366 27972 14418
rect 27916 14364 27972 14366
rect 28252 15036 28308 15092
rect 28140 13858 28196 13860
rect 28140 13806 28142 13858
rect 28142 13806 28194 13858
rect 28194 13806 28196 13858
rect 28140 13804 28196 13806
rect 27916 13356 27972 13412
rect 27804 12796 27860 12852
rect 28588 16156 28644 16212
rect 28588 15932 28644 15988
rect 28924 18508 28980 18564
rect 29148 20636 29204 20692
rect 29372 20188 29428 20244
rect 29484 20018 29540 20020
rect 29484 19966 29486 20018
rect 29486 19966 29538 20018
rect 29538 19966 29540 20018
rect 29484 19964 29540 19966
rect 29260 19740 29316 19796
rect 29036 17836 29092 17892
rect 29148 19628 29204 19684
rect 29260 19404 29316 19460
rect 29932 21644 29988 21700
rect 29708 19404 29764 19460
rect 29484 19180 29540 19236
rect 29372 19068 29428 19124
rect 30044 21532 30100 21588
rect 30604 25116 30660 25172
rect 30492 24108 30548 24164
rect 30716 24444 30772 24500
rect 30268 23100 30324 23156
rect 30268 22652 30324 22708
rect 30604 22876 30660 22932
rect 31200 33738 31256 33740
rect 31200 33686 31202 33738
rect 31202 33686 31254 33738
rect 31254 33686 31256 33738
rect 31200 33684 31256 33686
rect 31304 33738 31360 33740
rect 31304 33686 31306 33738
rect 31306 33686 31358 33738
rect 31358 33686 31360 33738
rect 31304 33684 31360 33686
rect 31408 33738 31464 33740
rect 31408 33686 31410 33738
rect 31410 33686 31462 33738
rect 31462 33686 31464 33738
rect 31408 33684 31464 33686
rect 32956 33404 33012 33460
rect 33740 33628 33796 33684
rect 31836 32562 31892 32564
rect 31836 32510 31838 32562
rect 31838 32510 31890 32562
rect 31890 32510 31892 32562
rect 31836 32508 31892 32510
rect 31724 32338 31780 32340
rect 31724 32286 31726 32338
rect 31726 32286 31778 32338
rect 31778 32286 31780 32338
rect 31724 32284 31780 32286
rect 31052 32172 31108 32228
rect 31200 32170 31256 32172
rect 31200 32118 31202 32170
rect 31202 32118 31254 32170
rect 31254 32118 31256 32170
rect 31200 32116 31256 32118
rect 31304 32170 31360 32172
rect 31304 32118 31306 32170
rect 31306 32118 31358 32170
rect 31358 32118 31360 32170
rect 31304 32116 31360 32118
rect 31408 32170 31464 32172
rect 31408 32118 31410 32170
rect 31410 32118 31462 32170
rect 31462 32118 31464 32170
rect 31408 32116 31464 32118
rect 31388 31612 31444 31668
rect 31052 30994 31108 30996
rect 31052 30942 31054 30994
rect 31054 30942 31106 30994
rect 31106 30942 31108 30994
rect 31052 30940 31108 30942
rect 31724 31106 31780 31108
rect 31724 31054 31726 31106
rect 31726 31054 31778 31106
rect 31778 31054 31780 31106
rect 31724 31052 31780 31054
rect 32172 31836 32228 31892
rect 31388 30828 31444 30884
rect 31200 30602 31256 30604
rect 31200 30550 31202 30602
rect 31202 30550 31254 30602
rect 31254 30550 31256 30602
rect 31200 30548 31256 30550
rect 31304 30602 31360 30604
rect 31304 30550 31306 30602
rect 31306 30550 31358 30602
rect 31358 30550 31360 30602
rect 31304 30548 31360 30550
rect 31408 30602 31464 30604
rect 31408 30550 31410 30602
rect 31410 30550 31462 30602
rect 31462 30550 31464 30602
rect 31408 30548 31464 30550
rect 31200 29034 31256 29036
rect 31200 28982 31202 29034
rect 31202 28982 31254 29034
rect 31254 28982 31256 29034
rect 31200 28980 31256 28982
rect 31304 29034 31360 29036
rect 31304 28982 31306 29034
rect 31306 28982 31358 29034
rect 31358 28982 31360 29034
rect 31304 28980 31360 28982
rect 31408 29034 31464 29036
rect 31408 28982 31410 29034
rect 31410 28982 31462 29034
rect 31462 28982 31464 29034
rect 31408 28980 31464 28982
rect 31276 27746 31332 27748
rect 31276 27694 31278 27746
rect 31278 27694 31330 27746
rect 31330 27694 31332 27746
rect 31276 27692 31332 27694
rect 31612 27580 31668 27636
rect 31200 27466 31256 27468
rect 31200 27414 31202 27466
rect 31202 27414 31254 27466
rect 31254 27414 31256 27466
rect 31200 27412 31256 27414
rect 31304 27466 31360 27468
rect 31304 27414 31306 27466
rect 31306 27414 31358 27466
rect 31358 27414 31360 27466
rect 31304 27412 31360 27414
rect 31408 27466 31464 27468
rect 31408 27414 31410 27466
rect 31410 27414 31462 27466
rect 31462 27414 31464 27466
rect 31408 27412 31464 27414
rect 32060 30994 32116 30996
rect 32060 30942 32062 30994
rect 32062 30942 32114 30994
rect 32114 30942 32116 30994
rect 32060 30940 32116 30942
rect 32284 32620 32340 32676
rect 32732 31948 32788 32004
rect 32284 31724 32340 31780
rect 32396 30940 32452 30996
rect 32396 30770 32452 30772
rect 32396 30718 32398 30770
rect 32398 30718 32450 30770
rect 32450 30718 32452 30770
rect 32396 30716 32452 30718
rect 32508 30322 32564 30324
rect 32508 30270 32510 30322
rect 32510 30270 32562 30322
rect 32562 30270 32564 30322
rect 32508 30268 32564 30270
rect 32620 29932 32676 29988
rect 32284 29596 32340 29652
rect 32508 29484 32564 29540
rect 32060 28140 32116 28196
rect 32172 27970 32228 27972
rect 32172 27918 32174 27970
rect 32174 27918 32226 27970
rect 32226 27918 32228 27970
rect 32172 27916 32228 27918
rect 32060 27746 32116 27748
rect 32060 27694 32062 27746
rect 32062 27694 32114 27746
rect 32114 27694 32116 27746
rect 32060 27692 32116 27694
rect 32172 27580 32228 27636
rect 31200 25898 31256 25900
rect 31200 25846 31202 25898
rect 31202 25846 31254 25898
rect 31254 25846 31256 25898
rect 31200 25844 31256 25846
rect 31304 25898 31360 25900
rect 31304 25846 31306 25898
rect 31306 25846 31358 25898
rect 31358 25846 31360 25898
rect 31304 25844 31360 25846
rect 31408 25898 31464 25900
rect 31408 25846 31410 25898
rect 31410 25846 31462 25898
rect 31462 25846 31464 25898
rect 31408 25844 31464 25846
rect 31052 25004 31108 25060
rect 30940 24892 30996 24948
rect 30828 22876 30884 22932
rect 30828 22258 30884 22260
rect 30828 22206 30830 22258
rect 30830 22206 30882 22258
rect 30882 22206 30884 22258
rect 30828 22204 30884 22206
rect 30940 22316 30996 22372
rect 31164 24556 31220 24612
rect 31612 25452 31668 25508
rect 31200 24330 31256 24332
rect 31200 24278 31202 24330
rect 31202 24278 31254 24330
rect 31254 24278 31256 24330
rect 31200 24276 31256 24278
rect 31304 24330 31360 24332
rect 31304 24278 31306 24330
rect 31306 24278 31358 24330
rect 31358 24278 31360 24330
rect 31304 24276 31360 24278
rect 31408 24330 31464 24332
rect 31408 24278 31410 24330
rect 31410 24278 31462 24330
rect 31462 24278 31464 24330
rect 31612 24332 31668 24388
rect 31408 24276 31464 24278
rect 32396 27858 32452 27860
rect 32396 27806 32398 27858
rect 32398 27806 32450 27858
rect 32450 27806 32452 27858
rect 32396 27804 32452 27806
rect 32172 24892 32228 24948
rect 31836 23100 31892 23156
rect 31724 22988 31780 23044
rect 31200 22762 31256 22764
rect 31200 22710 31202 22762
rect 31202 22710 31254 22762
rect 31254 22710 31256 22762
rect 31200 22708 31256 22710
rect 31304 22762 31360 22764
rect 31304 22710 31306 22762
rect 31306 22710 31358 22762
rect 31358 22710 31360 22762
rect 31304 22708 31360 22710
rect 31408 22762 31464 22764
rect 31408 22710 31410 22762
rect 31410 22710 31462 22762
rect 31462 22710 31464 22762
rect 31408 22708 31464 22710
rect 31612 22540 31668 22596
rect 31388 22370 31444 22372
rect 31388 22318 31390 22370
rect 31390 22318 31442 22370
rect 31442 22318 31444 22370
rect 31388 22316 31444 22318
rect 31052 21644 31108 21700
rect 30492 21532 30548 21588
rect 30380 21420 30436 21476
rect 30268 20636 30324 20692
rect 30156 19628 30212 19684
rect 30156 19404 30212 19460
rect 30044 19180 30100 19236
rect 29932 19122 29988 19124
rect 29932 19070 29934 19122
rect 29934 19070 29986 19122
rect 29986 19070 29988 19122
rect 29932 19068 29988 19070
rect 29148 17276 29204 17332
rect 29148 16268 29204 16324
rect 29260 16210 29316 16212
rect 29260 16158 29262 16210
rect 29262 16158 29314 16210
rect 29314 16158 29316 16210
rect 29260 16156 29316 16158
rect 28700 15820 28756 15876
rect 28476 15090 28532 15092
rect 28476 15038 28478 15090
rect 28478 15038 28530 15090
rect 28530 15038 28532 15090
rect 28476 15036 28532 15038
rect 28588 14812 28644 14868
rect 28588 13244 28644 13300
rect 28364 13020 28420 13076
rect 28924 14924 28980 14980
rect 28812 14700 28868 14756
rect 28364 12796 28420 12852
rect 28252 11676 28308 11732
rect 28476 11618 28532 11620
rect 28476 11566 28478 11618
rect 28478 11566 28530 11618
rect 28530 11566 28532 11618
rect 28476 11564 28532 11566
rect 28364 10668 28420 10724
rect 28028 9548 28084 9604
rect 26916 9434 26972 9436
rect 26916 9382 26918 9434
rect 26918 9382 26970 9434
rect 26970 9382 26972 9434
rect 26916 9380 26972 9382
rect 27020 9434 27076 9436
rect 27020 9382 27022 9434
rect 27022 9382 27074 9434
rect 27074 9382 27076 9434
rect 27020 9380 27076 9382
rect 27124 9434 27180 9436
rect 27124 9382 27126 9434
rect 27126 9382 27178 9434
rect 27178 9382 27180 9434
rect 27124 9380 27180 9382
rect 26012 9266 26068 9268
rect 26012 9214 26014 9266
rect 26014 9214 26066 9266
rect 26066 9214 26068 9266
rect 26012 9212 26068 9214
rect 25788 8204 25844 8260
rect 27356 9042 27412 9044
rect 27356 8990 27358 9042
rect 27358 8990 27410 9042
rect 27410 8990 27412 9042
rect 27356 8988 27412 8990
rect 26684 8092 26740 8148
rect 26796 8204 26852 8260
rect 25900 7756 25956 7812
rect 24220 7474 24276 7476
rect 24220 7422 24222 7474
rect 24222 7422 24274 7474
rect 24274 7422 24276 7474
rect 24220 7420 24276 7422
rect 24556 6578 24612 6580
rect 24556 6526 24558 6578
rect 24558 6526 24610 6578
rect 24610 6526 24612 6578
rect 24556 6524 24612 6526
rect 24332 6412 24388 6468
rect 24556 6300 24612 6356
rect 24444 5964 24500 6020
rect 24108 5068 24164 5124
rect 23212 4562 23268 4564
rect 23212 4510 23214 4562
rect 23214 4510 23266 4562
rect 23266 4510 23268 4562
rect 23212 4508 23268 4510
rect 22632 3946 22688 3948
rect 22632 3894 22634 3946
rect 22634 3894 22686 3946
rect 22686 3894 22688 3946
rect 22632 3892 22688 3894
rect 22736 3946 22792 3948
rect 22736 3894 22738 3946
rect 22738 3894 22790 3946
rect 22790 3894 22792 3946
rect 22736 3892 22792 3894
rect 22840 3946 22896 3948
rect 22840 3894 22842 3946
rect 22842 3894 22894 3946
rect 22894 3894 22896 3946
rect 22840 3892 22896 3894
rect 21868 3666 21924 3668
rect 21868 3614 21870 3666
rect 21870 3614 21922 3666
rect 21922 3614 21924 3666
rect 21868 3612 21924 3614
rect 22204 3612 22260 3668
rect 20748 3554 20804 3556
rect 20748 3502 20750 3554
rect 20750 3502 20802 3554
rect 20802 3502 20804 3554
rect 20748 3500 20804 3502
rect 24780 6466 24836 6468
rect 24780 6414 24782 6466
rect 24782 6414 24834 6466
rect 24834 6414 24836 6466
rect 24780 6412 24836 6414
rect 25228 6300 25284 6356
rect 25788 7474 25844 7476
rect 25788 7422 25790 7474
rect 25790 7422 25842 7474
rect 25842 7422 25844 7474
rect 25788 7420 25844 7422
rect 25340 5964 25396 6020
rect 25452 6748 25508 6804
rect 25116 5852 25172 5908
rect 25676 6748 25732 6804
rect 24556 5292 24612 5348
rect 25452 5628 25508 5684
rect 25564 5516 25620 5572
rect 25340 5180 25396 5236
rect 25788 5292 25844 5348
rect 25564 5068 25620 5124
rect 24780 4396 24836 4452
rect 26572 7420 26628 7476
rect 27244 8092 27300 8148
rect 28028 8146 28084 8148
rect 28028 8094 28030 8146
rect 28030 8094 28082 8146
rect 28082 8094 28084 8146
rect 28028 8092 28084 8094
rect 26916 7866 26972 7868
rect 26916 7814 26918 7866
rect 26918 7814 26970 7866
rect 26970 7814 26972 7866
rect 26916 7812 26972 7814
rect 27020 7866 27076 7868
rect 27020 7814 27022 7866
rect 27022 7814 27074 7866
rect 27074 7814 27076 7866
rect 27020 7812 27076 7814
rect 27124 7866 27180 7868
rect 27124 7814 27126 7866
rect 27126 7814 27178 7866
rect 27178 7814 27180 7866
rect 27124 7812 27180 7814
rect 26460 6690 26516 6692
rect 26460 6638 26462 6690
rect 26462 6638 26514 6690
rect 26514 6638 26516 6690
rect 26460 6636 26516 6638
rect 26684 6524 26740 6580
rect 27020 6524 27076 6580
rect 26916 6298 26972 6300
rect 26916 6246 26918 6298
rect 26918 6246 26970 6298
rect 26970 6246 26972 6298
rect 26916 6244 26972 6246
rect 27020 6298 27076 6300
rect 27020 6246 27022 6298
rect 27022 6246 27074 6298
rect 27074 6246 27076 6298
rect 27020 6244 27076 6246
rect 27124 6298 27180 6300
rect 27124 6246 27126 6298
rect 27126 6246 27178 6298
rect 27178 6246 27180 6298
rect 27124 6244 27180 6246
rect 27580 7586 27636 7588
rect 27580 7534 27582 7586
rect 27582 7534 27634 7586
rect 27634 7534 27636 7586
rect 27580 7532 27636 7534
rect 27916 7980 27972 8036
rect 27580 6748 27636 6804
rect 27356 6524 27412 6580
rect 27356 5964 27412 6020
rect 26460 5906 26516 5908
rect 26460 5854 26462 5906
rect 26462 5854 26514 5906
rect 26514 5854 26516 5906
rect 26460 5852 26516 5854
rect 26012 5404 26068 5460
rect 26460 5068 26516 5124
rect 26916 4730 26972 4732
rect 26916 4678 26918 4730
rect 26918 4678 26970 4730
rect 26970 4678 26972 4730
rect 26916 4676 26972 4678
rect 27020 4730 27076 4732
rect 27020 4678 27022 4730
rect 27022 4678 27074 4730
rect 27074 4678 27076 4730
rect 27020 4676 27076 4678
rect 27124 4730 27180 4732
rect 27124 4678 27126 4730
rect 27126 4678 27178 4730
rect 27178 4678 27180 4730
rect 27124 4676 27180 4678
rect 26236 4508 26292 4564
rect 28140 7474 28196 7476
rect 28140 7422 28142 7474
rect 28142 7422 28194 7474
rect 28194 7422 28196 7474
rect 28140 7420 28196 7422
rect 28028 7196 28084 7252
rect 27916 7084 27972 7140
rect 28140 6748 28196 6804
rect 28588 9714 28644 9716
rect 28588 9662 28590 9714
rect 28590 9662 28642 9714
rect 28642 9662 28644 9714
rect 28588 9660 28644 9662
rect 28812 8988 28868 9044
rect 28364 8034 28420 8036
rect 28364 7982 28366 8034
rect 28366 7982 28418 8034
rect 28418 7982 28420 8034
rect 28364 7980 28420 7982
rect 28476 7474 28532 7476
rect 28476 7422 28478 7474
rect 28478 7422 28530 7474
rect 28530 7422 28532 7474
rect 28476 7420 28532 7422
rect 28588 7308 28644 7364
rect 28364 7084 28420 7140
rect 27356 5292 27412 5348
rect 28140 6412 28196 6468
rect 27916 6018 27972 6020
rect 27916 5966 27918 6018
rect 27918 5966 27970 6018
rect 27970 5966 27972 6018
rect 27916 5964 27972 5966
rect 27468 5628 27524 5684
rect 28028 5346 28084 5348
rect 28028 5294 28030 5346
rect 28030 5294 28082 5346
rect 28082 5294 28084 5346
rect 28028 5292 28084 5294
rect 27356 4898 27412 4900
rect 27356 4846 27358 4898
rect 27358 4846 27410 4898
rect 27410 4846 27412 4898
rect 27356 4844 27412 4846
rect 27244 4508 27300 4564
rect 28028 4508 28084 4564
rect 24668 4226 24724 4228
rect 24668 4174 24670 4226
rect 24670 4174 24722 4226
rect 24722 4174 24724 4226
rect 24668 4172 24724 4174
rect 24220 3724 24276 3780
rect 25340 4338 25396 4340
rect 25340 4286 25342 4338
rect 25342 4286 25394 4338
rect 25394 4286 25396 4338
rect 25340 4284 25396 4286
rect 27468 4172 27524 4228
rect 28140 4396 28196 4452
rect 28588 6860 28644 6916
rect 28588 6636 28644 6692
rect 29148 13692 29204 13748
rect 29036 13244 29092 13300
rect 29148 13132 29204 13188
rect 29036 12124 29092 12180
rect 29148 11676 29204 11732
rect 29820 17948 29876 18004
rect 29372 15820 29428 15876
rect 30044 18620 30100 18676
rect 30268 19292 30324 19348
rect 30156 18060 30212 18116
rect 31164 21586 31220 21588
rect 31164 21534 31166 21586
rect 31166 21534 31218 21586
rect 31218 21534 31220 21586
rect 31164 21532 31220 21534
rect 30492 19964 30548 20020
rect 30604 19292 30660 19348
rect 30716 19234 30772 19236
rect 30716 19182 30718 19234
rect 30718 19182 30770 19234
rect 30770 19182 30772 19234
rect 30716 19180 30772 19182
rect 30604 18562 30660 18564
rect 30604 18510 30606 18562
rect 30606 18510 30658 18562
rect 30658 18510 30660 18562
rect 30604 18508 30660 18510
rect 30940 21308 30996 21364
rect 31200 21194 31256 21196
rect 31200 21142 31202 21194
rect 31202 21142 31254 21194
rect 31254 21142 31256 21194
rect 31200 21140 31256 21142
rect 31304 21194 31360 21196
rect 31304 21142 31306 21194
rect 31306 21142 31358 21194
rect 31358 21142 31360 21194
rect 31304 21140 31360 21142
rect 31408 21194 31464 21196
rect 31408 21142 31410 21194
rect 31410 21142 31462 21194
rect 31462 21142 31464 21194
rect 31408 21140 31464 21142
rect 31948 23212 32004 23268
rect 32060 23100 32116 23156
rect 32060 22316 32116 22372
rect 32172 23884 32228 23940
rect 33404 31554 33460 31556
rect 33404 31502 33406 31554
rect 33406 31502 33458 31554
rect 33458 31502 33460 31554
rect 33404 31500 33460 31502
rect 35196 34524 35252 34580
rect 35196 33628 35252 33684
rect 34412 32732 34468 32788
rect 34076 31948 34132 32004
rect 33964 31106 34020 31108
rect 33964 31054 33966 31106
rect 33966 31054 34018 31106
rect 34018 31054 34020 31106
rect 33964 31052 34020 31054
rect 32956 30994 33012 30996
rect 32956 30942 32958 30994
rect 32958 30942 33010 30994
rect 33010 30942 33012 30994
rect 32956 30940 33012 30942
rect 33404 30994 33460 30996
rect 33404 30942 33406 30994
rect 33406 30942 33458 30994
rect 33458 30942 33460 30994
rect 33404 30940 33460 30942
rect 32956 30492 33012 30548
rect 34860 32674 34916 32676
rect 34860 32622 34862 32674
rect 34862 32622 34914 32674
rect 34914 32622 34916 32674
rect 34860 32620 34916 32622
rect 35980 33292 36036 33348
rect 35484 32954 35540 32956
rect 35484 32902 35486 32954
rect 35486 32902 35538 32954
rect 35538 32902 35540 32954
rect 35484 32900 35540 32902
rect 35588 32954 35644 32956
rect 35588 32902 35590 32954
rect 35590 32902 35642 32954
rect 35642 32902 35644 32954
rect 35588 32900 35644 32902
rect 35692 32954 35748 32956
rect 35692 32902 35694 32954
rect 35694 32902 35746 32954
rect 35746 32902 35748 32954
rect 35692 32900 35748 32902
rect 34300 30828 34356 30884
rect 34412 30268 34468 30324
rect 33180 29708 33236 29764
rect 33292 29202 33348 29204
rect 33292 29150 33294 29202
rect 33294 29150 33346 29202
rect 33346 29150 33348 29202
rect 33292 29148 33348 29150
rect 33068 28364 33124 28420
rect 33404 28364 33460 28420
rect 33180 28140 33236 28196
rect 32732 27132 32788 27188
rect 32844 26460 32900 26516
rect 33852 29596 33908 29652
rect 33852 29372 33908 29428
rect 33628 28252 33684 28308
rect 34188 29932 34244 29988
rect 34412 29650 34468 29652
rect 34412 29598 34414 29650
rect 34414 29598 34466 29650
rect 34466 29598 34468 29650
rect 34412 29596 34468 29598
rect 34300 29484 34356 29540
rect 34636 30994 34692 30996
rect 34636 30942 34638 30994
rect 34638 30942 34690 30994
rect 34690 30942 34692 30994
rect 34636 30940 34692 30942
rect 34748 30268 34804 30324
rect 34636 29986 34692 29988
rect 34636 29934 34638 29986
rect 34638 29934 34690 29986
rect 34690 29934 34692 29986
rect 34636 29932 34692 29934
rect 34860 29708 34916 29764
rect 34524 29372 34580 29428
rect 34076 28364 34132 28420
rect 35484 31386 35540 31388
rect 35484 31334 35486 31386
rect 35486 31334 35538 31386
rect 35538 31334 35540 31386
rect 35484 31332 35540 31334
rect 35588 31386 35644 31388
rect 35588 31334 35590 31386
rect 35590 31334 35642 31386
rect 35642 31334 35644 31386
rect 35588 31332 35644 31334
rect 35692 31386 35748 31388
rect 35692 31334 35694 31386
rect 35694 31334 35746 31386
rect 35746 31334 35748 31386
rect 35692 31332 35748 31334
rect 35084 30828 35140 30884
rect 35084 30492 35140 30548
rect 35484 29818 35540 29820
rect 35484 29766 35486 29818
rect 35486 29766 35538 29818
rect 35538 29766 35540 29818
rect 35484 29764 35540 29766
rect 35588 29818 35644 29820
rect 35588 29766 35590 29818
rect 35590 29766 35642 29818
rect 35642 29766 35644 29818
rect 35588 29764 35644 29766
rect 35692 29818 35748 29820
rect 35692 29766 35694 29818
rect 35694 29766 35746 29818
rect 35746 29766 35748 29818
rect 35692 29764 35748 29766
rect 35084 29426 35140 29428
rect 35084 29374 35086 29426
rect 35086 29374 35138 29426
rect 35138 29374 35140 29426
rect 35084 29372 35140 29374
rect 33180 26460 33236 26516
rect 33180 26236 33236 26292
rect 33068 25900 33124 25956
rect 32844 25394 32900 25396
rect 32844 25342 32846 25394
rect 32846 25342 32898 25394
rect 32898 25342 32900 25394
rect 32844 25340 32900 25342
rect 33180 25564 33236 25620
rect 33180 25228 33236 25284
rect 32732 23884 32788 23940
rect 32844 24780 32900 24836
rect 32284 23548 32340 23604
rect 32172 22146 32228 22148
rect 32172 22094 32174 22146
rect 32174 22094 32226 22146
rect 32226 22094 32228 22146
rect 32172 22092 32228 22094
rect 31836 21420 31892 21476
rect 32060 21698 32116 21700
rect 32060 21646 32062 21698
rect 32062 21646 32114 21698
rect 32114 21646 32116 21698
rect 32060 21644 32116 21646
rect 32172 21532 32228 21588
rect 32508 21362 32564 21364
rect 32508 21310 32510 21362
rect 32510 21310 32562 21362
rect 32562 21310 32564 21362
rect 32508 21308 32564 21310
rect 32396 21196 32452 21252
rect 32284 20748 32340 20804
rect 32956 24556 33012 24612
rect 33180 24722 33236 24724
rect 33180 24670 33182 24722
rect 33182 24670 33234 24722
rect 33234 24670 33236 24722
rect 33180 24668 33236 24670
rect 34636 28140 34692 28196
rect 33404 25618 33460 25620
rect 33404 25566 33406 25618
rect 33406 25566 33458 25618
rect 33458 25566 33460 25618
rect 33404 25564 33460 25566
rect 34076 26796 34132 26852
rect 34188 26684 34244 26740
rect 33964 26402 34020 26404
rect 33964 26350 33966 26402
rect 33966 26350 34018 26402
rect 34018 26350 34020 26402
rect 33964 26348 34020 26350
rect 33740 25900 33796 25956
rect 33628 25116 33684 25172
rect 33404 24610 33460 24612
rect 33404 24558 33406 24610
rect 33406 24558 33458 24610
rect 33458 24558 33460 24610
rect 33404 24556 33460 24558
rect 33180 23548 33236 23604
rect 33292 23266 33348 23268
rect 33292 23214 33294 23266
rect 33294 23214 33346 23266
rect 33346 23214 33348 23266
rect 33292 23212 33348 23214
rect 33068 22370 33124 22372
rect 33068 22318 33070 22370
rect 33070 22318 33122 22370
rect 33122 22318 33124 22370
rect 33068 22316 33124 22318
rect 32844 21084 32900 21140
rect 32396 20524 32452 20580
rect 31612 20130 31668 20132
rect 31612 20078 31614 20130
rect 31614 20078 31666 20130
rect 31666 20078 31668 20130
rect 31612 20076 31668 20078
rect 31836 20018 31892 20020
rect 31836 19966 31838 20018
rect 31838 19966 31890 20018
rect 31890 19966 31892 20018
rect 31836 19964 31892 19966
rect 31200 19626 31256 19628
rect 31200 19574 31202 19626
rect 31202 19574 31254 19626
rect 31254 19574 31256 19626
rect 31200 19572 31256 19574
rect 31304 19626 31360 19628
rect 31304 19574 31306 19626
rect 31306 19574 31358 19626
rect 31358 19574 31360 19626
rect 31304 19572 31360 19574
rect 31408 19626 31464 19628
rect 31408 19574 31410 19626
rect 31410 19574 31462 19626
rect 31462 19574 31464 19626
rect 31408 19572 31464 19574
rect 30380 17724 30436 17780
rect 31052 19068 31108 19124
rect 30156 17554 30212 17556
rect 30156 17502 30158 17554
rect 30158 17502 30210 17554
rect 30210 17502 30212 17554
rect 30156 17500 30212 17502
rect 29484 16380 29540 16436
rect 29372 14812 29428 14868
rect 30044 16268 30100 16324
rect 29932 14252 29988 14308
rect 29708 13580 29764 13636
rect 29708 13020 29764 13076
rect 30828 18172 30884 18228
rect 30940 17890 30996 17892
rect 30940 17838 30942 17890
rect 30942 17838 30994 17890
rect 30994 17838 30996 17890
rect 30940 17836 30996 17838
rect 30716 17164 30772 17220
rect 31500 18732 31556 18788
rect 32284 19794 32340 19796
rect 32284 19742 32286 19794
rect 32286 19742 32338 19794
rect 32338 19742 32340 19794
rect 32284 19740 32340 19742
rect 32284 19346 32340 19348
rect 32284 19294 32286 19346
rect 32286 19294 32338 19346
rect 32338 19294 32340 19346
rect 32284 19292 32340 19294
rect 33068 20130 33124 20132
rect 33068 20078 33070 20130
rect 33070 20078 33122 20130
rect 33122 20078 33124 20130
rect 33068 20076 33124 20078
rect 33292 21868 33348 21924
rect 31948 18508 32004 18564
rect 31836 18450 31892 18452
rect 31836 18398 31838 18450
rect 31838 18398 31890 18450
rect 31890 18398 31892 18450
rect 31836 18396 31892 18398
rect 31200 18058 31256 18060
rect 31200 18006 31202 18058
rect 31202 18006 31254 18058
rect 31254 18006 31256 18058
rect 31200 18004 31256 18006
rect 31304 18058 31360 18060
rect 31304 18006 31306 18058
rect 31306 18006 31358 18058
rect 31358 18006 31360 18058
rect 31304 18004 31360 18006
rect 31408 18058 31464 18060
rect 31408 18006 31410 18058
rect 31410 18006 31462 18058
rect 31462 18006 31464 18058
rect 31408 18004 31464 18006
rect 32508 17948 32564 18004
rect 32172 17836 32228 17892
rect 31276 17778 31332 17780
rect 31276 17726 31278 17778
rect 31278 17726 31330 17778
rect 31330 17726 31332 17778
rect 31276 17724 31332 17726
rect 31724 17388 31780 17444
rect 32620 17388 32676 17444
rect 30380 16492 30436 16548
rect 30716 16716 30772 16772
rect 30940 16770 30996 16772
rect 30940 16718 30942 16770
rect 30942 16718 30994 16770
rect 30994 16718 30996 16770
rect 30940 16716 30996 16718
rect 31200 16490 31256 16492
rect 31200 16438 31202 16490
rect 31202 16438 31254 16490
rect 31254 16438 31256 16490
rect 31200 16436 31256 16438
rect 31304 16490 31360 16492
rect 31304 16438 31306 16490
rect 31306 16438 31358 16490
rect 31358 16438 31360 16490
rect 31304 16436 31360 16438
rect 31408 16490 31464 16492
rect 31408 16438 31410 16490
rect 31410 16438 31462 16490
rect 31462 16438 31464 16490
rect 31408 16436 31464 16438
rect 30492 15036 30548 15092
rect 30156 14924 30212 14980
rect 30268 12962 30324 12964
rect 30268 12910 30270 12962
rect 30270 12910 30322 12962
rect 30322 12910 30324 12962
rect 30268 12908 30324 12910
rect 29932 12684 29988 12740
rect 29596 10668 29652 10724
rect 32396 16882 32452 16884
rect 32396 16830 32398 16882
rect 32398 16830 32450 16882
rect 32450 16830 32452 16882
rect 32396 16828 32452 16830
rect 32172 16604 32228 16660
rect 31724 15932 31780 15988
rect 31500 15036 31556 15092
rect 31200 14922 31256 14924
rect 31200 14870 31202 14922
rect 31202 14870 31254 14922
rect 31254 14870 31256 14922
rect 31200 14868 31256 14870
rect 31304 14922 31360 14924
rect 31304 14870 31306 14922
rect 31306 14870 31358 14922
rect 31358 14870 31360 14922
rect 31304 14868 31360 14870
rect 31408 14922 31464 14924
rect 31408 14870 31410 14922
rect 31410 14870 31462 14922
rect 31462 14870 31464 14922
rect 31408 14868 31464 14870
rect 30940 13580 30996 13636
rect 31052 14252 31108 14308
rect 30940 12738 30996 12740
rect 30940 12686 30942 12738
rect 30942 12686 30994 12738
rect 30994 12686 30996 12738
rect 30940 12684 30996 12686
rect 30380 12236 30436 12292
rect 33180 17836 33236 17892
rect 33740 24444 33796 24500
rect 33964 24498 34020 24500
rect 33964 24446 33966 24498
rect 33966 24446 34018 24498
rect 34018 24446 34020 24498
rect 33964 24444 34020 24446
rect 33852 24332 33908 24388
rect 33628 23042 33684 23044
rect 33628 22990 33630 23042
rect 33630 22990 33682 23042
rect 33682 22990 33684 23042
rect 33628 22988 33684 22990
rect 33628 21586 33684 21588
rect 33628 21534 33630 21586
rect 33630 21534 33682 21586
rect 33682 21534 33684 21586
rect 33628 21532 33684 21534
rect 34412 28028 34468 28084
rect 34748 28082 34804 28084
rect 34748 28030 34750 28082
rect 34750 28030 34802 28082
rect 34802 28030 34804 28082
rect 34748 28028 34804 28030
rect 34412 27804 34468 27860
rect 34412 26402 34468 26404
rect 34412 26350 34414 26402
rect 34414 26350 34466 26402
rect 34466 26350 34468 26402
rect 34412 26348 34468 26350
rect 34300 26290 34356 26292
rect 34300 26238 34302 26290
rect 34302 26238 34354 26290
rect 34354 26238 34356 26290
rect 34300 26236 34356 26238
rect 34188 25788 34244 25844
rect 34188 25282 34244 25284
rect 34188 25230 34190 25282
rect 34190 25230 34242 25282
rect 34242 25230 34244 25282
rect 34188 25228 34244 25230
rect 34188 24892 34244 24948
rect 34188 23324 34244 23380
rect 34300 22876 34356 22932
rect 34860 26684 34916 26740
rect 35484 28250 35540 28252
rect 35484 28198 35486 28250
rect 35486 28198 35538 28250
rect 35538 28198 35540 28250
rect 35484 28196 35540 28198
rect 35588 28250 35644 28252
rect 35588 28198 35590 28250
rect 35590 28198 35642 28250
rect 35642 28198 35644 28250
rect 35588 28196 35644 28198
rect 35692 28250 35748 28252
rect 35692 28198 35694 28250
rect 35694 28198 35746 28250
rect 35746 28198 35748 28250
rect 35692 28196 35748 28198
rect 35084 28028 35140 28084
rect 35084 27858 35140 27860
rect 35084 27806 35086 27858
rect 35086 27806 35138 27858
rect 35138 27806 35140 27858
rect 35084 27804 35140 27806
rect 34972 26460 35028 26516
rect 35084 26796 35140 26852
rect 34860 26402 34916 26404
rect 34860 26350 34862 26402
rect 34862 26350 34914 26402
rect 34914 26350 34916 26402
rect 34860 26348 34916 26350
rect 34860 25676 34916 25732
rect 35484 26682 35540 26684
rect 35484 26630 35486 26682
rect 35486 26630 35538 26682
rect 35538 26630 35540 26682
rect 35484 26628 35540 26630
rect 35588 26682 35644 26684
rect 35588 26630 35590 26682
rect 35590 26630 35642 26682
rect 35642 26630 35644 26682
rect 35588 26628 35644 26630
rect 35692 26682 35748 26684
rect 35692 26630 35694 26682
rect 35694 26630 35746 26682
rect 35746 26630 35748 26682
rect 35692 26628 35748 26630
rect 35196 26348 35252 26404
rect 35484 25114 35540 25116
rect 35484 25062 35486 25114
rect 35486 25062 35538 25114
rect 35538 25062 35540 25114
rect 35484 25060 35540 25062
rect 35588 25114 35644 25116
rect 35588 25062 35590 25114
rect 35590 25062 35642 25114
rect 35642 25062 35644 25114
rect 35588 25060 35644 25062
rect 35692 25114 35748 25116
rect 35692 25062 35694 25114
rect 35694 25062 35746 25114
rect 35746 25062 35748 25114
rect 35692 25060 35748 25062
rect 34860 24668 34916 24724
rect 34412 24556 34468 24612
rect 34636 24444 34692 24500
rect 34412 22428 34468 22484
rect 34300 22092 34356 22148
rect 34076 21644 34132 21700
rect 34412 21868 34468 21924
rect 33964 21474 34020 21476
rect 33964 21422 33966 21474
rect 33966 21422 34018 21474
rect 34018 21422 34020 21474
rect 33964 21420 34020 21422
rect 33516 18284 33572 18340
rect 33404 18060 33460 18116
rect 33404 17612 33460 17668
rect 33628 17500 33684 17556
rect 33516 17276 33572 17332
rect 32732 16098 32788 16100
rect 32732 16046 32734 16098
rect 32734 16046 32786 16098
rect 32786 16046 32788 16098
rect 32732 16044 32788 16046
rect 32620 15484 32676 15540
rect 32172 15092 32228 15148
rect 31836 14252 31892 14308
rect 31948 14812 32004 14868
rect 31612 13804 31668 13860
rect 31724 13468 31780 13524
rect 31200 13354 31256 13356
rect 31200 13302 31202 13354
rect 31202 13302 31254 13354
rect 31254 13302 31256 13354
rect 31200 13300 31256 13302
rect 31304 13354 31360 13356
rect 31304 13302 31306 13354
rect 31306 13302 31358 13354
rect 31358 13302 31360 13354
rect 31304 13300 31360 13302
rect 31408 13354 31464 13356
rect 31408 13302 31410 13354
rect 31410 13302 31462 13354
rect 31462 13302 31464 13354
rect 31408 13300 31464 13302
rect 31164 13132 31220 13188
rect 32396 14812 32452 14868
rect 32620 14812 32676 14868
rect 32732 15036 32788 15092
rect 32172 14700 32228 14756
rect 31948 13020 32004 13076
rect 32060 14476 32116 14532
rect 31836 12572 31892 12628
rect 32396 13468 32452 13524
rect 31724 11900 31780 11956
rect 29820 10444 29876 10500
rect 29932 9714 29988 9716
rect 29932 9662 29934 9714
rect 29934 9662 29986 9714
rect 29986 9662 29988 9714
rect 29932 9660 29988 9662
rect 29932 9436 29988 9492
rect 28924 7644 28980 7700
rect 29372 8764 29428 8820
rect 29484 8428 29540 8484
rect 31200 11786 31256 11788
rect 31200 11734 31202 11786
rect 31202 11734 31254 11786
rect 31254 11734 31256 11786
rect 31200 11732 31256 11734
rect 31304 11786 31360 11788
rect 31304 11734 31306 11786
rect 31306 11734 31358 11786
rect 31358 11734 31360 11786
rect 31304 11732 31360 11734
rect 31408 11786 31464 11788
rect 31408 11734 31410 11786
rect 31410 11734 31462 11786
rect 31462 11734 31464 11786
rect 31408 11732 31464 11734
rect 32508 11900 32564 11956
rect 32396 11564 32452 11620
rect 32732 11564 32788 11620
rect 31052 11452 31108 11508
rect 31276 11340 31332 11396
rect 32284 11340 32340 11396
rect 32620 10780 32676 10836
rect 30828 10722 30884 10724
rect 30828 10670 30830 10722
rect 30830 10670 30882 10722
rect 30882 10670 30884 10722
rect 30828 10668 30884 10670
rect 31836 10722 31892 10724
rect 31836 10670 31838 10722
rect 31838 10670 31890 10722
rect 31890 10670 31892 10722
rect 31836 10668 31892 10670
rect 30940 10498 30996 10500
rect 30940 10446 30942 10498
rect 30942 10446 30994 10498
rect 30994 10446 30996 10498
rect 30940 10444 30996 10446
rect 31200 10218 31256 10220
rect 31200 10166 31202 10218
rect 31202 10166 31254 10218
rect 31254 10166 31256 10218
rect 31200 10164 31256 10166
rect 31304 10218 31360 10220
rect 31304 10166 31306 10218
rect 31306 10166 31358 10218
rect 31358 10166 31360 10218
rect 31304 10164 31360 10166
rect 31408 10218 31464 10220
rect 31408 10166 31410 10218
rect 31410 10166 31462 10218
rect 31462 10166 31464 10218
rect 31408 10164 31464 10166
rect 30828 9660 30884 9716
rect 30716 9602 30772 9604
rect 30716 9550 30718 9602
rect 30718 9550 30770 9602
rect 30770 9550 30772 9602
rect 30716 9548 30772 9550
rect 30604 9436 30660 9492
rect 30044 8988 30100 9044
rect 30380 8988 30436 9044
rect 30716 9042 30772 9044
rect 30716 8990 30718 9042
rect 30718 8990 30770 9042
rect 30770 8990 30772 9042
rect 30716 8988 30772 8990
rect 31164 8764 31220 8820
rect 32396 9154 32452 9156
rect 32396 9102 32398 9154
rect 32398 9102 32450 9154
rect 32450 9102 32452 9154
rect 32396 9100 32452 9102
rect 31612 9042 31668 9044
rect 31612 8990 31614 9042
rect 31614 8990 31666 9042
rect 31666 8990 31668 9042
rect 31612 8988 31668 8990
rect 30044 8316 30100 8372
rect 29820 8258 29876 8260
rect 29820 8206 29822 8258
rect 29822 8206 29874 8258
rect 29874 8206 29876 8258
rect 29820 8204 29876 8206
rect 30716 8258 30772 8260
rect 30716 8206 30718 8258
rect 30718 8206 30770 8258
rect 30770 8206 30772 8258
rect 30716 8204 30772 8206
rect 29372 7698 29428 7700
rect 29372 7646 29374 7698
rect 29374 7646 29426 7698
rect 29426 7646 29428 7698
rect 29372 7644 29428 7646
rect 29932 7980 29988 8036
rect 30492 7868 30548 7924
rect 29260 7532 29316 7588
rect 29260 6860 29316 6916
rect 30044 7586 30100 7588
rect 30044 7534 30046 7586
rect 30046 7534 30098 7586
rect 30098 7534 30100 7586
rect 30044 7532 30100 7534
rect 29932 7474 29988 7476
rect 29932 7422 29934 7474
rect 29934 7422 29986 7474
rect 29986 7422 29988 7474
rect 29932 7420 29988 7422
rect 29484 6748 29540 6804
rect 29484 6466 29540 6468
rect 29484 6414 29486 6466
rect 29486 6414 29538 6466
rect 29538 6414 29540 6466
rect 29484 6412 29540 6414
rect 30940 8034 30996 8036
rect 30940 7982 30942 8034
rect 30942 7982 30994 8034
rect 30994 7982 30996 8034
rect 30940 7980 30996 7982
rect 31200 8650 31256 8652
rect 31200 8598 31202 8650
rect 31202 8598 31254 8650
rect 31254 8598 31256 8650
rect 31200 8596 31256 8598
rect 31304 8650 31360 8652
rect 31304 8598 31306 8650
rect 31306 8598 31358 8650
rect 31358 8598 31360 8650
rect 31304 8596 31360 8598
rect 31408 8650 31464 8652
rect 31408 8598 31410 8650
rect 31410 8598 31462 8650
rect 31462 8598 31464 8650
rect 31408 8596 31464 8598
rect 31276 8316 31332 8372
rect 31164 8092 31220 8148
rect 31612 7980 31668 8036
rect 32060 8146 32116 8148
rect 32060 8094 32062 8146
rect 32062 8094 32114 8146
rect 32114 8094 32116 8146
rect 32060 8092 32116 8094
rect 32060 7868 32116 7924
rect 32172 7644 32228 7700
rect 31836 7586 31892 7588
rect 31836 7534 31838 7586
rect 31838 7534 31890 7586
rect 31890 7534 31892 7586
rect 31836 7532 31892 7534
rect 31276 7474 31332 7476
rect 31276 7422 31278 7474
rect 31278 7422 31330 7474
rect 31330 7422 31332 7474
rect 31276 7420 31332 7422
rect 31200 7082 31256 7084
rect 31200 7030 31202 7082
rect 31202 7030 31254 7082
rect 31254 7030 31256 7082
rect 31200 7028 31256 7030
rect 31304 7082 31360 7084
rect 31304 7030 31306 7082
rect 31306 7030 31358 7082
rect 31358 7030 31360 7082
rect 31304 7028 31360 7030
rect 31408 7082 31464 7084
rect 31408 7030 31410 7082
rect 31410 7030 31462 7082
rect 31462 7030 31464 7082
rect 31408 7028 31464 7030
rect 31164 6690 31220 6692
rect 31164 6638 31166 6690
rect 31166 6638 31218 6690
rect 31218 6638 31220 6690
rect 31164 6636 31220 6638
rect 31052 5740 31108 5796
rect 31724 5740 31780 5796
rect 31200 5514 31256 5516
rect 31200 5462 31202 5514
rect 31202 5462 31254 5514
rect 31254 5462 31256 5514
rect 31200 5460 31256 5462
rect 31304 5514 31360 5516
rect 31304 5462 31306 5514
rect 31306 5462 31358 5514
rect 31358 5462 31360 5514
rect 31304 5460 31360 5462
rect 31408 5514 31464 5516
rect 31408 5462 31410 5514
rect 31410 5462 31462 5514
rect 31462 5462 31464 5514
rect 31408 5460 31464 5462
rect 29036 4956 29092 5012
rect 28924 4396 28980 4452
rect 27244 3836 27300 3892
rect 25564 3666 25620 3668
rect 25564 3614 25566 3666
rect 25566 3614 25618 3666
rect 25618 3614 25620 3666
rect 25564 3612 25620 3614
rect 25340 3388 25396 3444
rect 26916 3162 26972 3164
rect 26916 3110 26918 3162
rect 26918 3110 26970 3162
rect 26970 3110 26972 3162
rect 26916 3108 26972 3110
rect 27020 3162 27076 3164
rect 27020 3110 27022 3162
rect 27022 3110 27074 3162
rect 27074 3110 27076 3162
rect 27020 3108 27076 3110
rect 27124 3162 27180 3164
rect 27124 3110 27126 3162
rect 27126 3110 27178 3162
rect 27178 3110 27180 3162
rect 27124 3108 27180 3110
rect 28700 3836 28756 3892
rect 28364 3724 28420 3780
rect 27804 3442 27860 3444
rect 27804 3390 27806 3442
rect 27806 3390 27858 3442
rect 27858 3390 27860 3442
rect 27804 3388 27860 3390
rect 28476 3500 28532 3556
rect 29036 4284 29092 4340
rect 31276 4956 31332 5012
rect 29372 4172 29428 4228
rect 30604 4844 30660 4900
rect 32396 8818 32452 8820
rect 32396 8766 32398 8818
rect 32398 8766 32450 8818
rect 32450 8766 32452 8818
rect 32396 8764 32452 8766
rect 32284 6748 32340 6804
rect 29820 3836 29876 3892
rect 30268 4172 30324 4228
rect 29372 3554 29428 3556
rect 29372 3502 29374 3554
rect 29374 3502 29426 3554
rect 29426 3502 29428 3554
rect 29372 3500 29428 3502
rect 29820 3442 29876 3444
rect 29820 3390 29822 3442
rect 29822 3390 29874 3442
rect 29874 3390 29876 3442
rect 29820 3388 29876 3390
rect 30044 3388 30100 3444
rect 31200 3946 31256 3948
rect 31200 3894 31202 3946
rect 31202 3894 31254 3946
rect 31254 3894 31256 3946
rect 31200 3892 31256 3894
rect 31304 3946 31360 3948
rect 31304 3894 31306 3946
rect 31306 3894 31358 3946
rect 31358 3894 31360 3946
rect 31304 3892 31360 3894
rect 31408 3946 31464 3948
rect 31408 3894 31410 3946
rect 31410 3894 31462 3946
rect 31462 3894 31464 3946
rect 31408 3892 31464 3894
rect 31052 3554 31108 3556
rect 31052 3502 31054 3554
rect 31054 3502 31106 3554
rect 31106 3502 31108 3554
rect 31052 3500 31108 3502
rect 31612 3500 31668 3556
rect 30604 3442 30660 3444
rect 30604 3390 30606 3442
rect 30606 3390 30658 3442
rect 30658 3390 30660 3442
rect 30604 3388 30660 3390
rect 31500 3442 31556 3444
rect 31500 3390 31502 3442
rect 31502 3390 31554 3442
rect 31554 3390 31556 3442
rect 31500 3388 31556 3390
rect 32396 3554 32452 3556
rect 32396 3502 32398 3554
rect 32398 3502 32450 3554
rect 32450 3502 32452 3554
rect 32396 3500 32452 3502
rect 32284 3276 32340 3332
rect 33292 15986 33348 15988
rect 33292 15934 33294 15986
rect 33294 15934 33346 15986
rect 33346 15934 33348 15986
rect 33292 15932 33348 15934
rect 34076 21308 34132 21364
rect 33852 19740 33908 19796
rect 33852 18956 33908 19012
rect 35196 23042 35252 23044
rect 35196 22990 35198 23042
rect 35198 22990 35250 23042
rect 35250 22990 35252 23042
rect 35196 22988 35252 22990
rect 35484 23546 35540 23548
rect 35484 23494 35486 23546
rect 35486 23494 35538 23546
rect 35538 23494 35540 23546
rect 35484 23492 35540 23494
rect 35588 23546 35644 23548
rect 35588 23494 35590 23546
rect 35590 23494 35642 23546
rect 35642 23494 35644 23546
rect 35588 23492 35644 23494
rect 35692 23546 35748 23548
rect 35692 23494 35694 23546
rect 35694 23494 35746 23546
rect 35746 23494 35748 23546
rect 35692 23492 35748 23494
rect 34748 22540 34804 22596
rect 34972 22594 35028 22596
rect 34972 22542 34974 22594
rect 34974 22542 35026 22594
rect 35026 22542 35028 22594
rect 34972 22540 35028 22542
rect 34860 22428 34916 22484
rect 35484 21978 35540 21980
rect 35484 21926 35486 21978
rect 35486 21926 35538 21978
rect 35538 21926 35540 21978
rect 35484 21924 35540 21926
rect 35588 21978 35644 21980
rect 35588 21926 35590 21978
rect 35590 21926 35642 21978
rect 35642 21926 35644 21978
rect 35588 21924 35644 21926
rect 35692 21978 35748 21980
rect 35692 21926 35694 21978
rect 35694 21926 35746 21978
rect 35746 21926 35748 21978
rect 35692 21924 35748 21926
rect 35196 21756 35252 21812
rect 35084 21532 35140 21588
rect 34748 21026 34804 21028
rect 34748 20974 34750 21026
rect 34750 20974 34802 21026
rect 34802 20974 34804 21026
rect 34748 20972 34804 20974
rect 34412 20076 34468 20132
rect 34300 19458 34356 19460
rect 34300 19406 34302 19458
rect 34302 19406 34354 19458
rect 34354 19406 34356 19458
rect 34300 19404 34356 19406
rect 34636 19404 34692 19460
rect 34076 18450 34132 18452
rect 34076 18398 34078 18450
rect 34078 18398 34130 18450
rect 34130 18398 34132 18450
rect 34076 18396 34132 18398
rect 34076 18060 34132 18116
rect 33964 17276 34020 17332
rect 33180 15426 33236 15428
rect 33180 15374 33182 15426
rect 33182 15374 33234 15426
rect 33234 15374 33236 15426
rect 33180 15372 33236 15374
rect 33516 15090 33572 15092
rect 33516 15038 33518 15090
rect 33518 15038 33570 15090
rect 33570 15038 33572 15090
rect 33516 15036 33572 15038
rect 33180 14364 33236 14420
rect 33516 13522 33572 13524
rect 33516 13470 33518 13522
rect 33518 13470 33570 13522
rect 33570 13470 33572 13522
rect 33516 13468 33572 13470
rect 33180 12402 33236 12404
rect 33180 12350 33182 12402
rect 33182 12350 33234 12402
rect 33234 12350 33236 12402
rect 33180 12348 33236 12350
rect 33852 16604 33908 16660
rect 33852 15820 33908 15876
rect 33964 15932 34020 15988
rect 34412 17554 34468 17556
rect 34412 17502 34414 17554
rect 34414 17502 34466 17554
rect 34466 17502 34468 17554
rect 34412 17500 34468 17502
rect 34860 18172 34916 18228
rect 34636 18060 34692 18116
rect 35084 18956 35140 19012
rect 34188 16716 34244 16772
rect 33740 15708 33796 15764
rect 33740 13468 33796 13524
rect 33964 13020 34020 13076
rect 33628 12124 33684 12180
rect 33516 11954 33572 11956
rect 33516 11902 33518 11954
rect 33518 11902 33570 11954
rect 33570 11902 33572 11954
rect 33516 11900 33572 11902
rect 32956 11506 33012 11508
rect 32956 11454 32958 11506
rect 32958 11454 33010 11506
rect 33010 11454 33012 11506
rect 32956 11452 33012 11454
rect 33516 11676 33572 11732
rect 33516 11506 33572 11508
rect 33516 11454 33518 11506
rect 33518 11454 33570 11506
rect 33570 11454 33572 11506
rect 33516 11452 33572 11454
rect 34188 12796 34244 12852
rect 34076 12290 34132 12292
rect 34076 12238 34078 12290
rect 34078 12238 34130 12290
rect 34130 12238 34132 12290
rect 34076 12236 34132 12238
rect 33180 10332 33236 10388
rect 34076 11676 34132 11732
rect 34188 11452 34244 11508
rect 34636 15820 34692 15876
rect 34748 15538 34804 15540
rect 34748 15486 34750 15538
rect 34750 15486 34802 15538
rect 34802 15486 34804 15538
rect 34748 15484 34804 15486
rect 34748 13858 34804 13860
rect 34748 13806 34750 13858
rect 34750 13806 34802 13858
rect 34802 13806 34804 13858
rect 34748 13804 34804 13806
rect 34412 12850 34468 12852
rect 34412 12798 34414 12850
rect 34414 12798 34466 12850
rect 34466 12798 34468 12850
rect 34412 12796 34468 12798
rect 34412 11452 34468 11508
rect 34188 10332 34244 10388
rect 34412 10556 34468 10612
rect 35084 17276 35140 17332
rect 35484 20410 35540 20412
rect 35484 20358 35486 20410
rect 35486 20358 35538 20410
rect 35538 20358 35540 20410
rect 35484 20356 35540 20358
rect 35588 20410 35644 20412
rect 35588 20358 35590 20410
rect 35590 20358 35642 20410
rect 35642 20358 35644 20410
rect 35588 20356 35644 20358
rect 35692 20410 35748 20412
rect 35692 20358 35694 20410
rect 35694 20358 35746 20410
rect 35746 20358 35748 20410
rect 35692 20356 35748 20358
rect 35484 18842 35540 18844
rect 35484 18790 35486 18842
rect 35486 18790 35538 18842
rect 35538 18790 35540 18842
rect 35484 18788 35540 18790
rect 35588 18842 35644 18844
rect 35588 18790 35590 18842
rect 35590 18790 35642 18842
rect 35642 18790 35644 18842
rect 35588 18788 35644 18790
rect 35692 18842 35748 18844
rect 35692 18790 35694 18842
rect 35694 18790 35746 18842
rect 35746 18790 35748 18842
rect 35692 18788 35748 18790
rect 35308 18396 35364 18452
rect 35196 16098 35252 16100
rect 35196 16046 35198 16098
rect 35198 16046 35250 16098
rect 35250 16046 35252 16098
rect 35196 16044 35252 16046
rect 35084 15986 35140 15988
rect 35084 15934 35086 15986
rect 35086 15934 35138 15986
rect 35138 15934 35140 15986
rect 35084 15932 35140 15934
rect 35484 17274 35540 17276
rect 35484 17222 35486 17274
rect 35486 17222 35538 17274
rect 35538 17222 35540 17274
rect 35484 17220 35540 17222
rect 35588 17274 35644 17276
rect 35588 17222 35590 17274
rect 35590 17222 35642 17274
rect 35642 17222 35644 17274
rect 35588 17220 35644 17222
rect 35692 17274 35748 17276
rect 35692 17222 35694 17274
rect 35694 17222 35746 17274
rect 35746 17222 35748 17274
rect 35692 17220 35748 17222
rect 36204 31612 36260 31668
rect 36204 22540 36260 22596
rect 35980 20972 36036 21028
rect 35868 16044 35924 16100
rect 35084 15538 35140 15540
rect 35084 15486 35086 15538
rect 35086 15486 35138 15538
rect 35138 15486 35140 15538
rect 35084 15484 35140 15486
rect 35084 13468 35140 13524
rect 34636 11676 34692 11732
rect 34636 11506 34692 11508
rect 34636 11454 34638 11506
rect 34638 11454 34690 11506
rect 34690 11454 34692 11506
rect 34636 11452 34692 11454
rect 35484 15706 35540 15708
rect 35484 15654 35486 15706
rect 35486 15654 35538 15706
rect 35538 15654 35540 15706
rect 35484 15652 35540 15654
rect 35588 15706 35644 15708
rect 35588 15654 35590 15706
rect 35590 15654 35642 15706
rect 35642 15654 35644 15706
rect 35588 15652 35644 15654
rect 35692 15706 35748 15708
rect 35692 15654 35694 15706
rect 35694 15654 35746 15706
rect 35746 15654 35748 15706
rect 35692 15652 35748 15654
rect 34860 12124 34916 12180
rect 33964 9772 34020 9828
rect 34412 9436 34468 9492
rect 33852 9100 33908 9156
rect 34188 8204 34244 8260
rect 35308 15484 35364 15540
rect 35084 11394 35140 11396
rect 35084 11342 35086 11394
rect 35086 11342 35138 11394
rect 35138 11342 35140 11394
rect 35084 11340 35140 11342
rect 35196 10668 35252 10724
rect 35084 10610 35140 10612
rect 35084 10558 35086 10610
rect 35086 10558 35138 10610
rect 35138 10558 35140 10610
rect 35084 10556 35140 10558
rect 34860 9436 34916 9492
rect 35484 14138 35540 14140
rect 35484 14086 35486 14138
rect 35486 14086 35538 14138
rect 35538 14086 35540 14138
rect 35484 14084 35540 14086
rect 35588 14138 35644 14140
rect 35588 14086 35590 14138
rect 35590 14086 35642 14138
rect 35642 14086 35644 14138
rect 35588 14084 35644 14086
rect 35692 14138 35748 14140
rect 35692 14086 35694 14138
rect 35694 14086 35746 14138
rect 35746 14086 35748 14138
rect 35692 14084 35748 14086
rect 35484 12570 35540 12572
rect 35484 12518 35486 12570
rect 35486 12518 35538 12570
rect 35538 12518 35540 12570
rect 35484 12516 35540 12518
rect 35588 12570 35644 12572
rect 35588 12518 35590 12570
rect 35590 12518 35642 12570
rect 35642 12518 35644 12570
rect 35588 12516 35644 12518
rect 35692 12570 35748 12572
rect 35692 12518 35694 12570
rect 35694 12518 35746 12570
rect 35746 12518 35748 12570
rect 35692 12516 35748 12518
rect 35484 11002 35540 11004
rect 35484 10950 35486 11002
rect 35486 10950 35538 11002
rect 35538 10950 35540 11002
rect 35484 10948 35540 10950
rect 35588 11002 35644 11004
rect 35588 10950 35590 11002
rect 35590 10950 35642 11002
rect 35642 10950 35644 11002
rect 35588 10948 35644 10950
rect 35692 11002 35748 11004
rect 35692 10950 35694 11002
rect 35694 10950 35746 11002
rect 35746 10950 35748 11002
rect 35692 10948 35748 10950
rect 35196 9826 35252 9828
rect 35196 9774 35198 9826
rect 35198 9774 35250 9826
rect 35250 9774 35252 9826
rect 35196 9772 35252 9774
rect 35484 9434 35540 9436
rect 35484 9382 35486 9434
rect 35486 9382 35538 9434
rect 35538 9382 35540 9434
rect 35484 9380 35540 9382
rect 35588 9434 35644 9436
rect 35588 9382 35590 9434
rect 35590 9382 35642 9434
rect 35642 9382 35644 9434
rect 35588 9380 35644 9382
rect 35692 9434 35748 9436
rect 35692 9382 35694 9434
rect 35694 9382 35746 9434
rect 35746 9382 35748 9434
rect 35692 9380 35748 9382
rect 34972 8428 35028 8484
rect 34636 5122 34692 5124
rect 34636 5070 34638 5122
rect 34638 5070 34690 5122
rect 34690 5070 34692 5122
rect 34636 5068 34692 5070
rect 35484 7866 35540 7868
rect 35484 7814 35486 7866
rect 35486 7814 35538 7866
rect 35538 7814 35540 7866
rect 35484 7812 35540 7814
rect 35588 7866 35644 7868
rect 35588 7814 35590 7866
rect 35590 7814 35642 7866
rect 35642 7814 35644 7866
rect 35588 7812 35644 7814
rect 35692 7866 35748 7868
rect 35692 7814 35694 7866
rect 35694 7814 35746 7866
rect 35746 7814 35748 7866
rect 35692 7812 35748 7814
rect 35308 7698 35364 7700
rect 35308 7646 35310 7698
rect 35310 7646 35362 7698
rect 35362 7646 35364 7698
rect 35308 7644 35364 7646
rect 35484 6298 35540 6300
rect 35484 6246 35486 6298
rect 35486 6246 35538 6298
rect 35538 6246 35540 6298
rect 35484 6244 35540 6246
rect 35588 6298 35644 6300
rect 35588 6246 35590 6298
rect 35590 6246 35642 6298
rect 35642 6246 35644 6298
rect 35588 6244 35644 6246
rect 35692 6298 35748 6300
rect 35692 6246 35694 6298
rect 35694 6246 35746 6298
rect 35746 6246 35748 6298
rect 35692 6244 35748 6246
rect 35196 5122 35252 5124
rect 35196 5070 35198 5122
rect 35198 5070 35250 5122
rect 35250 5070 35252 5122
rect 35196 5068 35252 5070
rect 35484 4730 35540 4732
rect 35484 4678 35486 4730
rect 35486 4678 35538 4730
rect 35538 4678 35540 4730
rect 35484 4676 35540 4678
rect 35588 4730 35644 4732
rect 35588 4678 35590 4730
rect 35590 4678 35642 4730
rect 35642 4678 35644 4730
rect 35588 4676 35644 4678
rect 35692 4730 35748 4732
rect 35692 4678 35694 4730
rect 35694 4678 35746 4730
rect 35746 4678 35748 4730
rect 35692 4676 35748 4678
rect 32956 3554 33012 3556
rect 32956 3502 32958 3554
rect 32958 3502 33010 3554
rect 33010 3502 33012 3554
rect 32956 3500 33012 3502
rect 32620 2268 32676 2324
rect 33404 3330 33460 3332
rect 33404 3278 33406 3330
rect 33406 3278 33458 3330
rect 33458 3278 33460 3330
rect 33404 3276 33460 3278
rect 35484 3162 35540 3164
rect 35484 3110 35486 3162
rect 35486 3110 35538 3162
rect 35538 3110 35540 3162
rect 35484 3108 35540 3110
rect 35588 3162 35644 3164
rect 35588 3110 35590 3162
rect 35590 3110 35642 3162
rect 35642 3110 35644 3162
rect 35588 3108 35644 3110
rect 35692 3162 35748 3164
rect 35692 3110 35694 3162
rect 35694 3110 35746 3162
rect 35746 3110 35748 3162
rect 35692 3108 35748 3110
<< metal3 >>
rect 36200 34580 37000 34608
rect 35186 34524 35196 34580
rect 35252 34524 37000 34580
rect 36200 34496 37000 34524
rect 5486 33684 5496 33740
rect 5552 33684 5600 33740
rect 5656 33684 5704 33740
rect 5760 33684 5770 33740
rect 14054 33684 14064 33740
rect 14120 33684 14168 33740
rect 14224 33684 14272 33740
rect 14328 33684 14338 33740
rect 22622 33684 22632 33740
rect 22688 33684 22736 33740
rect 22792 33684 22840 33740
rect 22896 33684 22906 33740
rect 31190 33684 31200 33740
rect 31256 33684 31304 33740
rect 31360 33684 31408 33740
rect 31464 33684 31474 33740
rect 33730 33628 33740 33684
rect 33796 33628 35196 33684
rect 35252 33628 35262 33684
rect 8194 33516 8204 33572
rect 8260 33516 10556 33572
rect 10612 33516 10622 33572
rect 12338 33516 12348 33572
rect 12404 33516 13916 33572
rect 13972 33516 13982 33572
rect 20626 33516 20636 33572
rect 20692 33516 25564 33572
rect 25620 33516 25630 33572
rect 16034 33404 16044 33460
rect 16100 33404 25228 33460
rect 25284 33404 25294 33460
rect 30146 33404 30156 33460
rect 30212 33404 32956 33460
rect 33012 33404 33022 33460
rect 8978 33292 8988 33348
rect 9044 33292 9996 33348
rect 10052 33292 10062 33348
rect 27346 33292 27356 33348
rect 27412 33292 35980 33348
rect 36036 33292 36046 33348
rect 9770 32900 9780 32956
rect 9836 32900 9884 32956
rect 9940 32900 9988 32956
rect 10044 32900 10054 32956
rect 18338 32900 18348 32956
rect 18404 32900 18452 32956
rect 18508 32900 18556 32956
rect 18612 32900 18622 32956
rect 26906 32900 26916 32956
rect 26972 32900 27020 32956
rect 27076 32900 27124 32956
rect 27180 32900 27190 32956
rect 35474 32900 35484 32956
rect 35540 32900 35588 32956
rect 35644 32900 35692 32956
rect 35748 32900 35758 32956
rect 28466 32844 28476 32900
rect 28532 32844 30380 32900
rect 30436 32844 30446 32900
rect 8306 32732 8316 32788
rect 8372 32732 9548 32788
rect 9604 32732 9614 32788
rect 15810 32732 15820 32788
rect 15876 32732 19852 32788
rect 19908 32732 19918 32788
rect 28578 32732 28588 32788
rect 28644 32732 34412 32788
rect 34468 32732 34478 32788
rect 16818 32620 16828 32676
rect 16884 32620 18284 32676
rect 18340 32620 18350 32676
rect 32274 32620 32284 32676
rect 32340 32620 34860 32676
rect 34916 32620 34926 32676
rect 17490 32508 17500 32564
rect 17556 32508 20524 32564
rect 20580 32508 20972 32564
rect 21028 32508 23324 32564
rect 23380 32508 23884 32564
rect 23940 32508 23950 32564
rect 27794 32508 27804 32564
rect 27860 32508 31836 32564
rect 31892 32508 31902 32564
rect 6850 32396 6860 32452
rect 6916 32396 7868 32452
rect 7924 32396 7934 32452
rect 15362 32396 15372 32452
rect 15428 32396 16268 32452
rect 16324 32396 17612 32452
rect 17668 32396 17678 32452
rect 21746 32396 21756 32452
rect 21812 32396 26236 32452
rect 26292 32396 26302 32452
rect 28018 32396 28028 32452
rect 28084 32396 29148 32452
rect 29204 32396 29214 32452
rect 22418 32284 22428 32340
rect 22484 32284 23436 32340
rect 23492 32284 23502 32340
rect 28242 32284 28252 32340
rect 28308 32284 31724 32340
rect 31780 32284 31790 32340
rect 26674 32172 26684 32228
rect 26740 32172 31052 32228
rect 31108 32172 31118 32228
rect 5486 32116 5496 32172
rect 5552 32116 5600 32172
rect 5656 32116 5704 32172
rect 5760 32116 5770 32172
rect 14054 32116 14064 32172
rect 14120 32116 14168 32172
rect 14224 32116 14272 32172
rect 14328 32116 14338 32172
rect 22622 32116 22632 32172
rect 22688 32116 22736 32172
rect 22792 32116 22840 32172
rect 22896 32116 22906 32172
rect 31190 32116 31200 32172
rect 31256 32116 31304 32172
rect 31360 32116 31408 32172
rect 31464 32116 31474 32172
rect 22530 31948 22540 32004
rect 22596 31948 23772 32004
rect 23828 31948 23838 32004
rect 32722 31948 32732 32004
rect 32788 31948 34076 32004
rect 34132 31948 34142 32004
rect 36200 31892 37000 31920
rect 6290 31836 6300 31892
rect 6356 31836 6524 31892
rect 6580 31836 8652 31892
rect 8708 31836 10220 31892
rect 10276 31836 11900 31892
rect 11956 31836 11966 31892
rect 17378 31836 17388 31892
rect 17444 31836 20412 31892
rect 20468 31836 24780 31892
rect 24836 31836 24846 31892
rect 28466 31836 28476 31892
rect 28532 31836 29260 31892
rect 29316 31836 29708 31892
rect 29764 31836 32172 31892
rect 32228 31836 32238 31892
rect 35980 31836 37000 31892
rect 8082 31724 8092 31780
rect 8148 31724 14588 31780
rect 14644 31724 14654 31780
rect 17714 31724 17724 31780
rect 17780 31724 18844 31780
rect 18900 31724 18910 31780
rect 21186 31724 21196 31780
rect 21252 31724 21756 31780
rect 21812 31724 21822 31780
rect 26898 31724 26908 31780
rect 26964 31724 32284 31780
rect 32340 31724 32350 31780
rect 35980 31668 36036 31836
rect 36200 31808 37000 31836
rect 8194 31612 8204 31668
rect 8260 31612 9212 31668
rect 9268 31612 9278 31668
rect 20066 31612 20076 31668
rect 20132 31612 21420 31668
rect 21476 31612 23548 31668
rect 23604 31612 23614 31668
rect 28242 31612 28252 31668
rect 28308 31612 31388 31668
rect 31444 31612 31454 31668
rect 35980 31612 36204 31668
rect 36260 31612 36270 31668
rect 12114 31500 12124 31556
rect 12180 31500 12460 31556
rect 12516 31500 13244 31556
rect 13300 31500 13804 31556
rect 13860 31500 13870 31556
rect 20626 31500 20636 31556
rect 20692 31500 22988 31556
rect 23044 31500 25340 31556
rect 25396 31500 25406 31556
rect 26450 31500 26460 31556
rect 26516 31500 33404 31556
rect 33460 31500 33470 31556
rect 22082 31388 22092 31444
rect 22148 31388 26348 31444
rect 26404 31388 26414 31444
rect 9770 31332 9780 31388
rect 9836 31332 9884 31388
rect 9940 31332 9988 31388
rect 10044 31332 10054 31388
rect 18338 31332 18348 31388
rect 18404 31332 18452 31388
rect 18508 31332 18556 31388
rect 18612 31332 18622 31388
rect 26906 31332 26916 31388
rect 26972 31332 27020 31388
rect 27076 31332 27124 31388
rect 27180 31332 27190 31388
rect 35474 31332 35484 31388
rect 35540 31332 35588 31388
rect 35644 31332 35692 31388
rect 35748 31332 35758 31388
rect 16146 31276 16156 31332
rect 16212 31276 17500 31332
rect 17556 31276 17566 31332
rect 22642 31276 22652 31332
rect 22708 31276 23212 31332
rect 23268 31276 23278 31332
rect 15362 31164 15372 31220
rect 15428 31164 15708 31220
rect 15764 31164 17948 31220
rect 18004 31164 18014 31220
rect 19506 31164 19516 31220
rect 19572 31164 20748 31220
rect 20804 31164 20814 31220
rect 28018 31164 28028 31220
rect 28084 31164 29260 31220
rect 29316 31164 30828 31220
rect 30884 31164 30894 31220
rect 15820 31052 16324 31108
rect 16706 31052 16716 31108
rect 16772 31052 17388 31108
rect 17444 31052 17454 31108
rect 17602 31052 17612 31108
rect 17668 31052 18732 31108
rect 18788 31052 18798 31108
rect 19058 31052 19068 31108
rect 19124 31052 25452 31108
rect 25508 31052 25518 31108
rect 27458 31052 27468 31108
rect 27524 31052 28476 31108
rect 28532 31052 28542 31108
rect 30604 31052 31724 31108
rect 31780 31052 31790 31108
rect 33058 31052 33068 31108
rect 33124 31052 33964 31108
rect 34020 31052 34030 31108
rect 7298 30940 7308 30996
rect 7364 30940 7980 30996
rect 8036 30940 10444 30996
rect 10500 30940 10510 30996
rect 11554 30940 11564 30996
rect 11620 30940 14588 30996
rect 14644 30940 15596 30996
rect 15652 30940 15662 30996
rect 15820 30884 15876 31052
rect 16268 30996 16324 31052
rect 30604 30996 30660 31052
rect 16034 30940 16044 30996
rect 16100 30940 16110 30996
rect 16258 30940 16268 30996
rect 16324 30940 17500 30996
rect 17556 30940 17566 30996
rect 18386 30940 18396 30996
rect 18452 30940 19404 30996
rect 19460 30940 20188 30996
rect 20244 30940 20254 30996
rect 21522 30940 21532 30996
rect 21588 30940 22764 30996
rect 22820 30940 23436 30996
rect 23492 30940 23502 30996
rect 29138 30940 29148 30996
rect 29204 30940 30604 30996
rect 30660 30940 30670 30996
rect 31042 30940 31052 30996
rect 31108 30940 32060 30996
rect 32116 30940 32126 30996
rect 32386 30940 32396 30996
rect 32452 30940 32956 30996
rect 33012 30940 33022 30996
rect 33394 30940 33404 30996
rect 33460 30940 34636 30996
rect 34692 30940 34702 30996
rect 14914 30828 14924 30884
rect 14980 30828 15876 30884
rect 16044 30772 16100 30940
rect 32396 30884 32452 30940
rect 20514 30828 20524 30884
rect 20580 30828 23548 30884
rect 23604 30828 23614 30884
rect 24210 30828 24220 30884
rect 24276 30828 25900 30884
rect 25956 30828 27692 30884
rect 27748 30828 27758 30884
rect 29922 30828 29932 30884
rect 29988 30828 30828 30884
rect 30884 30828 30894 30884
rect 31378 30828 31388 30884
rect 31444 30828 32452 30884
rect 34290 30828 34300 30884
rect 34356 30828 35084 30884
rect 35140 30828 35150 30884
rect 11218 30716 11228 30772
rect 11284 30716 16100 30772
rect 23548 30772 23604 30828
rect 23548 30716 25340 30772
rect 25396 30716 25406 30772
rect 30370 30716 30380 30772
rect 30436 30716 32396 30772
rect 32452 30716 32462 30772
rect 24658 30604 24668 30660
rect 24724 30604 26236 30660
rect 26292 30604 26302 30660
rect 5486 30548 5496 30604
rect 5552 30548 5600 30604
rect 5656 30548 5704 30604
rect 5760 30548 5770 30604
rect 14054 30548 14064 30604
rect 14120 30548 14168 30604
rect 14224 30548 14272 30604
rect 14328 30548 14338 30604
rect 22622 30548 22632 30604
rect 22688 30548 22736 30604
rect 22792 30548 22840 30604
rect 22896 30548 22906 30604
rect 31190 30548 31200 30604
rect 31256 30548 31304 30604
rect 31360 30548 31408 30604
rect 31464 30548 31474 30604
rect 32946 30492 32956 30548
rect 33012 30492 35084 30548
rect 35140 30492 35150 30548
rect 12562 30380 12572 30436
rect 12628 30380 14028 30436
rect 14084 30380 14094 30436
rect 15092 30380 17724 30436
rect 17780 30380 17790 30436
rect 15092 30324 15148 30380
rect 7532 30268 8932 30324
rect 9510 30268 9548 30324
rect 9604 30268 9614 30324
rect 12684 30268 15148 30324
rect 19394 30268 19404 30324
rect 19460 30268 20412 30324
rect 20468 30268 20478 30324
rect 21532 30268 21868 30324
rect 21924 30268 21934 30324
rect 25330 30268 25340 30324
rect 25396 30268 27804 30324
rect 27860 30268 27870 30324
rect 32498 30268 32508 30324
rect 32564 30268 34412 30324
rect 34468 30268 34748 30324
rect 34804 30268 34814 30324
rect 7532 30212 7588 30268
rect 6402 30156 6412 30212
rect 6468 30156 7084 30212
rect 7140 30156 7588 30212
rect 8876 30212 8932 30268
rect 12684 30212 12740 30268
rect 21532 30212 21588 30268
rect 8876 30156 10668 30212
rect 10724 30156 10734 30212
rect 12562 30156 12572 30212
rect 12628 30156 12740 30212
rect 20738 30156 20748 30212
rect 20804 30156 21588 30212
rect 21746 30156 21756 30212
rect 21812 30156 23884 30212
rect 23940 30156 23950 30212
rect 28578 30156 28588 30212
rect 28644 30156 29260 30212
rect 29316 30156 29326 30212
rect 8194 30044 8204 30100
rect 8260 30044 13020 30100
rect 13076 30044 13086 30100
rect 15092 30044 21532 30100
rect 21588 30044 21598 30100
rect 22082 30044 22092 30100
rect 22148 30044 24892 30100
rect 24948 30044 24958 30100
rect 15092 29988 15148 30044
rect 4610 29932 4620 29988
rect 4676 29932 5628 29988
rect 5684 29932 5694 29988
rect 7298 29932 7308 29988
rect 7364 29932 8316 29988
rect 8372 29932 8382 29988
rect 9986 29932 9996 29988
rect 10052 29932 10892 29988
rect 10948 29932 10958 29988
rect 11564 29932 15148 29988
rect 21970 29932 21980 29988
rect 22036 29932 23212 29988
rect 23268 29932 23278 29988
rect 32610 29932 32620 29988
rect 32676 29932 34188 29988
rect 34244 29932 34254 29988
rect 34598 29932 34636 29988
rect 34692 29932 34702 29988
rect 11564 29876 11620 29932
rect 10322 29820 10332 29876
rect 10388 29820 11620 29876
rect 13906 29820 13916 29876
rect 13972 29820 16380 29876
rect 16436 29820 16446 29876
rect 20402 29820 20412 29876
rect 20468 29820 21196 29876
rect 21252 29820 23324 29876
rect 23380 29820 23390 29876
rect 9770 29764 9780 29820
rect 9836 29764 9884 29820
rect 9940 29764 9988 29820
rect 10044 29764 10054 29820
rect 18338 29764 18348 29820
rect 18404 29764 18452 29820
rect 18508 29764 18556 29820
rect 18612 29764 18622 29820
rect 26906 29764 26916 29820
rect 26972 29764 27020 29820
rect 27076 29764 27124 29820
rect 27180 29764 27190 29820
rect 35474 29764 35484 29820
rect 35540 29764 35588 29820
rect 35644 29764 35692 29820
rect 35748 29764 35758 29820
rect 6738 29708 6748 29764
rect 6804 29708 8204 29764
rect 8260 29708 8270 29764
rect 9202 29708 9212 29764
rect 9268 29708 9548 29764
rect 9604 29708 9614 29764
rect 33170 29708 33180 29764
rect 33236 29708 34860 29764
rect 34916 29708 34926 29764
rect 34860 29652 34916 29708
rect 7858 29596 7868 29652
rect 7924 29596 8876 29652
rect 8932 29596 10108 29652
rect 10164 29596 10174 29652
rect 11106 29596 11116 29652
rect 11172 29596 11452 29652
rect 11508 29596 12572 29652
rect 12628 29596 12638 29652
rect 16818 29596 16828 29652
rect 16884 29596 19068 29652
rect 19124 29596 19134 29652
rect 23650 29596 23660 29652
rect 23716 29596 24108 29652
rect 24164 29596 24668 29652
rect 24724 29596 26908 29652
rect 28466 29596 28476 29652
rect 28532 29596 32284 29652
rect 32340 29596 32350 29652
rect 33842 29596 33852 29652
rect 33908 29596 34412 29652
rect 34468 29596 34478 29652
rect 34860 29596 35364 29652
rect 26852 29540 26908 29596
rect 5730 29484 5740 29540
rect 5796 29484 9996 29540
rect 10052 29484 10062 29540
rect 16930 29484 16940 29540
rect 16996 29484 18844 29540
rect 18900 29484 18910 29540
rect 21186 29484 21196 29540
rect 21252 29484 22204 29540
rect 22260 29484 22270 29540
rect 26852 29484 27132 29540
rect 27188 29484 32508 29540
rect 32564 29484 32574 29540
rect 34290 29484 34300 29540
rect 34356 29484 35140 29540
rect 35084 29428 35140 29484
rect 6514 29372 6524 29428
rect 6580 29372 7532 29428
rect 7588 29372 7756 29428
rect 7812 29372 8652 29428
rect 8708 29372 8718 29428
rect 9314 29372 9324 29428
rect 9380 29372 9884 29428
rect 9940 29372 9950 29428
rect 16258 29372 16268 29428
rect 16324 29372 17276 29428
rect 17332 29372 17342 29428
rect 17826 29372 17836 29428
rect 17892 29372 18620 29428
rect 18676 29372 18686 29428
rect 22754 29372 22764 29428
rect 22820 29372 25228 29428
rect 25284 29372 25294 29428
rect 33842 29372 33852 29428
rect 33908 29372 34524 29428
rect 34580 29372 34590 29428
rect 35046 29372 35084 29428
rect 35140 29372 35150 29428
rect 9538 29260 9548 29316
rect 9604 29260 11620 29316
rect 16594 29260 16604 29316
rect 16660 29260 17724 29316
rect 17780 29260 17790 29316
rect 18022 29260 18060 29316
rect 18116 29260 18126 29316
rect 23762 29260 23772 29316
rect 23828 29260 28924 29316
rect 28980 29260 28990 29316
rect 11564 29204 11620 29260
rect 35308 29204 35364 29596
rect 36200 29204 37000 29232
rect 8978 29148 8988 29204
rect 9044 29148 10780 29204
rect 10836 29148 10846 29204
rect 11554 29148 11564 29204
rect 11620 29148 16268 29204
rect 16324 29148 17164 29204
rect 17220 29148 17230 29204
rect 17378 29148 17388 29204
rect 17444 29148 17836 29204
rect 17892 29148 21980 29204
rect 22036 29148 22876 29204
rect 22932 29148 23212 29204
rect 23268 29148 23278 29204
rect 28802 29148 28812 29204
rect 28868 29148 33292 29204
rect 33348 29148 33358 29204
rect 35308 29148 37000 29204
rect 36200 29120 37000 29148
rect 16594 29036 16604 29092
rect 16660 29036 17052 29092
rect 17108 29036 17118 29092
rect 5486 28980 5496 29036
rect 5552 28980 5600 29036
rect 5656 28980 5704 29036
rect 5760 28980 5770 29036
rect 14054 28980 14064 29036
rect 14120 28980 14168 29036
rect 14224 28980 14272 29036
rect 14328 28980 14338 29036
rect 22622 28980 22632 29036
rect 22688 28980 22736 29036
rect 22792 28980 22840 29036
rect 22896 28980 22906 29036
rect 31190 28980 31200 29036
rect 31256 28980 31304 29036
rect 31360 28980 31408 29036
rect 31464 28980 31474 29036
rect 8754 28924 8764 28980
rect 8820 28924 9324 28980
rect 9380 28924 10892 28980
rect 10948 28924 13692 28980
rect 13748 28924 13758 28980
rect 16370 28924 16380 28980
rect 16436 28924 17836 28980
rect 17892 28924 17902 28980
rect 18918 28924 18956 28980
rect 19012 28924 19022 28980
rect 5170 28812 5180 28868
rect 5236 28812 6860 28868
rect 6916 28812 6926 28868
rect 11218 28812 11228 28868
rect 11284 28812 19740 28868
rect 19796 28812 19806 28868
rect 6626 28700 6636 28756
rect 6692 28700 7308 28756
rect 7364 28700 7644 28756
rect 7700 28700 7710 28756
rect 11778 28700 11788 28756
rect 11844 28700 12236 28756
rect 12292 28700 15372 28756
rect 15428 28700 15438 28756
rect 15922 28700 15932 28756
rect 15988 28700 17500 28756
rect 17556 28700 17566 28756
rect 19282 28700 19292 28756
rect 19348 28700 21308 28756
rect 21364 28700 21374 28756
rect 26562 28700 26572 28756
rect 26628 28700 28476 28756
rect 28532 28700 28542 28756
rect 6850 28588 6860 28644
rect 6916 28588 12460 28644
rect 12516 28588 12684 28644
rect 12740 28588 12750 28644
rect 15026 28588 15036 28644
rect 15092 28588 15820 28644
rect 15876 28588 15886 28644
rect 16940 28588 18732 28644
rect 18788 28588 18798 28644
rect 21186 28588 21196 28644
rect 21252 28588 23772 28644
rect 23828 28588 23838 28644
rect 9986 28476 9996 28532
rect 10052 28476 11340 28532
rect 11396 28476 11406 28532
rect 12684 28308 12740 28588
rect 16940 28532 16996 28588
rect 13794 28476 13804 28532
rect 13860 28476 14588 28532
rect 14644 28476 14654 28532
rect 16930 28476 16940 28532
rect 16996 28476 17006 28532
rect 19954 28476 19964 28532
rect 20020 28476 21308 28532
rect 21364 28476 21374 28532
rect 27570 28476 27580 28532
rect 27636 28476 28700 28532
rect 28756 28476 28766 28532
rect 13682 28364 13692 28420
rect 13748 28364 14700 28420
rect 14756 28364 14766 28420
rect 18946 28364 18956 28420
rect 19012 28364 19852 28420
rect 19908 28364 19918 28420
rect 20290 28364 20300 28420
rect 20356 28364 21420 28420
rect 21476 28364 21486 28420
rect 26226 28364 26236 28420
rect 26292 28364 28364 28420
rect 28420 28364 28430 28420
rect 30258 28364 30268 28420
rect 30324 28364 33068 28420
rect 33124 28364 33134 28420
rect 33394 28364 33404 28420
rect 33460 28364 34076 28420
rect 34132 28364 34142 28420
rect 8530 28252 8540 28308
rect 8596 28252 9324 28308
rect 9380 28252 9390 28308
rect 12684 28252 17500 28308
rect 17556 28252 17566 28308
rect 17714 28252 17724 28308
rect 17780 28252 18172 28308
rect 18228 28252 18238 28308
rect 18834 28252 18844 28308
rect 18900 28252 19292 28308
rect 19348 28252 22316 28308
rect 22372 28252 22382 28308
rect 24546 28252 24556 28308
rect 24612 28252 25228 28308
rect 25284 28252 25294 28308
rect 27346 28252 27356 28308
rect 27412 28252 33628 28308
rect 33684 28252 33694 28308
rect 9770 28196 9780 28252
rect 9836 28196 9884 28252
rect 9940 28196 9988 28252
rect 10044 28196 10054 28252
rect 18338 28196 18348 28252
rect 18404 28196 18452 28252
rect 18508 28196 18556 28252
rect 18612 28196 18622 28252
rect 24556 28196 24612 28252
rect 26906 28196 26916 28252
rect 26972 28196 27020 28252
rect 27076 28196 27124 28252
rect 27180 28196 27190 28252
rect 35474 28196 35484 28252
rect 35540 28196 35588 28252
rect 35644 28196 35692 28252
rect 35748 28196 35758 28252
rect 15586 28140 15596 28196
rect 15652 28140 17612 28196
rect 17668 28140 17678 28196
rect 19506 28140 19516 28196
rect 19572 28140 22204 28196
rect 22260 28140 24612 28196
rect 27346 28140 27356 28196
rect 27412 28140 32060 28196
rect 32116 28140 32126 28196
rect 33170 28140 33180 28196
rect 33236 28140 34636 28196
rect 34692 28140 34702 28196
rect 32060 28084 32116 28140
rect 7410 28028 7420 28084
rect 7476 28028 8540 28084
rect 8596 28028 8764 28084
rect 8820 28028 8830 28084
rect 18050 28028 18060 28084
rect 18116 28028 21756 28084
rect 21812 28028 21822 28084
rect 29250 28028 29260 28084
rect 29316 28028 30380 28084
rect 30436 28028 30446 28084
rect 32060 28028 34412 28084
rect 34468 28028 34478 28084
rect 34738 28028 34748 28084
rect 34804 28028 35084 28084
rect 35140 28028 35150 28084
rect 9090 27916 9100 27972
rect 9156 27916 10332 27972
rect 10388 27916 10398 27972
rect 13682 27916 13692 27972
rect 13748 27916 14252 27972
rect 14308 27916 14318 27972
rect 15138 27916 15148 27972
rect 15204 27916 17388 27972
rect 17444 27916 19516 27972
rect 19572 27916 19582 27972
rect 20738 27916 20748 27972
rect 20804 27916 23212 27972
rect 23268 27916 25564 27972
rect 25620 27916 25630 27972
rect 30706 27916 30716 27972
rect 30772 27916 32172 27972
rect 32228 27916 32238 27972
rect 8978 27804 8988 27860
rect 9044 27804 10892 27860
rect 10948 27804 10958 27860
rect 12002 27804 12012 27860
rect 12068 27804 13692 27860
rect 13748 27804 14812 27860
rect 14868 27804 14878 27860
rect 17714 27804 17724 27860
rect 17780 27804 19404 27860
rect 19460 27804 19470 27860
rect 20962 27804 20972 27860
rect 21028 27804 21868 27860
rect 21924 27804 21934 27860
rect 22418 27804 22428 27860
rect 22484 27804 26236 27860
rect 26292 27804 26302 27860
rect 30482 27804 30492 27860
rect 30548 27804 32396 27860
rect 32452 27804 32462 27860
rect 34402 27804 34412 27860
rect 34468 27804 35084 27860
rect 35140 27804 35150 27860
rect 10892 27748 10948 27804
rect 5954 27692 5964 27748
rect 6020 27692 6972 27748
rect 7028 27692 7038 27748
rect 9538 27692 9548 27748
rect 9604 27692 9884 27748
rect 9940 27692 9950 27748
rect 10892 27692 15036 27748
rect 15092 27636 15148 27748
rect 15474 27692 15484 27748
rect 15540 27692 16044 27748
rect 16100 27692 18956 27748
rect 19012 27692 19068 27748
rect 19124 27692 19134 27748
rect 20514 27692 20524 27748
rect 20580 27692 21308 27748
rect 21364 27692 21374 27748
rect 31266 27692 31276 27748
rect 31332 27692 32060 27748
rect 32116 27692 32126 27748
rect 32284 27636 32340 27804
rect 6514 27580 6524 27636
rect 6580 27580 8092 27636
rect 8148 27580 10892 27636
rect 10948 27580 10958 27636
rect 12786 27580 12796 27636
rect 12852 27580 13804 27636
rect 13860 27580 13870 27636
rect 15092 27580 18452 27636
rect 19702 27580 19740 27636
rect 19796 27580 19806 27636
rect 20402 27580 20412 27636
rect 20468 27580 24892 27636
rect 24948 27580 24958 27636
rect 27122 27580 27132 27636
rect 27188 27580 27804 27636
rect 27860 27580 31612 27636
rect 31668 27580 31678 27636
rect 32162 27580 32172 27636
rect 32228 27580 32340 27636
rect 18396 27524 18452 27580
rect 18396 27468 19852 27524
rect 19908 27468 19918 27524
rect 30044 27468 30268 27524
rect 30324 27468 30334 27524
rect 5486 27412 5496 27468
rect 5552 27412 5600 27468
rect 5656 27412 5704 27468
rect 5760 27412 5770 27468
rect 14054 27412 14064 27468
rect 14120 27412 14168 27468
rect 14224 27412 14272 27468
rect 14328 27412 14338 27468
rect 22622 27412 22632 27468
rect 22688 27412 22736 27468
rect 22792 27412 22840 27468
rect 22896 27412 22906 27468
rect 30044 27412 30100 27468
rect 31190 27412 31200 27468
rect 31256 27412 31304 27468
rect 31360 27412 31408 27468
rect 31464 27412 31474 27468
rect 6290 27356 6300 27412
rect 6356 27356 7196 27412
rect 7252 27356 12908 27412
rect 12964 27356 13468 27412
rect 13524 27356 13534 27412
rect 16370 27356 16380 27412
rect 16436 27356 17836 27412
rect 17892 27356 20076 27412
rect 20132 27356 20142 27412
rect 30034 27356 30044 27412
rect 30100 27356 30110 27412
rect 4274 27244 4284 27300
rect 4340 27244 5628 27300
rect 5684 27244 5694 27300
rect 10322 27244 10332 27300
rect 10388 27244 11900 27300
rect 11956 27244 14588 27300
rect 14644 27244 14654 27300
rect 15698 27244 15708 27300
rect 15764 27244 18284 27300
rect 18340 27244 18350 27300
rect 18498 27244 18508 27300
rect 18564 27244 18956 27300
rect 19012 27244 19022 27300
rect 21746 27244 21756 27300
rect 21812 27244 22652 27300
rect 22708 27244 23100 27300
rect 23156 27244 23166 27300
rect 23426 27244 23436 27300
rect 23492 27244 23502 27300
rect 23436 27188 23492 27244
rect 6962 27132 6972 27188
rect 7028 27132 7420 27188
rect 7476 27132 7486 27188
rect 9874 27132 9884 27188
rect 9940 27132 11452 27188
rect 11508 27132 11518 27188
rect 14690 27132 14700 27188
rect 14756 27132 15260 27188
rect 15316 27132 18844 27188
rect 18900 27132 23492 27188
rect 25890 27132 25900 27188
rect 25956 27132 26572 27188
rect 26628 27132 26638 27188
rect 29922 27132 29932 27188
rect 29988 27132 32732 27188
rect 32788 27132 32798 27188
rect 6850 27020 6860 27076
rect 6916 27020 7868 27076
rect 7924 27020 7934 27076
rect 8194 27020 8204 27076
rect 8260 27020 8540 27076
rect 8596 27020 8606 27076
rect 10098 27020 10108 27076
rect 10164 27020 11004 27076
rect 11060 27020 11070 27076
rect 12562 27020 12572 27076
rect 12628 27020 14980 27076
rect 14924 26964 14980 27020
rect 16828 27020 17500 27076
rect 17556 27020 17566 27076
rect 17798 27020 17836 27076
rect 17892 27020 17902 27076
rect 18722 27020 18732 27076
rect 18788 27020 19852 27076
rect 19908 27020 19918 27076
rect 20066 27020 20076 27076
rect 20132 27020 20142 27076
rect 20514 27020 20524 27076
rect 20580 27020 22428 27076
rect 22484 27020 22494 27076
rect 16828 26964 16884 27020
rect 20076 26964 20132 27020
rect 12338 26908 12348 26964
rect 12404 26908 14700 26964
rect 14756 26908 14766 26964
rect 14924 26908 16828 26964
rect 16884 26908 16894 26964
rect 17266 26908 17276 26964
rect 17332 26908 18284 26964
rect 18340 26908 18350 26964
rect 19730 26908 19740 26964
rect 19796 26908 20132 26964
rect 20188 26908 20860 26964
rect 20916 26908 20926 26964
rect 22530 26908 22540 26964
rect 22596 26908 24444 26964
rect 24500 26908 24510 26964
rect 14924 26852 14980 26908
rect 7868 26796 9884 26852
rect 9940 26796 9950 26852
rect 13878 26796 13916 26852
rect 13972 26796 13982 26852
rect 14802 26796 14812 26852
rect 14868 26796 14980 26852
rect 19618 26796 19628 26852
rect 19684 26796 19740 26852
rect 19796 26796 19806 26852
rect 7868 26740 7924 26796
rect 20188 26740 20244 26908
rect 21410 26796 21420 26852
rect 21476 26796 22652 26852
rect 22708 26796 22718 26852
rect 23650 26796 23660 26852
rect 23716 26796 26796 26852
rect 26852 26796 26862 26852
rect 34066 26796 34076 26852
rect 34132 26796 35084 26852
rect 35140 26796 35150 26852
rect 7858 26684 7868 26740
rect 7924 26684 7934 26740
rect 15092 26684 16940 26740
rect 16996 26684 17388 26740
rect 17444 26684 17454 26740
rect 20150 26684 20188 26740
rect 20244 26684 22540 26740
rect 22596 26684 25564 26740
rect 25620 26684 25630 26740
rect 34178 26684 34188 26740
rect 34244 26684 34860 26740
rect 34916 26684 34926 26740
rect 9770 26628 9780 26684
rect 9836 26628 9884 26684
rect 9940 26628 9988 26684
rect 10044 26628 10054 26684
rect 15092 26628 15148 26684
rect 18338 26628 18348 26684
rect 18404 26628 18452 26684
rect 18508 26628 18556 26684
rect 18612 26628 18622 26684
rect 26906 26628 26916 26684
rect 26972 26628 27020 26684
rect 27076 26628 27124 26684
rect 27180 26628 27190 26684
rect 35474 26628 35484 26684
rect 35540 26628 35588 26684
rect 35644 26628 35692 26684
rect 35748 26628 35758 26684
rect 6850 26572 6860 26628
rect 6916 26572 7308 26628
rect 7364 26572 7374 26628
rect 7606 26572 7644 26628
rect 7700 26572 7710 26628
rect 8166 26572 8204 26628
rect 8260 26572 8270 26628
rect 8530 26572 8540 26628
rect 8596 26572 8932 26628
rect 10770 26572 10780 26628
rect 10836 26572 15148 26628
rect 18050 26572 18060 26628
rect 18116 26572 18228 26628
rect 19730 26572 19740 26628
rect 19796 26572 20076 26628
rect 20132 26572 20142 26628
rect 20626 26572 20636 26628
rect 20692 26572 21756 26628
rect 21812 26572 21822 26628
rect 8876 26516 8932 26572
rect 18172 26516 18228 26572
rect 36200 26516 37000 26544
rect 5730 26460 5740 26516
rect 5796 26460 8428 26516
rect 8484 26460 8494 26516
rect 8876 26460 9772 26516
rect 9828 26460 13356 26516
rect 13412 26460 15708 26516
rect 15764 26460 15774 26516
rect 18172 26460 18396 26516
rect 18452 26460 18462 26516
rect 20850 26460 20860 26516
rect 20916 26460 22092 26516
rect 22148 26460 22158 26516
rect 24658 26460 24668 26516
rect 24724 26460 25564 26516
rect 25620 26460 25630 26516
rect 27570 26460 27580 26516
rect 27636 26460 28812 26516
rect 28868 26460 28878 26516
rect 32834 26460 32844 26516
rect 32900 26460 33180 26516
rect 33236 26460 33246 26516
rect 34962 26460 34972 26516
rect 35028 26460 37000 26516
rect 36200 26432 37000 26460
rect 7410 26348 7420 26404
rect 7476 26348 7644 26404
rect 7700 26348 7710 26404
rect 8194 26348 8204 26404
rect 8260 26348 9884 26404
rect 9940 26348 9950 26404
rect 11554 26348 11564 26404
rect 11620 26348 12460 26404
rect 12516 26348 12526 26404
rect 14914 26348 14924 26404
rect 14980 26348 15820 26404
rect 15876 26348 15886 26404
rect 17154 26348 17164 26404
rect 17220 26348 19068 26404
rect 19124 26348 19134 26404
rect 22418 26348 22428 26404
rect 22484 26348 23212 26404
rect 23268 26348 23884 26404
rect 23940 26348 23950 26404
rect 33954 26348 33964 26404
rect 34020 26348 34412 26404
rect 34468 26348 34478 26404
rect 34850 26348 34860 26404
rect 34916 26348 35196 26404
rect 35252 26348 35262 26404
rect 9426 26236 9436 26292
rect 9492 26236 15148 26292
rect 15250 26236 15260 26292
rect 15316 26236 16156 26292
rect 16212 26236 16716 26292
rect 16772 26236 16782 26292
rect 17714 26236 17724 26292
rect 17780 26236 18060 26292
rect 18116 26236 18126 26292
rect 18284 26236 20412 26292
rect 20468 26236 20478 26292
rect 21858 26236 21868 26292
rect 21924 26236 22764 26292
rect 22820 26236 25340 26292
rect 25396 26236 25406 26292
rect 26674 26236 26684 26292
rect 26740 26236 28140 26292
rect 28196 26236 28206 26292
rect 33170 26236 33180 26292
rect 33236 26236 34300 26292
rect 34356 26236 34366 26292
rect 15092 26180 15148 26236
rect 18284 26180 18340 26236
rect 4386 26124 4396 26180
rect 4452 26124 6188 26180
rect 6244 26124 6254 26180
rect 12114 26124 12124 26180
rect 12180 26124 13132 26180
rect 13188 26124 13198 26180
rect 15092 26124 16492 26180
rect 16548 26124 18340 26180
rect 19730 26124 19740 26180
rect 19796 26124 21756 26180
rect 21812 26124 21822 26180
rect 10434 26012 10444 26068
rect 10500 26012 11900 26068
rect 11956 26012 11966 26068
rect 12684 26012 14700 26068
rect 14756 26012 14924 26068
rect 14980 26012 14990 26068
rect 21410 26012 21420 26068
rect 21476 26012 22204 26068
rect 22260 26012 22270 26068
rect 22428 26012 27916 26068
rect 27972 26012 27982 26068
rect 12684 25956 12740 26012
rect 22428 25956 22484 26012
rect 8530 25900 8540 25956
rect 8596 25900 9884 25956
rect 9940 25900 12740 25956
rect 15026 25900 15036 25956
rect 15092 25900 22484 25956
rect 33058 25900 33068 25956
rect 33124 25900 33740 25956
rect 33796 25900 33806 25956
rect 5486 25844 5496 25900
rect 5552 25844 5600 25900
rect 5656 25844 5704 25900
rect 5760 25844 5770 25900
rect 14054 25844 14064 25900
rect 14120 25844 14168 25900
rect 14224 25844 14272 25900
rect 14328 25844 14338 25900
rect 22622 25844 22632 25900
rect 22688 25844 22736 25900
rect 22792 25844 22840 25900
rect 22896 25844 22906 25900
rect 31190 25844 31200 25900
rect 31256 25844 31304 25900
rect 31360 25844 31408 25900
rect 31464 25844 31474 25900
rect 15474 25788 15484 25844
rect 15540 25788 16268 25844
rect 16324 25788 16334 25844
rect 18498 25788 18508 25844
rect 18564 25788 20412 25844
rect 20468 25788 21308 25844
rect 21364 25788 21374 25844
rect 21858 25788 21868 25844
rect 21924 25788 22036 25844
rect 34150 25788 34188 25844
rect 34244 25788 34254 25844
rect 16706 25676 16716 25732
rect 16772 25676 19628 25732
rect 19684 25676 19694 25732
rect 19842 25676 19852 25732
rect 19908 25676 21756 25732
rect 21812 25676 21822 25732
rect 21980 25620 22036 25788
rect 27458 25676 27468 25732
rect 27524 25676 28028 25732
rect 28084 25676 29428 25732
rect 29586 25676 29596 25732
rect 29652 25676 34860 25732
rect 34916 25676 34926 25732
rect 29372 25620 29428 25676
rect 13682 25564 13692 25620
rect 13748 25564 14028 25620
rect 14084 25564 17724 25620
rect 17780 25564 17790 25620
rect 19170 25564 19180 25620
rect 19236 25564 22036 25620
rect 23874 25564 23884 25620
rect 23940 25564 26460 25620
rect 26516 25564 29148 25620
rect 29204 25564 29214 25620
rect 29372 25564 33180 25620
rect 33236 25564 33404 25620
rect 33460 25564 33470 25620
rect 12898 25452 12908 25508
rect 12964 25452 15036 25508
rect 15092 25452 15102 25508
rect 17378 25452 17388 25508
rect 17444 25452 19404 25508
rect 19460 25452 19740 25508
rect 19796 25452 19806 25508
rect 27122 25452 27132 25508
rect 27188 25452 27692 25508
rect 27748 25452 27758 25508
rect 29474 25452 29484 25508
rect 29540 25452 31612 25508
rect 31668 25452 31678 25508
rect 6290 25340 6300 25396
rect 6356 25340 10220 25396
rect 10276 25340 10286 25396
rect 15092 25340 18508 25396
rect 18564 25340 18574 25396
rect 18834 25340 18844 25396
rect 18900 25340 19516 25396
rect 19572 25340 22092 25396
rect 22148 25340 22158 25396
rect 22978 25340 22988 25396
rect 23044 25340 24220 25396
rect 24276 25340 24286 25396
rect 28466 25340 28476 25396
rect 28532 25340 32844 25396
rect 32900 25340 32910 25396
rect 15092 25284 15148 25340
rect 3602 25228 3612 25284
rect 3668 25228 6860 25284
rect 6916 25228 6926 25284
rect 8082 25228 8092 25284
rect 8148 25228 12236 25284
rect 12292 25228 15148 25284
rect 18386 25228 18396 25284
rect 18452 25228 20188 25284
rect 20244 25228 20972 25284
rect 21028 25228 21038 25284
rect 23090 25228 23100 25284
rect 23156 25228 23436 25284
rect 23492 25228 23502 25284
rect 26002 25228 26012 25284
rect 26068 25228 33180 25284
rect 33236 25228 33246 25284
rect 34178 25228 34188 25284
rect 34244 25228 34254 25284
rect 13654 25116 13692 25172
rect 13748 25116 13758 25172
rect 21746 25116 21756 25172
rect 21812 25116 23660 25172
rect 23716 25116 23726 25172
rect 30594 25116 30604 25172
rect 30660 25116 33628 25172
rect 33684 25116 33694 25172
rect 9770 25060 9780 25116
rect 9836 25060 9884 25116
rect 9940 25060 9988 25116
rect 10044 25060 10054 25116
rect 18338 25060 18348 25116
rect 18404 25060 18452 25116
rect 18508 25060 18556 25116
rect 18612 25060 18622 25116
rect 26906 25060 26916 25116
rect 26972 25060 27020 25116
rect 27076 25060 27124 25116
rect 27180 25060 27190 25116
rect 34188 25060 34244 25228
rect 35474 25060 35484 25116
rect 35540 25060 35588 25116
rect 35644 25060 35692 25116
rect 35748 25060 35758 25116
rect 13234 25004 13244 25060
rect 13300 25004 14252 25060
rect 14308 25004 15092 25060
rect 29362 25004 29372 25060
rect 29428 25004 30044 25060
rect 30100 25004 30110 25060
rect 31042 25004 31052 25060
rect 31108 25004 34244 25060
rect 15036 24948 15092 25004
rect 12226 24892 12236 24948
rect 12292 24892 12796 24948
rect 12852 24892 14812 24948
rect 14868 24892 14878 24948
rect 15036 24892 19852 24948
rect 19908 24892 19918 24948
rect 24210 24892 24220 24948
rect 24276 24892 25228 24948
rect 25284 24892 25294 24948
rect 25442 24892 25452 24948
rect 25508 24892 30940 24948
rect 30996 24892 31006 24948
rect 32162 24892 32172 24948
rect 32228 24892 32238 24948
rect 34150 24892 34188 24948
rect 34244 24892 34254 24948
rect 11554 24780 11564 24836
rect 11620 24780 12012 24836
rect 12068 24780 12348 24836
rect 12404 24780 12414 24836
rect 14812 24724 14868 24892
rect 28354 24780 28364 24836
rect 28420 24780 29372 24836
rect 29428 24780 29438 24836
rect 32172 24724 32228 24892
rect 32834 24780 32844 24836
rect 32900 24780 35084 24836
rect 35140 24780 35150 24836
rect 6626 24668 6636 24724
rect 6692 24668 7196 24724
rect 7252 24668 7756 24724
rect 7812 24668 8316 24724
rect 8372 24668 9548 24724
rect 9604 24668 9614 24724
rect 14812 24668 15596 24724
rect 15652 24668 15662 24724
rect 16706 24668 16716 24724
rect 16772 24668 17052 24724
rect 17108 24668 20412 24724
rect 20468 24668 20478 24724
rect 23762 24668 23772 24724
rect 23828 24668 25228 24724
rect 25284 24668 25294 24724
rect 29026 24668 29036 24724
rect 29092 24668 33180 24724
rect 33236 24668 34860 24724
rect 34916 24668 34926 24724
rect 16716 24500 16772 24668
rect 17154 24556 17164 24612
rect 17220 24556 17724 24612
rect 17780 24556 18172 24612
rect 18228 24556 18844 24612
rect 18900 24556 18910 24612
rect 27458 24556 27468 24612
rect 27524 24556 31164 24612
rect 31220 24556 32956 24612
rect 33012 24556 33022 24612
rect 33394 24556 33404 24612
rect 33460 24556 34412 24612
rect 34468 24556 34478 24612
rect 32956 24500 33012 24556
rect 9090 24444 9100 24500
rect 9156 24444 9884 24500
rect 9940 24444 11116 24500
rect 11172 24444 13132 24500
rect 13188 24444 13580 24500
rect 13636 24444 14476 24500
rect 14532 24444 16772 24500
rect 29586 24444 29596 24500
rect 29652 24444 30716 24500
rect 30772 24444 30782 24500
rect 32956 24444 33740 24500
rect 33796 24444 33806 24500
rect 33954 24444 33964 24500
rect 34020 24444 34636 24500
rect 34692 24444 34702 24500
rect 26786 24332 26796 24388
rect 26852 24332 27804 24388
rect 27860 24332 28868 24388
rect 31602 24332 31612 24388
rect 31668 24332 33852 24388
rect 33908 24332 33918 24388
rect 5486 24276 5496 24332
rect 5552 24276 5600 24332
rect 5656 24276 5704 24332
rect 5760 24276 5770 24332
rect 14054 24276 14064 24332
rect 14120 24276 14168 24332
rect 14224 24276 14272 24332
rect 14328 24276 14338 24332
rect 22622 24276 22632 24332
rect 22688 24276 22736 24332
rect 22792 24276 22840 24332
rect 22896 24276 22906 24332
rect 28812 24276 28868 24332
rect 31190 24276 31200 24332
rect 31256 24276 31304 24332
rect 31360 24276 31408 24332
rect 31464 24276 31474 24332
rect 23986 24220 23996 24276
rect 24052 24220 27132 24276
rect 27188 24220 28364 24276
rect 28420 24220 28430 24276
rect 28802 24220 28812 24276
rect 28868 24220 29820 24276
rect 29876 24220 29886 24276
rect 25554 24108 25564 24164
rect 25620 24108 28588 24164
rect 28644 24108 30492 24164
rect 30548 24108 30558 24164
rect 23874 23996 23884 24052
rect 23940 23996 24332 24052
rect 24388 23996 26012 24052
rect 26068 23996 26078 24052
rect 12898 23884 12908 23940
rect 12964 23884 13580 23940
rect 13636 23884 14252 23940
rect 14308 23884 15148 23940
rect 19170 23884 19180 23940
rect 19236 23884 19852 23940
rect 19908 23884 19918 23940
rect 21522 23884 21532 23940
rect 21588 23884 22316 23940
rect 22372 23884 22764 23940
rect 22820 23884 22830 23940
rect 32162 23884 32172 23940
rect 32228 23884 32732 23940
rect 32788 23884 32798 23940
rect 7298 23772 7308 23828
rect 7364 23772 7756 23828
rect 7812 23772 10220 23828
rect 10276 23772 10286 23828
rect 15092 23716 15148 23884
rect 36200 23828 37000 23856
rect 17938 23772 17948 23828
rect 18004 23772 18956 23828
rect 19012 23772 19022 23828
rect 19506 23772 19516 23828
rect 19572 23772 20636 23828
rect 20692 23772 20702 23828
rect 27794 23772 27804 23828
rect 27860 23772 37000 23828
rect 36200 23744 37000 23772
rect 6738 23660 6748 23716
rect 6804 23660 7420 23716
rect 7476 23660 7868 23716
rect 7924 23660 7934 23716
rect 15092 23660 19740 23716
rect 19796 23660 20860 23716
rect 20916 23660 21084 23716
rect 21140 23660 21150 23716
rect 25442 23660 25452 23716
rect 25508 23660 26236 23716
rect 26292 23660 26302 23716
rect 26450 23660 26460 23716
rect 26516 23660 27580 23716
rect 27636 23660 27646 23716
rect 28242 23660 28252 23716
rect 28308 23660 29260 23716
rect 29316 23660 29326 23716
rect 12002 23548 12012 23604
rect 12068 23548 13356 23604
rect 13412 23548 13422 23604
rect 18722 23548 18732 23604
rect 18788 23548 19292 23604
rect 19348 23548 21308 23604
rect 21364 23548 21374 23604
rect 24322 23548 24332 23604
rect 24388 23548 24398 23604
rect 25106 23548 25116 23604
rect 25172 23548 26740 23604
rect 28018 23548 28028 23604
rect 28084 23548 28588 23604
rect 28644 23548 28654 23604
rect 32274 23548 32284 23604
rect 32340 23548 33180 23604
rect 33236 23548 33246 23604
rect 9770 23492 9780 23548
rect 9836 23492 9884 23548
rect 9940 23492 9988 23548
rect 10044 23492 10054 23548
rect 18338 23492 18348 23548
rect 18404 23492 18452 23548
rect 18508 23492 18556 23548
rect 18612 23492 18622 23548
rect 24332 23492 24388 23548
rect 6962 23436 6972 23492
rect 7028 23436 7980 23492
rect 8036 23436 8046 23492
rect 23538 23436 23548 23492
rect 23604 23436 24388 23492
rect 26114 23436 26124 23492
rect 26180 23436 26460 23492
rect 26516 23436 26526 23492
rect 17154 23324 17164 23380
rect 17220 23324 17724 23380
rect 17780 23324 17790 23380
rect 24658 23324 24668 23380
rect 24724 23324 26348 23380
rect 26404 23324 26414 23380
rect 26684 23268 26740 23548
rect 26906 23492 26916 23548
rect 26972 23492 27020 23548
rect 27076 23492 27124 23548
rect 27180 23492 27190 23548
rect 35474 23492 35484 23548
rect 35540 23492 35588 23548
rect 35644 23492 35692 23548
rect 35748 23492 35758 23548
rect 28354 23436 28364 23492
rect 28420 23436 29036 23492
rect 29092 23436 29102 23492
rect 27346 23324 27356 23380
rect 27412 23324 34188 23380
rect 34244 23324 34748 23380
rect 34804 23324 34814 23380
rect 24434 23212 24444 23268
rect 24500 23212 24510 23268
rect 26684 23212 27132 23268
rect 27188 23212 27198 23268
rect 28242 23212 28252 23268
rect 28308 23212 31948 23268
rect 32004 23212 33292 23268
rect 33348 23212 33358 23268
rect 8418 23100 8428 23156
rect 8484 23100 9436 23156
rect 9492 23100 9502 23156
rect 10546 23100 10556 23156
rect 10612 23100 13804 23156
rect 13860 23100 13870 23156
rect 19954 23100 19964 23156
rect 20020 23100 23212 23156
rect 23268 23100 23278 23156
rect 24444 23044 24500 23212
rect 26460 23100 28924 23156
rect 28980 23100 29148 23156
rect 29204 23100 29214 23156
rect 29922 23100 29932 23156
rect 29988 23100 29998 23156
rect 30258 23100 30268 23156
rect 30324 23100 31836 23156
rect 31892 23100 31902 23156
rect 32050 23100 32060 23156
rect 32116 23100 35252 23156
rect 4722 22988 4732 23044
rect 4788 22988 7308 23044
rect 7364 22988 7374 23044
rect 20626 22988 20636 23044
rect 20692 22988 21644 23044
rect 21700 22988 21710 23044
rect 23650 22988 23660 23044
rect 23716 22988 25228 23044
rect 25284 22988 25294 23044
rect 26460 22932 26516 23100
rect 29932 23044 29988 23100
rect 35196 23044 35252 23100
rect 26674 22988 26684 23044
rect 26740 22988 29988 23044
rect 31714 22988 31724 23044
rect 31780 22988 33628 23044
rect 33684 22988 33694 23044
rect 35186 22988 35196 23044
rect 35252 22988 35262 23044
rect 19394 22876 19404 22932
rect 19460 22876 21532 22932
rect 21588 22876 21598 22932
rect 21756 22876 26516 22932
rect 27010 22876 27020 22932
rect 27076 22876 27804 22932
rect 27860 22876 27870 22932
rect 28802 22876 28812 22932
rect 28868 22876 29820 22932
rect 29876 22876 30604 22932
rect 30660 22876 30670 22932
rect 30818 22876 30828 22932
rect 30884 22876 34300 22932
rect 34356 22876 34366 22932
rect 21756 22820 21812 22876
rect 19730 22764 19740 22820
rect 19796 22764 21812 22820
rect 26226 22764 26236 22820
rect 26292 22764 26302 22820
rect 27990 22764 28028 22820
rect 28084 22764 28094 22820
rect 5486 22708 5496 22764
rect 5552 22708 5600 22764
rect 5656 22708 5704 22764
rect 5760 22708 5770 22764
rect 14054 22708 14064 22764
rect 14120 22708 14168 22764
rect 14224 22708 14272 22764
rect 14328 22708 14338 22764
rect 22622 22708 22632 22764
rect 22688 22708 22736 22764
rect 22792 22708 22840 22764
rect 22896 22708 22906 22764
rect 26236 22708 26292 22764
rect 31190 22708 31200 22764
rect 31256 22708 31304 22764
rect 31360 22708 31408 22764
rect 31464 22708 31474 22764
rect 8194 22652 8204 22708
rect 8260 22652 9660 22708
rect 9716 22652 9726 22708
rect 26236 22652 30268 22708
rect 30324 22652 30334 22708
rect 7074 22540 7084 22596
rect 7140 22540 7756 22596
rect 7812 22540 10108 22596
rect 10164 22540 11564 22596
rect 11620 22540 11630 22596
rect 18050 22540 18060 22596
rect 18116 22540 19404 22596
rect 19460 22540 19470 22596
rect 23538 22540 23548 22596
rect 23604 22540 31612 22596
rect 31668 22540 31678 22596
rect 34710 22540 34748 22596
rect 34804 22540 34814 22596
rect 34962 22540 34972 22596
rect 35028 22540 36204 22596
rect 36260 22540 36270 22596
rect 8866 22428 8876 22484
rect 8932 22428 10332 22484
rect 10388 22428 10398 22484
rect 13794 22428 13804 22484
rect 13860 22428 16100 22484
rect 24658 22428 24668 22484
rect 24724 22428 29148 22484
rect 29204 22428 29820 22484
rect 29876 22428 29886 22484
rect 34402 22428 34412 22484
rect 34468 22428 34860 22484
rect 34916 22428 34926 22484
rect 16044 22372 16100 22428
rect 16034 22316 16044 22372
rect 16100 22316 17500 22372
rect 17556 22316 17566 22372
rect 27234 22316 27244 22372
rect 27300 22316 27916 22372
rect 27972 22316 29036 22372
rect 29092 22316 29102 22372
rect 29250 22316 29260 22372
rect 29316 22316 30940 22372
rect 30996 22316 31006 22372
rect 31378 22316 31388 22372
rect 31444 22316 32060 22372
rect 32116 22316 32126 22372
rect 33030 22316 33068 22372
rect 33124 22316 33134 22372
rect 11554 22204 11564 22260
rect 11620 22204 12460 22260
rect 12516 22204 12526 22260
rect 12898 22204 12908 22260
rect 12964 22204 20748 22260
rect 20804 22204 21308 22260
rect 21364 22204 22316 22260
rect 22372 22204 22382 22260
rect 30034 22204 30044 22260
rect 30100 22204 30828 22260
rect 30884 22204 30894 22260
rect 4386 22092 4396 22148
rect 4452 22092 6636 22148
rect 6692 22092 6702 22148
rect 10098 22092 10108 22148
rect 10164 22092 11900 22148
rect 11956 22092 11966 22148
rect 13570 22092 13580 22148
rect 13636 22092 15260 22148
rect 15316 22092 19964 22148
rect 20020 22092 20030 22148
rect 25218 22092 25228 22148
rect 25284 22092 26460 22148
rect 26516 22092 26526 22148
rect 29922 22092 29932 22148
rect 29988 22092 32172 22148
rect 32228 22092 32238 22148
rect 34290 22092 34300 22148
rect 34356 22092 34636 22148
rect 34692 22092 34702 22148
rect 34300 22036 34356 22092
rect 16818 21980 16828 22036
rect 16884 21980 18172 22036
rect 18228 21980 18238 22036
rect 25778 21980 25788 22036
rect 25844 21980 26684 22036
rect 26740 21980 26750 22036
rect 28466 21980 28476 22036
rect 28532 21980 28588 22036
rect 28644 21980 34356 22036
rect 9770 21924 9780 21980
rect 9836 21924 9884 21980
rect 9940 21924 9988 21980
rect 10044 21924 10054 21980
rect 18338 21924 18348 21980
rect 18404 21924 18452 21980
rect 18508 21924 18556 21980
rect 18612 21924 18622 21980
rect 26906 21924 26916 21980
rect 26972 21924 27020 21980
rect 27076 21924 27124 21980
rect 27180 21924 27190 21980
rect 35474 21924 35484 21980
rect 35540 21924 35588 21980
rect 35644 21924 35692 21980
rect 35748 21924 35758 21980
rect 11890 21868 11900 21924
rect 11956 21868 13356 21924
rect 13412 21868 13422 21924
rect 33282 21868 33292 21924
rect 33348 21868 34412 21924
rect 34468 21868 34478 21924
rect 10434 21756 10444 21812
rect 10500 21756 12908 21812
rect 12964 21756 12974 21812
rect 14466 21756 14476 21812
rect 14532 21756 15484 21812
rect 15540 21756 15550 21812
rect 18722 21756 18732 21812
rect 18788 21756 21084 21812
rect 21140 21756 21150 21812
rect 23650 21756 23660 21812
rect 23716 21756 25340 21812
rect 25396 21756 25406 21812
rect 27458 21756 27468 21812
rect 27524 21756 35196 21812
rect 35252 21756 35262 21812
rect 11900 21644 15372 21700
rect 15428 21644 15438 21700
rect 15810 21644 15820 21700
rect 15876 21644 19180 21700
rect 19236 21644 19246 21700
rect 24770 21644 24780 21700
rect 24836 21644 26684 21700
rect 26740 21644 26750 21700
rect 29250 21644 29260 21700
rect 29316 21644 29932 21700
rect 29988 21644 31052 21700
rect 31108 21644 31118 21700
rect 32050 21644 32060 21700
rect 32116 21644 34076 21700
rect 34132 21644 34142 21700
rect 11900 21588 11956 21644
rect 8418 21532 8428 21588
rect 8484 21532 10332 21588
rect 10388 21532 10398 21588
rect 10770 21532 10780 21588
rect 10836 21532 11956 21588
rect 27458 21532 27468 21588
rect 27524 21532 30044 21588
rect 30100 21532 30110 21588
rect 30482 21532 30492 21588
rect 30548 21532 31164 21588
rect 31220 21532 31230 21588
rect 32162 21532 32172 21588
rect 32228 21532 33628 21588
rect 33684 21532 35084 21588
rect 35140 21532 35150 21588
rect 6514 21420 6524 21476
rect 6580 21420 7196 21476
rect 7252 21420 7262 21476
rect 7522 21420 7532 21476
rect 7588 21420 8876 21476
rect 8932 21420 10892 21476
rect 10948 21420 10958 21476
rect 14690 21420 14700 21476
rect 14756 21420 16604 21476
rect 16660 21420 16670 21476
rect 17826 21420 17836 21476
rect 17892 21420 19404 21476
rect 19460 21420 19470 21476
rect 20738 21420 20748 21476
rect 20804 21420 21868 21476
rect 21924 21420 22876 21476
rect 22932 21420 24220 21476
rect 24276 21420 26236 21476
rect 26292 21420 26302 21476
rect 26646 21420 26684 21476
rect 26740 21420 26750 21476
rect 27010 21420 27020 21476
rect 27076 21420 30380 21476
rect 30436 21420 30446 21476
rect 31826 21420 31836 21476
rect 31892 21420 33964 21476
rect 34020 21420 34030 21476
rect 9314 21308 9324 21364
rect 9380 21308 15260 21364
rect 15316 21308 15326 21364
rect 17042 21308 17052 21364
rect 17108 21308 17948 21364
rect 18004 21308 18014 21364
rect 22530 21308 22540 21364
rect 22596 21308 30940 21364
rect 30996 21308 32228 21364
rect 32498 21308 32508 21364
rect 32564 21308 34076 21364
rect 34132 21308 34142 21364
rect 32172 21252 32228 21308
rect 23986 21196 23996 21252
rect 24052 21196 28812 21252
rect 28868 21196 28878 21252
rect 32172 21196 32396 21252
rect 32452 21196 32462 21252
rect 5486 21140 5496 21196
rect 5552 21140 5600 21196
rect 5656 21140 5704 21196
rect 5760 21140 5770 21196
rect 14054 21140 14064 21196
rect 14120 21140 14168 21196
rect 14224 21140 14272 21196
rect 14328 21140 14338 21196
rect 22622 21140 22632 21196
rect 22688 21140 22736 21196
rect 22792 21140 22840 21196
rect 22896 21140 22906 21196
rect 31190 21140 31200 21196
rect 31256 21140 31304 21196
rect 31360 21140 31408 21196
rect 31464 21140 31474 21196
rect 36200 21140 37000 21168
rect 26852 21084 28476 21140
rect 28532 21084 28542 21140
rect 32834 21084 32844 21140
rect 32900 21084 37000 21140
rect 26852 20916 26908 21084
rect 36200 21056 37000 21084
rect 27570 20972 27580 21028
rect 27636 20972 28252 21028
rect 28308 20972 28318 21028
rect 34738 20972 34748 21028
rect 34804 20972 35980 21028
rect 36036 20972 36046 21028
rect 10892 20860 11564 20916
rect 11620 20860 11630 20916
rect 22754 20860 22764 20916
rect 22820 20860 23996 20916
rect 24052 20860 24062 20916
rect 25218 20860 25228 20916
rect 25284 20860 26908 20916
rect 8530 20748 8540 20804
rect 8596 20748 9324 20804
rect 9380 20748 9390 20804
rect 10892 20692 10948 20860
rect 13234 20748 13244 20804
rect 13300 20748 13804 20804
rect 13860 20748 14588 20804
rect 14644 20748 14654 20804
rect 23492 20748 26796 20804
rect 26852 20748 26862 20804
rect 28242 20748 28252 20804
rect 28308 20748 32284 20804
rect 32340 20748 32350 20804
rect 8754 20636 8764 20692
rect 8820 20636 9548 20692
rect 9604 20636 10948 20692
rect 14914 20636 14924 20692
rect 14980 20636 15708 20692
rect 15764 20636 16940 20692
rect 16996 20636 17836 20692
rect 17892 20636 17902 20692
rect 18050 20636 18060 20692
rect 18116 20636 18620 20692
rect 18676 20636 18686 20692
rect 6514 20524 6524 20580
rect 6580 20524 7420 20580
rect 7476 20524 7486 20580
rect 10892 20468 10948 20636
rect 23492 20580 23548 20748
rect 24434 20636 24444 20692
rect 24500 20636 27356 20692
rect 27412 20636 28588 20692
rect 28644 20636 28654 20692
rect 28802 20636 28812 20692
rect 28868 20636 29148 20692
rect 29204 20636 30268 20692
rect 30324 20636 30334 20692
rect 18274 20524 18284 20580
rect 18340 20524 19964 20580
rect 20020 20524 20030 20580
rect 22866 20524 22876 20580
rect 22932 20524 23548 20580
rect 27570 20524 27580 20580
rect 27636 20524 32396 20580
rect 32452 20524 32462 20580
rect 10882 20412 10892 20468
rect 10948 20412 10958 20468
rect 11442 20412 11452 20468
rect 11508 20412 12236 20468
rect 12292 20412 12302 20468
rect 18834 20412 18844 20468
rect 18900 20412 19404 20468
rect 19460 20412 19470 20468
rect 9770 20356 9780 20412
rect 9836 20356 9884 20412
rect 9940 20356 9988 20412
rect 10044 20356 10054 20412
rect 18338 20356 18348 20412
rect 18404 20356 18452 20412
rect 18508 20356 18556 20412
rect 18612 20356 18622 20412
rect 26906 20356 26916 20412
rect 26972 20356 27020 20412
rect 27076 20356 27124 20412
rect 27180 20356 27190 20412
rect 35474 20356 35484 20412
rect 35540 20356 35588 20412
rect 35644 20356 35692 20412
rect 35748 20356 35758 20412
rect 20738 20300 20748 20356
rect 20804 20300 26684 20356
rect 26740 20300 26750 20356
rect 3714 20188 3724 20244
rect 3780 20188 5068 20244
rect 5124 20188 6300 20244
rect 6356 20188 6366 20244
rect 7858 20188 7868 20244
rect 7924 20188 8204 20244
rect 8260 20188 10332 20244
rect 10388 20188 10398 20244
rect 12898 20188 12908 20244
rect 12964 20188 13468 20244
rect 13524 20188 13534 20244
rect 15250 20188 15260 20244
rect 15316 20188 21420 20244
rect 21476 20188 23548 20244
rect 23604 20188 23614 20244
rect 26226 20188 26236 20244
rect 26292 20188 27132 20244
rect 27188 20188 27198 20244
rect 27794 20188 27804 20244
rect 27860 20188 28588 20244
rect 28644 20188 29372 20244
rect 29428 20188 29438 20244
rect 7970 20076 7980 20132
rect 8036 20076 9772 20132
rect 9828 20076 9838 20132
rect 16146 20076 16156 20132
rect 16212 20076 16604 20132
rect 16660 20076 17388 20132
rect 17444 20076 18284 20132
rect 18340 20076 19068 20132
rect 19124 20076 19134 20132
rect 24994 20076 25004 20132
rect 25060 20076 25900 20132
rect 25956 20076 26236 20132
rect 26292 20076 26302 20132
rect 28242 20076 28252 20132
rect 28308 20076 31612 20132
rect 31668 20076 31678 20132
rect 33058 20076 33068 20132
rect 33124 20076 34412 20132
rect 34468 20076 34478 20132
rect 8530 19964 8540 20020
rect 8596 19964 9436 20020
rect 9492 19964 9502 20020
rect 11218 19964 11228 20020
rect 11284 19964 12572 20020
rect 12628 19964 12638 20020
rect 15922 19964 15932 20020
rect 15988 19964 16716 20020
rect 16772 19964 16782 20020
rect 27346 19964 27356 20020
rect 27412 19964 29484 20020
rect 29540 19964 30492 20020
rect 30548 19964 30558 20020
rect 31826 19964 31836 20020
rect 31892 19964 35084 20020
rect 35140 19964 35150 20020
rect 5730 19852 5740 19908
rect 5796 19852 8652 19908
rect 8708 19852 8718 19908
rect 10210 19852 10220 19908
rect 10276 19852 12796 19908
rect 12852 19852 12862 19908
rect 20626 19852 20636 19908
rect 20692 19852 22092 19908
rect 22148 19852 22158 19908
rect 22978 19852 22988 19908
rect 23044 19852 23660 19908
rect 23716 19852 23726 19908
rect 25778 19852 25788 19908
rect 25844 19852 26572 19908
rect 26628 19852 26638 19908
rect 6850 19740 6860 19796
rect 6916 19740 7868 19796
rect 7924 19740 8428 19796
rect 8484 19740 9660 19796
rect 9716 19740 9726 19796
rect 10994 19740 11004 19796
rect 11060 19740 12348 19796
rect 12404 19740 14700 19796
rect 14756 19740 14766 19796
rect 25526 19740 25564 19796
rect 25620 19740 25630 19796
rect 25788 19740 26684 19796
rect 26740 19740 28364 19796
rect 28420 19740 29260 19796
rect 29316 19740 29326 19796
rect 31052 19740 32284 19796
rect 32340 19740 33852 19796
rect 33908 19740 33918 19796
rect 25788 19684 25844 19740
rect 25778 19628 25788 19684
rect 25844 19628 25854 19684
rect 26786 19628 26796 19684
rect 26852 19628 29148 19684
rect 29204 19628 30156 19684
rect 30212 19628 30222 19684
rect 5486 19572 5496 19628
rect 5552 19572 5600 19628
rect 5656 19572 5704 19628
rect 5760 19572 5770 19628
rect 14054 19572 14064 19628
rect 14120 19572 14168 19628
rect 14224 19572 14272 19628
rect 14328 19572 14338 19628
rect 22622 19572 22632 19628
rect 22688 19572 22736 19628
rect 22792 19572 22840 19628
rect 22896 19572 22906 19628
rect 31052 19572 31108 19740
rect 31190 19572 31200 19628
rect 31256 19572 31304 19628
rect 31360 19572 31408 19628
rect 31464 19572 31474 19628
rect 25218 19516 25228 19572
rect 25284 19516 26012 19572
rect 26068 19516 26078 19572
rect 26852 19516 31108 19572
rect 26852 19460 26908 19516
rect 13682 19404 13692 19460
rect 13748 19404 14812 19460
rect 14868 19404 14878 19460
rect 15922 19404 15932 19460
rect 15988 19404 16268 19460
rect 16324 19404 19404 19460
rect 19460 19404 24892 19460
rect 24948 19404 24958 19460
rect 25330 19404 25340 19460
rect 25396 19404 26908 19460
rect 27570 19404 27580 19460
rect 27636 19404 28028 19460
rect 28084 19404 29260 19460
rect 29316 19404 29708 19460
rect 29764 19404 29774 19460
rect 30146 19404 30156 19460
rect 30212 19404 34300 19460
rect 34356 19404 34366 19460
rect 34626 19404 34636 19460
rect 34692 19404 34702 19460
rect 29708 19348 29764 19404
rect 7522 19292 7532 19348
rect 7588 19292 8540 19348
rect 8596 19292 8988 19348
rect 9044 19292 9054 19348
rect 10994 19292 11004 19348
rect 11060 19292 25228 19348
rect 25284 19292 27020 19348
rect 27076 19292 27086 19348
rect 28242 19292 28252 19348
rect 28308 19292 28364 19348
rect 28420 19292 28430 19348
rect 29708 19292 30268 19348
rect 30324 19292 30334 19348
rect 30594 19292 30604 19348
rect 30660 19292 32284 19348
rect 32340 19292 32350 19348
rect 12674 19180 12684 19236
rect 12740 19180 13468 19236
rect 13524 19180 14140 19236
rect 14196 19180 14206 19236
rect 15026 19180 15036 19236
rect 15092 19180 15932 19236
rect 15988 19180 15998 19236
rect 20514 19180 20524 19236
rect 20580 19180 21756 19236
rect 21812 19180 21822 19236
rect 26012 19180 28700 19236
rect 28756 19180 29484 19236
rect 29540 19180 29550 19236
rect 30034 19180 30044 19236
rect 30100 19180 30716 19236
rect 30772 19180 30782 19236
rect 12786 19068 12796 19124
rect 12852 19068 13692 19124
rect 13748 19068 13758 19124
rect 16492 19068 24780 19124
rect 24836 19068 24846 19124
rect 9770 18788 9780 18844
rect 9836 18788 9884 18844
rect 9940 18788 9988 18844
rect 10044 18788 10054 18844
rect 13020 18788 13076 19068
rect 16492 19012 16548 19068
rect 14690 18956 14700 19012
rect 14756 18956 15148 19012
rect 15204 18956 15214 19012
rect 16370 18956 16380 19012
rect 16436 18956 16548 19012
rect 18722 18956 18732 19012
rect 18788 18956 22652 19012
rect 22708 18956 22718 19012
rect 23202 18956 23212 19012
rect 23268 18956 24108 19012
rect 24164 18956 25228 19012
rect 25284 18956 25294 19012
rect 26012 18900 26068 19180
rect 34636 19124 34692 19404
rect 26562 19068 26572 19124
rect 26628 19068 29372 19124
rect 29428 19068 29438 19124
rect 29922 19068 29932 19124
rect 29988 19068 31052 19124
rect 31108 19068 34692 19124
rect 26572 18956 28028 19012
rect 28084 18956 28094 19012
rect 28578 18956 28588 19012
rect 28644 18956 33852 19012
rect 33908 18956 35084 19012
rect 35140 18956 35150 19012
rect 26572 18900 26628 18956
rect 13794 18844 13804 18900
rect 13860 18844 14588 18900
rect 14644 18844 14924 18900
rect 14980 18844 14990 18900
rect 26002 18844 26012 18900
rect 26068 18844 26078 18900
rect 26338 18844 26348 18900
rect 26404 18844 26628 18900
rect 18338 18788 18348 18844
rect 18404 18788 18452 18844
rect 18508 18788 18556 18844
rect 18612 18788 18622 18844
rect 26906 18788 26916 18844
rect 26972 18788 27020 18844
rect 27076 18788 27124 18844
rect 27180 18788 27190 18844
rect 35474 18788 35484 18844
rect 35540 18788 35588 18844
rect 35644 18788 35692 18844
rect 35748 18788 35758 18844
rect 6962 18732 6972 18788
rect 7028 18732 8204 18788
rect 8260 18732 9100 18788
rect 9156 18732 9166 18788
rect 13010 18732 13020 18788
rect 13076 18732 13086 18788
rect 22418 18732 22428 18788
rect 22484 18732 24668 18788
rect 24724 18732 26404 18788
rect 28018 18732 28028 18788
rect 28084 18732 31500 18788
rect 31556 18732 31566 18788
rect 7298 18620 7308 18676
rect 7364 18620 7868 18676
rect 7924 18620 7934 18676
rect 24546 18620 24556 18676
rect 24612 18620 26124 18676
rect 26180 18620 26190 18676
rect 26348 18564 26404 18732
rect 26562 18620 26572 18676
rect 26628 18620 30044 18676
rect 30100 18620 30110 18676
rect 6066 18508 6076 18564
rect 6132 18508 6804 18564
rect 7410 18508 7420 18564
rect 7476 18508 7980 18564
rect 8036 18508 8046 18564
rect 12674 18508 12684 18564
rect 12740 18508 13468 18564
rect 13524 18508 13534 18564
rect 21634 18508 21644 18564
rect 21700 18508 26012 18564
rect 26068 18508 26078 18564
rect 26348 18508 27916 18564
rect 27972 18508 27982 18564
rect 28914 18508 28924 18564
rect 28980 18508 30604 18564
rect 30660 18508 30670 18564
rect 31910 18508 31948 18564
rect 32004 18508 32014 18564
rect 6748 18452 6804 18508
rect 36200 18452 37000 18480
rect 6748 18396 7308 18452
rect 7364 18396 8876 18452
rect 8932 18396 9548 18452
rect 9604 18396 10556 18452
rect 10612 18396 13580 18452
rect 13636 18396 13646 18452
rect 16258 18396 16268 18452
rect 16324 18396 17612 18452
rect 17668 18396 17678 18452
rect 23202 18396 23212 18452
rect 23268 18396 25340 18452
rect 25396 18396 25406 18452
rect 25554 18396 25564 18452
rect 25620 18396 26124 18452
rect 26180 18396 26190 18452
rect 26562 18396 26572 18452
rect 26628 18396 27020 18452
rect 27076 18396 27086 18452
rect 27318 18396 27356 18452
rect 27412 18396 27422 18452
rect 27570 18396 27580 18452
rect 27636 18396 27674 18452
rect 31826 18396 31836 18452
rect 31892 18396 34076 18452
rect 34132 18396 34142 18452
rect 35298 18396 35308 18452
rect 35364 18396 37000 18452
rect 27580 18340 27636 18396
rect 36200 18368 37000 18396
rect 8082 18284 8092 18340
rect 8148 18284 10220 18340
rect 10276 18284 10286 18340
rect 10434 18284 10444 18340
rect 10500 18284 13132 18340
rect 13188 18284 13198 18340
rect 15586 18284 15596 18340
rect 15652 18284 17836 18340
rect 17892 18284 17902 18340
rect 20850 18284 20860 18340
rect 20916 18284 21644 18340
rect 21700 18284 21710 18340
rect 23650 18284 23660 18340
rect 23716 18284 24220 18340
rect 24276 18284 27636 18340
rect 27692 18284 33516 18340
rect 33572 18284 33582 18340
rect 27692 18228 27748 18284
rect 25218 18172 25228 18228
rect 25284 18172 27132 18228
rect 27188 18172 27356 18228
rect 27412 18172 27748 18228
rect 28102 18172 28140 18228
rect 28196 18172 28206 18228
rect 30818 18172 30828 18228
rect 30884 18172 34860 18228
rect 34916 18172 34926 18228
rect 15586 18060 15596 18116
rect 15652 18060 18060 18116
rect 18116 18060 18844 18116
rect 18900 18060 19404 18116
rect 19460 18060 20748 18116
rect 20804 18060 21420 18116
rect 21476 18060 21486 18116
rect 26338 18060 26348 18116
rect 26404 18060 30156 18116
rect 30212 18060 30222 18116
rect 33394 18060 33404 18116
rect 33460 18060 34076 18116
rect 34132 18060 34636 18116
rect 34692 18060 34702 18116
rect 5486 18004 5496 18060
rect 5552 18004 5600 18060
rect 5656 18004 5704 18060
rect 5760 18004 5770 18060
rect 14054 18004 14064 18060
rect 14120 18004 14168 18060
rect 14224 18004 14272 18060
rect 14328 18004 14338 18060
rect 22622 18004 22632 18060
rect 22688 18004 22736 18060
rect 22792 18004 22840 18060
rect 22896 18004 22906 18060
rect 31190 18004 31200 18060
rect 31256 18004 31304 18060
rect 31360 18004 31408 18060
rect 31464 18004 31474 18060
rect 22978 17948 22988 18004
rect 23044 17948 25340 18004
rect 25396 17948 29820 18004
rect 29876 17948 29886 18004
rect 32470 17948 32508 18004
rect 32564 17948 32574 18004
rect 8978 17836 8988 17892
rect 9044 17836 9884 17892
rect 9940 17836 17724 17892
rect 17780 17836 23548 17892
rect 23604 17836 23614 17892
rect 26786 17836 26796 17892
rect 26852 17836 28028 17892
rect 28084 17836 28094 17892
rect 28690 17836 28700 17892
rect 28756 17836 29036 17892
rect 29092 17836 29102 17892
rect 30930 17836 30940 17892
rect 30996 17836 32172 17892
rect 32228 17836 33180 17892
rect 33236 17836 33246 17892
rect 15250 17724 15260 17780
rect 15316 17724 16156 17780
rect 16212 17724 17052 17780
rect 17108 17724 17118 17780
rect 25778 17724 25788 17780
rect 25844 17724 26348 17780
rect 26404 17724 26414 17780
rect 30370 17724 30380 17780
rect 30436 17724 31276 17780
rect 31332 17724 31342 17780
rect 12898 17612 12908 17668
rect 12964 17612 14028 17668
rect 14084 17612 14094 17668
rect 18274 17612 18284 17668
rect 18340 17612 19292 17668
rect 19348 17612 19628 17668
rect 19684 17612 20076 17668
rect 20132 17612 20142 17668
rect 21970 17612 21980 17668
rect 22036 17612 22988 17668
rect 23044 17612 23054 17668
rect 24322 17612 24332 17668
rect 24388 17612 25676 17668
rect 25732 17612 25742 17668
rect 28578 17612 28588 17668
rect 28644 17612 33404 17668
rect 33460 17612 33470 17668
rect 18284 17556 18340 17612
rect 13794 17500 13804 17556
rect 13860 17500 14252 17556
rect 14308 17500 14318 17556
rect 17826 17500 17836 17556
rect 17892 17500 18340 17556
rect 18610 17500 18620 17556
rect 18676 17500 19068 17556
rect 19124 17500 22428 17556
rect 22484 17500 22494 17556
rect 22642 17500 22652 17556
rect 22708 17500 25004 17556
rect 25060 17500 26012 17556
rect 26068 17500 26078 17556
rect 27570 17500 27580 17556
rect 27636 17500 30156 17556
rect 30212 17500 30222 17556
rect 33618 17500 33628 17556
rect 33684 17500 34412 17556
rect 34468 17500 34478 17556
rect 10882 17388 10892 17444
rect 10948 17388 12460 17444
rect 12516 17388 12526 17444
rect 17714 17388 17724 17444
rect 17780 17388 19516 17444
rect 19572 17388 23996 17444
rect 24052 17388 25452 17444
rect 25508 17388 25518 17444
rect 26674 17388 26684 17444
rect 26740 17388 27468 17444
rect 27524 17388 27534 17444
rect 28018 17388 28028 17444
rect 28084 17388 28476 17444
rect 28532 17388 31724 17444
rect 31780 17388 32620 17444
rect 32676 17388 32686 17444
rect 29138 17276 29148 17332
rect 29204 17276 33516 17332
rect 33572 17276 33964 17332
rect 34020 17276 34030 17332
rect 35046 17276 35084 17332
rect 35140 17276 35150 17332
rect 9770 17220 9780 17276
rect 9836 17220 9884 17276
rect 9940 17220 9988 17276
rect 10044 17220 10054 17276
rect 18338 17220 18348 17276
rect 18404 17220 18452 17276
rect 18508 17220 18556 17276
rect 18612 17220 18622 17276
rect 26906 17220 26916 17276
rect 26972 17220 27020 17276
rect 27076 17220 27124 17276
rect 27180 17220 27190 17276
rect 35474 17220 35484 17276
rect 35540 17220 35588 17276
rect 35644 17220 35692 17276
rect 35748 17220 35758 17276
rect 20850 17164 20860 17220
rect 20916 17164 25620 17220
rect 30706 17164 30716 17220
rect 30772 17164 34972 17220
rect 35028 17164 35038 17220
rect 25564 17108 25620 17164
rect 10322 17052 10332 17108
rect 10388 17052 10780 17108
rect 10836 17052 12796 17108
rect 12852 17052 12862 17108
rect 16818 17052 16828 17108
rect 16884 17052 17836 17108
rect 17892 17052 17902 17108
rect 18834 17052 18844 17108
rect 18900 17052 19292 17108
rect 19348 17052 19358 17108
rect 19842 17052 19852 17108
rect 19908 17052 24444 17108
rect 24500 17052 24510 17108
rect 25554 17052 25564 17108
rect 25620 17052 25630 17108
rect 26226 17052 26236 17108
rect 26292 17052 27356 17108
rect 27412 17052 27422 17108
rect 12674 16940 12684 16996
rect 12740 16940 13580 16996
rect 13636 16940 13646 16996
rect 19394 16940 19404 16996
rect 19460 16940 21980 16996
rect 22036 16940 22046 16996
rect 22306 16940 22316 16996
rect 22372 16940 25228 16996
rect 25284 16940 25294 16996
rect 25778 16940 25788 16996
rect 25844 16940 26684 16996
rect 26740 16940 28364 16996
rect 28420 16940 28430 16996
rect 9762 16828 9772 16884
rect 9828 16828 10444 16884
rect 10500 16828 10510 16884
rect 12002 16828 12012 16884
rect 12068 16828 13244 16884
rect 13300 16828 13916 16884
rect 13972 16828 15260 16884
rect 15316 16828 15326 16884
rect 20626 16828 20636 16884
rect 20692 16828 22204 16884
rect 22260 16828 22270 16884
rect 22530 16828 22540 16884
rect 22596 16828 23436 16884
rect 23492 16828 23502 16884
rect 26002 16828 26012 16884
rect 26068 16828 32396 16884
rect 32452 16828 32462 16884
rect 12012 16772 12068 16828
rect 10098 16716 10108 16772
rect 10164 16716 12068 16772
rect 21186 16716 21196 16772
rect 21252 16716 25788 16772
rect 25844 16716 25854 16772
rect 26674 16716 26684 16772
rect 26740 16716 27692 16772
rect 27748 16716 28028 16772
rect 28084 16716 30716 16772
rect 30772 16716 30782 16772
rect 30930 16716 30940 16772
rect 30996 16716 34188 16772
rect 34244 16716 34254 16772
rect 33852 16660 33908 16716
rect 8306 16604 8316 16660
rect 8372 16604 11004 16660
rect 11060 16604 11070 16660
rect 20290 16604 20300 16660
rect 20356 16604 26572 16660
rect 26628 16604 26638 16660
rect 26786 16604 26796 16660
rect 26852 16604 27244 16660
rect 27300 16604 27310 16660
rect 28466 16604 28476 16660
rect 28532 16604 32172 16660
rect 32228 16604 32238 16660
rect 33842 16604 33852 16660
rect 33908 16604 33918 16660
rect 20402 16492 20412 16548
rect 20468 16492 21420 16548
rect 21476 16492 21486 16548
rect 28018 16492 28028 16548
rect 28084 16492 30380 16548
rect 30436 16492 30446 16548
rect 5486 16436 5496 16492
rect 5552 16436 5600 16492
rect 5656 16436 5704 16492
rect 5760 16436 5770 16492
rect 14054 16436 14064 16492
rect 14120 16436 14168 16492
rect 14224 16436 14272 16492
rect 14328 16436 14338 16492
rect 22622 16436 22632 16492
rect 22688 16436 22736 16492
rect 22792 16436 22840 16492
rect 22896 16436 22906 16492
rect 31190 16436 31200 16492
rect 31256 16436 31304 16492
rect 31360 16436 31408 16492
rect 31464 16436 31474 16492
rect 18162 16380 18172 16436
rect 18228 16380 19628 16436
rect 19684 16380 19694 16436
rect 25330 16380 25340 16436
rect 25396 16380 25900 16436
rect 25956 16380 25966 16436
rect 28466 16380 28476 16436
rect 28532 16380 29484 16436
rect 29540 16380 29550 16436
rect 13794 16268 13804 16324
rect 13860 16268 15260 16324
rect 15316 16268 15326 16324
rect 18050 16268 18060 16324
rect 18116 16268 27468 16324
rect 27524 16268 28364 16324
rect 28420 16268 28430 16324
rect 29138 16268 29148 16324
rect 29204 16268 30044 16324
rect 30100 16268 30110 16324
rect 9202 16156 9212 16212
rect 9268 16156 11676 16212
rect 11732 16156 11742 16212
rect 15362 16156 15372 16212
rect 15428 16156 18732 16212
rect 18788 16156 18798 16212
rect 22082 16156 22092 16212
rect 22148 16156 25900 16212
rect 25956 16156 25966 16212
rect 28578 16156 28588 16212
rect 28644 16156 29260 16212
rect 29316 16156 29326 16212
rect 20738 16044 20748 16100
rect 20804 16044 21756 16100
rect 21812 16044 23884 16100
rect 23940 16044 23950 16100
rect 24210 16044 24220 16100
rect 24276 16044 25452 16100
rect 25508 16044 32732 16100
rect 32788 16044 32798 16100
rect 35186 16044 35196 16100
rect 35252 16044 35868 16100
rect 35924 16044 35934 16100
rect 23426 15932 23436 15988
rect 23492 15932 24556 15988
rect 24612 15932 24622 15988
rect 26898 15932 26908 15988
rect 26964 15932 28588 15988
rect 28644 15932 28654 15988
rect 31714 15932 31724 15988
rect 31780 15932 33292 15988
rect 33348 15932 33358 15988
rect 33954 15932 33964 15988
rect 34020 15932 35084 15988
rect 35140 15932 35150 15988
rect 19730 15820 19740 15876
rect 19796 15820 24668 15876
rect 24724 15820 25676 15876
rect 25732 15820 25742 15876
rect 26674 15820 26684 15876
rect 26740 15820 26796 15876
rect 26852 15820 26862 15876
rect 27010 15820 27020 15876
rect 27076 15820 27692 15876
rect 27748 15820 27758 15876
rect 28690 15820 28700 15876
rect 28756 15820 29372 15876
rect 29428 15820 29438 15876
rect 9770 15652 9780 15708
rect 9836 15652 9884 15708
rect 9940 15652 9988 15708
rect 10044 15652 10054 15708
rect 18338 15652 18348 15708
rect 18404 15652 18452 15708
rect 18508 15652 18556 15708
rect 18612 15652 18622 15708
rect 25676 15540 25732 15820
rect 33292 15764 33348 15932
rect 33842 15820 33852 15876
rect 33908 15820 34636 15876
rect 34692 15820 34702 15876
rect 36200 15764 37000 15792
rect 33292 15708 33740 15764
rect 33796 15708 33806 15764
rect 35868 15708 37000 15764
rect 26906 15652 26916 15708
rect 26972 15652 27020 15708
rect 27076 15652 27124 15708
rect 27180 15652 27190 15708
rect 35474 15652 35484 15708
rect 35540 15652 35588 15708
rect 35644 15652 35692 15708
rect 35748 15652 35758 15708
rect 26114 15596 26124 15652
rect 26180 15596 26348 15652
rect 26404 15596 26414 15652
rect 35868 15540 35924 15708
rect 36200 15680 37000 15708
rect 13458 15484 13468 15540
rect 13524 15484 14812 15540
rect 14868 15484 14878 15540
rect 25676 15484 27468 15540
rect 27524 15484 27534 15540
rect 32610 15484 32620 15540
rect 32676 15484 34748 15540
rect 34804 15484 34814 15540
rect 34962 15484 34972 15540
rect 35028 15484 35084 15540
rect 35140 15484 35150 15540
rect 35298 15484 35308 15540
rect 35364 15484 35924 15540
rect 14130 15372 14140 15428
rect 14196 15372 15148 15428
rect 24434 15372 24444 15428
rect 24500 15372 33180 15428
rect 33236 15372 33246 15428
rect 15092 15316 15148 15372
rect 15092 15260 16716 15316
rect 16772 15260 16782 15316
rect 21746 15260 21756 15316
rect 21812 15260 25676 15316
rect 25732 15260 25742 15316
rect 25900 15260 27132 15316
rect 27188 15260 27198 15316
rect 27766 15260 27804 15316
rect 27860 15260 27870 15316
rect 28214 15260 28252 15316
rect 28308 15260 28318 15316
rect 25900 15204 25956 15260
rect 17042 15148 17052 15204
rect 17108 15148 25228 15204
rect 25284 15148 25294 15204
rect 25442 15148 25452 15204
rect 25508 15148 25564 15204
rect 25620 15148 25956 15204
rect 26338 15148 26348 15204
rect 26404 15148 27412 15204
rect 27356 15092 27412 15148
rect 32162 15092 32172 15148
rect 32228 15092 32238 15148
rect 14354 15036 14364 15092
rect 14420 15036 14644 15092
rect 16930 15036 16940 15092
rect 16996 15036 25116 15092
rect 25172 15036 25182 15092
rect 26562 15036 26572 15092
rect 26628 15036 26908 15092
rect 26964 15036 26974 15092
rect 27356 15036 28252 15092
rect 28308 15036 28476 15092
rect 28532 15036 28542 15092
rect 30482 15036 30492 15092
rect 30548 15036 31500 15092
rect 31556 15036 31566 15092
rect 14588 14980 14644 15036
rect 32172 14980 32228 15092
rect 32722 15036 32732 15092
rect 32788 15036 33516 15092
rect 33572 15036 33582 15092
rect 14588 14924 14812 14980
rect 14868 14924 14878 14980
rect 26852 14924 27356 14980
rect 27412 14924 27422 14980
rect 27570 14924 27580 14980
rect 27636 14924 28644 14980
rect 28914 14924 28924 14980
rect 28980 14924 30156 14980
rect 30212 14924 30222 14980
rect 32162 14924 32172 14980
rect 32228 14924 32238 14980
rect 5486 14868 5496 14924
rect 5552 14868 5600 14924
rect 5656 14868 5704 14924
rect 5760 14868 5770 14924
rect 14054 14868 14064 14924
rect 14120 14868 14168 14924
rect 14224 14868 14272 14924
rect 14328 14868 14338 14924
rect 22622 14868 22632 14924
rect 22688 14868 22736 14924
rect 22792 14868 22840 14924
rect 22896 14868 22906 14924
rect 26852 14756 26908 14924
rect 28588 14868 28644 14924
rect 31190 14868 31200 14924
rect 31256 14868 31304 14924
rect 31360 14868 31408 14924
rect 31464 14868 31474 14924
rect 27654 14812 27692 14868
rect 27748 14812 27758 14868
rect 28578 14812 28588 14868
rect 28644 14812 29372 14868
rect 29428 14812 29438 14868
rect 31938 14812 31948 14868
rect 32004 14812 32396 14868
rect 32452 14812 32462 14868
rect 32610 14812 32620 14868
rect 32676 14812 32686 14868
rect 32620 14756 32676 14812
rect 9202 14700 9212 14756
rect 9268 14700 16828 14756
rect 16884 14700 16894 14756
rect 20738 14700 20748 14756
rect 20804 14700 24108 14756
rect 24164 14700 24174 14756
rect 24332 14700 26908 14756
rect 27906 14700 27916 14756
rect 27972 14700 28812 14756
rect 28868 14700 28878 14756
rect 32162 14700 32172 14756
rect 32228 14700 32676 14756
rect 24332 14644 24388 14700
rect 11218 14588 11228 14644
rect 11284 14588 11788 14644
rect 11844 14588 16940 14644
rect 16996 14588 17006 14644
rect 19058 14588 19068 14644
rect 19124 14588 24388 14644
rect 24658 14588 24668 14644
rect 24724 14588 33236 14644
rect 25778 14476 25788 14532
rect 25844 14476 27580 14532
rect 27636 14476 27646 14532
rect 32050 14476 32060 14532
rect 32116 14476 32508 14532
rect 32564 14476 32574 14532
rect 33180 14420 33236 14588
rect 17938 14364 17948 14420
rect 18004 14364 19852 14420
rect 19908 14364 23492 14420
rect 23986 14364 23996 14420
rect 24052 14364 27916 14420
rect 27972 14364 27982 14420
rect 33170 14364 33180 14420
rect 33236 14364 33246 14420
rect 23436 14308 23492 14364
rect 19394 14252 19404 14308
rect 19460 14252 20412 14308
rect 20468 14252 20478 14308
rect 21410 14252 21420 14308
rect 21476 14252 23212 14308
rect 23268 14252 23278 14308
rect 23436 14252 27412 14308
rect 29922 14252 29932 14308
rect 29988 14252 31052 14308
rect 31108 14252 31836 14308
rect 31892 14252 31902 14308
rect 20066 14140 20076 14196
rect 20132 14140 22316 14196
rect 22372 14140 26348 14196
rect 26404 14140 26414 14196
rect 9770 14084 9780 14140
rect 9836 14084 9884 14140
rect 9940 14084 9988 14140
rect 10044 14084 10054 14140
rect 18338 14084 18348 14140
rect 18404 14084 18452 14140
rect 18508 14084 18556 14140
rect 18612 14084 18622 14140
rect 26906 14084 26916 14140
rect 26972 14084 27020 14140
rect 27076 14084 27124 14140
rect 27180 14084 27190 14140
rect 19506 14028 19516 14084
rect 19572 14028 20748 14084
rect 20804 14028 21980 14084
rect 22036 14028 22046 14084
rect 25890 14028 25900 14084
rect 25956 14028 26460 14084
rect 26516 14028 26526 14084
rect 16594 13916 16604 13972
rect 16660 13916 17388 13972
rect 17444 13916 17454 13972
rect 23314 13916 23324 13972
rect 23380 13916 25228 13972
rect 25284 13916 26684 13972
rect 26740 13916 26750 13972
rect 19954 13804 19964 13860
rect 20020 13804 25788 13860
rect 25844 13804 25854 13860
rect 27356 13748 27412 14252
rect 35474 14084 35484 14140
rect 35540 14084 35588 14140
rect 35644 14084 35692 14140
rect 35748 14084 35758 14140
rect 27570 13804 27580 13860
rect 27636 13804 28140 13860
rect 28196 13804 28252 13860
rect 28308 13804 28318 13860
rect 31602 13804 31612 13860
rect 31668 13804 34748 13860
rect 34804 13804 34814 13860
rect 6850 13692 6860 13748
rect 6916 13692 7868 13748
rect 7924 13692 7934 13748
rect 13804 13692 15596 13748
rect 15652 13692 16716 13748
rect 16772 13692 16782 13748
rect 27356 13692 29148 13748
rect 29204 13692 29214 13748
rect 13804 13636 13860 13692
rect 27580 13636 27636 13692
rect 13346 13580 13356 13636
rect 13412 13580 13804 13636
rect 13860 13580 13870 13636
rect 14690 13580 14700 13636
rect 14756 13580 15036 13636
rect 15092 13580 15372 13636
rect 15428 13580 16156 13636
rect 16212 13580 16222 13636
rect 16482 13580 16492 13636
rect 16548 13580 18620 13636
rect 18676 13580 21868 13636
rect 21924 13580 21934 13636
rect 27570 13580 27580 13636
rect 27636 13580 27646 13636
rect 29698 13580 29708 13636
rect 29764 13580 30940 13636
rect 30996 13580 33796 13636
rect 16492 13524 16548 13580
rect 33740 13524 33796 13580
rect 12898 13468 12908 13524
rect 12964 13468 16548 13524
rect 27122 13468 27132 13524
rect 27188 13468 31724 13524
rect 31780 13468 31790 13524
rect 32386 13468 32396 13524
rect 32452 13468 33516 13524
rect 33572 13468 33582 13524
rect 33730 13468 33740 13524
rect 33796 13468 35084 13524
rect 35140 13468 35150 13524
rect 23202 13356 23212 13412
rect 23268 13356 27244 13412
rect 27300 13356 27310 13412
rect 27458 13356 27468 13412
rect 27524 13356 27916 13412
rect 27972 13356 27982 13412
rect 5486 13300 5496 13356
rect 5552 13300 5600 13356
rect 5656 13300 5704 13356
rect 5760 13300 5770 13356
rect 14054 13300 14064 13356
rect 14120 13300 14168 13356
rect 14224 13300 14272 13356
rect 14328 13300 14338 13356
rect 22622 13300 22632 13356
rect 22688 13300 22736 13356
rect 22792 13300 22840 13356
rect 22896 13300 22906 13356
rect 31190 13300 31200 13356
rect 31256 13300 31304 13356
rect 31360 13300 31408 13356
rect 31464 13300 31474 13356
rect 8306 13244 8316 13300
rect 8372 13244 11340 13300
rect 11396 13244 11788 13300
rect 11844 13244 11854 13300
rect 23090 13244 23100 13300
rect 23156 13244 23996 13300
rect 24052 13244 24062 13300
rect 28578 13244 28588 13300
rect 28644 13244 29036 13300
rect 29092 13244 29102 13300
rect 7186 13132 7196 13188
rect 7252 13132 7262 13188
rect 7410 13132 7420 13188
rect 7476 13132 8540 13188
rect 8596 13132 8606 13188
rect 23202 13132 23212 13188
rect 23268 13132 24668 13188
rect 24724 13132 26684 13188
rect 26740 13132 26750 13188
rect 29138 13132 29148 13188
rect 29204 13132 31164 13188
rect 31220 13132 31230 13188
rect 32162 13132 32172 13188
rect 32228 13132 32238 13188
rect 7196 12852 7252 13132
rect 11554 13020 11564 13076
rect 11620 13020 12796 13076
rect 12852 13020 12862 13076
rect 24322 13020 24332 13076
rect 24388 13020 25452 13076
rect 25508 13020 25518 13076
rect 26338 13020 26348 13076
rect 26404 13020 26796 13076
rect 26852 13020 26862 13076
rect 28354 13020 28364 13076
rect 28420 13020 29708 13076
rect 29764 13020 31948 13076
rect 32004 13020 32014 13076
rect 8082 12908 8092 12964
rect 8148 12908 8876 12964
rect 8932 12908 8942 12964
rect 10322 12908 10332 12964
rect 10388 12908 12460 12964
rect 12516 12908 12526 12964
rect 22978 12908 22988 12964
rect 23044 12908 27804 12964
rect 27860 12908 27870 12964
rect 28130 12908 28140 12964
rect 28196 12908 30268 12964
rect 30324 12908 30334 12964
rect 32172 12852 32228 13132
rect 36200 13076 37000 13104
rect 33954 13020 33964 13076
rect 34020 13020 37000 13076
rect 36200 12992 37000 13020
rect 6962 12796 6972 12852
rect 7028 12796 8764 12852
rect 8820 12796 9996 12852
rect 10052 12796 10062 12852
rect 10770 12796 10780 12852
rect 10836 12796 12236 12852
rect 12292 12796 12302 12852
rect 27794 12796 27804 12852
rect 27860 12796 28364 12852
rect 28420 12796 28430 12852
rect 29484 12796 32228 12852
rect 34178 12796 34188 12852
rect 34244 12796 34412 12852
rect 34468 12796 34478 12852
rect 29484 12740 29540 12796
rect 7522 12684 7532 12740
rect 7588 12684 8428 12740
rect 8484 12684 10444 12740
rect 10500 12684 10510 12740
rect 18946 12684 18956 12740
rect 19012 12684 19516 12740
rect 19572 12684 19582 12740
rect 19730 12684 19740 12740
rect 19796 12684 20300 12740
rect 20356 12684 20366 12740
rect 25442 12684 25452 12740
rect 25508 12684 29540 12740
rect 29922 12684 29932 12740
rect 29988 12684 30940 12740
rect 30996 12684 31006 12740
rect 6290 12572 6300 12628
rect 6356 12572 8316 12628
rect 8372 12572 8382 12628
rect 10332 12572 11564 12628
rect 11620 12572 11630 12628
rect 22306 12572 22316 12628
rect 22372 12572 23212 12628
rect 23268 12572 23278 12628
rect 27458 12572 27468 12628
rect 27524 12572 31836 12628
rect 31892 12572 31902 12628
rect 9770 12516 9780 12572
rect 9836 12516 9884 12572
rect 9940 12516 9988 12572
rect 10044 12516 10054 12572
rect 6178 12460 6188 12516
rect 6244 12460 8428 12516
rect 8484 12460 8494 12516
rect 4834 12348 4844 12404
rect 4900 12348 7756 12404
rect 7812 12348 7822 12404
rect 10332 12180 10388 12572
rect 18338 12516 18348 12572
rect 18404 12516 18452 12572
rect 18508 12516 18556 12572
rect 18612 12516 18622 12572
rect 26906 12516 26916 12572
rect 26972 12516 27020 12572
rect 27076 12516 27124 12572
rect 27180 12516 27190 12572
rect 35474 12516 35484 12572
rect 35540 12516 35588 12572
rect 35644 12516 35692 12572
rect 35748 12516 35758 12572
rect 22530 12460 22540 12516
rect 22596 12460 24220 12516
rect 24276 12460 25620 12516
rect 25564 12404 25620 12460
rect 13570 12348 13580 12404
rect 13636 12348 15148 12404
rect 15204 12348 15214 12404
rect 16482 12348 16492 12404
rect 16548 12348 17164 12404
rect 17220 12348 20524 12404
rect 20580 12348 21196 12404
rect 21252 12348 21262 12404
rect 21746 12348 21756 12404
rect 21812 12348 23660 12404
rect 23716 12348 25340 12404
rect 25396 12348 25406 12404
rect 25564 12348 33180 12404
rect 33236 12348 33246 12404
rect 30370 12236 30380 12292
rect 30436 12236 34076 12292
rect 34132 12236 34142 12292
rect 7634 12124 7644 12180
rect 7700 12124 8540 12180
rect 8596 12124 9100 12180
rect 9156 12124 9166 12180
rect 10322 12124 10332 12180
rect 10388 12124 10398 12180
rect 12450 12124 12460 12180
rect 12516 12124 13916 12180
rect 13972 12124 17948 12180
rect 18004 12124 18014 12180
rect 24658 12124 24668 12180
rect 24724 12124 25900 12180
rect 25956 12124 27580 12180
rect 27636 12124 29036 12180
rect 29092 12124 29102 12180
rect 33618 12124 33628 12180
rect 33684 12124 34860 12180
rect 34916 12124 34926 12180
rect 10098 12012 10108 12068
rect 10164 12012 11564 12068
rect 11620 12012 11630 12068
rect 25890 11900 25900 11956
rect 25956 11900 26908 11956
rect 26964 11900 31724 11956
rect 31780 11900 31790 11956
rect 32498 11900 32508 11956
rect 32564 11900 33516 11956
rect 33572 11900 33582 11956
rect 15138 11788 15148 11844
rect 15204 11788 16156 11844
rect 16212 11788 16222 11844
rect 5486 11732 5496 11788
rect 5552 11732 5600 11788
rect 5656 11732 5704 11788
rect 5760 11732 5770 11788
rect 14054 11732 14064 11788
rect 14120 11732 14168 11788
rect 14224 11732 14272 11788
rect 14328 11732 14338 11788
rect 22622 11732 22632 11788
rect 22688 11732 22736 11788
rect 22792 11732 22840 11788
rect 22896 11732 22906 11788
rect 31190 11732 31200 11788
rect 31256 11732 31304 11788
rect 31360 11732 31408 11788
rect 31464 11732 31474 11788
rect 25666 11676 25676 11732
rect 25732 11676 28252 11732
rect 28308 11676 29148 11732
rect 29204 11676 29214 11732
rect 31938 11676 31948 11732
rect 32004 11676 32014 11732
rect 33506 11676 33516 11732
rect 33572 11676 34076 11732
rect 34132 11676 34636 11732
rect 34692 11676 34702 11732
rect 31948 11620 32004 11676
rect 7970 11564 7980 11620
rect 8036 11564 8988 11620
rect 9044 11564 9884 11620
rect 9940 11564 9950 11620
rect 20290 11564 20300 11620
rect 20356 11564 20972 11620
rect 21028 11564 23100 11620
rect 23156 11564 25564 11620
rect 25620 11564 25630 11620
rect 28466 11564 28476 11620
rect 28532 11564 32004 11620
rect 32386 11564 32396 11620
rect 32452 11564 32732 11620
rect 32788 11564 33572 11620
rect 33516 11508 33572 11564
rect 9762 11452 9772 11508
rect 9828 11452 10556 11508
rect 10612 11452 10622 11508
rect 15922 11452 15932 11508
rect 15988 11452 16828 11508
rect 16884 11452 19516 11508
rect 19572 11452 19582 11508
rect 19954 11452 19964 11508
rect 20020 11452 20636 11508
rect 20692 11452 20702 11508
rect 31042 11452 31052 11508
rect 31108 11452 32956 11508
rect 33012 11452 33022 11508
rect 33506 11452 33516 11508
rect 33572 11452 34188 11508
rect 34244 11452 34412 11508
rect 34468 11452 34478 11508
rect 34598 11452 34636 11508
rect 34692 11452 34702 11508
rect 10994 11340 11004 11396
rect 11060 11340 11452 11396
rect 11508 11340 11900 11396
rect 11956 11340 12796 11396
rect 12852 11340 31276 11396
rect 31332 11340 32284 11396
rect 32340 11340 32350 11396
rect 34962 11340 34972 11396
rect 35028 11340 35084 11396
rect 35140 11340 35150 11396
rect 9650 11228 9660 11284
rect 9716 11228 10668 11284
rect 10724 11228 10734 11284
rect 20188 11228 22764 11284
rect 22820 11228 22830 11284
rect 23202 11228 23212 11284
rect 23268 11228 23660 11284
rect 23716 11228 23726 11284
rect 20188 11172 20244 11228
rect 9426 11116 9436 11172
rect 9492 11116 10332 11172
rect 10388 11116 10398 11172
rect 15250 11116 15260 11172
rect 15316 11116 16156 11172
rect 16212 11116 20188 11172
rect 20244 11116 20254 11172
rect 20738 11116 20748 11172
rect 20804 11116 21868 11172
rect 21924 11116 21934 11172
rect 24994 11116 25004 11172
rect 25060 11116 25676 11172
rect 25732 11116 25742 11172
rect 22306 11004 22316 11060
rect 22372 11004 23772 11060
rect 23828 11004 24892 11060
rect 24948 11004 24958 11060
rect 9770 10948 9780 11004
rect 9836 10948 9884 11004
rect 9940 10948 9988 11004
rect 10044 10948 10054 11004
rect 18338 10948 18348 11004
rect 18404 10948 18452 11004
rect 18508 10948 18556 11004
rect 18612 10948 18622 11004
rect 26906 10948 26916 11004
rect 26972 10948 27020 11004
rect 27076 10948 27124 11004
rect 27180 10948 27190 11004
rect 35474 10948 35484 11004
rect 35540 10948 35588 11004
rect 35644 10948 35692 11004
rect 35748 10948 35758 11004
rect 20738 10892 20748 10948
rect 20804 10892 21644 10948
rect 21700 10892 21710 10948
rect 19282 10780 19292 10836
rect 19348 10780 21420 10836
rect 21476 10780 21486 10836
rect 22754 10780 22764 10836
rect 22820 10780 23324 10836
rect 23380 10780 23390 10836
rect 23538 10780 23548 10836
rect 23604 10780 32620 10836
rect 32676 10780 32686 10836
rect 20636 10724 20692 10780
rect 20626 10668 20636 10724
rect 20692 10668 20702 10724
rect 21074 10668 21084 10724
rect 21140 10668 22428 10724
rect 22484 10668 22494 10724
rect 25106 10668 25116 10724
rect 25172 10668 26908 10724
rect 26964 10668 28364 10724
rect 28420 10668 28430 10724
rect 29586 10668 29596 10724
rect 29652 10668 30828 10724
rect 30884 10668 30894 10724
rect 31826 10668 31836 10724
rect 31892 10668 35196 10724
rect 35252 10668 35262 10724
rect 15558 10556 15596 10612
rect 15652 10556 15662 10612
rect 20514 10556 20524 10612
rect 20580 10556 21532 10612
rect 21588 10556 21598 10612
rect 24210 10556 24220 10612
rect 24276 10556 25228 10612
rect 25284 10556 25294 10612
rect 34402 10556 34412 10612
rect 34468 10556 35084 10612
rect 35140 10556 35150 10612
rect 10882 10444 10892 10500
rect 10948 10444 13244 10500
rect 13300 10444 13310 10500
rect 14578 10444 14588 10500
rect 14644 10444 15708 10500
rect 15764 10444 15774 10500
rect 29810 10444 29820 10500
rect 29876 10444 30940 10500
rect 30996 10444 31006 10500
rect 36200 10388 37000 10416
rect 8418 10332 8428 10388
rect 8484 10332 9660 10388
rect 9716 10332 9726 10388
rect 16454 10332 16492 10388
rect 16548 10332 16558 10388
rect 16706 10332 16716 10388
rect 16772 10332 25060 10388
rect 33170 10332 33180 10388
rect 33236 10332 34188 10388
rect 34244 10332 37000 10388
rect 5486 10164 5496 10220
rect 5552 10164 5600 10220
rect 5656 10164 5704 10220
rect 5760 10164 5770 10220
rect 14054 10164 14064 10220
rect 14120 10164 14168 10220
rect 14224 10164 14272 10220
rect 14328 10164 14338 10220
rect 22622 10164 22632 10220
rect 22688 10164 22736 10220
rect 22792 10164 22840 10220
rect 22896 10164 22906 10220
rect 7634 10108 7644 10164
rect 7700 10108 9436 10164
rect 9492 10108 9502 10164
rect 23100 10108 24108 10164
rect 24164 10108 24174 10164
rect 23100 10052 23156 10108
rect 14466 9996 14476 10052
rect 14532 9996 15036 10052
rect 15092 9996 16940 10052
rect 16996 9996 17006 10052
rect 21410 9996 21420 10052
rect 21476 9996 22540 10052
rect 22596 9996 23156 10052
rect 25004 10052 25060 10332
rect 36200 10304 37000 10332
rect 31190 10164 31200 10220
rect 31256 10164 31304 10220
rect 31360 10164 31408 10220
rect 31464 10164 31474 10220
rect 25004 9996 25228 10052
rect 25284 9996 25294 10052
rect 6738 9884 6748 9940
rect 6804 9884 8204 9940
rect 8260 9884 8270 9940
rect 13122 9884 13132 9940
rect 13188 9884 14140 9940
rect 14196 9884 14206 9940
rect 12898 9772 12908 9828
rect 12964 9772 14924 9828
rect 14980 9772 16156 9828
rect 16212 9772 16222 9828
rect 20290 9772 20300 9828
rect 20356 9772 24556 9828
rect 24612 9772 24622 9828
rect 33954 9772 33964 9828
rect 34020 9772 35196 9828
rect 35252 9772 35262 9828
rect 28578 9660 28588 9716
rect 28644 9660 29932 9716
rect 29988 9660 30828 9716
rect 30884 9660 30894 9716
rect 12226 9548 12236 9604
rect 12292 9548 13580 9604
rect 13636 9548 13646 9604
rect 14690 9548 14700 9604
rect 14756 9548 15372 9604
rect 15428 9548 15438 9604
rect 15922 9548 15932 9604
rect 15988 9548 15998 9604
rect 28018 9548 28028 9604
rect 28084 9548 30716 9604
rect 30772 9548 30782 9604
rect 15932 9492 15988 9548
rect 14802 9436 14812 9492
rect 14868 9436 15988 9492
rect 29922 9436 29932 9492
rect 29988 9436 30604 9492
rect 30660 9436 30670 9492
rect 34402 9436 34412 9492
rect 34468 9436 34860 9492
rect 34916 9436 34926 9492
rect 9770 9380 9780 9436
rect 9836 9380 9884 9436
rect 9940 9380 9988 9436
rect 10044 9380 10054 9436
rect 18338 9380 18348 9436
rect 18404 9380 18452 9436
rect 18508 9380 18556 9436
rect 18612 9380 18622 9436
rect 26906 9380 26916 9436
rect 26972 9380 27020 9436
rect 27076 9380 27124 9436
rect 27180 9380 27190 9436
rect 35474 9380 35484 9436
rect 35540 9380 35588 9436
rect 35644 9380 35692 9436
rect 35748 9380 35758 9436
rect 15474 9212 15484 9268
rect 15540 9212 15596 9268
rect 15652 9212 16604 9268
rect 16660 9212 16670 9268
rect 25218 9212 25228 9268
rect 25284 9212 26012 9268
rect 26068 9212 26078 9268
rect 15810 9100 15820 9156
rect 15876 9100 17388 9156
rect 17444 9100 17836 9156
rect 17892 9100 18284 9156
rect 18340 9100 18350 9156
rect 19730 9100 19740 9156
rect 19796 9100 21532 9156
rect 21588 9100 21598 9156
rect 22764 9100 24108 9156
rect 24164 9100 24332 9156
rect 24388 9100 24398 9156
rect 24546 9100 24556 9156
rect 24612 9100 32396 9156
rect 32452 9100 33852 9156
rect 33908 9100 33918 9156
rect 22764 9044 22820 9100
rect 18610 8988 18620 9044
rect 18676 8988 20188 9044
rect 20244 8988 22764 9044
rect 22820 8988 22830 9044
rect 24210 8988 24220 9044
rect 24276 8988 27356 9044
rect 27412 8988 28812 9044
rect 28868 8988 30044 9044
rect 30100 8988 30110 9044
rect 30370 8988 30380 9044
rect 30436 8988 30716 9044
rect 30772 8988 31612 9044
rect 31668 8988 31678 9044
rect 7074 8876 7084 8932
rect 7140 8876 8540 8932
rect 8596 8876 12124 8932
rect 12180 8876 12190 8932
rect 13570 8876 13580 8932
rect 13636 8876 15708 8932
rect 15764 8876 17052 8932
rect 17108 8876 17118 8932
rect 15026 8764 15036 8820
rect 15092 8764 16380 8820
rect 16436 8764 17612 8820
rect 17668 8764 17678 8820
rect 23986 8764 23996 8820
rect 24052 8764 29372 8820
rect 29428 8764 29438 8820
rect 31154 8764 31164 8820
rect 31220 8764 32396 8820
rect 32452 8764 32462 8820
rect 5486 8596 5496 8652
rect 5552 8596 5600 8652
rect 5656 8596 5704 8652
rect 5760 8596 5770 8652
rect 14054 8596 14064 8652
rect 14120 8596 14168 8652
rect 14224 8596 14272 8652
rect 14328 8596 14338 8652
rect 22622 8596 22632 8652
rect 22688 8596 22736 8652
rect 22792 8596 22840 8652
rect 22896 8596 22906 8652
rect 31190 8596 31200 8652
rect 31256 8596 31304 8652
rect 31360 8596 31408 8652
rect 31464 8596 31474 8652
rect 4162 8428 4172 8484
rect 4228 8428 6748 8484
rect 6804 8428 7644 8484
rect 7700 8428 7710 8484
rect 13906 8428 13916 8484
rect 13972 8428 13982 8484
rect 14130 8428 14140 8484
rect 14196 8428 17500 8484
rect 17556 8428 17566 8484
rect 17714 8428 17724 8484
rect 17780 8428 23772 8484
rect 23828 8428 24444 8484
rect 24500 8428 24510 8484
rect 29474 8428 29484 8484
rect 29540 8428 34972 8484
rect 35028 8428 35038 8484
rect 9538 8316 9548 8372
rect 9604 8316 9772 8372
rect 9828 8316 9838 8372
rect 8082 8204 8092 8260
rect 8148 8204 9100 8260
rect 9156 8204 10332 8260
rect 10388 8204 10398 8260
rect 8540 8148 8596 8204
rect 13916 8148 13972 8428
rect 17938 8316 17948 8372
rect 18004 8316 19292 8372
rect 19348 8316 19358 8372
rect 30034 8316 30044 8372
rect 30100 8316 31276 8372
rect 31332 8316 31342 8372
rect 15250 8204 15260 8260
rect 15316 8204 16716 8260
rect 16772 8204 21308 8260
rect 21364 8204 21374 8260
rect 25778 8204 25788 8260
rect 25844 8204 26796 8260
rect 26852 8204 27300 8260
rect 29810 8204 29820 8260
rect 29876 8204 30716 8260
rect 30772 8204 34188 8260
rect 34244 8204 34254 8260
rect 27244 8148 27300 8204
rect 8530 8092 8540 8148
rect 8596 8092 8606 8148
rect 13916 8092 15708 8148
rect 15764 8092 15774 8148
rect 16258 8092 16268 8148
rect 16324 8092 20748 8148
rect 20804 8092 20814 8148
rect 26674 8092 26684 8148
rect 26740 8092 26908 8148
rect 27234 8092 27244 8148
rect 27300 8092 28028 8148
rect 28084 8092 28094 8148
rect 31154 8092 31164 8148
rect 31220 8092 32060 8148
rect 32116 8092 32126 8148
rect 26852 8036 26908 8092
rect 5954 7980 5964 8036
rect 6020 7980 9996 8036
rect 10052 7980 10062 8036
rect 12898 7980 12908 8036
rect 12964 7980 14252 8036
rect 14308 7980 14318 8036
rect 16482 7980 16492 8036
rect 16548 7980 26180 8036
rect 26852 7980 27916 8036
rect 27972 7980 27982 8036
rect 28354 7980 28364 8036
rect 28420 7980 29932 8036
rect 29988 7980 29998 8036
rect 30930 7980 30940 8036
rect 30996 7980 31612 8036
rect 31668 7980 31678 8036
rect 9770 7812 9780 7868
rect 9836 7812 9884 7868
rect 9940 7812 9988 7868
rect 10044 7812 10054 7868
rect 18338 7812 18348 7868
rect 18404 7812 18452 7868
rect 18508 7812 18556 7868
rect 18612 7812 18622 7868
rect 15092 7756 17388 7812
rect 17444 7756 17454 7812
rect 19404 7756 23884 7812
rect 23940 7756 25900 7812
rect 25956 7756 25966 7812
rect 9090 7644 9100 7700
rect 9156 7644 10780 7700
rect 10836 7644 12236 7700
rect 12292 7644 12302 7700
rect 7410 7532 7420 7588
rect 7476 7532 7980 7588
rect 8036 7532 8428 7588
rect 8484 7532 9548 7588
rect 9604 7532 9614 7588
rect 15092 7476 15148 7756
rect 19404 7700 19460 7756
rect 26124 7700 26180 7980
rect 27916 7924 27972 7980
rect 27916 7868 30492 7924
rect 30548 7868 32060 7924
rect 32116 7868 32126 7924
rect 26906 7812 26916 7868
rect 26972 7812 27020 7868
rect 27076 7812 27124 7868
rect 27180 7812 27190 7868
rect 35474 7812 35484 7868
rect 35540 7812 35588 7868
rect 35644 7812 35692 7868
rect 35748 7812 35758 7868
rect 36200 7700 37000 7728
rect 15250 7644 15260 7700
rect 15316 7644 15820 7700
rect 15876 7644 15886 7700
rect 18386 7644 18396 7700
rect 18452 7644 19460 7700
rect 19516 7644 20524 7700
rect 20580 7644 21084 7700
rect 21140 7644 21150 7700
rect 26124 7644 28924 7700
rect 28980 7644 28990 7700
rect 29362 7644 29372 7700
rect 29428 7644 32172 7700
rect 32228 7644 32238 7700
rect 35298 7644 35308 7700
rect 35364 7644 37000 7700
rect 19516 7588 19572 7644
rect 36200 7616 37000 7644
rect 18498 7532 18508 7588
rect 18564 7532 19516 7588
rect 19572 7532 19582 7588
rect 19842 7532 19852 7588
rect 19908 7532 20412 7588
rect 20468 7532 20478 7588
rect 20962 7532 20972 7588
rect 21028 7532 21038 7588
rect 21522 7532 21532 7588
rect 21588 7532 24500 7588
rect 27570 7532 27580 7588
rect 27636 7532 29260 7588
rect 29316 7532 29326 7588
rect 30034 7532 30044 7588
rect 30100 7532 31836 7588
rect 31892 7532 31902 7588
rect 6290 7420 6300 7476
rect 6356 7420 7196 7476
rect 7252 7420 7262 7476
rect 10210 7420 10220 7476
rect 10276 7420 11452 7476
rect 11508 7420 13580 7476
rect 13636 7420 13916 7476
rect 13972 7420 15148 7476
rect 16258 7420 16268 7476
rect 16324 7420 18172 7476
rect 18228 7420 18238 7476
rect 6514 7308 6524 7364
rect 6580 7308 8092 7364
rect 8148 7308 8158 7364
rect 9314 7308 9324 7364
rect 9380 7308 9996 7364
rect 10052 7308 10062 7364
rect 18050 7308 18060 7364
rect 18116 7308 20188 7364
rect 20244 7308 20254 7364
rect 20972 7252 21028 7532
rect 23426 7420 23436 7476
rect 23492 7420 24220 7476
rect 24276 7420 24286 7476
rect 24444 7364 24500 7532
rect 25778 7420 25788 7476
rect 25844 7420 26572 7476
rect 26628 7420 28140 7476
rect 28196 7420 28476 7476
rect 28532 7420 28542 7476
rect 29922 7420 29932 7476
rect 29988 7420 31276 7476
rect 31332 7420 31342 7476
rect 22082 7308 22092 7364
rect 22148 7308 23548 7364
rect 23604 7308 23614 7364
rect 24444 7308 28588 7364
rect 28644 7308 28654 7364
rect 20972 7196 28028 7252
rect 28084 7196 28094 7252
rect 19170 7084 19180 7140
rect 19236 7084 20860 7140
rect 20916 7084 20926 7140
rect 27906 7084 27916 7140
rect 27972 7084 28364 7140
rect 28420 7084 28430 7140
rect 5486 7028 5496 7084
rect 5552 7028 5600 7084
rect 5656 7028 5704 7084
rect 5760 7028 5770 7084
rect 14054 7028 14064 7084
rect 14120 7028 14168 7084
rect 14224 7028 14272 7084
rect 14328 7028 14338 7084
rect 22622 7028 22632 7084
rect 22688 7028 22736 7084
rect 22792 7028 22840 7084
rect 22896 7028 22906 7084
rect 31190 7028 31200 7084
rect 31256 7028 31304 7084
rect 31360 7028 31408 7084
rect 31464 7028 31474 7084
rect 8642 6972 8652 7028
rect 8708 6972 9660 7028
rect 9716 6972 9726 7028
rect 9426 6860 9436 6916
rect 9492 6860 12460 6916
rect 12516 6860 12526 6916
rect 28578 6860 28588 6916
rect 28644 6860 29260 6916
rect 29316 6860 29326 6916
rect 6066 6748 6076 6804
rect 6132 6748 7308 6804
rect 7364 6748 8540 6804
rect 8596 6748 8606 6804
rect 23762 6748 23772 6804
rect 23828 6748 25452 6804
rect 25508 6748 25676 6804
rect 25732 6748 25742 6804
rect 27570 6748 27580 6804
rect 27636 6748 28140 6804
rect 28196 6748 28206 6804
rect 29474 6748 29484 6804
rect 29540 6748 32284 6804
rect 32340 6748 32350 6804
rect 31164 6692 31220 6748
rect 19282 6636 19292 6692
rect 19348 6636 20300 6692
rect 20356 6636 20366 6692
rect 21298 6636 21308 6692
rect 21364 6636 21756 6692
rect 21812 6636 26460 6692
rect 26516 6636 28588 6692
rect 28644 6636 28654 6692
rect 31154 6636 31164 6692
rect 31220 6636 31230 6692
rect 16482 6524 16492 6580
rect 16548 6524 18172 6580
rect 18228 6524 18238 6580
rect 18610 6524 18620 6580
rect 18676 6524 19516 6580
rect 19572 6524 19582 6580
rect 24546 6524 24556 6580
rect 24612 6524 26684 6580
rect 26740 6524 26750 6580
rect 27010 6524 27020 6580
rect 27076 6524 27356 6580
rect 27412 6524 27422 6580
rect 14802 6412 14812 6468
rect 14868 6412 15820 6468
rect 15876 6412 15886 6468
rect 9770 6244 9780 6300
rect 9836 6244 9884 6300
rect 9940 6244 9988 6300
rect 10044 6244 10054 6300
rect 16492 6132 16548 6524
rect 17154 6412 17164 6468
rect 17220 6412 18396 6468
rect 18452 6412 20748 6468
rect 20804 6412 20814 6468
rect 24322 6412 24332 6468
rect 24388 6412 24780 6468
rect 24836 6412 24846 6468
rect 28130 6412 28140 6468
rect 28196 6412 29484 6468
rect 29540 6412 29550 6468
rect 24546 6300 24556 6356
rect 24612 6300 25228 6356
rect 25284 6300 25294 6356
rect 18338 6244 18348 6300
rect 18404 6244 18452 6300
rect 18508 6244 18556 6300
rect 18612 6244 18622 6300
rect 26906 6244 26916 6300
rect 26972 6244 27020 6300
rect 27076 6244 27124 6300
rect 27180 6244 27190 6300
rect 35474 6244 35484 6300
rect 35540 6244 35588 6300
rect 35644 6244 35692 6300
rect 35748 6244 35758 6300
rect 13234 6076 13244 6132
rect 13300 6076 14476 6132
rect 14532 6076 16548 6132
rect 5954 5964 5964 6020
rect 6020 5964 10780 6020
rect 10836 5964 10846 6020
rect 11330 5964 11340 6020
rect 11396 5964 13468 6020
rect 13524 5964 13534 6020
rect 14242 5964 14252 6020
rect 14308 5964 16156 6020
rect 16212 5964 16222 6020
rect 20402 5964 20412 6020
rect 20468 5964 24444 6020
rect 24500 5964 25340 6020
rect 25396 5964 25406 6020
rect 27346 5964 27356 6020
rect 27412 5964 27916 6020
rect 27972 5964 27982 6020
rect 9538 5852 9548 5908
rect 9604 5852 11004 5908
rect 11060 5852 11070 5908
rect 12786 5852 12796 5908
rect 12852 5852 17388 5908
rect 17444 5852 17454 5908
rect 25106 5852 25116 5908
rect 25172 5852 26460 5908
rect 26516 5852 26526 5908
rect 6962 5740 6972 5796
rect 7028 5740 10108 5796
rect 10164 5740 10174 5796
rect 12450 5740 12460 5796
rect 12516 5740 13580 5796
rect 13636 5740 13646 5796
rect 16482 5740 16492 5796
rect 16548 5740 18060 5796
rect 18116 5740 19292 5796
rect 19348 5740 19358 5796
rect 22978 5740 22988 5796
rect 23044 5740 31052 5796
rect 31108 5740 31724 5796
rect 31780 5740 31790 5796
rect 11554 5628 11564 5684
rect 11620 5628 13020 5684
rect 13076 5628 13086 5684
rect 15362 5628 15372 5684
rect 15428 5628 17836 5684
rect 17892 5628 17902 5684
rect 20626 5628 20636 5684
rect 20692 5628 21868 5684
rect 21924 5628 21934 5684
rect 25442 5628 25452 5684
rect 25508 5628 27468 5684
rect 27524 5628 27534 5684
rect 8194 5516 8204 5572
rect 8260 5516 8988 5572
rect 9044 5516 10108 5572
rect 10164 5516 10174 5572
rect 25554 5516 25564 5572
rect 25620 5516 25630 5572
rect 5486 5460 5496 5516
rect 5552 5460 5600 5516
rect 5656 5460 5704 5516
rect 5760 5460 5770 5516
rect 14054 5460 14064 5516
rect 14120 5460 14168 5516
rect 14224 5460 14272 5516
rect 14328 5460 14338 5516
rect 22622 5460 22632 5516
rect 22688 5460 22736 5516
rect 22792 5460 22840 5516
rect 22896 5460 22906 5516
rect 25564 5460 25620 5516
rect 31190 5460 31200 5516
rect 31256 5460 31304 5516
rect 31360 5460 31408 5516
rect 31464 5460 31474 5516
rect 25564 5404 26012 5460
rect 26068 5404 26078 5460
rect 13458 5292 13468 5348
rect 13524 5292 14028 5348
rect 14084 5292 14094 5348
rect 24546 5292 24556 5348
rect 24612 5292 25788 5348
rect 25844 5292 25854 5348
rect 26460 5292 27356 5348
rect 27412 5292 27422 5348
rect 27990 5292 28028 5348
rect 28084 5292 28094 5348
rect 5730 5180 5740 5236
rect 5796 5180 9772 5236
rect 9828 5180 12796 5236
rect 12852 5180 12862 5236
rect 14578 5180 14588 5236
rect 14644 5180 15484 5236
rect 15540 5180 17052 5236
rect 17108 5180 17118 5236
rect 22530 5180 22540 5236
rect 22596 5180 25340 5236
rect 25396 5180 25406 5236
rect 26460 5124 26516 5292
rect 6066 5068 6076 5124
rect 6132 5068 9884 5124
rect 9940 5068 11788 5124
rect 11844 5068 11854 5124
rect 12012 5068 13468 5124
rect 13524 5068 13534 5124
rect 17378 5068 17388 5124
rect 17444 5068 19180 5124
rect 19236 5068 19246 5124
rect 24098 5068 24108 5124
rect 24164 5068 25564 5124
rect 25620 5068 26460 5124
rect 26516 5068 26526 5124
rect 34626 5068 34636 5124
rect 34692 5068 35196 5124
rect 35252 5068 35262 5124
rect 12012 5012 12068 5068
rect 35196 5012 35252 5068
rect 36200 5012 37000 5040
rect 6178 4956 6188 5012
rect 6244 4956 12068 5012
rect 16818 4956 16828 5012
rect 16884 4956 17500 5012
rect 17556 4956 17948 5012
rect 18004 4956 19292 5012
rect 19348 4956 19358 5012
rect 20066 4956 20076 5012
rect 20132 4956 22876 5012
rect 22932 4956 22942 5012
rect 29026 4956 29036 5012
rect 29092 4956 31276 5012
rect 31332 4956 31342 5012
rect 35196 4956 37000 5012
rect 36200 4928 37000 4956
rect 9650 4844 9660 4900
rect 9716 4844 12684 4900
rect 12740 4844 12750 4900
rect 14578 4844 14588 4900
rect 14644 4844 19068 4900
rect 19124 4844 19134 4900
rect 27346 4844 27356 4900
rect 27412 4844 30604 4900
rect 30660 4844 30670 4900
rect 10434 4732 10444 4788
rect 10500 4732 11676 4788
rect 11732 4732 11742 4788
rect 9770 4676 9780 4732
rect 9836 4676 9884 4732
rect 9940 4676 9988 4732
rect 10044 4676 10054 4732
rect 18338 4676 18348 4732
rect 18404 4676 18452 4732
rect 18508 4676 18556 4732
rect 18612 4676 18622 4732
rect 26906 4676 26916 4732
rect 26972 4676 27020 4732
rect 27076 4676 27124 4732
rect 27180 4676 27190 4732
rect 35474 4676 35484 4732
rect 35540 4676 35588 4732
rect 35644 4676 35692 4732
rect 35748 4676 35758 4732
rect 5394 4508 5404 4564
rect 5460 4508 5964 4564
rect 6020 4508 9324 4564
rect 9380 4508 11116 4564
rect 11172 4508 11182 4564
rect 16706 4508 16716 4564
rect 16772 4508 17500 4564
rect 17556 4508 17566 4564
rect 17826 4508 17836 4564
rect 17892 4508 18956 4564
rect 19012 4508 22764 4564
rect 22820 4508 23212 4564
rect 23268 4508 23278 4564
rect 26226 4508 26236 4564
rect 26292 4508 27244 4564
rect 27300 4508 28028 4564
rect 28084 4508 28094 4564
rect 15698 4396 15708 4452
rect 15764 4396 17612 4452
rect 17668 4396 17678 4452
rect 22642 4396 22652 4452
rect 22708 4396 24780 4452
rect 24836 4396 24846 4452
rect 28130 4396 28140 4452
rect 28196 4396 28924 4452
rect 28980 4396 28990 4452
rect 12450 4284 12460 4340
rect 12516 4284 16828 4340
rect 16884 4284 16894 4340
rect 25330 4284 25340 4340
rect 25396 4284 29036 4340
rect 29092 4284 29102 4340
rect 6402 4172 6412 4228
rect 6468 4172 9548 4228
rect 9604 4172 10444 4228
rect 10500 4172 10510 4228
rect 11666 4172 11676 4228
rect 11732 4172 12908 4228
rect 12964 4172 12974 4228
rect 17042 4172 17052 4228
rect 17108 4172 18396 4228
rect 18452 4172 18462 4228
rect 24658 4172 24668 4228
rect 24724 4172 27468 4228
rect 27524 4172 27534 4228
rect 29362 4172 29372 4228
rect 29428 4172 30268 4228
rect 30324 4172 30334 4228
rect 17042 3948 17052 4004
rect 17108 3948 17836 4004
rect 17892 3948 17902 4004
rect 5486 3892 5496 3948
rect 5552 3892 5600 3948
rect 5656 3892 5704 3948
rect 5760 3892 5770 3948
rect 14054 3892 14064 3948
rect 14120 3892 14168 3948
rect 14224 3892 14272 3948
rect 14328 3892 14338 3948
rect 22622 3892 22632 3948
rect 22688 3892 22736 3948
rect 22792 3892 22840 3948
rect 22896 3892 22906 3948
rect 31190 3892 31200 3948
rect 31256 3892 31304 3948
rect 31360 3892 31408 3948
rect 31464 3892 31474 3948
rect 27234 3836 27244 3892
rect 27300 3836 28700 3892
rect 28756 3836 29820 3892
rect 29876 3836 29886 3892
rect 7186 3724 7196 3780
rect 7252 3724 9212 3780
rect 9268 3724 9278 3780
rect 13580 3724 17276 3780
rect 17332 3724 17342 3780
rect 24210 3724 24220 3780
rect 24276 3724 28364 3780
rect 28420 3724 28430 3780
rect 13580 3556 13636 3724
rect 17490 3612 17500 3668
rect 17556 3612 18620 3668
rect 18676 3612 18686 3668
rect 19058 3612 19068 3668
rect 19124 3612 21868 3668
rect 21924 3612 21934 3668
rect 22194 3612 22204 3668
rect 22260 3612 25564 3668
rect 25620 3612 25630 3668
rect 13570 3500 13580 3556
rect 13636 3500 13646 3556
rect 13906 3500 13916 3556
rect 13972 3500 17612 3556
rect 17668 3500 17678 3556
rect 18386 3500 18396 3556
rect 18452 3500 20748 3556
rect 20804 3500 20814 3556
rect 28466 3500 28476 3556
rect 28532 3500 29372 3556
rect 29428 3500 31052 3556
rect 31108 3500 31118 3556
rect 31602 3500 31612 3556
rect 31668 3500 32396 3556
rect 32452 3500 32956 3556
rect 33012 3500 33022 3556
rect 13916 3444 13972 3500
rect 3938 3388 3948 3444
rect 4004 3388 4956 3444
rect 5012 3388 5022 3444
rect 8306 3388 8316 3444
rect 8372 3388 9716 3444
rect 13346 3388 13356 3444
rect 13412 3388 13972 3444
rect 25330 3388 25340 3444
rect 25396 3388 27804 3444
rect 27860 3388 29820 3444
rect 29876 3388 29886 3444
rect 30034 3388 30044 3444
rect 30100 3388 30604 3444
rect 30660 3388 31500 3444
rect 31556 3388 31566 3444
rect 9650 3332 9660 3388
rect 9716 3332 9726 3388
rect 32274 3276 32284 3332
rect 32340 3276 33404 3332
rect 33460 3276 33470 3332
rect 9770 3108 9780 3164
rect 9836 3108 9884 3164
rect 9940 3108 9988 3164
rect 10044 3108 10054 3164
rect 18338 3108 18348 3164
rect 18404 3108 18452 3164
rect 18508 3108 18556 3164
rect 18612 3108 18622 3164
rect 26906 3108 26916 3164
rect 26972 3108 27020 3164
rect 27076 3108 27124 3164
rect 27180 3108 27190 3164
rect 35474 3108 35484 3164
rect 35540 3108 35588 3164
rect 35644 3108 35692 3164
rect 35748 3108 35758 3164
rect 36200 2324 37000 2352
rect 32610 2268 32620 2324
rect 32676 2268 37000 2324
rect 36200 2240 37000 2268
<< via3 >>
rect 5496 33684 5552 33740
rect 5600 33684 5656 33740
rect 5704 33684 5760 33740
rect 14064 33684 14120 33740
rect 14168 33684 14224 33740
rect 14272 33684 14328 33740
rect 22632 33684 22688 33740
rect 22736 33684 22792 33740
rect 22840 33684 22896 33740
rect 31200 33684 31256 33740
rect 31304 33684 31360 33740
rect 31408 33684 31464 33740
rect 9780 32900 9836 32956
rect 9884 32900 9940 32956
rect 9988 32900 10044 32956
rect 18348 32900 18404 32956
rect 18452 32900 18508 32956
rect 18556 32900 18612 32956
rect 26916 32900 26972 32956
rect 27020 32900 27076 32956
rect 27124 32900 27180 32956
rect 35484 32900 35540 32956
rect 35588 32900 35644 32956
rect 35692 32900 35748 32956
rect 5496 32116 5552 32172
rect 5600 32116 5656 32172
rect 5704 32116 5760 32172
rect 14064 32116 14120 32172
rect 14168 32116 14224 32172
rect 14272 32116 14328 32172
rect 22632 32116 22688 32172
rect 22736 32116 22792 32172
rect 22840 32116 22896 32172
rect 31200 32116 31256 32172
rect 31304 32116 31360 32172
rect 31408 32116 31464 32172
rect 9780 31332 9836 31388
rect 9884 31332 9940 31388
rect 9988 31332 10044 31388
rect 18348 31332 18404 31388
rect 18452 31332 18508 31388
rect 18556 31332 18612 31388
rect 26916 31332 26972 31388
rect 27020 31332 27076 31388
rect 27124 31332 27180 31388
rect 35484 31332 35540 31388
rect 35588 31332 35644 31388
rect 35692 31332 35748 31388
rect 33068 31052 33124 31108
rect 5496 30548 5552 30604
rect 5600 30548 5656 30604
rect 5704 30548 5760 30604
rect 14064 30548 14120 30604
rect 14168 30548 14224 30604
rect 14272 30548 14328 30604
rect 22632 30548 22688 30604
rect 22736 30548 22792 30604
rect 22840 30548 22896 30604
rect 31200 30548 31256 30604
rect 31304 30548 31360 30604
rect 31408 30548 31464 30604
rect 9548 30268 9604 30324
rect 34636 29932 34692 29988
rect 13916 29820 13972 29876
rect 9780 29764 9836 29820
rect 9884 29764 9940 29820
rect 9988 29764 10044 29820
rect 18348 29764 18404 29820
rect 18452 29764 18508 29820
rect 18556 29764 18612 29820
rect 26916 29764 26972 29820
rect 27020 29764 27076 29820
rect 27124 29764 27180 29820
rect 35484 29764 35540 29820
rect 35588 29764 35644 29820
rect 35692 29764 35748 29820
rect 35084 29372 35140 29428
rect 18060 29260 18116 29316
rect 5496 28980 5552 29036
rect 5600 28980 5656 29036
rect 5704 28980 5760 29036
rect 14064 28980 14120 29036
rect 14168 28980 14224 29036
rect 14272 28980 14328 29036
rect 22632 28980 22688 29036
rect 22736 28980 22792 29036
rect 22840 28980 22896 29036
rect 31200 28980 31256 29036
rect 31304 28980 31360 29036
rect 31408 28980 31464 29036
rect 13692 28924 13748 28980
rect 18956 28924 19012 28980
rect 27580 28476 27636 28532
rect 19852 28364 19908 28420
rect 27356 28252 27412 28308
rect 9780 28196 9836 28252
rect 9884 28196 9940 28252
rect 9988 28196 10044 28252
rect 18348 28196 18404 28252
rect 18452 28196 18508 28252
rect 18556 28196 18612 28252
rect 26916 28196 26972 28252
rect 27020 28196 27076 28252
rect 27124 28196 27180 28252
rect 35484 28196 35540 28252
rect 35588 28196 35644 28252
rect 35692 28196 35748 28252
rect 18060 28028 18116 28084
rect 13692 27916 13748 27972
rect 9548 27692 9604 27748
rect 18956 27692 19012 27748
rect 19740 27580 19796 27636
rect 5496 27412 5552 27468
rect 5600 27412 5656 27468
rect 5704 27412 5760 27468
rect 14064 27412 14120 27468
rect 14168 27412 14224 27468
rect 14272 27412 14328 27468
rect 22632 27412 22688 27468
rect 22736 27412 22792 27468
rect 22840 27412 22896 27468
rect 31200 27412 31256 27468
rect 31304 27412 31360 27468
rect 31408 27412 31464 27468
rect 17836 27356 17892 27412
rect 8204 27020 8260 27076
rect 17836 27020 17892 27076
rect 13916 26796 13972 26852
rect 19740 26796 19796 26852
rect 9780 26628 9836 26684
rect 9884 26628 9940 26684
rect 9988 26628 10044 26684
rect 18348 26628 18404 26684
rect 18452 26628 18508 26684
rect 18556 26628 18612 26684
rect 26916 26628 26972 26684
rect 27020 26628 27076 26684
rect 27124 26628 27180 26684
rect 35484 26628 35540 26684
rect 35588 26628 35644 26684
rect 35692 26628 35748 26684
rect 7644 26572 7700 26628
rect 8204 26572 8260 26628
rect 18060 26572 18116 26628
rect 7644 26348 7700 26404
rect 5496 25844 5552 25900
rect 5600 25844 5656 25900
rect 5704 25844 5760 25900
rect 14064 25844 14120 25900
rect 14168 25844 14224 25900
rect 14272 25844 14328 25900
rect 22632 25844 22688 25900
rect 22736 25844 22792 25900
rect 22840 25844 22896 25900
rect 31200 25844 31256 25900
rect 31304 25844 31360 25900
rect 31408 25844 31464 25900
rect 34188 25788 34244 25844
rect 19852 25676 19908 25732
rect 13692 25116 13748 25172
rect 9780 25060 9836 25116
rect 9884 25060 9940 25116
rect 9988 25060 10044 25116
rect 18348 25060 18404 25116
rect 18452 25060 18508 25116
rect 18556 25060 18612 25116
rect 26916 25060 26972 25116
rect 27020 25060 27076 25116
rect 27124 25060 27180 25116
rect 35484 25060 35540 25116
rect 35588 25060 35644 25116
rect 35692 25060 35748 25116
rect 19852 24892 19908 24948
rect 34188 24892 34244 24948
rect 35084 24780 35140 24836
rect 5496 24276 5552 24332
rect 5600 24276 5656 24332
rect 5704 24276 5760 24332
rect 14064 24276 14120 24332
rect 14168 24276 14224 24332
rect 14272 24276 14328 24332
rect 22632 24276 22688 24332
rect 22736 24276 22792 24332
rect 22840 24276 22896 24332
rect 31200 24276 31256 24332
rect 31304 24276 31360 24332
rect 31408 24276 31464 24332
rect 26236 23660 26292 23716
rect 9780 23492 9836 23548
rect 9884 23492 9940 23548
rect 9988 23492 10044 23548
rect 18348 23492 18404 23548
rect 18452 23492 18508 23548
rect 18556 23492 18612 23548
rect 26916 23492 26972 23548
rect 27020 23492 27076 23548
rect 27124 23492 27180 23548
rect 35484 23492 35540 23548
rect 35588 23492 35644 23548
rect 35692 23492 35748 23548
rect 34748 23324 34804 23380
rect 25228 22988 25284 23044
rect 26236 22764 26292 22820
rect 28028 22764 28084 22820
rect 5496 22708 5552 22764
rect 5600 22708 5656 22764
rect 5704 22708 5760 22764
rect 14064 22708 14120 22764
rect 14168 22708 14224 22764
rect 14272 22708 14328 22764
rect 22632 22708 22688 22764
rect 22736 22708 22792 22764
rect 22840 22708 22896 22764
rect 31200 22708 31256 22764
rect 31304 22708 31360 22764
rect 31408 22708 31464 22764
rect 34748 22540 34804 22596
rect 33068 22316 33124 22372
rect 15260 22092 15316 22148
rect 34636 22092 34692 22148
rect 26684 21980 26740 22036
rect 28476 21980 28532 22036
rect 9780 21924 9836 21980
rect 9884 21924 9940 21980
rect 9988 21924 10044 21980
rect 18348 21924 18404 21980
rect 18452 21924 18508 21980
rect 18556 21924 18612 21980
rect 26916 21924 26972 21980
rect 27020 21924 27076 21980
rect 27124 21924 27180 21980
rect 35484 21924 35540 21980
rect 35588 21924 35644 21980
rect 35692 21924 35748 21980
rect 15372 21644 15428 21700
rect 15820 21644 15876 21700
rect 26684 21420 26740 21476
rect 5496 21140 5552 21196
rect 5600 21140 5656 21196
rect 5704 21140 5760 21196
rect 14064 21140 14120 21196
rect 14168 21140 14224 21196
rect 14272 21140 14328 21196
rect 22632 21140 22688 21196
rect 22736 21140 22792 21196
rect 22840 21140 22896 21196
rect 31200 21140 31256 21196
rect 31304 21140 31360 21196
rect 31408 21140 31464 21196
rect 28476 21084 28532 21140
rect 28252 20972 28308 21028
rect 9780 20356 9836 20412
rect 9884 20356 9940 20412
rect 9988 20356 10044 20412
rect 18348 20356 18404 20412
rect 18452 20356 18508 20412
rect 18556 20356 18612 20412
rect 26916 20356 26972 20412
rect 27020 20356 27076 20412
rect 27124 20356 27180 20412
rect 35484 20356 35540 20412
rect 35588 20356 35644 20412
rect 35692 20356 35748 20412
rect 26684 20300 26740 20356
rect 26236 20188 26292 20244
rect 28252 20076 28308 20132
rect 35084 19964 35140 20020
rect 25564 19740 25620 19796
rect 5496 19572 5552 19628
rect 5600 19572 5656 19628
rect 5704 19572 5760 19628
rect 14064 19572 14120 19628
rect 14168 19572 14224 19628
rect 14272 19572 14328 19628
rect 22632 19572 22688 19628
rect 22736 19572 22792 19628
rect 22840 19572 22896 19628
rect 31200 19572 31256 19628
rect 31304 19572 31360 19628
rect 31408 19572 31464 19628
rect 25228 19292 25284 19348
rect 28252 19292 28308 19348
rect 9780 18788 9836 18844
rect 9884 18788 9940 18844
rect 9988 18788 10044 18844
rect 18348 18788 18404 18844
rect 18452 18788 18508 18844
rect 18556 18788 18612 18844
rect 26916 18788 26972 18844
rect 27020 18788 27076 18844
rect 27124 18788 27180 18844
rect 35484 18788 35540 18844
rect 35588 18788 35644 18844
rect 35692 18788 35748 18844
rect 26124 18620 26180 18676
rect 26572 18620 26628 18676
rect 31948 18508 32004 18564
rect 26572 18396 26628 18452
rect 27356 18396 27412 18452
rect 27580 18396 27636 18452
rect 28140 18172 28196 18228
rect 5496 18004 5552 18060
rect 5600 18004 5656 18060
rect 5704 18004 5760 18060
rect 14064 18004 14120 18060
rect 14168 18004 14224 18060
rect 14272 18004 14328 18060
rect 22632 18004 22688 18060
rect 22736 18004 22792 18060
rect 22840 18004 22896 18060
rect 31200 18004 31256 18060
rect 31304 18004 31360 18060
rect 31408 18004 31464 18060
rect 32508 17948 32564 18004
rect 25788 17724 25844 17780
rect 28028 17388 28084 17444
rect 35084 17276 35140 17332
rect 9780 17220 9836 17276
rect 9884 17220 9940 17276
rect 9988 17220 10044 17276
rect 18348 17220 18404 17276
rect 18452 17220 18508 17276
rect 18556 17220 18612 17276
rect 26916 17220 26972 17276
rect 27020 17220 27076 17276
rect 27124 17220 27180 17276
rect 35484 17220 35540 17276
rect 35588 17220 35644 17276
rect 35692 17220 35748 17276
rect 34972 17164 35028 17220
rect 25564 17052 25620 17108
rect 25788 16716 25844 16772
rect 26684 16716 26740 16772
rect 27692 16716 27748 16772
rect 26572 16604 26628 16660
rect 28476 16604 28532 16660
rect 5496 16436 5552 16492
rect 5600 16436 5656 16492
rect 5704 16436 5760 16492
rect 14064 16436 14120 16492
rect 14168 16436 14224 16492
rect 14272 16436 14328 16492
rect 22632 16436 22688 16492
rect 22736 16436 22792 16492
rect 22840 16436 22896 16492
rect 31200 16436 31256 16492
rect 31304 16436 31360 16492
rect 31408 16436 31464 16492
rect 15260 16268 15316 16324
rect 26684 15820 26740 15876
rect 9780 15652 9836 15708
rect 9884 15652 9940 15708
rect 9988 15652 10044 15708
rect 18348 15652 18404 15708
rect 18452 15652 18508 15708
rect 18556 15652 18612 15708
rect 26916 15652 26972 15708
rect 27020 15652 27076 15708
rect 27124 15652 27180 15708
rect 35484 15652 35540 15708
rect 35588 15652 35644 15708
rect 35692 15652 35748 15708
rect 26348 15596 26404 15652
rect 34972 15484 35028 15540
rect 27804 15260 27860 15316
rect 28252 15260 28308 15316
rect 25564 15148 25620 15204
rect 26348 15148 26404 15204
rect 26572 15036 26628 15092
rect 28476 15036 28532 15092
rect 32172 14924 32228 14980
rect 5496 14868 5552 14924
rect 5600 14868 5656 14924
rect 5704 14868 5760 14924
rect 14064 14868 14120 14924
rect 14168 14868 14224 14924
rect 14272 14868 14328 14924
rect 22632 14868 22688 14924
rect 22736 14868 22792 14924
rect 22840 14868 22896 14924
rect 31200 14868 31256 14924
rect 31304 14868 31360 14924
rect 31408 14868 31464 14924
rect 27692 14812 27748 14868
rect 32508 14476 32564 14532
rect 9780 14084 9836 14140
rect 9884 14084 9940 14140
rect 9988 14084 10044 14140
rect 18348 14084 18404 14140
rect 18452 14084 18508 14140
rect 18556 14084 18612 14140
rect 26916 14084 26972 14140
rect 27020 14084 27076 14140
rect 27124 14084 27180 14140
rect 26684 13916 26740 13972
rect 35484 14084 35540 14140
rect 35588 14084 35644 14140
rect 35692 14084 35748 14140
rect 28252 13804 28308 13860
rect 5496 13300 5552 13356
rect 5600 13300 5656 13356
rect 5704 13300 5760 13356
rect 14064 13300 14120 13356
rect 14168 13300 14224 13356
rect 14272 13300 14328 13356
rect 22632 13300 22688 13356
rect 22736 13300 22792 13356
rect 22840 13300 22896 13356
rect 31200 13300 31256 13356
rect 31304 13300 31360 13356
rect 31408 13300 31464 13356
rect 32172 13132 32228 13188
rect 27804 12908 27860 12964
rect 28140 12908 28196 12964
rect 9780 12516 9836 12572
rect 9884 12516 9940 12572
rect 9988 12516 10044 12572
rect 18348 12516 18404 12572
rect 18452 12516 18508 12572
rect 18556 12516 18612 12572
rect 26916 12516 26972 12572
rect 27020 12516 27076 12572
rect 27124 12516 27180 12572
rect 35484 12516 35540 12572
rect 35588 12516 35644 12572
rect 35692 12516 35748 12572
rect 5496 11732 5552 11788
rect 5600 11732 5656 11788
rect 5704 11732 5760 11788
rect 14064 11732 14120 11788
rect 14168 11732 14224 11788
rect 14272 11732 14328 11788
rect 22632 11732 22688 11788
rect 22736 11732 22792 11788
rect 22840 11732 22896 11788
rect 31200 11732 31256 11788
rect 31304 11732 31360 11788
rect 31408 11732 31464 11788
rect 31948 11676 32004 11732
rect 34636 11452 34692 11508
rect 34972 11340 35028 11396
rect 9780 10948 9836 11004
rect 9884 10948 9940 11004
rect 9988 10948 10044 11004
rect 18348 10948 18404 11004
rect 18452 10948 18508 11004
rect 18556 10948 18612 11004
rect 26916 10948 26972 11004
rect 27020 10948 27076 11004
rect 27124 10948 27180 11004
rect 35484 10948 35540 11004
rect 35588 10948 35644 11004
rect 35692 10948 35748 11004
rect 15596 10556 15652 10612
rect 16492 10332 16548 10388
rect 5496 10164 5552 10220
rect 5600 10164 5656 10220
rect 5704 10164 5760 10220
rect 14064 10164 14120 10220
rect 14168 10164 14224 10220
rect 14272 10164 14328 10220
rect 22632 10164 22688 10220
rect 22736 10164 22792 10220
rect 22840 10164 22896 10220
rect 31200 10164 31256 10220
rect 31304 10164 31360 10220
rect 31408 10164 31464 10220
rect 9780 9380 9836 9436
rect 9884 9380 9940 9436
rect 9988 9380 10044 9436
rect 18348 9380 18404 9436
rect 18452 9380 18508 9436
rect 18556 9380 18612 9436
rect 26916 9380 26972 9436
rect 27020 9380 27076 9436
rect 27124 9380 27180 9436
rect 35484 9380 35540 9436
rect 35588 9380 35644 9436
rect 35692 9380 35748 9436
rect 15596 9212 15652 9268
rect 5496 8596 5552 8652
rect 5600 8596 5656 8652
rect 5704 8596 5760 8652
rect 14064 8596 14120 8652
rect 14168 8596 14224 8652
rect 14272 8596 14328 8652
rect 22632 8596 22688 8652
rect 22736 8596 22792 8652
rect 22840 8596 22896 8652
rect 31200 8596 31256 8652
rect 31304 8596 31360 8652
rect 31408 8596 31464 8652
rect 16492 7980 16548 8036
rect 9780 7812 9836 7868
rect 9884 7812 9940 7868
rect 9988 7812 10044 7868
rect 18348 7812 18404 7868
rect 18452 7812 18508 7868
rect 18556 7812 18612 7868
rect 26916 7812 26972 7868
rect 27020 7812 27076 7868
rect 27124 7812 27180 7868
rect 35484 7812 35540 7868
rect 35588 7812 35644 7868
rect 35692 7812 35748 7868
rect 28028 7196 28084 7252
rect 5496 7028 5552 7084
rect 5600 7028 5656 7084
rect 5704 7028 5760 7084
rect 14064 7028 14120 7084
rect 14168 7028 14224 7084
rect 14272 7028 14328 7084
rect 22632 7028 22688 7084
rect 22736 7028 22792 7084
rect 22840 7028 22896 7084
rect 31200 7028 31256 7084
rect 31304 7028 31360 7084
rect 31408 7028 31464 7084
rect 9780 6244 9836 6300
rect 9884 6244 9940 6300
rect 9988 6244 10044 6300
rect 18348 6244 18404 6300
rect 18452 6244 18508 6300
rect 18556 6244 18612 6300
rect 26916 6244 26972 6300
rect 27020 6244 27076 6300
rect 27124 6244 27180 6300
rect 35484 6244 35540 6300
rect 35588 6244 35644 6300
rect 35692 6244 35748 6300
rect 5496 5460 5552 5516
rect 5600 5460 5656 5516
rect 5704 5460 5760 5516
rect 14064 5460 14120 5516
rect 14168 5460 14224 5516
rect 14272 5460 14328 5516
rect 22632 5460 22688 5516
rect 22736 5460 22792 5516
rect 22840 5460 22896 5516
rect 31200 5460 31256 5516
rect 31304 5460 31360 5516
rect 31408 5460 31464 5516
rect 28028 5292 28084 5348
rect 9780 4676 9836 4732
rect 9884 4676 9940 4732
rect 9988 4676 10044 4732
rect 18348 4676 18404 4732
rect 18452 4676 18508 4732
rect 18556 4676 18612 4732
rect 26916 4676 26972 4732
rect 27020 4676 27076 4732
rect 27124 4676 27180 4732
rect 35484 4676 35540 4732
rect 35588 4676 35644 4732
rect 35692 4676 35748 4732
rect 5496 3892 5552 3948
rect 5600 3892 5656 3948
rect 5704 3892 5760 3948
rect 14064 3892 14120 3948
rect 14168 3892 14224 3948
rect 14272 3892 14328 3948
rect 22632 3892 22688 3948
rect 22736 3892 22792 3948
rect 22840 3892 22896 3948
rect 31200 3892 31256 3948
rect 31304 3892 31360 3948
rect 31408 3892 31464 3948
rect 9780 3108 9836 3164
rect 9884 3108 9940 3164
rect 9988 3108 10044 3164
rect 18348 3108 18404 3164
rect 18452 3108 18508 3164
rect 18556 3108 18612 3164
rect 26916 3108 26972 3164
rect 27020 3108 27076 3164
rect 27124 3108 27180 3164
rect 35484 3108 35540 3164
rect 35588 3108 35644 3164
rect 35692 3108 35748 3164
<< metal4 >>
rect 5468 33740 5788 33772
rect 5468 33684 5496 33740
rect 5552 33684 5600 33740
rect 5656 33684 5704 33740
rect 5760 33684 5788 33740
rect 5468 32172 5788 33684
rect 5468 32116 5496 32172
rect 5552 32116 5600 32172
rect 5656 32116 5704 32172
rect 5760 32116 5788 32172
rect 5468 30604 5788 32116
rect 5468 30548 5496 30604
rect 5552 30548 5600 30604
rect 5656 30548 5704 30604
rect 5760 30548 5788 30604
rect 5468 29036 5788 30548
rect 9752 32956 10072 33772
rect 9752 32900 9780 32956
rect 9836 32900 9884 32956
rect 9940 32900 9988 32956
rect 10044 32900 10072 32956
rect 9752 31388 10072 32900
rect 9752 31332 9780 31388
rect 9836 31332 9884 31388
rect 9940 31332 9988 31388
rect 10044 31332 10072 31388
rect 5468 28980 5496 29036
rect 5552 28980 5600 29036
rect 5656 28980 5704 29036
rect 5760 28980 5788 29036
rect 5468 27468 5788 28980
rect 9548 30324 9604 30334
rect 9548 27748 9604 30268
rect 9548 27682 9604 27692
rect 9752 29820 10072 31332
rect 14036 33740 14356 33772
rect 14036 33684 14064 33740
rect 14120 33684 14168 33740
rect 14224 33684 14272 33740
rect 14328 33684 14356 33740
rect 14036 32172 14356 33684
rect 14036 32116 14064 32172
rect 14120 32116 14168 32172
rect 14224 32116 14272 32172
rect 14328 32116 14356 32172
rect 14036 30604 14356 32116
rect 14036 30548 14064 30604
rect 14120 30548 14168 30604
rect 14224 30548 14272 30604
rect 14328 30548 14356 30604
rect 9752 29764 9780 29820
rect 9836 29764 9884 29820
rect 9940 29764 9988 29820
rect 10044 29764 10072 29820
rect 9752 28252 10072 29764
rect 13916 29876 13972 29886
rect 9752 28196 9780 28252
rect 9836 28196 9884 28252
rect 9940 28196 9988 28252
rect 10044 28196 10072 28252
rect 5468 27412 5496 27468
rect 5552 27412 5600 27468
rect 5656 27412 5704 27468
rect 5760 27412 5788 27468
rect 5468 25900 5788 27412
rect 8204 27076 8260 27086
rect 7644 26628 7700 26638
rect 7644 26404 7700 26572
rect 8204 26628 8260 27020
rect 8204 26562 8260 26572
rect 9752 26684 10072 28196
rect 9752 26628 9780 26684
rect 9836 26628 9884 26684
rect 9940 26628 9988 26684
rect 10044 26628 10072 26684
rect 7644 26338 7700 26348
rect 5468 25844 5496 25900
rect 5552 25844 5600 25900
rect 5656 25844 5704 25900
rect 5760 25844 5788 25900
rect 5468 24332 5788 25844
rect 5468 24276 5496 24332
rect 5552 24276 5600 24332
rect 5656 24276 5704 24332
rect 5760 24276 5788 24332
rect 5468 22764 5788 24276
rect 5468 22708 5496 22764
rect 5552 22708 5600 22764
rect 5656 22708 5704 22764
rect 5760 22708 5788 22764
rect 5468 21196 5788 22708
rect 5468 21140 5496 21196
rect 5552 21140 5600 21196
rect 5656 21140 5704 21196
rect 5760 21140 5788 21196
rect 5468 19628 5788 21140
rect 5468 19572 5496 19628
rect 5552 19572 5600 19628
rect 5656 19572 5704 19628
rect 5760 19572 5788 19628
rect 5468 18060 5788 19572
rect 5468 18004 5496 18060
rect 5552 18004 5600 18060
rect 5656 18004 5704 18060
rect 5760 18004 5788 18060
rect 5468 16492 5788 18004
rect 5468 16436 5496 16492
rect 5552 16436 5600 16492
rect 5656 16436 5704 16492
rect 5760 16436 5788 16492
rect 5468 14924 5788 16436
rect 5468 14868 5496 14924
rect 5552 14868 5600 14924
rect 5656 14868 5704 14924
rect 5760 14868 5788 14924
rect 5468 13356 5788 14868
rect 5468 13300 5496 13356
rect 5552 13300 5600 13356
rect 5656 13300 5704 13356
rect 5760 13300 5788 13356
rect 5468 11788 5788 13300
rect 5468 11732 5496 11788
rect 5552 11732 5600 11788
rect 5656 11732 5704 11788
rect 5760 11732 5788 11788
rect 5468 10220 5788 11732
rect 5468 10164 5496 10220
rect 5552 10164 5600 10220
rect 5656 10164 5704 10220
rect 5760 10164 5788 10220
rect 5468 8652 5788 10164
rect 5468 8596 5496 8652
rect 5552 8596 5600 8652
rect 5656 8596 5704 8652
rect 5760 8596 5788 8652
rect 5468 7084 5788 8596
rect 5468 7028 5496 7084
rect 5552 7028 5600 7084
rect 5656 7028 5704 7084
rect 5760 7028 5788 7084
rect 5468 5516 5788 7028
rect 5468 5460 5496 5516
rect 5552 5460 5600 5516
rect 5656 5460 5704 5516
rect 5760 5460 5788 5516
rect 5468 3948 5788 5460
rect 5468 3892 5496 3948
rect 5552 3892 5600 3948
rect 5656 3892 5704 3948
rect 5760 3892 5788 3948
rect 5468 3076 5788 3892
rect 9752 25116 10072 26628
rect 9752 25060 9780 25116
rect 9836 25060 9884 25116
rect 9940 25060 9988 25116
rect 10044 25060 10072 25116
rect 13692 28980 13748 28990
rect 13692 27972 13748 28924
rect 13692 25172 13748 27916
rect 13916 26852 13972 29820
rect 13916 26786 13972 26796
rect 14036 29036 14356 30548
rect 18320 32956 18640 33772
rect 18320 32900 18348 32956
rect 18404 32900 18452 32956
rect 18508 32900 18556 32956
rect 18612 32900 18640 32956
rect 18320 31388 18640 32900
rect 18320 31332 18348 31388
rect 18404 31332 18452 31388
rect 18508 31332 18556 31388
rect 18612 31332 18640 31388
rect 18320 29820 18640 31332
rect 18320 29764 18348 29820
rect 18404 29764 18452 29820
rect 18508 29764 18556 29820
rect 18612 29764 18640 29820
rect 14036 28980 14064 29036
rect 14120 28980 14168 29036
rect 14224 28980 14272 29036
rect 14328 28980 14356 29036
rect 14036 27468 14356 28980
rect 14036 27412 14064 27468
rect 14120 27412 14168 27468
rect 14224 27412 14272 27468
rect 14328 27412 14356 27468
rect 18060 29316 18116 29326
rect 18060 28084 18116 29260
rect 13692 25106 13748 25116
rect 14036 25900 14356 27412
rect 17836 27412 17892 27422
rect 17836 27076 17892 27356
rect 17836 27010 17892 27020
rect 18060 26628 18116 28028
rect 18060 26562 18116 26572
rect 18320 28252 18640 29764
rect 22604 33740 22924 33772
rect 22604 33684 22632 33740
rect 22688 33684 22736 33740
rect 22792 33684 22840 33740
rect 22896 33684 22924 33740
rect 22604 32172 22924 33684
rect 22604 32116 22632 32172
rect 22688 32116 22736 32172
rect 22792 32116 22840 32172
rect 22896 32116 22924 32172
rect 22604 30604 22924 32116
rect 22604 30548 22632 30604
rect 22688 30548 22736 30604
rect 22792 30548 22840 30604
rect 22896 30548 22924 30604
rect 22604 29036 22924 30548
rect 18320 28196 18348 28252
rect 18404 28196 18452 28252
rect 18508 28196 18556 28252
rect 18612 28196 18640 28252
rect 18320 26684 18640 28196
rect 18956 28980 19012 28990
rect 18956 27748 19012 28924
rect 22604 28980 22632 29036
rect 22688 28980 22736 29036
rect 22792 28980 22840 29036
rect 22896 28980 22924 29036
rect 18956 27682 19012 27692
rect 19852 28420 19908 28430
rect 19740 27636 19796 27646
rect 19740 26852 19796 27580
rect 19740 26786 19796 26796
rect 18320 26628 18348 26684
rect 18404 26628 18452 26684
rect 18508 26628 18556 26684
rect 18612 26628 18640 26684
rect 14036 25844 14064 25900
rect 14120 25844 14168 25900
rect 14224 25844 14272 25900
rect 14328 25844 14356 25900
rect 9752 23548 10072 25060
rect 9752 23492 9780 23548
rect 9836 23492 9884 23548
rect 9940 23492 9988 23548
rect 10044 23492 10072 23548
rect 9752 21980 10072 23492
rect 9752 21924 9780 21980
rect 9836 21924 9884 21980
rect 9940 21924 9988 21980
rect 10044 21924 10072 21980
rect 9752 20412 10072 21924
rect 9752 20356 9780 20412
rect 9836 20356 9884 20412
rect 9940 20356 9988 20412
rect 10044 20356 10072 20412
rect 9752 18844 10072 20356
rect 9752 18788 9780 18844
rect 9836 18788 9884 18844
rect 9940 18788 9988 18844
rect 10044 18788 10072 18844
rect 9752 17276 10072 18788
rect 9752 17220 9780 17276
rect 9836 17220 9884 17276
rect 9940 17220 9988 17276
rect 10044 17220 10072 17276
rect 9752 15708 10072 17220
rect 9752 15652 9780 15708
rect 9836 15652 9884 15708
rect 9940 15652 9988 15708
rect 10044 15652 10072 15708
rect 9752 14140 10072 15652
rect 9752 14084 9780 14140
rect 9836 14084 9884 14140
rect 9940 14084 9988 14140
rect 10044 14084 10072 14140
rect 9752 12572 10072 14084
rect 9752 12516 9780 12572
rect 9836 12516 9884 12572
rect 9940 12516 9988 12572
rect 10044 12516 10072 12572
rect 9752 11004 10072 12516
rect 9752 10948 9780 11004
rect 9836 10948 9884 11004
rect 9940 10948 9988 11004
rect 10044 10948 10072 11004
rect 9752 9436 10072 10948
rect 9752 9380 9780 9436
rect 9836 9380 9884 9436
rect 9940 9380 9988 9436
rect 10044 9380 10072 9436
rect 9752 7868 10072 9380
rect 9752 7812 9780 7868
rect 9836 7812 9884 7868
rect 9940 7812 9988 7868
rect 10044 7812 10072 7868
rect 9752 6300 10072 7812
rect 9752 6244 9780 6300
rect 9836 6244 9884 6300
rect 9940 6244 9988 6300
rect 10044 6244 10072 6300
rect 9752 4732 10072 6244
rect 9752 4676 9780 4732
rect 9836 4676 9884 4732
rect 9940 4676 9988 4732
rect 10044 4676 10072 4732
rect 9752 3164 10072 4676
rect 9752 3108 9780 3164
rect 9836 3108 9884 3164
rect 9940 3108 9988 3164
rect 10044 3108 10072 3164
rect 9752 3076 10072 3108
rect 14036 24332 14356 25844
rect 14036 24276 14064 24332
rect 14120 24276 14168 24332
rect 14224 24276 14272 24332
rect 14328 24276 14356 24332
rect 14036 22764 14356 24276
rect 14036 22708 14064 22764
rect 14120 22708 14168 22764
rect 14224 22708 14272 22764
rect 14328 22708 14356 22764
rect 14036 21196 14356 22708
rect 18320 25116 18640 26628
rect 18320 25060 18348 25116
rect 18404 25060 18452 25116
rect 18508 25060 18556 25116
rect 18612 25060 18640 25116
rect 18320 23548 18640 25060
rect 19852 25732 19908 28364
rect 19852 24948 19908 25676
rect 19852 24882 19908 24892
rect 22604 27468 22924 28980
rect 22604 27412 22632 27468
rect 22688 27412 22736 27468
rect 22792 27412 22840 27468
rect 22896 27412 22924 27468
rect 22604 25900 22924 27412
rect 22604 25844 22632 25900
rect 22688 25844 22736 25900
rect 22792 25844 22840 25900
rect 22896 25844 22924 25900
rect 18320 23492 18348 23548
rect 18404 23492 18452 23548
rect 18508 23492 18556 23548
rect 18612 23492 18640 23548
rect 14036 21140 14064 21196
rect 14120 21140 14168 21196
rect 14224 21140 14272 21196
rect 14328 21140 14356 21196
rect 14036 19628 14356 21140
rect 14036 19572 14064 19628
rect 14120 19572 14168 19628
rect 14224 19572 14272 19628
rect 14328 19572 14356 19628
rect 14036 18060 14356 19572
rect 14036 18004 14064 18060
rect 14120 18004 14168 18060
rect 14224 18004 14272 18060
rect 14328 18004 14356 18060
rect 14036 16492 14356 18004
rect 14036 16436 14064 16492
rect 14120 16436 14168 16492
rect 14224 16436 14272 16492
rect 14328 16436 14356 16492
rect 14036 14924 14356 16436
rect 15260 22148 15316 22158
rect 15260 16324 15316 22092
rect 18320 21980 18640 23492
rect 18320 21924 18348 21980
rect 18404 21924 18452 21980
rect 18508 21924 18556 21980
rect 18612 21924 18640 21980
rect 15372 21700 15876 21718
rect 15428 21662 15820 21700
rect 15372 21634 15428 21644
rect 15820 21634 15876 21644
rect 15260 16258 15316 16268
rect 18320 20412 18640 21924
rect 18320 20356 18348 20412
rect 18404 20356 18452 20412
rect 18508 20356 18556 20412
rect 18612 20356 18640 20412
rect 18320 18844 18640 20356
rect 18320 18788 18348 18844
rect 18404 18788 18452 18844
rect 18508 18788 18556 18844
rect 18612 18788 18640 18844
rect 18320 17276 18640 18788
rect 18320 17220 18348 17276
rect 18404 17220 18452 17276
rect 18508 17220 18556 17276
rect 18612 17220 18640 17276
rect 14036 14868 14064 14924
rect 14120 14868 14168 14924
rect 14224 14868 14272 14924
rect 14328 14868 14356 14924
rect 14036 13356 14356 14868
rect 14036 13300 14064 13356
rect 14120 13300 14168 13356
rect 14224 13300 14272 13356
rect 14328 13300 14356 13356
rect 14036 11788 14356 13300
rect 14036 11732 14064 11788
rect 14120 11732 14168 11788
rect 14224 11732 14272 11788
rect 14328 11732 14356 11788
rect 14036 10220 14356 11732
rect 18320 15708 18640 17220
rect 18320 15652 18348 15708
rect 18404 15652 18452 15708
rect 18508 15652 18556 15708
rect 18612 15652 18640 15708
rect 18320 14140 18640 15652
rect 18320 14084 18348 14140
rect 18404 14084 18452 14140
rect 18508 14084 18556 14140
rect 18612 14084 18640 14140
rect 18320 12572 18640 14084
rect 18320 12516 18348 12572
rect 18404 12516 18452 12572
rect 18508 12516 18556 12572
rect 18612 12516 18640 12572
rect 18320 11004 18640 12516
rect 18320 10948 18348 11004
rect 18404 10948 18452 11004
rect 18508 10948 18556 11004
rect 18612 10948 18640 11004
rect 14036 10164 14064 10220
rect 14120 10164 14168 10220
rect 14224 10164 14272 10220
rect 14328 10164 14356 10220
rect 14036 8652 14356 10164
rect 15596 10612 15652 10622
rect 15596 9268 15652 10556
rect 15596 9202 15652 9212
rect 16492 10388 16548 10398
rect 14036 8596 14064 8652
rect 14120 8596 14168 8652
rect 14224 8596 14272 8652
rect 14328 8596 14356 8652
rect 14036 7084 14356 8596
rect 16492 8036 16548 10332
rect 16492 7970 16548 7980
rect 18320 9436 18640 10948
rect 18320 9380 18348 9436
rect 18404 9380 18452 9436
rect 18508 9380 18556 9436
rect 18612 9380 18640 9436
rect 14036 7028 14064 7084
rect 14120 7028 14168 7084
rect 14224 7028 14272 7084
rect 14328 7028 14356 7084
rect 14036 5516 14356 7028
rect 14036 5460 14064 5516
rect 14120 5460 14168 5516
rect 14224 5460 14272 5516
rect 14328 5460 14356 5516
rect 14036 3948 14356 5460
rect 14036 3892 14064 3948
rect 14120 3892 14168 3948
rect 14224 3892 14272 3948
rect 14328 3892 14356 3948
rect 14036 3076 14356 3892
rect 18320 7868 18640 9380
rect 18320 7812 18348 7868
rect 18404 7812 18452 7868
rect 18508 7812 18556 7868
rect 18612 7812 18640 7868
rect 18320 6300 18640 7812
rect 18320 6244 18348 6300
rect 18404 6244 18452 6300
rect 18508 6244 18556 6300
rect 18612 6244 18640 6300
rect 18320 4732 18640 6244
rect 18320 4676 18348 4732
rect 18404 4676 18452 4732
rect 18508 4676 18556 4732
rect 18612 4676 18640 4732
rect 18320 3164 18640 4676
rect 18320 3108 18348 3164
rect 18404 3108 18452 3164
rect 18508 3108 18556 3164
rect 18612 3108 18640 3164
rect 18320 3076 18640 3108
rect 22604 24332 22924 25844
rect 22604 24276 22632 24332
rect 22688 24276 22736 24332
rect 22792 24276 22840 24332
rect 22896 24276 22924 24332
rect 22604 22764 22924 24276
rect 26888 32956 27208 33772
rect 26888 32900 26916 32956
rect 26972 32900 27020 32956
rect 27076 32900 27124 32956
rect 27180 32900 27208 32956
rect 26888 31388 27208 32900
rect 26888 31332 26916 31388
rect 26972 31332 27020 31388
rect 27076 31332 27124 31388
rect 27180 31332 27208 31388
rect 26888 29820 27208 31332
rect 26888 29764 26916 29820
rect 26972 29764 27020 29820
rect 27076 29764 27124 29820
rect 27180 29764 27208 29820
rect 26888 28252 27208 29764
rect 31172 33740 31492 33772
rect 31172 33684 31200 33740
rect 31256 33684 31304 33740
rect 31360 33684 31408 33740
rect 31464 33684 31492 33740
rect 31172 32172 31492 33684
rect 31172 32116 31200 32172
rect 31256 32116 31304 32172
rect 31360 32116 31408 32172
rect 31464 32116 31492 32172
rect 31172 30604 31492 32116
rect 35456 32956 35776 33772
rect 35456 32900 35484 32956
rect 35540 32900 35588 32956
rect 35644 32900 35692 32956
rect 35748 32900 35776 32956
rect 35456 31388 35776 32900
rect 35456 31332 35484 31388
rect 35540 31332 35588 31388
rect 35644 31332 35692 31388
rect 35748 31332 35776 31388
rect 31172 30548 31200 30604
rect 31256 30548 31304 30604
rect 31360 30548 31408 30604
rect 31464 30548 31492 30604
rect 31172 29036 31492 30548
rect 31172 28980 31200 29036
rect 31256 28980 31304 29036
rect 31360 28980 31408 29036
rect 31464 28980 31492 29036
rect 27580 28532 27636 28542
rect 26888 28196 26916 28252
rect 26972 28196 27020 28252
rect 27076 28196 27124 28252
rect 27180 28196 27208 28252
rect 26888 26684 27208 28196
rect 26888 26628 26916 26684
rect 26972 26628 27020 26684
rect 27076 26628 27124 26684
rect 27180 26628 27208 26684
rect 26888 25116 27208 26628
rect 26888 25060 26916 25116
rect 26972 25060 27020 25116
rect 27076 25060 27124 25116
rect 27180 25060 27208 25116
rect 26236 23716 26292 23726
rect 22604 22708 22632 22764
rect 22688 22708 22736 22764
rect 22792 22708 22840 22764
rect 22896 22708 22924 22764
rect 22604 21196 22924 22708
rect 22604 21140 22632 21196
rect 22688 21140 22736 21196
rect 22792 21140 22840 21196
rect 22896 21140 22924 21196
rect 22604 19628 22924 21140
rect 22604 19572 22632 19628
rect 22688 19572 22736 19628
rect 22792 19572 22840 19628
rect 22896 19572 22924 19628
rect 22604 18060 22924 19572
rect 25228 23044 25284 23054
rect 25228 19348 25284 22988
rect 26236 22820 26292 23660
rect 26236 20244 26292 22764
rect 26888 23548 27208 25060
rect 26888 23492 26916 23548
rect 26972 23492 27020 23548
rect 27076 23492 27124 23548
rect 27180 23492 27208 23548
rect 26684 22036 26740 22046
rect 26684 21476 26740 21980
rect 26684 21410 26740 21420
rect 26888 21980 27208 23492
rect 26888 21924 26916 21980
rect 26972 21924 27020 21980
rect 27076 21924 27124 21980
rect 27180 21924 27208 21980
rect 26888 20412 27208 21924
rect 26236 20178 26292 20188
rect 26684 20356 26740 20366
rect 25228 19282 25284 19292
rect 25564 19796 25620 19806
rect 22604 18004 22632 18060
rect 22688 18004 22736 18060
rect 22792 18004 22840 18060
rect 22896 18004 22924 18060
rect 22604 16492 22924 18004
rect 22604 16436 22632 16492
rect 22688 16436 22736 16492
rect 22792 16436 22840 16492
rect 22896 16436 22924 16492
rect 22604 14924 22924 16436
rect 25564 17108 25620 19740
rect 26124 18676 26180 18686
rect 26572 18676 26628 18686
rect 26180 18620 26572 18658
rect 26124 18602 26628 18620
rect 26572 18452 26628 18462
rect 25564 15204 25620 17052
rect 25788 17780 25844 17790
rect 25788 16772 25844 17724
rect 25788 16706 25844 16716
rect 26572 16660 26628 18396
rect 26684 16772 26740 20300
rect 26684 16706 26740 16716
rect 26888 20356 26916 20412
rect 26972 20356 27020 20412
rect 27076 20356 27124 20412
rect 27180 20356 27208 20412
rect 26888 18844 27208 20356
rect 26888 18788 26916 18844
rect 26972 18788 27020 18844
rect 27076 18788 27124 18844
rect 27180 18788 27208 18844
rect 26888 17276 27208 18788
rect 27356 28308 27412 28318
rect 27356 18452 27412 28252
rect 27356 18386 27412 18396
rect 27580 18452 27636 28476
rect 31172 27468 31492 28980
rect 31172 27412 31200 27468
rect 31256 27412 31304 27468
rect 31360 27412 31408 27468
rect 31464 27412 31492 27468
rect 31172 25900 31492 27412
rect 31172 25844 31200 25900
rect 31256 25844 31304 25900
rect 31360 25844 31408 25900
rect 31464 25844 31492 25900
rect 31172 24332 31492 25844
rect 31172 24276 31200 24332
rect 31256 24276 31304 24332
rect 31360 24276 31408 24332
rect 31464 24276 31492 24332
rect 27580 18386 27636 18396
rect 28028 22820 28084 22830
rect 28028 17444 28084 22764
rect 31172 22764 31492 24276
rect 31172 22708 31200 22764
rect 31256 22708 31304 22764
rect 31360 22708 31408 22764
rect 31464 22708 31492 22764
rect 28476 22036 28532 22046
rect 28476 21140 28532 21980
rect 28476 21074 28532 21084
rect 31172 21196 31492 22708
rect 33068 31108 33124 31118
rect 33068 22372 33124 31052
rect 34636 29988 34692 29998
rect 34188 25844 34244 25854
rect 34188 24948 34244 25788
rect 34188 24882 34244 24892
rect 33068 22306 33124 22316
rect 31172 21140 31200 21196
rect 31256 21140 31304 21196
rect 31360 21140 31408 21196
rect 31464 21140 31492 21196
rect 28252 21028 28308 21038
rect 28252 20132 28308 20972
rect 28252 19348 28308 20076
rect 28252 19282 28308 19292
rect 31172 19628 31492 21140
rect 31172 19572 31200 19628
rect 31256 19572 31304 19628
rect 31360 19572 31408 19628
rect 31464 19572 31492 19628
rect 28028 17378 28084 17388
rect 28140 18228 28196 18238
rect 26888 17220 26916 17276
rect 26972 17220 27020 17276
rect 27076 17220 27124 17276
rect 27180 17220 27208 17276
rect 25564 15138 25620 15148
rect 26348 15652 26404 15662
rect 26348 15204 26404 15596
rect 26348 15138 26404 15148
rect 26572 15092 26628 16604
rect 26572 15026 26628 15036
rect 26684 15876 26740 15886
rect 22604 14868 22632 14924
rect 22688 14868 22736 14924
rect 22792 14868 22840 14924
rect 22896 14868 22924 14924
rect 22604 13356 22924 14868
rect 26684 13972 26740 15820
rect 26684 13906 26740 13916
rect 26888 15708 27208 17220
rect 26888 15652 26916 15708
rect 26972 15652 27020 15708
rect 27076 15652 27124 15708
rect 27180 15652 27208 15708
rect 26888 14140 27208 15652
rect 27692 16772 27748 16782
rect 27692 14868 27748 16716
rect 27692 14802 27748 14812
rect 27804 15316 27860 15326
rect 26888 14084 26916 14140
rect 26972 14084 27020 14140
rect 27076 14084 27124 14140
rect 27180 14084 27208 14140
rect 22604 13300 22632 13356
rect 22688 13300 22736 13356
rect 22792 13300 22840 13356
rect 22896 13300 22924 13356
rect 22604 11788 22924 13300
rect 22604 11732 22632 11788
rect 22688 11732 22736 11788
rect 22792 11732 22840 11788
rect 22896 11732 22924 11788
rect 22604 10220 22924 11732
rect 22604 10164 22632 10220
rect 22688 10164 22736 10220
rect 22792 10164 22840 10220
rect 22896 10164 22924 10220
rect 22604 8652 22924 10164
rect 22604 8596 22632 8652
rect 22688 8596 22736 8652
rect 22792 8596 22840 8652
rect 22896 8596 22924 8652
rect 22604 7084 22924 8596
rect 22604 7028 22632 7084
rect 22688 7028 22736 7084
rect 22792 7028 22840 7084
rect 22896 7028 22924 7084
rect 22604 5516 22924 7028
rect 22604 5460 22632 5516
rect 22688 5460 22736 5516
rect 22792 5460 22840 5516
rect 22896 5460 22924 5516
rect 22604 3948 22924 5460
rect 22604 3892 22632 3948
rect 22688 3892 22736 3948
rect 22792 3892 22840 3948
rect 22896 3892 22924 3948
rect 22604 3076 22924 3892
rect 26888 12572 27208 14084
rect 27804 12964 27860 15260
rect 27804 12898 27860 12908
rect 28140 12964 28196 18172
rect 31172 18060 31492 19572
rect 34636 22148 34692 29932
rect 35456 29820 35776 31332
rect 35456 29764 35484 29820
rect 35540 29764 35588 29820
rect 35644 29764 35692 29820
rect 35748 29764 35776 29820
rect 35084 29428 35140 29438
rect 35084 24836 35140 29372
rect 35084 24770 35140 24780
rect 35456 28252 35776 29764
rect 35456 28196 35484 28252
rect 35540 28196 35588 28252
rect 35644 28196 35692 28252
rect 35748 28196 35776 28252
rect 35456 26684 35776 28196
rect 35456 26628 35484 26684
rect 35540 26628 35588 26684
rect 35644 26628 35692 26684
rect 35748 26628 35776 26684
rect 35456 25116 35776 26628
rect 35456 25060 35484 25116
rect 35540 25060 35588 25116
rect 35644 25060 35692 25116
rect 35748 25060 35776 25116
rect 35456 23548 35776 25060
rect 35456 23492 35484 23548
rect 35540 23492 35588 23548
rect 35644 23492 35692 23548
rect 35748 23492 35776 23548
rect 34748 23380 34804 23390
rect 34748 22596 34804 23324
rect 34748 22530 34804 22540
rect 31172 18004 31200 18060
rect 31256 18004 31304 18060
rect 31360 18004 31408 18060
rect 31464 18004 31492 18060
rect 28476 16660 28532 16670
rect 28252 15316 28308 15326
rect 28252 13860 28308 15260
rect 28476 15092 28532 16604
rect 28476 15026 28532 15036
rect 31172 16492 31492 18004
rect 31172 16436 31200 16492
rect 31256 16436 31304 16492
rect 31360 16436 31408 16492
rect 31464 16436 31492 16492
rect 28252 13794 28308 13804
rect 31172 14924 31492 16436
rect 31172 14868 31200 14924
rect 31256 14868 31304 14924
rect 31360 14868 31408 14924
rect 31464 14868 31492 14924
rect 28140 12898 28196 12908
rect 31172 13356 31492 14868
rect 31172 13300 31200 13356
rect 31256 13300 31304 13356
rect 31360 13300 31408 13356
rect 31464 13300 31492 13356
rect 26888 12516 26916 12572
rect 26972 12516 27020 12572
rect 27076 12516 27124 12572
rect 27180 12516 27208 12572
rect 26888 11004 27208 12516
rect 26888 10948 26916 11004
rect 26972 10948 27020 11004
rect 27076 10948 27124 11004
rect 27180 10948 27208 11004
rect 26888 9436 27208 10948
rect 26888 9380 26916 9436
rect 26972 9380 27020 9436
rect 27076 9380 27124 9436
rect 27180 9380 27208 9436
rect 26888 7868 27208 9380
rect 26888 7812 26916 7868
rect 26972 7812 27020 7868
rect 27076 7812 27124 7868
rect 27180 7812 27208 7868
rect 26888 6300 27208 7812
rect 31172 11788 31492 13300
rect 31172 11732 31200 11788
rect 31256 11732 31304 11788
rect 31360 11732 31408 11788
rect 31464 11732 31492 11788
rect 31172 10220 31492 11732
rect 31948 18564 32004 18574
rect 31948 11732 32004 18508
rect 32508 18004 32564 18014
rect 32172 14980 32228 14990
rect 32172 13188 32228 14924
rect 32508 14532 32564 17948
rect 32508 14466 32564 14476
rect 32172 13122 32228 13132
rect 31948 11666 32004 11676
rect 34636 11508 34692 22092
rect 35456 21980 35776 23492
rect 35456 21924 35484 21980
rect 35540 21924 35588 21980
rect 35644 21924 35692 21980
rect 35748 21924 35776 21980
rect 35456 20412 35776 21924
rect 35456 20356 35484 20412
rect 35540 20356 35588 20412
rect 35644 20356 35692 20412
rect 35748 20356 35776 20412
rect 35084 20020 35140 20030
rect 35084 17332 35140 19964
rect 35084 17266 35140 17276
rect 35456 18844 35776 20356
rect 35456 18788 35484 18844
rect 35540 18788 35588 18844
rect 35644 18788 35692 18844
rect 35748 18788 35776 18844
rect 35456 17276 35776 18788
rect 34636 11442 34692 11452
rect 34972 17220 35028 17230
rect 34972 15540 35028 17164
rect 34972 11396 35028 15484
rect 34972 11330 35028 11340
rect 35456 17220 35484 17276
rect 35540 17220 35588 17276
rect 35644 17220 35692 17276
rect 35748 17220 35776 17276
rect 35456 15708 35776 17220
rect 35456 15652 35484 15708
rect 35540 15652 35588 15708
rect 35644 15652 35692 15708
rect 35748 15652 35776 15708
rect 35456 14140 35776 15652
rect 35456 14084 35484 14140
rect 35540 14084 35588 14140
rect 35644 14084 35692 14140
rect 35748 14084 35776 14140
rect 35456 12572 35776 14084
rect 35456 12516 35484 12572
rect 35540 12516 35588 12572
rect 35644 12516 35692 12572
rect 35748 12516 35776 12572
rect 31172 10164 31200 10220
rect 31256 10164 31304 10220
rect 31360 10164 31408 10220
rect 31464 10164 31492 10220
rect 31172 8652 31492 10164
rect 31172 8596 31200 8652
rect 31256 8596 31304 8652
rect 31360 8596 31408 8652
rect 31464 8596 31492 8652
rect 26888 6244 26916 6300
rect 26972 6244 27020 6300
rect 27076 6244 27124 6300
rect 27180 6244 27208 6300
rect 26888 4732 27208 6244
rect 28028 7252 28084 7262
rect 28028 5348 28084 7196
rect 28028 5282 28084 5292
rect 31172 7084 31492 8596
rect 31172 7028 31200 7084
rect 31256 7028 31304 7084
rect 31360 7028 31408 7084
rect 31464 7028 31492 7084
rect 31172 5516 31492 7028
rect 31172 5460 31200 5516
rect 31256 5460 31304 5516
rect 31360 5460 31408 5516
rect 31464 5460 31492 5516
rect 26888 4676 26916 4732
rect 26972 4676 27020 4732
rect 27076 4676 27124 4732
rect 27180 4676 27208 4732
rect 26888 3164 27208 4676
rect 26888 3108 26916 3164
rect 26972 3108 27020 3164
rect 27076 3108 27124 3164
rect 27180 3108 27208 3164
rect 26888 3076 27208 3108
rect 31172 3948 31492 5460
rect 31172 3892 31200 3948
rect 31256 3892 31304 3948
rect 31360 3892 31408 3948
rect 31464 3892 31492 3948
rect 31172 3076 31492 3892
rect 35456 11004 35776 12516
rect 35456 10948 35484 11004
rect 35540 10948 35588 11004
rect 35644 10948 35692 11004
rect 35748 10948 35776 11004
rect 35456 9436 35776 10948
rect 35456 9380 35484 9436
rect 35540 9380 35588 9436
rect 35644 9380 35692 9436
rect 35748 9380 35776 9436
rect 35456 7868 35776 9380
rect 35456 7812 35484 7868
rect 35540 7812 35588 7868
rect 35644 7812 35692 7868
rect 35748 7812 35776 7868
rect 35456 6300 35776 7812
rect 35456 6244 35484 6300
rect 35540 6244 35588 6300
rect 35644 6244 35692 6300
rect 35748 6244 35776 6300
rect 35456 4732 35776 6244
rect 35456 4676 35484 4732
rect 35540 4676 35588 4732
rect 35644 4676 35692 4732
rect 35748 4676 35776 4732
rect 35456 3164 35776 4676
rect 35456 3108 35484 3164
rect 35540 3108 35588 3164
rect 35644 3108 35692 3164
rect 35748 3108 35776 3164
rect 35456 3076 35776 3108
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0511_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _0512_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30576 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0513_
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0514_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19264 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _0515_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24864 0 -1 15680
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0516_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20944 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0517_
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0518_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20048 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0519_
timestamp 1698431365
transform 1 0 32480 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0520_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20944 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  _0521_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21616 0 -1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _0522_
timestamp 1698431365
transform 1 0 23296 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0523_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32032 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0524_
timestamp 1698431365
transform -1 0 28224 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0525_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27216 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0526_
timestamp 1698431365
transform 1 0 23520 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0527_
timestamp 1698431365
transform 1 0 23856 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0528_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  _0529_
timestamp 1698431365
transform -1 0 24864 0 1 15680
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0530_
timestamp 1698431365
transform -1 0 20944 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0531_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26544 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0532_
timestamp 1698431365
transform -1 0 34496 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0533_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23744 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0534_
timestamp 1698431365
transform 1 0 26992 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0535_
timestamp 1698431365
transform 1 0 32256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0536_
timestamp 1698431365
transform 1 0 34496 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0537_
timestamp 1698431365
transform -1 0 34608 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0538_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 35392 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0539_
timestamp 1698431365
transform -1 0 34496 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0540_
timestamp 1698431365
transform -1 0 26992 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0541_
timestamp 1698431365
transform -1 0 32256 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0542_
timestamp 1698431365
transform -1 0 30016 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _0543_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 25872 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0544_
timestamp 1698431365
transform -1 0 34160 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _0545_
timestamp 1698431365
transform 1 0 17920 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0546_
timestamp 1698431365
transform -1 0 22512 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0547_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21504 0 1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _0548_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23072 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _0549_
timestamp 1698431365
transform 1 0 21728 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0550_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31248 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0551_
timestamp 1698431365
transform 1 0 26880 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0552_
timestamp 1698431365
transform 1 0 26880 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0553_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34160 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0554_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 34160 0 -1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0555_
timestamp 1698431365
transform -1 0 35280 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0556_
timestamp 1698431365
transform -1 0 32032 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0557_
timestamp 1698431365
transform -1 0 34832 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0558_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32480 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0559_
timestamp 1698431365
transform 1 0 24752 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0560_
timestamp 1698431365
transform -1 0 29456 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0561_
timestamp 1698431365
transform 1 0 29344 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0562_
timestamp 1698431365
transform 1 0 27776 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0563_
timestamp 1698431365
transform 1 0 34384 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0564_
timestamp 1698431365
transform -1 0 32592 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0565_
timestamp 1698431365
transform -1 0 31472 0 -1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0566_
timestamp 1698431365
transform 1 0 34160 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0567_
timestamp 1698431365
transform -1 0 34160 0 -1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0568_
timestamp 1698431365
transform 1 0 30128 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0569_
timestamp 1698431365
transform -1 0 28784 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0570_
timestamp 1698431365
transform 1 0 32704 0 1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0571_
timestamp 1698431365
transform -1 0 27776 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0572_
timestamp 1698431365
transform 1 0 24192 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0573_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26208 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0574_
timestamp 1698431365
transform 1 0 25984 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0575_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25984 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0576_
timestamp 1698431365
transform -1 0 25760 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0577_
timestamp 1698431365
transform 1 0 26432 0 1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0578_
timestamp 1698431365
transform -1 0 26320 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0579_
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0580_
timestamp 1698431365
transform -1 0 28784 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0581_
timestamp 1698431365
transform 1 0 26320 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0582_
timestamp 1698431365
transform 1 0 30464 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0583_
timestamp 1698431365
transform -1 0 29792 0 -1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0584_
timestamp 1698431365
transform 1 0 28672 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0585_
timestamp 1698431365
transform -1 0 28784 0 1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0586_
timestamp 1698431365
transform -1 0 32704 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0587_
timestamp 1698431365
transform -1 0 28784 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0588_
timestamp 1698431365
transform -1 0 28784 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0589_
timestamp 1698431365
transform -1 0 20272 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0590_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14448 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0591_
timestamp 1698431365
transform -1 0 14672 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0592_
timestamp 1698431365
transform -1 0 18368 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _0593_
timestamp 1698431365
transform -1 0 21616 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0594_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 25984 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0595_
timestamp 1698431365
transform -1 0 23520 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0596_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27104 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0597_
timestamp 1698431365
transform -1 0 35280 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0598_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28000 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0599_
timestamp 1698431365
transform -1 0 33824 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0600_
timestamp 1698431365
transform -1 0 28672 0 -1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0601_
timestamp 1698431365
transform 1 0 31584 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0602_
timestamp 1698431365
transform -1 0 31136 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0603_
timestamp 1698431365
transform 1 0 34496 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0604_
timestamp 1698431365
transform -1 0 27552 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0605_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28784 0 1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0606_
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0607_
timestamp 1698431365
transform -1 0 29792 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _0608_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33040 0 -1 23520
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0609_
timestamp 1698431365
transform -1 0 35392 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0610_
timestamp 1698431365
transform 1 0 34384 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0611_
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _0612_
timestamp 1698431365
transform -1 0 34832 0 -1 21952
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _0613_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30128 0 1 20384
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0614_
timestamp 1698431365
transform 1 0 30688 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0615_
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0616_
timestamp 1698431365
transform 1 0 28224 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0617_
timestamp 1698431365
transform -1 0 35056 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0618_
timestamp 1698431365
transform -1 0 32592 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0619_
timestamp 1698431365
transform -1 0 35392 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _0620_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32704 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0621_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32704 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0622_
timestamp 1698431365
transform -1 0 35168 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0623_
timestamp 1698431365
transform -1 0 30352 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _0624_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 34048 0 1 18816
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0625_
timestamp 1698431365
transform -1 0 29904 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0626_
timestamp 1698431365
transform -1 0 28448 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0627_
timestamp 1698431365
transform -1 0 30128 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0628_
timestamp 1698431365
transform -1 0 32704 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0629_
timestamp 1698431365
transform 1 0 26208 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0630_
timestamp 1698431365
transform -1 0 27328 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0631_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27328 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0632_
timestamp 1698431365
transform -1 0 28672 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0633_
timestamp 1698431365
transform -1 0 25984 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0634_
timestamp 1698431365
transform 1 0 26544 0 -1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0635_
timestamp 1698431365
transform 1 0 30016 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0636_
timestamp 1698431365
transform 1 0 28224 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0637_
timestamp 1698431365
transform -1 0 30800 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0638_
timestamp 1698431365
transform 1 0 21280 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0639_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _0640_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26208 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0641_
timestamp 1698431365
transform 1 0 18928 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _0642_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15904 0 1 15680
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0643_
timestamp 1698431365
transform -1 0 9184 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0644_
timestamp 1698431365
transform 1 0 11312 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0645_
timestamp 1698431365
transform -1 0 8512 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0646_
timestamp 1698431365
transform -1 0 9184 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0647_
timestamp 1698431365
transform 1 0 8288 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0648_
timestamp 1698431365
transform 1 0 6720 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0649_
timestamp 1698431365
transform -1 0 6496 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0650_
timestamp 1698431365
transform 1 0 7392 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0651_
timestamp 1698431365
transform 1 0 6496 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0652_
timestamp 1698431365
transform -1 0 28672 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0653_
timestamp 1698431365
transform -1 0 34496 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0654_
timestamp 1698431365
transform -1 0 26208 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0655_
timestamp 1698431365
transform 1 0 10640 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0656_
timestamp 1698431365
transform -1 0 13776 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0657_
timestamp 1698431365
transform 1 0 12096 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0658_
timestamp 1698431365
transform 1 0 11088 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0659_
timestamp 1698431365
transform -1 0 21280 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0660_
timestamp 1698431365
transform -1 0 23408 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0661_
timestamp 1698431365
transform -1 0 17920 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0662_
timestamp 1698431365
transform 1 0 11312 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0663_
timestamp 1698431365
transform 1 0 9184 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0664_
timestamp 1698431365
transform 1 0 15120 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0665_
timestamp 1698431365
transform -1 0 14000 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0666_
timestamp 1698431365
transform 1 0 12656 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0667_
timestamp 1698431365
transform -1 0 10080 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0668_
timestamp 1698431365
transform 1 0 5488 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0669_
timestamp 1698431365
transform 1 0 10640 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0670_
timestamp 1698431365
transform 1 0 13440 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0671_
timestamp 1698431365
transform 1 0 5488 0 1 3136
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0672_
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0673_
timestamp 1698431365
transform 1 0 13776 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0674_
timestamp 1698431365
transform -1 0 17024 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0675_
timestamp 1698431365
transform 1 0 14336 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0676_
timestamp 1698431365
transform 1 0 18592 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0677_
timestamp 1698431365
transform -1 0 19376 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0678_
timestamp 1698431365
transform 1 0 15792 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0679_
timestamp 1698431365
transform 1 0 15232 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0680_
timestamp 1698431365
transform 1 0 13104 0 1 3136
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0681_
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0682_
timestamp 1698431365
transform 1 0 16912 0 1 3136
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0683_
timestamp 1698431365
transform 1 0 18144 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0684_
timestamp 1698431365
transform 1 0 18704 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0685_
timestamp 1698431365
transform -1 0 22960 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0686_
timestamp 1698431365
transform 1 0 18144 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0687_
timestamp 1698431365
transform 1 0 19600 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0688_
timestamp 1698431365
transform -1 0 20272 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _0689_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23296 0 -1 20384
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0690_
timestamp 1698431365
transform -1 0 20944 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0691_
timestamp 1698431365
transform -1 0 16688 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0692_
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0693_
timestamp 1698431365
transform -1 0 20720 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0694_
timestamp 1698431365
transform -1 0 18816 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0695_
timestamp 1698431365
transform -1 0 18032 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0696_
timestamp 1698431365
transform -1 0 17360 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0697_
timestamp 1698431365
transform -1 0 16800 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0698_
timestamp 1698431365
transform -1 0 17472 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0699_
timestamp 1698431365
transform -1 0 24864 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0700_
timestamp 1698431365
transform -1 0 20048 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0701_
timestamp 1698431365
transform -1 0 20720 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0702_
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0703_
timestamp 1698431365
transform -1 0 15680 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0704_
timestamp 1698431365
transform 1 0 14000 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0705_
timestamp 1698431365
transform -1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0706_
timestamp 1698431365
transform -1 0 18704 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0707_
timestamp 1698431365
transform 1 0 15456 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0708_
timestamp 1698431365
transform 1 0 15456 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0709_
timestamp 1698431365
transform 1 0 13888 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0710_
timestamp 1698431365
transform -1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0711_
timestamp 1698431365
transform -1 0 21280 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0712_
timestamp 1698431365
transform 1 0 15680 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0713_
timestamp 1698431365
transform 1 0 15008 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0714_
timestamp 1698431365
transform 1 0 15568 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0715_
timestamp 1698431365
transform 1 0 14672 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0716_
timestamp 1698431365
transform -1 0 20832 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0717_
timestamp 1698431365
transform 1 0 20048 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0718_
timestamp 1698431365
transform -1 0 29568 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0719_
timestamp 1698431365
transform 1 0 21280 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0720_
timestamp 1698431365
transform 1 0 19152 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0721_
timestamp 1698431365
transform 1 0 21056 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0722_
timestamp 1698431365
transform -1 0 20944 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0723_
timestamp 1698431365
transform 1 0 19264 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0724_
timestamp 1698431365
transform -1 0 32032 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0725_
timestamp 1698431365
transform -1 0 22960 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0726_
timestamp 1698431365
transform 1 0 21280 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0727_
timestamp 1698431365
transform 1 0 22176 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0728_
timestamp 1698431365
transform 1 0 20384 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0729_
timestamp 1698431365
transform -1 0 32480 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0730_
timestamp 1698431365
transform -1 0 24304 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0731_
timestamp 1698431365
transform 1 0 22400 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0732_
timestamp 1698431365
transform -1 0 23968 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0733_
timestamp 1698431365
transform 1 0 22512 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0734_
timestamp 1698431365
transform -1 0 34272 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0735_
timestamp 1698431365
transform 1 0 24304 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0736_
timestamp 1698431365
transform 1 0 23968 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0737_
timestamp 1698431365
transform 1 0 15120 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0738_
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0739_
timestamp 1698431365
transform 1 0 24752 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0740_
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0741_
timestamp 1698431365
transform 1 0 26992 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0742_
timestamp 1698431365
transform -1 0 28784 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0743_
timestamp 1698431365
transform 1 0 26768 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0744_
timestamp 1698431365
transform 1 0 25312 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0745_
timestamp 1698431365
transform -1 0 28336 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0746_
timestamp 1698431365
transform 1 0 26992 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0747_
timestamp 1698431365
transform -1 0 27776 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0748_
timestamp 1698431365
transform -1 0 24752 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0749_
timestamp 1698431365
transform -1 0 27664 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0750_
timestamp 1698431365
transform 1 0 23968 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0751_
timestamp 1698431365
transform 1 0 23296 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0752_
timestamp 1698431365
transform -1 0 27104 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0753_
timestamp 1698431365
transform -1 0 25648 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0754_
timestamp 1698431365
transform 1 0 24416 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0755_
timestamp 1698431365
transform -1 0 25760 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0756_
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0757_
timestamp 1698431365
transform 1 0 25648 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0758_
timestamp 1698431365
transform -1 0 26880 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0759_
timestamp 1698431365
transform -1 0 26656 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0760_
timestamp 1698431365
transform -1 0 26208 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0761_
timestamp 1698431365
transform -1 0 28336 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0762_
timestamp 1698431365
transform 1 0 26880 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0763_
timestamp 1698431365
transform 1 0 26208 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0764_
timestamp 1698431365
transform 1 0 27776 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0765_
timestamp 1698431365
transform 1 0 26992 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0766_
timestamp 1698431365
transform 1 0 28112 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0767_
timestamp 1698431365
transform 1 0 27888 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0768_
timestamp 1698431365
transform 1 0 28336 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0769_
timestamp 1698431365
transform -1 0 29904 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0770_
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0771_
timestamp 1698431365
transform 1 0 31472 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0772_
timestamp 1698431365
transform 1 0 29904 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0773_
timestamp 1698431365
transform -1 0 31360 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0774_
timestamp 1698431365
transform 1 0 29680 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0775_
timestamp 1698431365
transform -1 0 31136 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0776_
timestamp 1698431365
transform -1 0 31472 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0777_
timestamp 1698431365
transform 1 0 29120 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0778_
timestamp 1698431365
transform -1 0 30240 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0779_
timestamp 1698431365
transform 1 0 31248 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0780_
timestamp 1698431365
transform 1 0 30464 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0781_
timestamp 1698431365
transform 1 0 32144 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0782_
timestamp 1698431365
transform 1 0 30352 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0783_
timestamp 1698431365
transform -1 0 13552 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0784_
timestamp 1698431365
transform 1 0 30688 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0785_
timestamp 1698431365
transform -1 0 30464 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0786_
timestamp 1698431365
transform -1 0 34944 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0787_
timestamp 1698431365
transform -1 0 35280 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0788_
timestamp 1698431365
transform -1 0 33824 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0789_
timestamp 1698431365
transform -1 0 34720 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0790_
timestamp 1698431365
transform -1 0 32704 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0791_
timestamp 1698431365
transform -1 0 20944 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _0792_
timestamp 1698431365
transform 1 0 20944 0 -1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0793_
timestamp 1698431365
transform 1 0 19264 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0794_
timestamp 1698431365
transform -1 0 25872 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0795_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22288 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0796_
timestamp 1698431365
transform 1 0 9968 0 -1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0797_
timestamp 1698431365
transform -1 0 16576 0 -1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0798_
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0799_
timestamp 1698431365
transform 1 0 19376 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0800_
timestamp 1698431365
transform 1 0 22400 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0801_
timestamp 1698431365
transform -1 0 20944 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0802_
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0803_
timestamp 1698431365
transform -1 0 20272 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0804_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21504 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0805_
timestamp 1698431365
transform -1 0 17360 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0806_
timestamp 1698431365
transform -1 0 14784 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _0807_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21280 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0808_
timestamp 1698431365
transform -1 0 27104 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0809_
timestamp 1698431365
transform 1 0 17920 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0810_
timestamp 1698431365
transform 1 0 23296 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0811_
timestamp 1698431365
transform -1 0 13776 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0812_
timestamp 1698431365
transform 1 0 12432 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0813_
timestamp 1698431365
transform -1 0 23408 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0814_
timestamp 1698431365
transform -1 0 28896 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0815_
timestamp 1698431365
transform 1 0 27216 0 1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0816_
timestamp 1698431365
transform -1 0 29456 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0817_
timestamp 1698431365
transform -1 0 31472 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0818_
timestamp 1698431365
transform 1 0 14672 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0819_
timestamp 1698431365
transform 1 0 23296 0 1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0820_
timestamp 1698431365
transform 1 0 9632 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0821_
timestamp 1698431365
transform 1 0 19152 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0822_
timestamp 1698431365
transform 1 0 23296 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0823_
timestamp 1698431365
transform -1 0 21616 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0824_
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0825_
timestamp 1698431365
transform -1 0 22064 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0826_
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0827_
timestamp 1698431365
transform -1 0 30464 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0828_
timestamp 1698431365
transform 1 0 31584 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0829_
timestamp 1698431365
transform 1 0 30464 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0830_
timestamp 1698431365
transform -1 0 24864 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0831_
timestamp 1698431365
transform -1 0 32032 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0832_
timestamp 1698431365
transform 1 0 27664 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0833_
timestamp 1698431365
transform -1 0 32032 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0834_
timestamp 1698431365
transform 1 0 26096 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0835_
timestamp 1698431365
transform 1 0 25760 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0836_
timestamp 1698431365
transform -1 0 9184 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0837_
timestamp 1698431365
transform 1 0 9632 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0838_
timestamp 1698431365
transform 1 0 8288 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0839_
timestamp 1698431365
transform -1 0 8736 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0840_
timestamp 1698431365
transform 1 0 7280 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0841_
timestamp 1698431365
transform -1 0 8400 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0842_
timestamp 1698431365
transform 1 0 7168 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0843_
timestamp 1698431365
transform -1 0 9968 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0844_
timestamp 1698431365
transform -1 0 9296 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0845_
timestamp 1698431365
transform -1 0 8960 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0846_
timestamp 1698431365
transform -1 0 7616 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0847_
timestamp 1698431365
transform -1 0 7168 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0848_
timestamp 1698431365
transform -1 0 12992 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0849_
timestamp 1698431365
transform 1 0 6384 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0850_
timestamp 1698431365
transform -1 0 8176 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0851_
timestamp 1698431365
transform -1 0 10640 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0852_
timestamp 1698431365
transform -1 0 7504 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0853_
timestamp 1698431365
transform 1 0 7056 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0854_
timestamp 1698431365
transform 1 0 9072 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0855_
timestamp 1698431365
transform 1 0 8624 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0856_
timestamp 1698431365
transform 1 0 7952 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0857_
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0858_
timestamp 1698431365
transform -1 0 11872 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0859_
timestamp 1698431365
transform 1 0 10192 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0860_
timestamp 1698431365
transform 1 0 10864 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0861_
timestamp 1698431365
transform 1 0 11648 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0862_
timestamp 1698431365
transform 1 0 11760 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0863_
timestamp 1698431365
transform -1 0 14000 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0864_
timestamp 1698431365
transform 1 0 11312 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0865_
timestamp 1698431365
transform 1 0 10752 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0866_
timestamp 1698431365
transform -1 0 13328 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0867_
timestamp 1698431365
transform -1 0 13664 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0868_
timestamp 1698431365
transform -1 0 13104 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0869_
timestamp 1698431365
transform -1 0 15456 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0870_
timestamp 1698431365
transform -1 0 14000 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0871_
timestamp 1698431365
transform -1 0 12656 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0872_
timestamp 1698431365
transform 1 0 12208 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0873_
timestamp 1698431365
transform -1 0 14784 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0874_
timestamp 1698431365
transform 1 0 12544 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0875_
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0876_
timestamp 1698431365
transform -1 0 16240 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0877_
timestamp 1698431365
transform 1 0 14000 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0878_
timestamp 1698431365
transform 1 0 14448 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0879_
timestamp 1698431365
transform 1 0 14896 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0880_
timestamp 1698431365
transform 1 0 15792 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0881_
timestamp 1698431365
transform -1 0 17920 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0882_
timestamp 1698431365
transform 1 0 16464 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0883_
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0884_
timestamp 1698431365
transform -1 0 18704 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0885_
timestamp 1698431365
transform 1 0 15792 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0886_
timestamp 1698431365
transform 1 0 16352 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0887_
timestamp 1698431365
transform -1 0 19152 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0888_
timestamp 1698431365
transform -1 0 18480 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0889_
timestamp 1698431365
transform -1 0 18592 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0890_
timestamp 1698431365
transform -1 0 19488 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0891_
timestamp 1698431365
transform 1 0 19152 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0892_
timestamp 1698431365
transform -1 0 17920 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0893_
timestamp 1698431365
transform -1 0 18144 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _0894_
timestamp 1698431365
transform -1 0 22176 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0895_
timestamp 1698431365
transform -1 0 16912 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0896_
timestamp 1698431365
transform -1 0 15456 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0897_
timestamp 1698431365
transform 1 0 6832 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0898_
timestamp 1698431365
transform -1 0 16352 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0899_
timestamp 1698431365
transform -1 0 19264 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0900_
timestamp 1698431365
transform 1 0 8176 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0901_
timestamp 1698431365
transform -1 0 8736 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0902_
timestamp 1698431365
transform 1 0 12432 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0903_
timestamp 1698431365
transform -1 0 14112 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0904_
timestamp 1698431365
transform 1 0 6720 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0905_
timestamp 1698431365
transform -1 0 6160 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0906_
timestamp 1698431365
transform -1 0 8176 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0907_
timestamp 1698431365
transform -1 0 8288 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0908_
timestamp 1698431365
transform -1 0 10080 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0909_
timestamp 1698431365
transform 1 0 6496 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0910_
timestamp 1698431365
transform -1 0 7840 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0911_
timestamp 1698431365
transform 1 0 7056 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0912_
timestamp 1698431365
transform -1 0 7392 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0913_
timestamp 1698431365
transform -1 0 11200 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0914_
timestamp 1698431365
transform -1 0 17024 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0915_
timestamp 1698431365
transform 1 0 6272 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0916_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6944 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0917_
timestamp 1698431365
transform 1 0 8176 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0918_
timestamp 1698431365
transform -1 0 12432 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0919_
timestamp 1698431365
transform 1 0 8176 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0920_
timestamp 1698431365
transform -1 0 10528 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0921_
timestamp 1698431365
transform -1 0 5936 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0922_
timestamp 1698431365
transform 1 0 8288 0 -1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0923_
timestamp 1698431365
transform -1 0 17920 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0924_
timestamp 1698431365
transform -1 0 11312 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0925_
timestamp 1698431365
transform -1 0 12768 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0926_
timestamp 1698431365
transform 1 0 7056 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0927_
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0928_
timestamp 1698431365
transform -1 0 10192 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0929_
timestamp 1698431365
transform -1 0 8400 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0930_
timestamp 1698431365
transform -1 0 11872 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0931_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10528 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0932_
timestamp 1698431365
transform 1 0 7616 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0933_
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0934_
timestamp 1698431365
transform -1 0 10416 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0935_
timestamp 1698431365
transform -1 0 9856 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0936_
timestamp 1698431365
transform -1 0 13328 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0937_
timestamp 1698431365
transform 1 0 10976 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0938_
timestamp 1698431365
transform -1 0 11536 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0939_
timestamp 1698431365
transform 1 0 11200 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0940_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9744 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0941_
timestamp 1698431365
transform 1 0 6160 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0942_
timestamp 1698431365
transform -1 0 6720 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0943_
timestamp 1698431365
transform 1 0 12096 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0944_
timestamp 1698431365
transform 1 0 11760 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0945_
timestamp 1698431365
transform 1 0 12096 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0946_
timestamp 1698431365
transform 1 0 12544 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0947_
timestamp 1698431365
transform 1 0 11984 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0948_
timestamp 1698431365
transform -1 0 14896 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0949_
timestamp 1698431365
transform -1 0 14000 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0950_
timestamp 1698431365
transform -1 0 13104 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0951_
timestamp 1698431365
transform 1 0 13328 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0952_
timestamp 1698431365
transform -1 0 13888 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0953_
timestamp 1698431365
transform -1 0 14112 0 -1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0954_
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0955_
timestamp 1698431365
transform -1 0 12992 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0956_
timestamp 1698431365
transform -1 0 18928 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0957_
timestamp 1698431365
transform 1 0 14784 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0958_
timestamp 1698431365
transform 1 0 15232 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0959_
timestamp 1698431365
transform 1 0 17472 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _0960_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17024 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _0961_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0962_
timestamp 1698431365
transform -1 0 19600 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0963_
timestamp 1698431365
transform 1 0 14672 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0964_
timestamp 1698431365
transform 1 0 17360 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0965_
timestamp 1698431365
transform 1 0 15680 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0966_
timestamp 1698431365
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0967_
timestamp 1698431365
transform 1 0 18480 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0968_
timestamp 1698431365
transform -1 0 17472 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0969_
timestamp 1698431365
transform 1 0 16352 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0970_
timestamp 1698431365
transform -1 0 19152 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0971_
timestamp 1698431365
transform -1 0 17920 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0972_
timestamp 1698431365
transform -1 0 15680 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0973_
timestamp 1698431365
transform -1 0 15792 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0974_
timestamp 1698431365
transform -1 0 15568 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0975_
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0976_
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0977_
timestamp 1698431365
transform 1 0 19824 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0978_
timestamp 1698431365
transform 1 0 19488 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0979_
timestamp 1698431365
transform 1 0 18032 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0980_
timestamp 1698431365
transform -1 0 19152 0 -1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0981_
timestamp 1698431365
transform 1 0 18704 0 1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0982_
timestamp 1698431365
transform 1 0 20272 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0983_
timestamp 1698431365
transform 1 0 22512 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0984_
timestamp 1698431365
transform -1 0 25648 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0985_
timestamp 1698431365
transform -1 0 24640 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0986_
timestamp 1698431365
transform 1 0 19712 0 1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0987_
timestamp 1698431365
transform -1 0 20832 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0988_
timestamp 1698431365
transform -1 0 21952 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0989_
timestamp 1698431365
transform 1 0 17248 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0990_
timestamp 1698431365
transform -1 0 19040 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0991_
timestamp 1698431365
transform 1 0 21392 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0992_
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0993_
timestamp 1698431365
transform -1 0 28672 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0994_
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0995_
timestamp 1698431365
transform 1 0 20048 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0996_
timestamp 1698431365
transform 1 0 20272 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0997_
timestamp 1698431365
transform -1 0 22848 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _0998_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19040 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0999_
timestamp 1698431365
transform 1 0 19488 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1000_
timestamp 1698431365
transform 1 0 22960 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1001_
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1002_
timestamp 1698431365
transform -1 0 11536 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1003_
timestamp 1698431365
transform 1 0 10416 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1004_
timestamp 1698431365
transform 1 0 10080 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1005_
timestamp 1698431365
transform 1 0 11984 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1006_
timestamp 1698431365
transform 1 0 10304 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1007_
timestamp 1698431365
transform -1 0 10416 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1008_
timestamp 1698431365
transform -1 0 7952 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1009_
timestamp 1698431365
transform -1 0 9632 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1010_
timestamp 1698431365
transform -1 0 9968 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1011_
timestamp 1698431365
transform -1 0 10304 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1012_
timestamp 1698431365
transform -1 0 10864 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1013_
timestamp 1698431365
transform 1 0 8288 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1014_
timestamp 1698431365
transform 1 0 7952 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1015_
timestamp 1698431365
transform -1 0 9744 0 1 3136
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1016_
timestamp 1698431365
transform 1 0 7840 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1017_
timestamp 1698431365
transform -1 0 7280 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1018_
timestamp 1698431365
transform -1 0 10640 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1019_
timestamp 1698431365
transform 1 0 6944 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1020_
timestamp 1698431365
transform -1 0 6944 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1021_
timestamp 1698431365
transform 1 0 5824 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1022_
timestamp 1698431365
transform 1 0 7280 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1023_
timestamp 1698431365
transform 1 0 6384 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1024_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8736 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1025_
timestamp 1698431365
transform -1 0 7952 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1026_
timestamp 1698431365
transform -1 0 12880 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1027_
timestamp 1698431365
transform -1 0 12656 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1028_
timestamp 1698431365
transform 1 0 9744 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1029_
timestamp 1698431365
transform 1 0 11536 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1030_
timestamp 1698431365
transform -1 0 17024 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1031_
timestamp 1698431365
transform -1 0 17696 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1032_
timestamp 1698431365
transform 1 0 17696 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1033_
timestamp 1698431365
transform 1 0 19152 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1034_
timestamp 1698431365
transform -1 0 18144 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1035_
timestamp 1698431365
transform 1 0 11984 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1036_
timestamp 1698431365
transform 1 0 12208 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1037_
timestamp 1698431365
transform 1 0 13776 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1038_
timestamp 1698431365
transform 1 0 17808 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1039_
timestamp 1698431365
transform 1 0 19152 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1040_
timestamp 1698431365
transform 1 0 21504 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1041_
timestamp 1698431365
transform 1 0 23856 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1042_
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1043_
timestamp 1698431365
transform 1 0 21616 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1044_
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1045_
timestamp 1698431365
transform -1 0 31584 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1046_
timestamp 1698431365
transform 1 0 28896 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1047_
timestamp 1698431365
transform 1 0 31136 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1048_
timestamp 1698431365
transform 1 0 27104 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1049_
timestamp 1698431365
transform 1 0 29904 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1050_
timestamp 1698431365
transform 1 0 32032 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1051_
timestamp 1698431365
transform 1 0 29456 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1052_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23296 0 1 25088
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1053_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1054_
timestamp 1698431365
transform -1 0 32480 0 1 15680
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1055_
timestamp 1698431365
transform -1 0 30688 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1056_
timestamp 1698431365
transform -1 0 35392 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1057_
timestamp 1698431365
transform 1 0 29456 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1058_
timestamp 1698431365
transform -1 0 35392 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1059_
timestamp 1698431365
transform -1 0 35392 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1060_
timestamp 1698431365
transform -1 0 20048 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1061_
timestamp 1698431365
transform 1 0 13552 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1062_
timestamp 1698431365
transform 1 0 22736 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1063_
timestamp 1698431365
transform -1 0 26544 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1064_
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1065_
timestamp 1698431365
transform 1 0 19712 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1066_
timestamp 1698431365
transform 1 0 29008 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1067_
timestamp 1698431365
transform 1 0 27216 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1068_
timestamp 1698431365
transform 1 0 32144 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1069_
timestamp 1698431365
transform -1 0 30240 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1070_
timestamp 1698431365
transform 1 0 32144 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1071_
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1072_
timestamp 1698431365
transform 1 0 28224 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1073_
timestamp 1698431365
transform -1 0 27776 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1074_
timestamp 1698431365
transform 1 0 7168 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1075_
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1076_
timestamp 1698431365
transform 1 0 4816 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1077_
timestamp 1698431365
transform 1 0 3472 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1078_
timestamp 1698431365
transform 1 0 3808 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1079_
timestamp 1698431365
transform 1 0 7280 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1080_
timestamp 1698431365
transform 1 0 10304 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1081_
timestamp 1698431365
transform 1 0 9744 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1082_
timestamp 1698431365
transform 1 0 9296 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1083_
timestamp 1698431365
transform 1 0 9856 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1084_
timestamp 1698431365
transform 1 0 11760 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1085_
timestamp 1698431365
transform 1 0 13776 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1086_
timestamp 1698431365
transform 1 0 16352 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1087_
timestamp 1698431365
transform 1 0 13776 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1088_
timestamp 1698431365
transform -1 0 20944 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1089_
timestamp 1698431365
transform 1 0 15904 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1090_
timestamp 1698431365
transform 1 0 3360 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1091_
timestamp 1698431365
transform 1 0 4256 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1092_
timestamp 1698431365
transform 1 0 3696 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1093_
timestamp 1698431365
transform 1 0 5936 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1094_
timestamp 1698431365
transform 1 0 8400 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1095_
timestamp 1698431365
transform 1 0 3472 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1096_
timestamp 1698431365
transform 1 0 11872 0 -1 31360
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1097_
timestamp 1698431365
transform 1 0 12208 0 -1 32928
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1098_
timestamp 1698431365
transform 1 0 16800 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1099_
timestamp 1698431365
transform 1 0 17360 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1100_
timestamp 1698431365
transform 1 0 12992 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1101_
timestamp 1698431365
transform 1 0 20384 0 -1 32928
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1102_
timestamp 1698431365
transform 1 0 20720 0 1 32928
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1103_
timestamp 1698431365
transform 1 0 23184 0 1 31360
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1104_
timestamp 1698431365
transform 1 0 23520 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1105_
timestamp 1698431365
transform 1 0 23968 0 1 29792
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1106_
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1107_
timestamp 1698431365
transform -1 0 12656 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1108_
timestamp 1698431365
transform 1 0 6832 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1109_
timestamp 1698431365
transform 1 0 5936 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1110_
timestamp 1698431365
transform 1 0 5712 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1111_
timestamp 1698431365
transform -1 0 7280 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0524__I $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 27440 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0532__I
timestamp 1698431365
transform 1 0 35168 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0533__I
timestamp 1698431365
transform 1 0 23520 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0535__I
timestamp 1698431365
transform -1 0 22624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0537__I
timestamp 1698431365
transform -1 0 33712 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0545__A1
timestamp 1698431365
transform -1 0 18928 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0545__A2
timestamp 1698431365
transform 1 0 18816 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0555__I
timestamp 1698431365
transform 1 0 35168 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0557__I
timestamp 1698431365
transform -1 0 34160 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0562__A3
timestamp 1698431365
transform 1 0 34160 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0572__A1
timestamp 1698431365
transform -1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0574__A1
timestamp 1698431365
transform 1 0 25088 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0576__A1
timestamp 1698431365
transform 1 0 23632 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0578__A1
timestamp 1698431365
transform -1 0 24416 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0590__I
timestamp 1698431365
transform -1 0 14448 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0592__B
timestamp 1698431365
transform 1 0 16800 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0592__C
timestamp 1698431365
transform -1 0 17920 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0597__I
timestamp 1698431365
transform -1 0 34944 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0598__A1
timestamp 1698431365
transform 1 0 23296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0602__A1
timestamp 1698431365
transform 1 0 31808 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0608__C
timestamp 1698431365
transform -1 0 34720 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0611__A1
timestamp 1698431365
transform -1 0 34160 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0618__A2
timestamp 1698431365
transform -1 0 32816 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0619__A1
timestamp 1698431365
transform -1 0 34720 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0622__A2
timestamp 1698431365
transform 1 0 33488 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0623__A2
timestamp 1698431365
transform 1 0 21504 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0636__B
timestamp 1698431365
transform -1 0 29568 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0640__A1
timestamp 1698431365
transform 1 0 23744 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0641__A1
timestamp 1698431365
transform 1 0 21392 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0641__A2
timestamp 1698431365
transform 1 0 19824 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0642__A1
timestamp 1698431365
transform 1 0 18592 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0643__I
timestamp 1698431365
transform 1 0 9856 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0644__I
timestamp 1698431365
transform 1 0 12768 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0646__I
timestamp 1698431365
transform 1 0 9184 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0647__B
timestamp 1698431365
transform 1 0 8064 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0650__B
timestamp 1698431365
transform 1 0 8288 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0653__A2
timestamp 1698431365
transform 1 0 33488 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0654__A2
timestamp 1698431365
transform 1 0 21168 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0654__A3
timestamp 1698431365
transform -1 0 26656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0655__I
timestamp 1698431365
transform -1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0657__A2
timestamp 1698431365
transform 1 0 13552 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0658__A1
timestamp 1698431365
transform 1 0 11984 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0659__I
timestamp 1698431365
transform 1 0 21392 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0660__A3
timestamp 1698431365
transform 1 0 24080 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0661__I
timestamp 1698431365
transform 1 0 18256 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0664__I
timestamp 1698431365
transform 1 0 14896 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0674__I
timestamp 1698431365
transform 1 0 15680 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0677__I
timestamp 1698431365
transform -1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0679__A2
timestamp 1698431365
transform -1 0 15232 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0682__A2
timestamp 1698431365
transform 1 0 18928 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0685__A2
timestamp 1698431365
transform 1 0 23184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0689__A2
timestamp 1698431365
transform 1 0 23632 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0692__A1
timestamp 1698431365
transform -1 0 22960 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0692__A3
timestamp 1698431365
transform -1 0 23072 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0737__I
timestamp 1698431365
transform -1 0 16240 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0738__I
timestamp 1698431365
transform -1 0 25088 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0743__A1
timestamp 1698431365
transform -1 0 26880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0743__A3
timestamp 1698431365
transform -1 0 21840 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0763__I
timestamp 1698431365
transform 1 0 25984 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0783__I
timestamp 1698431365
transform 1 0 13776 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0784__B
timestamp 1698431365
transform 1 0 32256 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0794__A1
timestamp 1698431365
transform 1 0 24640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0813__B
timestamp 1698431365
transform 1 0 22288 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0818__A1
timestamp 1698431365
transform 1 0 15568 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0825__B
timestamp 1698431365
transform 1 0 20720 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0829__A1
timestamp 1698431365
transform 1 0 28560 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0830__A1
timestamp 1698431365
transform 1 0 24080 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0832__A1
timestamp 1698431365
transform 1 0 29232 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0837__B
timestamp 1698431365
transform 1 0 10752 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0838__A1
timestamp 1698431365
transform 1 0 9184 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0842__B
timestamp 1698431365
transform 1 0 8400 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0845__B
timestamp 1698431365
transform -1 0 10416 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0892__I
timestamp 1698431365
transform 1 0 18144 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0895__I
timestamp 1698431365
transform -1 0 17136 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0904__B
timestamp 1698431365
transform 1 0 8512 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0908__I
timestamp 1698431365
transform -1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0920__C
timestamp 1698431365
transform 1 0 11536 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0928__C
timestamp 1698431365
transform -1 0 9072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0934__C
timestamp 1698431365
transform -1 0 10976 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0936__I
timestamp 1698431365
transform 1 0 11088 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0941__B
timestamp 1698431365
transform 1 0 7392 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0951__I
timestamp 1698431365
transform 1 0 14448 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0961__C
timestamp 1698431365
transform -1 0 22736 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0968__A1
timestamp 1698431365
transform 1 0 16128 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0975__C
timestamp 1698431365
transform 1 0 14224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1000__B
timestamp 1698431365
transform 1 0 24080 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1001__C
timestamp 1698431365
transform 1 0 23184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1002__A1
timestamp 1698431365
transform 1 0 11760 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1003__B
timestamp 1698431365
transform 1 0 11424 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1006__B
timestamp 1698431365
transform 1 0 11872 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1008__I
timestamp 1698431365
transform 1 0 7952 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1009__I
timestamp 1698431365
transform -1 0 10416 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1011__I
timestamp 1698431365
transform 1 0 9408 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1012__I
timestamp 1698431365
transform 1 0 10864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1040__CLK
timestamp 1698431365
transform 1 0 23632 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1042__CLK
timestamp 1698431365
transform 1 0 26432 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1043__CLK
timestamp 1698431365
transform 1 0 28560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1052__CLK
timestamp 1698431365
transform 1 0 23072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1062__CLK
timestamp 1698431365
transform 1 0 26208 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1063__CLK
timestamp 1698431365
transform 1 0 24192 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1064__CLK
timestamp 1698431365
transform 1 0 23744 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1065__CLK
timestamp 1698431365
transform 1 0 23184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1074__CLK
timestamp 1698431365
transform -1 0 10864 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1075__CLK
timestamp 1698431365
transform 1 0 10528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1076__CLK
timestamp 1698431365
transform 1 0 6384 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1077__CLK
timestamp 1698431365
transform 1 0 8848 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1078__CLK
timestamp 1698431365
transform 1 0 6720 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1079__CLK
timestamp 1698431365
transform 1 0 10864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1080__CLK
timestamp 1698431365
transform 1 0 13776 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1081__CLK
timestamp 1698431365
transform 1 0 14224 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1082__CLK
timestamp 1698431365
transform 1 0 13552 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1083__CLK
timestamp 1698431365
transform -1 0 13328 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1084__CLK
timestamp 1698431365
transform 1 0 15232 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1085__CLK
timestamp 1698431365
transform 1 0 17024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1086__CLK
timestamp 1698431365
transform 1 0 16128 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1087__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1088__CLK
timestamp 1698431365
transform 1 0 21840 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1089__CLK
timestamp 1698431365
transform 1 0 15680 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1090__CLK
timestamp 1698431365
transform 1 0 7616 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1091__CLK
timestamp 1698431365
transform 1 0 8400 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1092__CLK
timestamp 1698431365
transform 1 0 6496 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1093__CLK
timestamp 1698431365
transform -1 0 10304 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1094__CLK
timestamp 1698431365
transform 1 0 11872 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1095__CLK
timestamp 1698431365
transform 1 0 6944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1096__CLK
timestamp 1698431365
transform 1 0 14224 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1097__CLK
timestamp 1698431365
transform 1 0 14224 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1098__CLK
timestamp 1698431365
transform 1 0 24528 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1099__CLK
timestamp 1698431365
transform 1 0 24080 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1100__CLK
timestamp 1698431365
transform 1 0 13776 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1101__CLK
timestamp 1698431365
transform 1 0 25872 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1102__CLK
timestamp 1698431365
transform 1 0 27552 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1103__CLK
timestamp 1698431365
transform 1 0 27328 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1104__CLK
timestamp 1698431365
transform 1 0 23296 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1105__CLK
timestamp 1698431365
transform 1 0 27664 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_i_I
timestamp 1698431365
transform 1 0 23072 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_0__f_clk_i_I
timestamp 1698431365
transform 1 0 15232 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_1__f_clk_i_I
timestamp 1698431365
transform -1 0 21616 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_2__f_clk_i_I
timestamp 1698431365
transform 1 0 14224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_3__f_clk_i_I
timestamp 1698431365
transform 1 0 19712 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_4__f_clk_i_I
timestamp 1698431365
transform 1 0 21392 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_5__f_clk_i_I
timestamp 1698431365
transform 1 0 27328 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_6__f_clk_i_I
timestamp 1698431365
transform -1 0 23856 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_7__f_clk_i_I
timestamp 1698431365
transform -1 0 29008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 33264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 33824 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 35392 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 33264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 33712 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 34048 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 34496 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 34272 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform -1 0 34720 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform -1 0 34720 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform 1 0 23744 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform 1 0 29792 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform 1 0 29792 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform 1 0 31024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform 1 0 31472 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform 1 0 32928 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform -1 0 33376 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform -1 0 34720 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output33_I
timestamp 1698431365
transform 1 0 32480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output35_I
timestamp 1698431365
transform 1 0 28672 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24528 0 -1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_0__f_clk_i
timestamp 1698431365
transform -1 0 15008 0 -1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_1__f_clk_i
timestamp 1698431365
transform 1 0 15120 0 1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_2__f_clk_i
timestamp 1698431365
transform -1 0 13104 0 1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_3__f_clk_i
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_4__f_clk_i
timestamp 1698431365
transform 1 0 21616 0 1 14112
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_5__f_clk_i
timestamp 1698431365
transform 1 0 26432 0 -1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_6__f_clk_i
timestamp 1698431365
transform 1 0 22624 0 1 28224
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_7__f_clk_i
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout58
timestamp 1698431365
transform -1 0 15232 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout59
timestamp 1698431365
transform 1 0 15680 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout60
timestamp 1698431365
transform 1 0 7616 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout61
timestamp 1698431365
transform -1 0 8400 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout62
timestamp 1698431365
transform -1 0 30688 0 -1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout63
timestamp 1698431365
transform 1 0 34608 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout64
timestamp 1698431365
transform -1 0 32256 0 -1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout65
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout66
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_6 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_36 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_75
timestamp 1698431365
transform 1 0 9744 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_252
timestamp 1698431365
transform 1 0 29568 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_256
timestamp 1698431365
transform 1 0 30016 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_263
timestamp 1698431365
transform 1 0 30800 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_267
timestamp 1698431365
transform 1 0 31248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_271
timestamp 1698431365
transform 1 0 31696 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_280
timestamp 1698431365
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_284
timestamp 1698431365
transform 1 0 33152 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_291
timestamp 1698431365
transform 1 0 33936 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_295
timestamp 1698431365
transform 1 0 34384 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_10
timestamp 1698431365
transform 1 0 2464 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_12
timestamp 1698431365
transform 1 0 2688 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_68
timestamp 1698431365
transform 1 0 8960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_109
timestamp 1698431365
transform 1 0 13552 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_155
timestamp 1698431365
transform 1 0 18704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_193
timestamp 1698431365
transform 1 0 22960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_197
timestamp 1698431365
transform 1 0 23408 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_199
timestamp 1698431365
transform 1 0 23632 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698431365
transform 1 0 32480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_286 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33376 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_302
timestamp 1698431365
transform 1 0 35168 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_4
timestamp 1698431365
transform 1 0 1792 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_31
timestamp 1698431365
transform 1 0 4816 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_104
timestamp 1698431365
transform 1 0 12992 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_115
timestamp 1698431365
transform 1 0 14224 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_226
timestamp 1698431365
transform 1 0 26656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_228
timestamp 1698431365
transform 1 0 26880 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_241
timestamp 1698431365
transform 1 0 28336 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_252
timestamp 1698431365
transform 1 0 29568 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_256 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30016 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_288
timestamp 1698431365
transform 1 0 33600 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_34
timestamp 1698431365
transform 1 0 5152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_36
timestamp 1698431365
transform 1 0 5376 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_42
timestamp 1698431365
transform 1 0 6048 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_120
timestamp 1698431365
transform 1 0 14784 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_137
timestamp 1698431365
transform 1 0 16688 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_139
timestamp 1698431365
transform 1 0 16912 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_199
timestamp 1698431365
transform 1 0 23632 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_201
timestamp 1698431365
transform 1 0 23856 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_244
timestamp 1698431365
transform 1 0 28672 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_275
timestamp 1698431365
transform 1 0 32144 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_279
timestamp 1698431365
transform 1 0 32592 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_298
timestamp 1698431365
transform 1 0 34720 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_302
timestamp 1698431365
transform 1 0 35168 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_171
timestamp 1698431365
transform 1 0 20496 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_222
timestamp 1698431365
transform 1 0 26208 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_226
timestamp 1698431365
transform 1 0 26656 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698431365
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_268
timestamp 1698431365
transform 1 0 31360 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_300
timestamp 1698431365
transform 1 0 34944 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_34
timestamp 1698431365
transform 1 0 5152 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_80
timestamp 1698431365
transform 1 0 10304 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_82
timestamp 1698431365
transform 1 0 10528 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_94
timestamp 1698431365
transform 1 0 11872 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_124
timestamp 1698431365
transform 1 0 15232 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_148
timestamp 1698431365
transform 1 0 17920 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_183
timestamp 1698431365
transform 1 0 21840 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_191
timestamp 1698431365
transform 1 0 22736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_195
timestamp 1698431365
transform 1 0 23184 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_209
timestamp 1698431365
transform 1 0 24752 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_222
timestamp 1698431365
transform 1 0 26208 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_246
timestamp 1698431365
transform 1 0 28896 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_277
timestamp 1698431365
transform 1 0 32368 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_279
timestamp 1698431365
transform 1 0 32592 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_294
timestamp 1698431365
transform 1 0 34272 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_39
timestamp 1698431365
transform 1 0 5712 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_61
timestamp 1698431365
transform 1 0 8176 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_70
timestamp 1698431365
transform 1 0 9184 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_103
timestamp 1698431365
transform 1 0 12880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_121
timestamp 1698431365
transform 1 0 14896 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_173
timestamp 1698431365
transform 1 0 20720 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_181
timestamp 1698431365
transform 1 0 21616 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_197
timestamp 1698431365
transform 1 0 23408 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_205
timestamp 1698431365
transform 1 0 24304 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_209
timestamp 1698431365
transform 1 0 24752 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_212
timestamp 1698431365
transform 1 0 25088 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_228
timestamp 1698431365
transform 1 0 26880 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_235
timestamp 1698431365
transform 1 0 27664 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_243
timestamp 1698431365
transform 1 0 28560 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_249
timestamp 1698431365
transform 1 0 29232 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_295
timestamp 1698431365
transform 1 0 34384 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_297
timestamp 1698431365
transform 1 0 34608 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_18
timestamp 1698431365
transform 1 0 3360 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_22
timestamp 1698431365
transform 1 0 3808 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_67
timestamp 1698431365
transform 1 0 8848 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_69
timestamp 1698431365
transform 1 0 9072 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_122
timestamp 1698431365
transform 1 0 15008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_126
timestamp 1698431365
transform 1 0 15456 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_138
timestamp 1698431365
transform 1 0 16800 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_156
timestamp 1698431365
transform 1 0 18816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_158
timestamp 1698431365
transform 1 0 19040 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_193
timestamp 1698431365
transform 1 0 22960 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_197
timestamp 1698431365
transform 1 0 23408 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_199
timestamp 1698431365
transform 1 0 23632 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_218
timestamp 1698431365
transform 1 0 25760 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_228
timestamp 1698431365
transform 1 0 26880 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_292
timestamp 1698431365
transform 1 0 34048 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_296
timestamp 1698431365
transform 1 0 34496 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_300
timestamp 1698431365
transform 1 0 34944 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_45
timestamp 1698431365
transform 1 0 6384 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_78
timestamp 1698431365
transform 1 0 10080 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_85
timestamp 1698431365
transform 1 0 10864 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_95
timestamp 1698431365
transform 1 0 11984 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_104
timestamp 1698431365
transform 1 0 12992 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_111
timestamp 1698431365
transform 1 0 13776 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_149
timestamp 1698431365
transform 1 0 18032 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_153
timestamp 1698431365
transform 1 0 18480 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_161
timestamp 1698431365
transform 1 0 19376 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_165
timestamp 1698431365
transform 1 0 19824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_173
timestamp 1698431365
transform 1 0 20720 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_185
timestamp 1698431365
transform 1 0 22064 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_187
timestamp 1698431365
transform 1 0 22288 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_196
timestamp 1698431365
transform 1 0 23296 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_200
timestamp 1698431365
transform 1 0 23744 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_230
timestamp 1698431365
transform 1 0 27104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_234
timestamp 1698431365
transform 1 0 27552 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_238
timestamp 1698431365
transform 1 0 28000 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_249
timestamp 1698431365
transform 1 0 29232 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_268
timestamp 1698431365
transform 1 0 31360 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_276
timestamp 1698431365
transform 1 0 32256 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_278
timestamp 1698431365
transform 1 0 32480 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_281
timestamp 1698431365
transform 1 0 32816 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_285
timestamp 1698431365
transform 1 0 33264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_289
timestamp 1698431365
transform 1 0 33712 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_293
timestamp 1698431365
transform 1 0 34160 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_295
timestamp 1698431365
transform 1 0 34384 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_34
timestamp 1698431365
transform 1 0 5152 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_50
timestamp 1698431365
transform 1 0 6944 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_58
timestamp 1698431365
transform 1 0 7840 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_61
timestamp 1698431365
transform 1 0 8176 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_69
timestamp 1698431365
transform 1 0 9072 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_77
timestamp 1698431365
transform 1 0 9968 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_81
timestamp 1698431365
transform 1 0 10416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_87
timestamp 1698431365
transform 1 0 11088 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_134
timestamp 1698431365
transform 1 0 16352 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_138
timestamp 1698431365
transform 1 0 16800 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_158
timestamp 1698431365
transform 1 0 19040 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_166
timestamp 1698431365
transform 1 0 19936 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_220
timestamp 1698431365
transform 1 0 25984 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_226
timestamp 1698431365
transform 1 0 26656 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_230
timestamp 1698431365
transform 1 0 27104 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_270
timestamp 1698431365
transform 1 0 31584 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_274
timestamp 1698431365
transform 1 0 32032 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_278
timestamp 1698431365
transform 1 0 32480 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_286
timestamp 1698431365
transform 1 0 33376 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_303
timestamp 1698431365
transform 1 0 35280 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_66
timestamp 1698431365
transform 1 0 8736 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_74
timestamp 1698431365
transform 1 0 9632 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_78
timestamp 1698431365
transform 1 0 10080 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_88
timestamp 1698431365
transform 1 0 11200 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_92
timestamp 1698431365
transform 1 0 11648 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_96
timestamp 1698431365
transform 1 0 12096 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_104
timestamp 1698431365
transform 1 0 12992 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_115
timestamp 1698431365
transform 1 0 14224 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_143
timestamp 1698431365
transform 1 0 17360 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_179
timestamp 1698431365
transform 1 0 21392 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_217
timestamp 1698431365
transform 1 0 25648 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_224
timestamp 1698431365
transform 1 0 26432 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_228
timestamp 1698431365
transform 1 0 26880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_230
timestamp 1698431365
transform 1 0 27104 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_238
timestamp 1698431365
transform 1 0 28000 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_244
timestamp 1698431365
transform 1 0 28672 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_284
timestamp 1698431365
transform 1 0 33152 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_286
timestamp 1698431365
transform 1 0 33376 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_303
timestamp 1698431365
transform 1 0 35280 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_18
timestamp 1698431365
transform 1 0 3360 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_26
timestamp 1698431365
transform 1 0 4256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_101
timestamp 1698431365
transform 1 0 12656 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_146
timestamp 1698431365
transform 1 0 17696 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_184
timestamp 1698431365
transform 1 0 21952 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_197
timestamp 1698431365
transform 1 0 23408 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_222
timestamp 1698431365
transform 1 0 26208 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_279
timestamp 1698431365
transform 1 0 32592 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_297
timestamp 1698431365
transform 1 0 34608 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_70
timestamp 1698431365
transform 1 0 9184 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_72
timestamp 1698431365
transform 1 0 9408 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_100
timestamp 1698431365
transform 1 0 12544 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_104
timestamp 1698431365
transform 1 0 12992 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_115
timestamp 1698431365
transform 1 0 14224 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_119
timestamp 1698431365
transform 1 0 14672 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_121
timestamp 1698431365
transform 1 0 14896 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_128
timestamp 1698431365
transform 1 0 15680 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_130
timestamp 1698431365
transform 1 0 15904 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_137
timestamp 1698431365
transform 1 0 16688 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_153
timestamp 1698431365
transform 1 0 18480 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_157
timestamp 1698431365
transform 1 0 18928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_159
timestamp 1698431365
transform 1 0 19152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698431365
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_179
timestamp 1698431365
transform 1 0 21392 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698431365
transform 1 0 28672 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_274
timestamp 1698431365
transform 1 0 32032 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_34
timestamp 1698431365
transform 1 0 5152 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_42
timestamp 1698431365
transform 1 0 6048 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_46
timestamp 1698431365
transform 1 0 6496 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_56
timestamp 1698431365
transform 1 0 7616 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_109
timestamp 1698431365
transform 1 0 13552 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_113
timestamp 1698431365
transform 1 0 14000 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_129
timestamp 1698431365
transform 1 0 15792 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_133
timestamp 1698431365
transform 1 0 16240 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_137
timestamp 1698431365
transform 1 0 16688 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_139
timestamp 1698431365
transform 1 0 16912 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_150
timestamp 1698431365
transform 1 0 18144 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_156
timestamp 1698431365
transform 1 0 18816 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_175
timestamp 1698431365
transform 1 0 20944 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_177
timestamp 1698431365
transform 1 0 21168 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_220
timestamp 1698431365
transform 1 0 25984 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_303
timestamp 1698431365
transform 1 0 35280 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_53
timestamp 1698431365
transform 1 0 7280 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_61
timestamp 1698431365
transform 1 0 8176 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_64
timestamp 1698431365
transform 1 0 8512 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_68
timestamp 1698431365
transform 1 0 8960 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_72
timestamp 1698431365
transform 1 0 9408 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_76
timestamp 1698431365
transform 1 0 9856 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_91
timestamp 1698431365
transform 1 0 11536 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_95
timestamp 1698431365
transform 1 0 11984 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_103
timestamp 1698431365
transform 1 0 12880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_167
timestamp 1698431365
transform 1 0 20048 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_239
timestamp 1698431365
transform 1 0 28112 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698431365
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_104
timestamp 1698431365
transform 1 0 12992 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_125
timestamp 1698431365
transform 1 0 15344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_129
timestamp 1698431365
transform 1 0 15792 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_137
timestamp 1698431365
transform 1 0 16688 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698431365
transform 1 0 16912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_172
timestamp 1698431365
transform 1 0 20608 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_176
timestamp 1698431365
transform 1 0 21056 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_179
timestamp 1698431365
transform 1 0 21392 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_246
timestamp 1698431365
transform 1 0 28896 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_303
timestamp 1698431365
transform 1 0 35280 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_69
timestamp 1698431365
transform 1 0 9072 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_72
timestamp 1698431365
transform 1 0 9408 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_114
timestamp 1698431365
transform 1 0 14112 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_118
timestamp 1698431365
transform 1 0 14560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_120
timestamp 1698431365
transform 1 0 14784 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_127
timestamp 1698431365
transform 1 0 15568 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_129
timestamp 1698431365
transform 1 0 15792 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_160
timestamp 1698431365
transform 1 0 19264 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_164
timestamp 1698431365
transform 1 0 19712 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_186
timestamp 1698431365
transform 1 0 22176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_190
timestamp 1698431365
transform 1 0 22624 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_219
timestamp 1698431365
transform 1 0 25872 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_221
timestamp 1698431365
transform 1 0 26096 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_34
timestamp 1698431365
transform 1 0 5152 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_50
timestamp 1698431365
transform 1 0 6944 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_58
timestamp 1698431365
transform 1 0 7840 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_82
timestamp 1698431365
transform 1 0 10528 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_86
timestamp 1698431365
transform 1 0 10976 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_90
timestamp 1698431365
transform 1 0 11424 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_92
timestamp 1698431365
transform 1 0 11648 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_122
timestamp 1698431365
transform 1 0 15008 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_126
timestamp 1698431365
transform 1 0 15456 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_134
timestamp 1698431365
transform 1 0 16352 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_152
timestamp 1698431365
transform 1 0 18368 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_192
timestamp 1698431365
transform 1 0 22848 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_258
timestamp 1698431365
transform 1 0 30240 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_45
timestamp 1698431365
transform 1 0 6384 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_49
timestamp 1698431365
transform 1 0 6832 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_51
timestamp 1698431365
transform 1 0 7056 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_81
timestamp 1698431365
transform 1 0 10416 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_85
timestamp 1698431365
transform 1 0 10864 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_93
timestamp 1698431365
transform 1 0 11760 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_120
timestamp 1698431365
transform 1 0 14784 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_128
timestamp 1698431365
transform 1 0 15680 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_134
timestamp 1698431365
transform 1 0 16352 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_138
timestamp 1698431365
transform 1 0 16800 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_142
timestamp 1698431365
transform 1 0 17248 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_194
timestamp 1698431365
transform 1 0 23072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_210
timestamp 1698431365
transform 1 0 24864 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_274
timestamp 1698431365
transform 1 0 32032 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_34
timestamp 1698431365
transform 1 0 5152 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_50
timestamp 1698431365
transform 1 0 6944 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_52
timestamp 1698431365
transform 1 0 7168 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_63
timestamp 1698431365
transform 1 0 8400 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_80
timestamp 1698431365
transform 1 0 10304 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_84
timestamp 1698431365
transform 1 0 10752 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_92
timestamp 1698431365
transform 1 0 11648 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_107
timestamp 1698431365
transform 1 0 13328 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_150
timestamp 1698431365
transform 1 0 18144 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_154
timestamp 1698431365
transform 1 0 18592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_207
timestamp 1698431365
transform 1 0 24528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698431365
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_242
timestamp 1698431365
transform 1 0 28448 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_263
timestamp 1698431365
transform 1 0 30800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_301
timestamp 1698431365
transform 1 0 35056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_303
timestamp 1698431365
transform 1 0 35280 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_118
timestamp 1698431365
transform 1 0 14560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_120
timestamp 1698431365
transform 1 0 14784 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_163
timestamp 1698431365
transform 1 0 19600 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_181
timestamp 1698431365
transform 1 0 21616 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_183
timestamp 1698431365
transform 1 0 21840 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_197
timestamp 1698431365
transform 1 0 23408 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_201
timestamp 1698431365
transform 1 0 23856 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_205
timestamp 1698431365
transform 1 0 24304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_207
timestamp 1698431365
transform 1 0 24528 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_249
timestamp 1698431365
transform 1 0 29232 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_302
timestamp 1698431365
transform 1 0 35168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_18
timestamp 1698431365
transform 1 0 3360 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_26
timestamp 1698431365
transform 1 0 4256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_30
timestamp 1698431365
transform 1 0 4704 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1698431365
transform 1 0 8960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_77
timestamp 1698431365
transform 1 0 9968 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_81
timestamp 1698431365
transform 1 0 10416 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_83
timestamp 1698431365
transform 1 0 10640 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_110
timestamp 1698431365
transform 1 0 13664 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_118
timestamp 1698431365
transform 1 0 14560 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_126
timestamp 1698431365
transform 1 0 15456 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_133
timestamp 1698431365
transform 1 0 16240 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_153
timestamp 1698431365
transform 1 0 18480 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_161
timestamp 1698431365
transform 1 0 19376 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_169
timestamp 1698431365
transform 1 0 20272 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698431365
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_267
timestamp 1698431365
transform 1 0 31248 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_66
timestamp 1698431365
transform 1 0 8736 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_68
timestamp 1698431365
transform 1 0 8960 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_104
timestamp 1698431365
transform 1 0 12992 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_113
timestamp 1698431365
transform 1 0 14000 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_123
timestamp 1698431365
transform 1 0 15120 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_127
timestamp 1698431365
transform 1 0 15568 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_142
timestamp 1698431365
transform 1 0 17248 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_159
timestamp 1698431365
transform 1 0 19152 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_179
timestamp 1698431365
transform 1 0 21392 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_225
timestamp 1698431365
transform 1 0 26544 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_255
timestamp 1698431365
transform 1 0 29904 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_302
timestamp 1698431365
transform 1 0 35168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_18
timestamp 1698431365
transform 1 0 3360 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_48
timestamp 1698431365
transform 1 0 6720 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_50
timestamp 1698431365
transform 1 0 6944 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_61
timestamp 1698431365
transform 1 0 8176 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_65
timestamp 1698431365
transform 1 0 8624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_69
timestamp 1698431365
transform 1 0 9072 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_76
timestamp 1698431365
transform 1 0 9856 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_83
timestamp 1698431365
transform 1 0 10640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_87
timestamp 1698431365
transform 1 0 11088 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_91
timestamp 1698431365
transform 1 0 11536 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_97
timestamp 1698431365
transform 1 0 12208 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_181
timestamp 1698431365
transform 1 0 21616 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_185
timestamp 1698431365
transform 1 0 22064 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_187
timestamp 1698431365
transform 1 0 22288 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_190
timestamp 1698431365
transform 1 0 22624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_194
timestamp 1698431365
transform 1 0 23072 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_198
timestamp 1698431365
transform 1 0 23520 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_202
timestamp 1698431365
transform 1 0 23968 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_206
timestamp 1698431365
transform 1 0 24416 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_220
timestamp 1698431365
transform 1 0 25984 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_82
timestamp 1698431365
transform 1 0 10528 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_84
timestamp 1698431365
transform 1 0 10752 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_104
timestamp 1698431365
transform 1 0 12992 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_123
timestamp 1698431365
transform 1 0 15120 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_127
timestamp 1698431365
transform 1 0 15568 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_164
timestamp 1698431365
transform 1 0 19712 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_171
timestamp 1698431365
transform 1 0 20496 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_185
timestamp 1698431365
transform 1 0 22064 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_189
timestamp 1698431365
transform 1 0 22512 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_220
timestamp 1698431365
transform 1 0 25984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_277
timestamp 1698431365
transform 1 0 32368 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_18
timestamp 1698431365
transform 1 0 3360 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_64
timestamp 1698431365
transform 1 0 8512 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_109
timestamp 1698431365
transform 1 0 13552 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_113
timestamp 1698431365
transform 1 0 14000 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_117
timestamp 1698431365
transform 1 0 14448 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_133
timestamp 1698431365
transform 1 0 16240 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_137
timestamp 1698431365
transform 1 0 16688 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698431365
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_155
timestamp 1698431365
transform 1 0 18704 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_193
timestamp 1698431365
transform 1 0 22960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_197
timestamp 1698431365
transform 1 0 23408 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_201
timestamp 1698431365
transform 1 0 23856 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_218
timestamp 1698431365
transform 1 0 25760 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_234
timestamp 1698431365
transform 1 0 27552 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_236
timestamp 1698431365
transform 1 0 27776 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_45
timestamp 1698431365
transform 1 0 6384 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_47
timestamp 1698431365
transform 1 0 6608 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_162
timestamp 1698431365
transform 1 0 19488 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_166
timestamp 1698431365
transform 1 0 19936 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698431365
transform 1 0 20832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_184
timestamp 1698431365
transform 1 0 21952 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_186
timestamp 1698431365
transform 1 0 22176 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_189
timestamp 1698431365
transform 1 0 22512 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_197
timestamp 1698431365
transform 1 0 23408 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_247
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_34
timestamp 1698431365
transform 1 0 5152 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_42
timestamp 1698431365
transform 1 0 6048 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_66
timestamp 1698431365
transform 1 0 8736 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_78
timestamp 1698431365
transform 1 0 10080 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_84
timestamp 1698431365
transform 1 0 10752 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_86
timestamp 1698431365
transform 1 0 10976 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_94
timestamp 1698431365
transform 1 0 11872 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_115
timestamp 1698431365
transform 1 0 14224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_129
timestamp 1698431365
transform 1 0 15792 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698431365
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_148
timestamp 1698431365
transform 1 0 17920 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_152
timestamp 1698431365
transform 1 0 18368 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_160
timestamp 1698431365
transform 1 0 19264 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_170
timestamp 1698431365
transform 1 0 20384 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_174
timestamp 1698431365
transform 1 0 20832 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_197
timestamp 1698431365
transform 1 0 23408 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_199
timestamp 1698431365
transform 1 0 23632 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_202
timestamp 1698431365
transform 1 0 23968 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_206
timestamp 1698431365
transform 1 0 24416 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_241
timestamp 1698431365
transform 1 0 28336 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_303
timestamp 1698431365
transform 1 0 35280 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_41
timestamp 1698431365
transform 1 0 5936 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_48
timestamp 1698431365
transform 1 0 6720 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_52
timestamp 1698431365
transform 1 0 7168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_56
timestamp 1698431365
transform 1 0 7616 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_62
timestamp 1698431365
transform 1 0 8288 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_70
timestamp 1698431365
transform 1 0 9184 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_74
timestamp 1698431365
transform 1 0 9632 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_85
timestamp 1698431365
transform 1 0 10864 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_93
timestamp 1698431365
transform 1 0 11760 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_112
timestamp 1698431365
transform 1 0 13888 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_125
timestamp 1698431365
transform 1 0 15344 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_133
timestamp 1698431365
transform 1 0 16240 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_137
timestamp 1698431365
transform 1 0 16688 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_141
timestamp 1698431365
transform 1 0 17136 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_168
timestamp 1698431365
transform 1 0 20160 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_190
timestamp 1698431365
transform 1 0 22624 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_227
timestamp 1698431365
transform 1 0 26768 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_291
timestamp 1698431365
transform 1 0 33936 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_303
timestamp 1698431365
transform 1 0 35280 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_18
timestamp 1698431365
transform 1 0 3360 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_48
timestamp 1698431365
transform 1 0 6720 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698431365
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_82
timestamp 1698431365
transform 1 0 10528 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_86
timestamp 1698431365
transform 1 0 10976 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_114
timestamp 1698431365
transform 1 0 14112 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_160
timestamp 1698431365
transform 1 0 19264 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_162
timestamp 1698431365
transform 1 0 19488 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_179
timestamp 1698431365
transform 1 0 21392 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_203
timestamp 1698431365
transform 1 0 24080 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_207
timestamp 1698431365
transform 1 0 24528 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_271
timestamp 1698431365
transform 1 0 31696 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_278
timestamp 1698431365
transform 1 0 32480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_303
timestamp 1698431365
transform 1 0 35280 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_60
timestamp 1698431365
transform 1 0 8064 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_82
timestamp 1698431365
transform 1 0 10528 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_91
timestamp 1698431365
transform 1 0 11536 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_121
timestamp 1698431365
transform 1 0 14896 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_128
timestamp 1698431365
transform 1 0 15680 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_134
timestamp 1698431365
transform 1 0 16352 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_136
timestamp 1698431365
transform 1 0 16576 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_159
timestamp 1698431365
transform 1 0 19152 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_161
timestamp 1698431365
transform 1 0 19376 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_192
timestamp 1698431365
transform 1 0 22848 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_227
timestamp 1698431365
transform 1 0 26768 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698431365
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_273
timestamp 1698431365
transform 1 0 31920 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_47
timestamp 1698431365
transform 1 0 6608 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_62
timestamp 1698431365
transform 1 0 8288 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698431365
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_88
timestamp 1698431365
transform 1 0 11200 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_92
timestamp 1698431365
transform 1 0 11648 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_113
timestamp 1698431365
transform 1 0 14000 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_127
timestamp 1698431365
transform 1 0 15568 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_138
timestamp 1698431365
transform 1 0 16800 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_159
timestamp 1698431365
transform 1 0 19152 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_227
timestamp 1698431365
transform 1 0 26768 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_279
timestamp 1698431365
transform 1 0 32592 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_288
timestamp 1698431365
transform 1 0 33600 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_303
timestamp 1698431365
transform 1 0 35280 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_45
timestamp 1698431365
transform 1 0 6384 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_54
timestamp 1698431365
transform 1 0 7392 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_58
timestamp 1698431365
transform 1 0 7840 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_60
timestamp 1698431365
transform 1 0 8064 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_89
timestamp 1698431365
transform 1 0 11312 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_93
timestamp 1698431365
transform 1 0 11760 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_97
timestamp 1698431365
transform 1 0 12208 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_117
timestamp 1698431365
transform 1 0 14448 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_132
timestamp 1698431365
transform 1 0 16128 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_152
timestamp 1698431365
transform 1 0 18368 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_154
timestamp 1698431365
transform 1 0 18592 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_173
timestamp 1698431365
transform 1 0 20720 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_187
timestamp 1698431365
transform 1 0 22288 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_189
timestamp 1698431365
transform 1 0 22512 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_244
timestamp 1698431365
transform 1 0 28672 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_303
timestamp 1698431365
transform 1 0 35280 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_18
timestamp 1698431365
transform 1 0 3360 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_20
timestamp 1698431365
transform 1 0 3584 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_69
timestamp 1698431365
transform 1 0 9072 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_82
timestamp 1698431365
transform 1 0 10528 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_102
timestamp 1698431365
transform 1 0 12768 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_129
timestamp 1698431365
transform 1 0 15792 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_193
timestamp 1698431365
transform 1 0 22960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_197
timestamp 1698431365
transform 1 0 23408 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_201
timestamp 1698431365
transform 1 0 23856 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_205
timestamp 1698431365
transform 1 0 24304 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_209
timestamp 1698431365
transform 1 0 24752 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_238
timestamp 1698431365
transform 1 0 28000 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_242
timestamp 1698431365
transform 1 0 28448 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_244
timestamp 1698431365
transform 1 0 28672 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_276
timestamp 1698431365
transform 1 0 32256 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_41
timestamp 1698431365
transform 1 0 5936 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_43
timestamp 1698431365
transform 1 0 6160 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_55
timestamp 1698431365
transform 1 0 7504 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_63
timestamp 1698431365
transform 1 0 8400 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_111
timestamp 1698431365
transform 1 0 13776 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_187
timestamp 1698431365
transform 1 0 22288 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_191
timestamp 1698431365
transform 1 0 22736 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_201
timestamp 1698431365
transform 1 0 23856 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_233
timestamp 1698431365
transform 1 0 27440 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_237
timestamp 1698431365
transform 1 0 27888 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_241
timestamp 1698431365
transform 1 0 28336 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_280
timestamp 1698431365
transform 1 0 32704 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_282
timestamp 1698431365
transform 1 0 32928 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_285
timestamp 1698431365
transform 1 0 33264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_289
timestamp 1698431365
transform 1 0 33712 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_293
timestamp 1698431365
transform 1 0 34160 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_295
timestamp 1698431365
transform 1 0 34384 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_18
timestamp 1698431365
transform 1 0 3360 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_61
timestamp 1698431365
transform 1 0 8176 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_65
timestamp 1698431365
transform 1 0 8624 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_69
timestamp 1698431365
transform 1 0 9072 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_76
timestamp 1698431365
transform 1 0 9856 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_208
timestamp 1698431365
transform 1 0 24640 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_217
timestamp 1698431365
transform 1 0 25648 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_221
timestamp 1698431365
transform 1 0 26096 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_229
timestamp 1698431365
transform 1 0 26992 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_300
timestamp 1698431365
transform 1 0 34944 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_57
timestamp 1698431365
transform 1 0 7728 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_92
timestamp 1698431365
transform 1 0 11648 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_96
timestamp 1698431365
transform 1 0 12096 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_104
timestamp 1698431365
transform 1 0 12992 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_113
timestamp 1698431365
transform 1 0 14000 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_172
timestamp 1698431365
transform 1 0 20608 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_174
timestamp 1698431365
transform 1 0 20832 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_230
timestamp 1698431365
transform 1 0 27104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_234
timestamp 1698431365
transform 1 0 27552 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_302
timestamp 1698431365
transform 1 0 35168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_34
timestamp 1698431365
transform 1 0 5152 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_38
timestamp 1698431365
transform 1 0 5600 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_40
timestamp 1698431365
transform 1 0 5824 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_76
timestamp 1698431365
transform 1 0 9856 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_80
timestamp 1698431365
transform 1 0 10304 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_96
timestamp 1698431365
transform 1 0 12096 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_201
timestamp 1698431365
transform 1 0 23856 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_205
timestamp 1698431365
transform 1 0 24304 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_209
timestamp 1698431365
transform 1 0 24752 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_238
timestamp 1698431365
transform 1 0 28000 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_274
timestamp 1698431365
transform 1 0 32032 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_278
timestamp 1698431365
transform 1 0 32480 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_286
timestamp 1698431365
transform 1 0 33376 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_290
timestamp 1698431365
transform 1 0 33824 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_294
timestamp 1698431365
transform 1 0 34272 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_7
timestamp 1698431365
transform 1 0 2128 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_11
timestamp 1698431365
transform 1 0 2576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_17
timestamp 1698431365
transform 1 0 3248 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_21
timestamp 1698431365
transform 1 0 3696 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_27
timestamp 1698431365
transform 1 0 4368 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_29
timestamp 1698431365
transform 1 0 4592 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_36
timestamp 1698431365
transform 1 0 5376 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_70
timestamp 1698431365
transform 1 0 9184 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_133
timestamp 1698431365
transform 1 0 16240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_135
timestamp 1698431365
transform 1 0 16464 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_167
timestamp 1698431365
transform 1 0 20048 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_169
timestamp 1698431365
transform 1 0 20272 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_172
timestamp 1698431365
transform 1 0 20608 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_232
timestamp 1698431365
transform 1 0 27328 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_236
timestamp 1698431365
transform 1 0 27776 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_240
timestamp 1698431365
transform 1 0 28224 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_303
timestamp 1698431365
transform 1 0 35280 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform 1 0 34720 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform -1 0 35392 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform -1 0 35392 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform -1 0 34384 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform 1 0 33712 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform -1 0 35392 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform -1 0 35392 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input8
timestamp 1698431365
transform -1 0 35392 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input9
timestamp 1698431365
transform 1 0 26880 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input10
timestamp 1698431365
transform -1 0 35280 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform -1 0 35392 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform 1 0 23520 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform -1 0 28000 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform -1 0 28896 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform -1 0 29568 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform -1 0 30800 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698431365
transform -1 0 32704 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698431365
transform -1 0 33936 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform -1 0 35392 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12880 0 -1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698431365
transform 1 0 9856 0 1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698431365
transform 1 0 14448 0 1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698431365
transform 1 0 14448 0 1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698431365
transform 1 0 17360 0 1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698431365
transform 1 0 17472 0 -1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output26
timestamp 1698431365
transform 1 0 19600 0 -1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output27
timestamp 1698431365
transform 1 0 24416 0 1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output28
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output29
timestamp 1698431365
transform 1 0 21952 0 -1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output30
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output31
timestamp 1698431365
transform 1 0 29792 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output32
timestamp 1698431365
transform 1 0 32256 0 1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output33
timestamp 1698431365
transform 1 0 32256 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output34
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output35
timestamp 1698431365
transform 1 0 28896 0 1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output36
timestamp 1698431365
transform 1 0 29232 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output37
timestamp 1698431365
transform 1 0 29792 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output38
timestamp 1698431365
transform -1 0 32704 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output39
timestamp 1698431365
transform -1 0 31696 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output40
timestamp 1698431365
transform -1 0 28784 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output41
timestamp 1698431365
transform 1 0 6048 0 1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output42
timestamp 1698431365
transform 1 0 10192 0 1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output43
timestamp 1698431365
transform -1 0 4816 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output44
timestamp 1698431365
transform -1 0 5712 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output45
timestamp 1698431365
transform -1 0 5152 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output46
timestamp 1698431365
transform -1 0 9184 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output47
timestamp 1698431365
transform -1 0 8960 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output48
timestamp 1698431365
transform -1 0 10192 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output49
timestamp 1698431365
transform 1 0 32480 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output50
timestamp 1698431365
transform -1 0 13104 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output51
timestamp 1698431365
transform 1 0 9856 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output52
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output53
timestamp 1698431365
transform 1 0 13664 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output54
timestamp 1698431365
transform 1 0 17472 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output55
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output56
timestamp 1698431365
transform 1 0 20720 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output57
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_39 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_40
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 35616 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_41
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 35616 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_42
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 35616 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_43
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 35616 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_44
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 35616 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_45
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 35616 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_46
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 35616 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_47
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 35616 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_48
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 35616 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_49
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 35616 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_50
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 35616 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_51
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 35616 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_52
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 35616 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_53
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 35616 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_54
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 35616 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_55
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 35616 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_56
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 35616 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_57
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 35616 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_58
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 35616 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_59
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 35616 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_60
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 35616 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_61
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 35616 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_62
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 35616 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_63
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 35616 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_64
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 35616 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_65
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 35616 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_66
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 35616 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_67
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 35616 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_68
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 35616 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_69
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 35616 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_70
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 35616 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_71
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 35616 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_72
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 35616 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_73
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 35616 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_74
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 35616 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_75
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 35616 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_76
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 35616 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_77
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 35616 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer1
timestamp 1698431365
transform -1 0 23632 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  rebuffer2
timestamp 1698431365
transform -1 0 27104 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_78 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_79
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_80
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_81
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_82
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_83
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_84
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_85
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_86
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_87
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_88
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_89
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_90
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_91
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_92
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_93
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_94
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_95
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_96
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_97
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_98
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_99
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_100
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_101
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_102
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_103
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_104
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_105
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_106
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_107
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_108
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_109
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_110
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_111
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_112
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_113
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_114
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_115
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_116
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_117
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_118
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_119
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_120
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_121
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_122
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_123
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_124
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_125
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_126
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_127
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_128
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_129
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_130
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_131
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_132
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_133
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_134
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_135
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_136
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_137
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_138
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_139
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_140
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_141
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_142
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_143
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_144
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_145
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_146
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_147
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_148
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_149
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_150
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_151
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_152
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_153
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_154
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_155
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_156
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_157
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_158
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_159
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_160
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_161
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_162
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_163
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_164
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_165
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_166
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_167
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_168
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_169
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_170
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_171
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_172
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_173
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_174
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_175
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_176
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_177
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_178
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_179
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_180
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_181
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_182
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_183
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_184
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_185
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_186
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_187
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_188
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_189
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_190
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_191
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_192
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_193
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_194
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_195
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_196
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_197
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_198
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_199
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_200
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_201
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_202
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_203
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_204
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_205
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_206
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_207
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_208
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_209
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_210
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_211
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_212
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_213
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_214
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_215
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_216
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_217
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_218
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_219
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_220
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_221
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_222
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_223
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_224
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_225
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_226
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_227
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_228
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_229
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_230
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_231
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_232
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_233
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_234
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_235
timestamp 1698431365
transform 1 0 8960 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_236
timestamp 1698431365
transform 1 0 12768 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_237
timestamp 1698431365
transform 1 0 16576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_238
timestamp 1698431365
transform 1 0 20384 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_239
timestamp 1698431365
transform 1 0 24192 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_240
timestamp 1698431365
transform 1 0 28000 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_241
timestamp 1698431365
transform 1 0 31808 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_mc14500_67 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 2128 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_mc14500_68
timestamp 1698431365
transform -1 0 3248 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_mc14500_69
timestamp 1698431365
transform -1 0 4368 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_mc14500_70
timestamp 1698431365
transform 1 0 4704 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_mc14500_71
timestamp 1698431365
transform 1 0 5600 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_mc14500_72
timestamp 1698431365
transform -1 0 7728 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_mc14500_73
timestamp 1698431365
transform -1 0 9856 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_mc14500_74
timestamp 1698431365
transform -1 0 9856 0 1 32928
box -86 -86 534 870
<< labels >>
flabel metal3 s 36200 29120 37000 29232 0 FreeSans 448 0 0 0 SDI
port 0 nsew signal input
flabel metal3 s 36200 2240 37000 2352 0 FreeSans 448 0 0 0 clk_i
port 1 nsew signal input
flabel metal3 s 36200 34496 37000 34608 0 FreeSans 448 0 0 0 custom_setting
port 2 nsew signal input
flabel metal3 s 36200 7616 37000 7728 0 FreeSans 448 0 0 0 io_in[0]
port 3 nsew signal input
flabel metal3 s 36200 10304 37000 10416 0 FreeSans 448 0 0 0 io_in[1]
port 4 nsew signal input
flabel metal3 s 36200 12992 37000 13104 0 FreeSans 448 0 0 0 io_in[2]
port 5 nsew signal input
flabel metal3 s 36200 15680 37000 15792 0 FreeSans 448 0 0 0 io_in[3]
port 6 nsew signal input
flabel metal3 s 36200 18368 37000 18480 0 FreeSans 448 0 0 0 io_in[4]
port 7 nsew signal input
flabel metal3 s 36200 21056 37000 21168 0 FreeSans 448 0 0 0 io_in[5]
port 8 nsew signal input
flabel metal3 s 36200 23744 37000 23856 0 FreeSans 448 0 0 0 io_in[6]
port 9 nsew signal input
flabel metal3 s 36200 26432 37000 26544 0 FreeSans 448 0 0 0 io_in[7]
port 10 nsew signal input
flabel metal2 s 1568 36200 1680 37000 0 FreeSans 448 90 0 0 io_out[0]
port 11 nsew signal tristate
flabel metal2 s 12768 36200 12880 37000 0 FreeSans 448 90 0 0 io_out[10]
port 12 nsew signal tristate
flabel metal2 s 13888 36200 14000 37000 0 FreeSans 448 90 0 0 io_out[11]
port 13 nsew signal tristate
flabel metal2 s 15008 36200 15120 37000 0 FreeSans 448 90 0 0 io_out[12]
port 14 nsew signal tristate
flabel metal2 s 16128 36200 16240 37000 0 FreeSans 448 90 0 0 io_out[13]
port 15 nsew signal tristate
flabel metal2 s 17248 36200 17360 37000 0 FreeSans 448 90 0 0 io_out[14]
port 16 nsew signal tristate
flabel metal2 s 18368 36200 18480 37000 0 FreeSans 448 90 0 0 io_out[15]
port 17 nsew signal tristate
flabel metal2 s 19488 36200 19600 37000 0 FreeSans 448 90 0 0 io_out[16]
port 18 nsew signal tristate
flabel metal2 s 20608 36200 20720 37000 0 FreeSans 448 90 0 0 io_out[17]
port 19 nsew signal tristate
flabel metal2 s 21728 36200 21840 37000 0 FreeSans 448 90 0 0 io_out[18]
port 20 nsew signal tristate
flabel metal2 s 22848 36200 22960 37000 0 FreeSans 448 90 0 0 io_out[19]
port 21 nsew signal tristate
flabel metal2 s 2688 36200 2800 37000 0 FreeSans 448 90 0 0 io_out[1]
port 22 nsew signal tristate
flabel metal2 s 23968 36200 24080 37000 0 FreeSans 448 90 0 0 io_out[20]
port 23 nsew signal tristate
flabel metal2 s 25088 36200 25200 37000 0 FreeSans 448 90 0 0 io_out[21]
port 24 nsew signal tristate
flabel metal2 s 26208 36200 26320 37000 0 FreeSans 448 90 0 0 io_out[22]
port 25 nsew signal tristate
flabel metal2 s 27328 36200 27440 37000 0 FreeSans 448 90 0 0 io_out[23]
port 26 nsew signal tristate
flabel metal2 s 28448 36200 28560 37000 0 FreeSans 448 90 0 0 io_out[24]
port 27 nsew signal tristate
flabel metal2 s 29568 36200 29680 37000 0 FreeSans 448 90 0 0 io_out[25]
port 28 nsew signal tristate
flabel metal2 s 30688 36200 30800 37000 0 FreeSans 448 90 0 0 io_out[26]
port 29 nsew signal tristate
flabel metal2 s 31808 36200 31920 37000 0 FreeSans 448 90 0 0 io_out[27]
port 30 nsew signal tristate
flabel metal2 s 32928 36200 33040 37000 0 FreeSans 448 90 0 0 io_out[28]
port 31 nsew signal tristate
flabel metal2 s 34048 36200 34160 37000 0 FreeSans 448 90 0 0 io_out[29]
port 32 nsew signal tristate
flabel metal2 s 3808 36200 3920 37000 0 FreeSans 448 90 0 0 io_out[2]
port 33 nsew signal tristate
flabel metal2 s 35168 36200 35280 37000 0 FreeSans 448 90 0 0 io_out[30]
port 34 nsew signal tristate
flabel metal2 s 4928 36200 5040 37000 0 FreeSans 448 90 0 0 io_out[3]
port 35 nsew signal tristate
flabel metal2 s 6048 36200 6160 37000 0 FreeSans 448 90 0 0 io_out[4]
port 36 nsew signal tristate
flabel metal2 s 7168 36200 7280 37000 0 FreeSans 448 90 0 0 io_out[5]
port 37 nsew signal tristate
flabel metal2 s 8288 36200 8400 37000 0 FreeSans 448 90 0 0 io_out[6]
port 38 nsew signal tristate
flabel metal2 s 9408 36200 9520 37000 0 FreeSans 448 90 0 0 io_out[7]
port 39 nsew signal tristate
flabel metal2 s 10528 36200 10640 37000 0 FreeSans 448 90 0 0 io_out[8]
port 40 nsew signal tristate
flabel metal2 s 11648 36200 11760 37000 0 FreeSans 448 90 0 0 io_out[9]
port 41 nsew signal tristate
flabel metal3 s 36200 4928 37000 5040 0 FreeSans 448 0 0 0 rst_n
port 42 nsew signal input
flabel metal2 s 1792 0 1904 800 0 FreeSans 448 90 0 0 sram_addr[0]
port 43 nsew signal tristate
flabel metal2 s 3360 0 3472 800 0 FreeSans 448 90 0 0 sram_addr[1]
port 44 nsew signal tristate
flabel metal2 s 4928 0 5040 800 0 FreeSans 448 90 0 0 sram_addr[2]
port 45 nsew signal tristate
flabel metal2 s 6496 0 6608 800 0 FreeSans 448 90 0 0 sram_addr[3]
port 46 nsew signal tristate
flabel metal2 s 8064 0 8176 800 0 FreeSans 448 90 0 0 sram_addr[4]
port 47 nsew signal tristate
flabel metal2 s 9632 0 9744 800 0 FreeSans 448 90 0 0 sram_addr[5]
port 48 nsew signal tristate
flabel metal3 s 36200 31808 37000 31920 0 FreeSans 448 0 0 0 sram_gwe
port 49 nsew signal tristate
flabel metal2 s 11200 0 11312 800 0 FreeSans 448 90 0 0 sram_in[0]
port 50 nsew signal tristate
flabel metal2 s 12768 0 12880 800 0 FreeSans 448 90 0 0 sram_in[1]
port 51 nsew signal tristate
flabel metal2 s 14336 0 14448 800 0 FreeSans 448 90 0 0 sram_in[2]
port 52 nsew signal tristate
flabel metal2 s 15904 0 16016 800 0 FreeSans 448 90 0 0 sram_in[3]
port 53 nsew signal tristate
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 sram_in[4]
port 54 nsew signal tristate
flabel metal2 s 19040 0 19152 800 0 FreeSans 448 90 0 0 sram_in[5]
port 55 nsew signal tristate
flabel metal2 s 20608 0 20720 800 0 FreeSans 448 90 0 0 sram_in[6]
port 56 nsew signal tristate
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 sram_in[7]
port 57 nsew signal tristate
flabel metal2 s 23744 0 23856 800 0 FreeSans 448 90 0 0 sram_out[0]
port 58 nsew signal input
flabel metal2 s 25312 0 25424 800 0 FreeSans 448 90 0 0 sram_out[1]
port 59 nsew signal input
flabel metal2 s 26880 0 26992 800 0 FreeSans 448 90 0 0 sram_out[2]
port 60 nsew signal input
flabel metal2 s 28448 0 28560 800 0 FreeSans 448 90 0 0 sram_out[3]
port 61 nsew signal input
flabel metal2 s 30016 0 30128 800 0 FreeSans 448 90 0 0 sram_out[4]
port 62 nsew signal input
flabel metal2 s 31584 0 31696 800 0 FreeSans 448 90 0 0 sram_out[5]
port 63 nsew signal input
flabel metal2 s 33152 0 33264 800 0 FreeSans 448 90 0 0 sram_out[6]
port 64 nsew signal input
flabel metal2 s 34720 0 34832 800 0 FreeSans 448 90 0 0 sram_out[7]
port 65 nsew signal input
flabel metal4 s 5468 3076 5788 33772 0 FreeSans 1280 90 0 0 vdd
port 66 nsew power bidirectional
flabel metal4 s 14036 3076 14356 33772 0 FreeSans 1280 90 0 0 vdd
port 66 nsew power bidirectional
flabel metal4 s 22604 3076 22924 33772 0 FreeSans 1280 90 0 0 vdd
port 66 nsew power bidirectional
flabel metal4 s 31172 3076 31492 33772 0 FreeSans 1280 90 0 0 vdd
port 66 nsew power bidirectional
flabel metal4 s 9752 3076 10072 33772 0 FreeSans 1280 90 0 0 vss
port 67 nsew ground bidirectional
flabel metal4 s 18320 3076 18640 33772 0 FreeSans 1280 90 0 0 vss
port 67 nsew ground bidirectional
flabel metal4 s 26888 3076 27208 33772 0 FreeSans 1280 90 0 0 vss
port 67 nsew ground bidirectional
flabel metal4 s 35456 3076 35776 33772 0 FreeSans 1280 90 0 0 vss
port 67 nsew ground bidirectional
rlabel metal1 18480 33712 18480 33712 0 vdd
rlabel via1 18560 32928 18560 32928 0 vss
rlabel metal2 34888 29904 34888 29904 0 SDI
rlabel metal2 31192 15960 31192 15960 0 _0000_
rlabel metal3 21728 14616 21728 14616 0 _0001_
rlabel metal2 17976 16016 17976 16016 0 _0002_
rlabel metal3 24528 21784 24528 21784 0 _0003_
rlabel metal2 25592 21168 25592 21168 0 _0004_
rlabel metal2 26040 25032 26040 25032 0 _0005_
rlabel metal3 29848 28056 29848 28056 0 _0006_
rlabel metal2 33096 26712 33096 26712 0 _0007_
rlabel metal2 33096 24472 33096 24472 0 _0008_
rlabel metal2 28280 26236 28280 26236 0 _0009_
rlabel metal2 29680 25256 29680 25256 0 _0010_
rlabel metal2 7784 11704 7784 11704 0 _0011_
rlabel metal2 6944 12264 6944 12264 0 _0012_
rlabel metal2 11816 8344 11816 8344 0 _0013_
rlabel metal3 12320 4200 12320 4200 0 _0014_
rlabel metal2 10696 5264 10696 5264 0 _0015_
rlabel metal2 13608 5488 13608 5488 0 _0016_
rlabel metal2 16072 5096 16072 5096 0 _0017_
rlabel metal3 17136 4536 17136 4536 0 _0018_
rlabel metal2 18648 5488 18648 5488 0 _0019_
rlabel metal2 20048 4424 20048 4424 0 _0020_
rlabel metal2 17192 8120 17192 8120 0 _0021_
rlabel metal2 12936 7784 12936 7784 0 _0022_
rlabel metal3 13664 9912 13664 9912 0 _0023_
rlabel metal2 14952 11760 14952 11760 0 _0024_
rlabel metal2 18760 12488 18760 12488 0 _0025_
rlabel metal2 20104 9688 20104 9688 0 _0026_
rlabel metal2 22456 11760 22456 11760 0 _0027_
rlabel metal2 24808 10080 24808 10080 0 _0028_
rlabel metal2 22120 7000 22120 7000 0 _0029_
rlabel metal3 23968 5208 23968 5208 0 _0030_
rlabel metal2 25984 4424 25984 4424 0 _0031_
rlabel metal2 30632 4648 30632 4648 0 _0032_
rlabel metal2 29848 6048 29848 6048 0 _0033_
rlabel metal2 31192 7896 31192 7896 0 _0034_
rlabel metal2 28056 9352 28056 9352 0 _0035_
rlabel metal2 30184 10584 30184 10584 0 _0036_
rlabel metal2 33544 32200 33544 32200 0 _0037_
rlabel metal2 30408 30464 30408 30464 0 _0038_
rlabel metal2 23016 25144 23016 25144 0 _0039_
rlabel metal2 29792 10696 29792 10696 0 _0040_
rlabel metal2 14952 15148 14952 15148 0 _0041_
rlabel metal2 21672 22568 21672 22568 0 _0042_
rlabel metal2 29960 31248 29960 31248 0 _0043_
rlabel metal2 28056 32144 28056 32144 0 _0044_
rlabel metal2 26264 12152 26264 12152 0 _0045_
rlabel metal2 8568 17304 8568 17304 0 _0046_
rlabel metal2 6496 19320 6496 19320 0 _0047_
rlabel metal3 7224 19880 7224 19880 0 _0048_
rlabel metal2 4424 21896 4424 21896 0 _0049_
rlabel metal3 6048 23016 6048 23016 0 _0050_
rlabel metal2 8232 22568 8232 22568 0 _0051_
rlabel metal2 11256 22568 11256 22568 0 _0052_
rlabel metal2 11592 20440 11592 20440 0 _0053_
rlabel metal2 10248 19600 10248 19600 0 _0054_
rlabel metal2 10864 16184 10864 16184 0 _0055_
rlabel metal3 13160 16968 13160 16968 0 _0056_
rlabel metal2 14728 18704 14728 18704 0 _0057_
rlabel metal2 17528 18872 17528 18872 0 _0058_
rlabel metal2 16632 21168 16632 21168 0 _0059_
rlabel metal3 19152 20552 19152 20552 0 _0060_
rlabel metal2 16856 22904 16856 22904 0 _0061_
rlabel metal3 4984 27272 4984 27272 0 _0062_
rlabel metal3 6048 28840 6048 28840 0 _0063_
rlabel metal2 4648 29736 4648 29736 0 _0064_
rlabel metal2 8120 32200 8120 32200 0 _0065_
rlabel metal2 9576 31416 9576 31416 0 _0066_
rlabel metal2 6216 25928 6216 25928 0 _0067_
rlabel metal2 12824 29792 12824 29792 0 _0068_
rlabel metal2 12712 28112 12712 28112 0 _0069_
rlabel metal2 17864 31416 17864 31416 0 _0070_
rlabel metal2 18312 32256 18312 32256 0 _0071_
rlabel metal2 13608 31696 13608 31696 0 _0072_
rlabel metal2 20832 30408 20832 30408 0 _0073_
rlabel metal2 21616 33208 21616 33208 0 _0074_
rlabel metal2 21784 30072 21784 30072 0 _0075_
rlabel metal3 23520 26936 23520 26936 0 _0076_
rlabel metal2 22120 29232 22120 29232 0 _0077_
rlabel metal2 10360 14056 10360 14056 0 _0078_
rlabel metal2 11704 12096 11704 12096 0 _0079_
rlabel metal2 8232 9464 8232 9464 0 _0080_
rlabel metal2 6888 5824 6888 5824 0 _0081_
rlabel metal2 6608 4424 6608 4424 0 _0082_
rlabel metal2 6664 8624 6664 8624 0 _0083_
rlabel metal2 24248 12712 24248 12712 0 _0084_
rlabel metal3 32536 15960 32536 15960 0 _0085_
rlabel metal2 24584 15568 24584 15568 0 _0086_
rlabel metal2 20776 14000 20776 14000 0 _0087_
rlabel metal2 22064 15960 22064 15960 0 _0088_
rlabel metal2 24696 15904 24696 15904 0 _0089_
rlabel metal2 24472 16576 24472 16576 0 _0090_
rlabel metal2 25424 16968 25424 16968 0 _0091_
rlabel metal3 24864 16072 24864 16072 0 _0092_
rlabel metal3 21448 16856 21448 16856 0 _0093_
rlabel metal3 23016 16856 23016 16856 0 _0094_
rlabel metal2 21448 17920 21448 17920 0 _0095_
rlabel metal2 26824 18144 26824 18144 0 _0096_
rlabel metal2 24024 13608 24024 13608 0 _0097_
rlabel metal2 24360 13384 24360 13384 0 _0098_
rlabel metal2 24696 12096 24696 12096 0 _0099_
rlabel metal2 26824 17248 26824 17248 0 _0100_
rlabel metal3 22848 16072 22848 16072 0 _0101_
rlabel metal2 20328 16912 20328 16912 0 _0102_
rlabel metal2 27496 18368 27496 18368 0 _0103_
rlabel metal2 27160 24080 27160 24080 0 _0104_
rlabel metal2 33096 25256 33096 25256 0 _0105_
rlabel metal2 34104 19488 34104 19488 0 _0106_
rlabel metal2 35112 21448 35112 21448 0 _0107_
rlabel metal2 35336 23520 35336 23520 0 _0108_
rlabel metal2 34496 24808 34496 24808 0 _0109_
rlabel metal2 26824 19824 26824 19824 0 _0110_
rlabel metal3 25816 19712 25816 19712 0 _0111_
rlabel metal2 31360 21560 31360 21560 0 _0112_
rlabel metal2 27608 19320 27608 19320 0 _0113_
rlabel metal2 25088 16296 25088 16296 0 _0114_
rlabel metal2 19656 18984 19656 18984 0 _0115_
rlabel metal3 20552 17528 20552 17528 0 _0116_
rlabel metal2 22176 12376 22176 12376 0 _0117_
rlabel metal2 22344 17304 22344 17304 0 _0118_
rlabel metal2 21896 17080 21896 17080 0 _0119_
rlabel metal2 24024 20664 24024 20664 0 _0120_
rlabel metal2 27832 22344 27832 22344 0 _0121_
rlabel metal3 27776 25704 27776 25704 0 _0122_
rlabel metal2 34776 25480 34776 25480 0 _0123_
rlabel metal3 34216 26376 34216 26376 0 _0124_
rlabel metal3 28280 17416 28280 17416 0 _0125_
rlabel metal2 25144 23688 25144 23688 0 _0126_
rlabel metal2 33432 21000 33432 21000 0 _0127_
rlabel metal2 25480 23800 25480 23800 0 _0128_
rlabel metal2 28616 24024 28616 24024 0 _0129_
rlabel metal3 23856 18536 23856 18536 0 _0130_
rlabel metal2 15288 15904 15288 15904 0 _0131_
rlabel metal2 34328 25088 34328 25088 0 _0132_
rlabel metal3 31136 24696 31136 24696 0 _0133_
rlabel metal3 31696 27720 31696 27720 0 _0134_
rlabel metal3 34328 24472 34328 24472 0 _0135_
rlabel metal2 28280 23744 28280 23744 0 _0136_
rlabel metal2 28504 24696 28504 24696 0 _0137_
rlabel metal3 24472 23016 24472 23016 0 _0138_
rlabel metal3 25536 23352 25536 23352 0 _0139_
rlabel metal2 26432 21336 26432 21336 0 _0140_
rlabel metal2 26544 20104 26544 20104 0 _0141_
rlabel metal2 25480 22344 25480 22344 0 _0142_
rlabel metal3 25872 22120 25872 22120 0 _0143_
rlabel metal2 25928 22624 25928 22624 0 _0144_
rlabel metal3 27048 23688 27048 23688 0 _0145_
rlabel metal2 28840 23016 28840 23016 0 _0146_
rlabel metal2 30744 23464 30744 23464 0 _0147_
rlabel metal2 28672 25368 28672 25368 0 _0148_
rlabel metal2 29736 12992 29736 12992 0 _0149_
rlabel metal2 18088 16632 18088 16632 0 _0150_
rlabel metal3 22904 13832 22904 13832 0 _0151_
rlabel metal3 18928 16408 18928 16408 0 _0152_
rlabel metal2 15176 12544 15176 12544 0 _0153_
rlabel metal2 16800 17080 16800 17080 0 _0154_
rlabel metal3 25704 15176 25704 15176 0 _0155_
rlabel metal2 23352 13440 23352 13440 0 _0156_
rlabel metal3 25424 12936 25424 12936 0 _0157_
rlabel metal2 25424 18536 25424 18536 0 _0158_
rlabel metal2 28672 20888 28672 20888 0 _0159_
rlabel metal2 31976 22792 31976 22792 0 _0160_
rlabel metal2 28392 21280 28392 21280 0 _0161_
rlabel metal3 30296 20776 30296 20776 0 _0162_
rlabel metal3 32312 19096 32312 19096 0 _0163_
rlabel metal3 25928 20664 25928 20664 0 _0164_
rlabel metal2 27384 20888 27384 20888 0 _0165_
rlabel metal2 32424 19880 32424 19880 0 _0166_
rlabel metal2 33208 21616 33208 21616 0 _0167_
rlabel metal2 33936 23016 33936 23016 0 _0168_
rlabel metal2 31752 21952 31752 21952 0 _0169_
rlabel metal2 34664 22232 34664 22232 0 _0170_
rlabel metal2 33768 21616 33768 21616 0 _0171_
rlabel metal2 33152 23800 33152 23800 0 _0172_
rlabel metal2 31864 21224 31864 21224 0 _0173_
rlabel metal2 30632 19992 30632 19992 0 _0174_
rlabel metal2 32200 18144 32200 18144 0 _0175_
rlabel metal3 32984 18424 32984 18424 0 _0176_
rlabel metal2 31976 19264 31976 19264 0 _0177_
rlabel metal3 26124 19432 26124 19432 0 _0178_
rlabel metal2 32088 13440 32088 13440 0 _0179_
rlabel metal2 35112 16800 35112 16800 0 _0180_
rlabel metal2 31752 19096 31752 19096 0 _0181_
rlabel metal2 31416 18816 31416 18816 0 _0182_
rlabel via2 26376 18088 26376 18088 0 _0183_
rlabel via3 26600 18639 26600 18639 0 _0184_
rlabel metal2 28056 18704 28056 18704 0 _0185_
rlabel metal3 29008 16408 29008 16408 0 _0186_
rlabel metal3 29232 12936 29232 12936 0 _0187_
rlabel metal2 26600 19488 26600 19488 0 _0188_
rlabel metal2 26264 19096 26264 19096 0 _0189_
rlabel metal2 26488 17528 26488 17528 0 _0190_
rlabel metal3 27384 15848 27384 15848 0 _0191_
rlabel metal2 28056 16352 28056 16352 0 _0192_
rlabel metal2 27664 15624 27664 15624 0 _0193_
rlabel metal2 25816 18088 25816 18088 0 _0194_
rlabel metal2 27608 17304 27608 17304 0 _0195_
rlabel metal2 30464 16296 30464 16296 0 _0196_
rlabel metal2 30072 14616 30072 14616 0 _0197_
rlabel metal3 20272 13608 20272 13608 0 _0198_
rlabel metal2 25704 18088 25704 18088 0 _0199_
rlabel metal2 16408 17472 16408 17472 0 _0200_
rlabel metal3 18648 17416 18648 17416 0 _0201_
rlabel metal2 16856 15456 16856 15456 0 _0202_
rlabel metal2 10024 13104 10024 13104 0 _0203_
rlabel metal2 8344 12432 8344 12432 0 _0204_
rlabel metal2 7952 12376 7952 12376 0 _0205_
rlabel metal2 10528 12712 10528 12712 0 _0206_
rlabel metal2 8568 13104 8568 13104 0 _0207_
rlabel metal2 6216 13104 6216 13104 0 _0208_
rlabel metal2 7448 12936 7448 12936 0 _0209_
rlabel metal3 22456 25984 22456 25984 0 _0210_
rlabel metal3 24696 18984 24696 18984 0 _0211_
rlabel metal3 21168 15176 21168 15176 0 _0212_
rlabel metal2 11144 8736 11144 8736 0 _0213_
rlabel metal2 16184 9912 16184 9912 0 _0214_
rlabel metal2 12096 9800 12096 9800 0 _0215_
rlabel metal2 24640 19992 24640 19992 0 _0216_
rlabel metal2 18200 16072 18200 16072 0 _0217_
rlabel metal2 17416 7728 17416 7728 0 _0218_
rlabel metal2 13048 4984 13048 4984 0 _0219_
rlabel metal2 12712 4592 12712 4592 0 _0220_
rlabel metal2 13608 21896 13608 21896 0 _0221_
rlabel metal3 14168 15512 14168 15512 0 _0222_
rlabel metal3 10304 5880 10304 5880 0 _0223_
rlabel metal3 8400 5992 8400 5992 0 _0224_
rlabel metal2 13832 6552 13832 6552 0 _0225_
rlabel metal2 6104 3528 6104 3528 0 _0226_
rlabel metal2 16184 5936 16184 5936 0 _0227_
rlabel metal2 18256 6552 18256 6552 0 _0228_
rlabel metal2 15848 6160 15848 6160 0 _0229_
rlabel metal2 19152 15848 19152 15848 0 _0230_
rlabel metal2 16520 5824 16520 5824 0 _0231_
rlabel metal2 17640 4368 17640 4368 0 _0232_
rlabel metal2 17304 4032 17304 4032 0 _0233_
rlabel metal2 17416 4312 17416 4312 0 _0234_
rlabel metal2 18704 4536 18704 4536 0 _0235_
rlabel metal2 22792 4088 22792 4088 0 _0236_
rlabel metal2 19656 6608 19656 6608 0 _0237_
rlabel metal2 19824 20104 19824 20104 0 _0238_
rlabel metal3 21168 19208 21168 19208 0 _0239_
rlabel metal2 20608 18984 20608 18984 0 _0240_
rlabel metal2 16968 9912 16968 9912 0 _0241_
rlabel metal2 25032 18200 25032 18200 0 _0242_
rlabel metal2 20216 8344 20216 8344 0 _0243_
rlabel metal2 15848 9352 15848 9352 0 _0244_
rlabel metal2 17416 9688 17416 9688 0 _0245_
rlabel metal2 15512 9408 15512 9408 0 _0246_
rlabel metal2 16632 9016 16632 9016 0 _0247_
rlabel metal2 24528 4536 24528 4536 0 _0248_
rlabel metal3 19040 7560 19040 7560 0 _0249_
rlabel metal2 20216 6720 20216 6720 0 _0250_
rlabel metal2 17528 8680 17528 8680 0 _0251_
rlabel metal2 14728 8904 14728 8904 0 _0252_
rlabel metal2 25928 7728 25928 7728 0 _0253_
rlabel metal3 17248 7448 17248 7448 0 _0254_
rlabel metal2 15736 7896 15736 7896 0 _0255_
rlabel metal2 14616 10136 14616 10136 0 _0256_
rlabel metal3 21000 7392 21000 7392 0 _0257_
rlabel metal2 20776 7896 20776 7896 0 _0258_
rlabel metal3 15960 9520 15960 9520 0 _0259_
rlabel metal3 15736 11144 15736 11144 0 _0260_
rlabel metal2 15624 11368 15624 11368 0 _0261_
rlabel metal2 23072 12152 23072 12152 0 _0262_
rlabel metal3 20384 10808 20384 10808 0 _0263_
rlabel metal3 24472 7448 24472 7448 0 _0264_
rlabel metal2 21616 7224 21616 7224 0 _0265_
rlabel metal2 19432 12152 19432 12152 0 _0266_
rlabel metal2 23800 10920 23800 10920 0 _0267_
rlabel metal3 20328 11480 20328 11480 0 _0268_
rlabel metal2 23016 7280 23016 7280 0 _0269_
rlabel metal2 22400 9240 22400 9240 0 _0270_
rlabel metal3 21056 10584 21056 10584 0 _0271_
rlabel metal3 21784 10696 21784 10696 0 _0272_
rlabel metal2 24024 8960 24024 8960 0 _0273_
rlabel metal2 23800 9520 23800 9520 0 _0274_
rlabel metal2 22680 9968 22680 9968 0 _0275_
rlabel metal2 23688 11032 23688 11032 0 _0276_
rlabel metal2 33936 7672 33936 7672 0 _0277_
rlabel metal2 24752 9240 24752 9240 0 _0278_
rlabel metal3 24752 10584 24752 10584 0 _0279_
rlabel metal2 15624 13776 15624 13776 0 _0280_
rlabel metal2 25536 9240 25536 9240 0 _0281_
rlabel metal2 25704 10864 25704 10864 0 _0282_
rlabel metal2 28504 19712 28504 19712 0 _0283_
rlabel metal2 26264 18200 26264 18200 0 _0284_
rlabel metal2 26712 17640 26712 17640 0 _0285_
rlabel metal2 25648 13944 25648 13944 0 _0286_
rlabel metal2 25704 6720 25704 6720 0 _0287_
rlabel metal3 31192 6720 31192 6720 0 _0288_
rlabel metal2 24584 7000 24584 7000 0 _0289_
rlabel metal3 23856 7448 23856 7448 0 _0290_
rlabel metal2 25592 5040 25592 5040 0 _0291_
rlabel metal2 24192 6104 24192 6104 0 _0292_
rlabel metal2 26600 7504 26600 7504 0 _0293_
rlabel metal2 25144 7056 25144 7056 0 _0294_
rlabel metal2 25256 6048 25256 6048 0 _0295_
rlabel metal2 25480 5264 25480 5264 0 _0296_
rlabel metal2 26152 6664 26152 6664 0 _0297_
rlabel metal2 26600 5712 26600 5712 0 _0298_
rlabel metal2 26376 5320 26376 5320 0 _0299_
rlabel metal2 27720 6664 27720 6664 0 _0300_
rlabel metal2 27160 5432 27160 5432 0 _0301_
rlabel metal2 26712 8624 26712 8624 0 _0302_
rlabel metal2 27832 5096 27832 5096 0 _0303_
rlabel metal3 29288 9688 29288 9688 0 _0304_
rlabel metal2 30128 8120 30128 8120 0 _0305_
rlabel metal2 28952 6664 28952 6664 0 _0306_
rlabel metal2 29792 6664 29792 6664 0 _0307_
rlabel metal3 30240 10696 30240 10696 0 _0308_
rlabel metal2 30632 6776 30632 6776 0 _0309_
rlabel metal2 30576 6440 30576 6440 0 _0310_
rlabel metal3 30632 7448 30632 7448 0 _0311_
rlabel metal2 30856 7728 30856 7728 0 _0312_
rlabel metal2 29624 7840 29624 7840 0 _0313_
rlabel metal2 29960 8904 29960 8904 0 _0314_
rlabel metal2 31528 9464 31528 9464 0 _0315_
rlabel metal2 31192 8904 31192 8904 0 _0316_
rlabel metal2 30576 9240 30576 9240 0 _0317_
rlabel metal3 11816 17080 11816 17080 0 _0318_
rlabel metal2 29848 10136 29848 10136 0 _0319_
rlabel metal3 34048 30968 34048 30968 0 _0320_
rlabel metal2 32984 30744 32984 30744 0 _0321_
rlabel metal2 34216 29792 34216 29792 0 _0322_
rlabel metal2 21056 24696 21056 24696 0 _0323_
rlabel metal2 22008 25424 22008 25424 0 _0324_
rlabel metal2 19600 24920 19600 24920 0 _0325_
rlabel metal2 21896 25928 21896 25928 0 _0326_
rlabel metal3 21840 31528 21840 31528 0 _0327_
rlabel metal2 17752 30688 17752 30688 0 _0328_
rlabel metal3 16688 31192 16688 31192 0 _0329_
rlabel metal3 19824 30968 19824 30968 0 _0330_
rlabel metal2 22568 26600 22568 26600 0 _0331_
rlabel metal2 22680 26656 22680 26656 0 _0332_
rlabel metal2 20440 25592 20440 25592 0 _0333_
rlabel metal2 21672 26264 21672 26264 0 _0334_
rlabel metal3 18424 25480 18424 25480 0 _0335_
rlabel metal2 21448 25872 21448 25872 0 _0336_
rlabel metal3 17192 27048 17192 27048 0 _0337_
rlabel metal2 18984 28504 18984 28504 0 _0338_
rlabel metal2 22904 25200 22904 25200 0 _0339_
rlabel metal2 23688 25704 23688 25704 0 _0340_
rlabel metal3 18312 26488 18312 26488 0 _0341_
rlabel metal2 23352 25368 23352 25368 0 _0342_
rlabel metal3 14224 20776 14224 20776 0 _0343_
rlabel metal3 21056 22232 21056 22232 0 _0344_
rlabel metal2 27440 11368 27440 11368 0 _0345_
rlabel metal2 28000 11592 28000 11592 0 _0346_
rlabel metal2 31192 13048 31192 13048 0 _0347_
rlabel metal2 17752 18928 17752 18928 0 _0348_
rlabel via3 15400 21681 15400 21681 0 _0349_
rlabel metal2 21560 22624 21560 22624 0 _0350_
rlabel metal2 21448 20888 21448 20888 0 _0351_
rlabel metal2 18648 23128 18648 23128 0 _0352_
rlabel metal2 21896 23016 21896 23016 0 _0353_
rlabel metal2 24696 22792 24696 22792 0 _0354_
rlabel metal2 29400 24360 29400 24360 0 _0355_
rlabel metal3 31584 30968 31584 30968 0 _0356_
rlabel metal2 24304 23352 24304 23352 0 _0357_
rlabel metal2 28168 31976 28168 31976 0 _0358_
rlabel metal2 31752 13328 31752 13328 0 _0359_
rlabel metal2 26040 12432 26040 12432 0 _0360_
rlabel metal2 8232 18648 8232 18648 0 _0361_
rlabel metal2 9016 17024 9016 17024 0 _0362_
rlabel metal2 8232 20496 8232 20496 0 _0363_
rlabel metal2 7784 19544 7784 19544 0 _0364_
rlabel metal2 7896 18536 7896 18536 0 _0365_
rlabel metal3 9016 19992 9016 19992 0 _0366_
rlabel metal2 8792 19600 8792 19600 0 _0367_
rlabel metal2 7056 21784 7056 21784 0 _0368_
rlabel metal2 6664 21224 6664 21224 0 _0369_
rlabel metal3 12040 22232 12040 22232 0 _0370_
rlabel metal2 7672 22456 7672 22456 0 _0371_
rlabel metal2 10136 21952 10136 21952 0 _0372_
rlabel metal2 7112 23408 7112 23408 0 _0373_
rlabel metal2 11760 21672 11760 21672 0 _0374_
rlabel metal2 9464 23352 9464 23352 0 _0375_
rlabel metal3 8960 23128 8960 23128 0 _0376_
rlabel metal2 11368 23520 11368 23520 0 _0377_
rlabel metal2 10920 23520 10920 23520 0 _0378_
rlabel metal2 11704 20664 11704 20664 0 _0379_
rlabel metal2 11480 20272 11480 20272 0 _0380_
rlabel metal3 13496 17640 13496 17640 0 _0381_
rlabel metal3 11928 19992 11928 19992 0 _0382_
rlabel metal3 13832 19208 13832 19208 0 _0383_
rlabel metal2 13160 20048 13160 20048 0 _0384_
rlabel metal2 13832 18984 13832 18984 0 _0385_
rlabel metal2 12712 18088 12712 18088 0 _0386_
rlabel metal2 12376 17920 12376 17920 0 _0387_
rlabel metal3 14056 17528 14056 17528 0 _0388_
rlabel metal2 13440 17640 13440 17640 0 _0389_
rlabel metal2 15400 19600 15400 19600 0 _0390_
rlabel metal2 14728 19208 14728 19208 0 _0391_
rlabel metal2 15624 19488 15624 19488 0 _0392_
rlabel metal3 16968 18424 16968 18424 0 _0393_
rlabel metal3 18704 20104 18704 20104 0 _0394_
rlabel metal2 17136 18424 17136 18424 0 _0395_
rlabel metal2 16744 21392 16744 21392 0 _0396_
rlabel metal2 16408 20776 16408 20776 0 _0397_
rlabel metal3 18368 20664 18368 20664 0 _0398_
rlabel metal2 17976 20272 17976 20272 0 _0399_
rlabel metal2 17808 23128 17808 23128 0 _0400_
rlabel metal3 18760 22568 18760 22568 0 _0401_
rlabel metal2 17472 24920 17472 24920 0 _0402_
rlabel metal3 18592 24696 18592 24696 0 _0403_
rlabel metal2 16744 25984 16744 25984 0 _0404_
rlabel metal2 15848 27104 15848 27104 0 _0405_
rlabel metal2 8008 25704 8008 25704 0 _0406_
rlabel metal2 8344 26768 8344 26768 0 _0407_
rlabel metal3 19320 27048 19320 27048 0 _0408_
rlabel metal2 7784 26852 7784 26852 0 _0409_
rlabel metal3 7112 26488 7112 26488 0 _0410_
rlabel metal2 12936 27160 12936 27160 0 _0411_
rlabel metal2 7448 25648 7448 25648 0 _0412_
rlabel metal2 5992 27496 5992 27496 0 _0413_
rlabel metal2 7672 26712 7672 26712 0 _0414_
rlabel metal2 7784 25928 7784 25928 0 _0415_
rlabel metal3 8960 24696 8960 24696 0 _0416_
rlabel metal2 7056 24920 7056 24920 0 _0417_
rlabel metal2 7560 26600 7560 26600 0 _0418_
rlabel metal2 7560 28056 7560 28056 0 _0419_
rlabel metal2 21560 29344 21560 29344 0 _0420_
rlabel metal2 16520 26264 16520 26264 0 _0421_
rlabel metal2 6832 29960 6832 29960 0 _0422_
rlabel metal2 8344 28952 8344 28952 0 _0423_
rlabel metal2 8680 26712 8680 26712 0 _0424_
rlabel metal2 11928 27104 11928 27104 0 _0425_
rlabel metal2 9128 29064 9128 29064 0 _0426_
rlabel metal2 10024 29400 10024 29400 0 _0427_
rlabel metal2 10808 28896 10808 28896 0 _0428_
rlabel metal2 17416 26600 17416 26600 0 _0429_
rlabel metal2 11032 29344 11032 29344 0 _0430_
rlabel metal2 12264 29120 12264 29120 0 _0431_
rlabel metal2 7560 25088 7560 25088 0 _0432_
rlabel metal2 9576 30240 9576 30240 0 _0433_
rlabel metal2 9240 30968 9240 30968 0 _0434_
rlabel metal2 11368 30240 11368 30240 0 _0435_
rlabel metal2 9576 26880 9576 26880 0 _0436_
rlabel metal2 8120 24976 8120 24976 0 _0437_
rlabel metal2 9744 28392 9744 28392 0 _0438_
rlabel metal2 9912 28952 9912 28952 0 _0439_
rlabel via2 12264 24920 12264 24920 0 _0440_
rlabel metal3 12040 26376 12040 26376 0 _0441_
rlabel metal2 11368 26544 11368 26544 0 _0442_
rlabel metal2 10472 25872 10472 25872 0 _0443_
rlabel metal3 8288 25368 8288 25368 0 _0444_
rlabel metal2 6440 26264 6440 26264 0 _0445_
rlabel metal2 12600 25088 12600 25088 0 _0446_
rlabel metal2 12152 25872 12152 25872 0 _0447_
rlabel metal2 12712 25816 12712 25816 0 _0448_
rlabel metal2 13048 26180 13048 26180 0 _0449_
rlabel metal2 12320 25704 12320 25704 0 _0450_
rlabel metal2 14000 27048 14000 27048 0 _0451_
rlabel metal2 13272 28112 13272 28112 0 _0452_
rlabel metal2 18144 27048 18144 27048 0 _0453_
rlabel metal2 13608 25872 13608 25872 0 _0454_
rlabel metal2 13664 26824 13664 26824 0 _0455_
rlabel metal2 13832 27384 13832 27384 0 _0456_
rlabel metal2 18256 29512 18256 29512 0 _0457_
rlabel metal2 15344 25480 15344 25480 0 _0458_
rlabel metal3 16744 28728 16744 28728 0 _0459_
rlabel metal2 17752 29064 17752 29064 0 _0460_
rlabel metal3 16800 29400 16800 29400 0 _0461_
rlabel metal3 22288 31080 22288 31080 0 _0462_
rlabel metal2 15288 24696 15288 24696 0 _0463_
rlabel metal3 21504 31752 21504 31752 0 _0464_
rlabel metal2 17080 28840 17080 28840 0 _0465_
rlabel metal3 17976 29624 17976 29624 0 _0466_
rlabel metal3 16968 28560 16968 28560 0 _0467_
rlabel metal2 16520 30688 16520 30688 0 _0468_
rlabel metal2 18200 28056 18200 28056 0 _0469_
rlabel metal3 16296 27944 16296 27944 0 _0470_
rlabel metal2 15400 27496 15400 27496 0 _0471_
rlabel metal2 15232 24920 15232 24920 0 _0472_
rlabel metal2 14616 28112 14616 28112 0 _0473_
rlabel metal2 13496 29400 13496 29400 0 _0474_
rlabel metal2 20328 23576 20328 23576 0 _0475_
rlabel metal2 19712 27272 19712 27272 0 _0476_
rlabel metal2 18536 27160 18536 27160 0 _0477_
rlabel metal2 19096 28224 19096 28224 0 _0478_
rlabel metal2 19432 29512 19432 29512 0 _0479_
rlabel metal3 23128 30968 23128 30968 0 _0480_
rlabel metal3 22064 30856 22064 30856 0 _0481_
rlabel metal2 21448 31696 21448 31696 0 _0482_
rlabel metal2 20104 28056 20104 28056 0 _0483_
rlabel metal3 20944 27720 20944 27720 0 _0484_
rlabel metal2 18200 25536 18200 25536 0 _0485_
rlabel metal2 18872 25592 18872 25592 0 _0486_
rlabel metal2 21784 30968 21784 30968 0 _0487_
rlabel metal2 26264 28112 26264 28112 0 _0488_
rlabel metal2 25592 27832 25592 27832 0 _0489_
rlabel metal2 20608 26824 20608 26824 0 _0490_
rlabel metal3 21504 26488 21504 26488 0 _0491_
rlabel metal2 20104 25088 20104 25088 0 _0492_
rlabel metal2 19880 24920 19880 24920 0 _0493_
rlabel metal2 21896 29400 21896 29400 0 _0494_
rlabel metal2 10248 14616 10248 14616 0 _0495_
rlabel metal2 10696 13776 10696 13776 0 _0496_
rlabel metal3 11424 12936 11424 12936 0 _0497_
rlabel metal3 10192 11480 10192 11480 0 _0498_
rlabel metal2 7448 8960 7448 8960 0 _0499_
rlabel metal2 10472 5600 10472 5600 0 _0500_
rlabel metal2 8232 9016 8232 9016 0 _0501_
rlabel metal3 8792 7560 8792 7560 0 _0502_
rlabel metal3 9744 8232 9744 8232 0 _0503_
rlabel metal2 8624 8344 8624 8344 0 _0504_
rlabel metal2 9240 3640 9240 3640 0 _0505_
rlabel metal2 6552 7000 6552 7000 0 _0506_
rlabel metal2 10136 5824 10136 5824 0 _0507_
rlabel metal3 6776 7448 6776 7448 0 _0508_
rlabel metal2 6440 8120 6440 8120 0 _0509_
rlabel metal2 7336 8232 7336 8232 0 _0510_
rlabel metal3 34426 2296 34426 2296 0 clk_i
rlabel metal2 21672 17920 21672 17920 0 clknet_0_clk_i
rlabel metal2 6104 4704 6104 4704 0 clknet_3_0__leaf_clk_i
rlabel metal2 19320 8680 19320 8680 0 clknet_3_1__leaf_clk_i
rlabel metal3 12096 18424 12096 18424 0 clknet_3_2__leaf_clk_i
rlabel metal2 15736 23128 15736 23128 0 clknet_3_3__leaf_clk_i
rlabel metal2 26152 20776 26152 20776 0 clknet_3_4__leaf_clk_i
rlabel metal2 24248 9408 24248 9408 0 clknet_3_5__leaf_clk_i
rlabel metal3 21616 23128 21616 23128 0 clknet_3_6__leaf_clk_i
rlabel metal2 32424 25396 32424 25396 0 clknet_3_7__leaf_clk_i
rlabel metal2 35224 33600 35224 33600 0 custom_setting
rlabel metal2 8120 19264 8120 19264 0 dest\[0\]
rlabel metal2 15512 23296 15512 23296 0 dest\[10\]
rlabel metal2 16800 20104 16800 20104 0 dest\[11\]
rlabel metal2 19432 19376 19432 19376 0 dest\[12\]
rlabel metal2 18312 23352 18312 23352 0 dest\[13\]
rlabel metal2 19488 22232 19488 22232 0 dest\[14\]
rlabel metal2 19208 23856 19208 23856 0 dest\[15\]
rlabel metal3 21952 23912 21952 23912 0 dest\[16\]
rlabel metal2 7560 19712 7560 19712 0 dest\[1\]
rlabel metal2 7896 19824 7896 19824 0 dest\[2\]
rlabel metal2 7224 23912 7224 23912 0 dest\[3\]
rlabel metal2 8232 23408 8232 23408 0 dest\[4\]
rlabel metal2 8904 22848 8904 22848 0 dest\[5\]
rlabel metal3 11984 24808 11984 24808 0 dest\[6\]
rlabel metal2 12824 20720 12824 20720 0 dest\[7\]
rlabel metal2 12376 19544 12376 19544 0 dest\[8\]
rlabel metal2 13720 19264 13720 19264 0 dest\[9\]
rlabel metal2 16408 8904 16408 8904 0 dia\[0\]
rlabel metal2 15288 7840 15288 7840 0 dia\[1\]
rlabel metal2 15848 10192 15848 10192 0 dia\[2\]
rlabel metal2 16856 11760 16856 11760 0 dia\[3\]
rlabel metal2 20552 11032 20552 11032 0 dia\[4\]
rlabel metal2 22624 9576 22624 9576 0 dia\[5\]
rlabel metal2 24360 11144 24360 11144 0 dia\[6\]
rlabel metal2 25144 10920 25144 10920 0 dia\[7\]
rlabel metal2 24360 6216 24360 6216 0 dib\[0\]
rlabel metal2 25312 4984 25312 4984 0 dib\[1\]
rlabel metal2 26264 4704 26264 4704 0 dib\[2\]
rlabel metal2 28168 6272 28168 6272 0 dib\[3\]
rlabel metal3 30968 7560 30968 7560 0 dib\[4\]
rlabel metal3 32480 8232 32480 8232 0 dib\[5\]
rlabel metal3 31192 9016 31192 9016 0 dib\[6\]
rlabel metal2 33096 16072 33096 16072 0 dib\[7\]
rlabel metal3 35770 7672 35770 7672 0 io_in[0]
rlabel metal2 34216 10472 34216 10472 0 io_in[1]
rlabel metal2 33880 12208 33880 12208 0 io_in[2]
rlabel metal3 35616 15512 35616 15512 0 io_in[3]
rlabel metal2 35056 12152 35056 12152 0 io_in[4]
rlabel metal3 34538 21112 34538 21112 0 io_in[5]
rlabel metal3 25760 21672 25760 21672 0 io_in[6]
rlabel metal3 35602 26488 35602 26488 0 io_in[7]
rlabel metal2 12824 34482 12824 34482 0 io_out[10]
rlabel metal3 13160 33544 13160 33544 0 io_out[11]
rlabel metal2 15064 33306 15064 33306 0 io_out[12]
rlabel metal2 16072 32536 16072 32536 0 io_out[13]
rlabel metal2 17304 34818 17304 34818 0 io_out[14]
rlabel metal2 18424 34874 18424 34874 0 io_out[15]
rlabel metal2 19544 33698 19544 33698 0 io_out[16]
rlabel metal2 20664 34874 20664 34874 0 io_out[17]
rlabel metal3 24024 32424 24024 32424 0 io_out[18]
rlabel metal2 22904 35042 22904 35042 0 io_out[19]
rlabel metal2 26264 30128 26264 30128 0 io_out[20]
rlabel metal2 25368 30520 25368 30520 0 io_out[21]
rlabel metal2 26488 32088 26488 32088 0 io_out[22]
rlabel metal3 35392 21000 35392 21000 0 io_out[23]
rlabel metal2 30632 29008 30632 29008 0 io_out[24]
rlabel metal2 29624 34874 29624 34874 0 io_out[25]
rlabel metal2 30800 29736 30800 29736 0 io_out[26]
rlabel metal2 31304 36232 31304 36232 0 io_out[27]
rlabel metal2 30296 25732 30296 25732 0 io_out[28]
rlabel metal3 31360 27160 31360 27160 0 io_out[29]
rlabel metal3 28224 26488 28224 26488 0 io_out[30]
rlabel metal2 8232 33488 8232 33488 0 io_out[8]
rlabel metal2 11816 30968 11816 30968 0 io_out[9]
rlabel metal3 11536 12824 11536 12824 0 mar\[0\]
rlabel metal2 9688 11424 9688 11424 0 mar\[1\]
rlabel metal2 25144 16968 25144 16968 0 mc14500.DATA_OUT
rlabel metal2 27888 10472 27888 10472 0 mc14500.IEN_l
rlabel metal2 24696 13104 24696 13104 0 mc14500.OEN_l
rlabel metal2 16632 14280 16632 14280 0 mc14500.X1
rlabel metal2 32312 13272 32312 13272 0 mc14500.instr_l\[0\]
rlabel metal3 33040 11928 33040 11928 0 mc14500.instr_l\[1\]
rlabel metal3 33152 15064 33152 15064 0 mc14500.instr_l\[2\]
rlabel metal2 33096 16352 33096 16352 0 mc14500.instr_l\[3\]
rlabel metal2 20440 14392 20440 14392 0 mc14500.skip
rlabel metal3 35560 16072 35560 16072 0 net1
rlabel metal2 34552 19544 34552 19544 0 net10
rlabel metal2 29680 16968 29680 16968 0 net11
rlabel metal2 24472 8064 24472 8064 0 net12
rlabel metal2 27496 3808 27496 3808 0 net13
rlabel metal2 24248 3976 24248 3976 0 net14
rlabel metal2 29008 3416 29008 3416 0 net15
rlabel metal2 30296 3808 30296 3808 0 net16
rlabel metal2 32144 3416 32144 3416 0 net17
rlabel metal3 32872 3304 32872 3304 0 net18
rlabel metal2 34832 4648 34832 4648 0 net19
rlabel metal3 29624 31752 29624 31752 0 net2
rlabel metal3 10640 30072 10640 30072 0 net20
rlabel metal2 9016 32872 9016 32872 0 net21
rlabel metal2 11592 31416 11592 31416 0 net22
rlabel metal2 6552 26516 6552 26516 0 net23
rlabel metal2 16296 31024 16296 31024 0 net24
rlabel metal3 16520 32424 16520 32424 0 net25
rlabel metal2 19880 33096 19880 33096 0 net26
rlabel metal3 22624 31864 22624 31864 0 net27
rlabel metal3 20664 33432 20664 33432 0 net28
rlabel metal2 22456 32088 22456 32088 0 net29
rlabel metal2 34664 10360 34664 10360 0 net3
rlabel metal3 24024 29400 24024 29400 0 net30
rlabel metal2 26656 25704 26656 25704 0 net31
rlabel metal2 26600 27944 26600 27944 0 net32
rlabel metal3 25144 26488 25144 26488 0 net33
rlabel metal2 23912 25984 23912 25984 0 net34
rlabel metal2 28728 30800 28728 30800 0 net35
rlabel metal2 28616 17192 28616 17192 0 net36
rlabel metal2 29960 25312 29960 25312 0 net37
rlabel metal2 32088 23912 32088 23912 0 net38
rlabel metal2 31528 26572 31528 26572 0 net39
rlabel metal3 32256 12264 32256 12264 0 net4
rlabel metal2 26712 29232 26712 29232 0 net40
rlabel metal3 7336 30184 7336 30184 0 net41
rlabel metal2 10472 30576 10472 30576 0 net42
rlabel metal2 4872 8568 4872 8568 0 net43
rlabel metal2 5656 10920 5656 10920 0 net44
rlabel metal2 4200 6216 4200 6216 0 net45
rlabel metal2 8792 5040 8792 5040 0 net46
rlabel metal2 9016 5376 9016 5376 0 net47
rlabel metal2 9688 6160 9688 6160 0 net48
rlabel metal3 33544 31080 33544 31080 0 net49
rlabel metal2 34272 11256 34272 11256 0 net5
rlabel metal3 9688 8344 9688 8344 0 net50
rlabel metal2 10472 4144 10472 4144 0 net51
rlabel metal2 9800 5600 9800 5600 0 net52
rlabel metal2 14560 5768 14560 5768 0 net53
rlabel metal2 13944 3864 13944 3864 0 net54
rlabel metal2 18424 3976 18424 3976 0 net55
rlabel metal3 17808 6440 17808 6440 0 net56
rlabel metal3 23744 4424 23744 4424 0 net57
rlabel metal2 18872 27048 18872 27048 0 net58
rlabel metal2 17640 31192 17640 31192 0 net59
rlabel metal2 33656 16744 33656 16744 0 net6
rlabel metal3 16072 30856 16072 30856 0 net60
rlabel metal2 10192 29624 10192 29624 0 net61
rlabel metal2 33768 12880 33768 12880 0 net62
rlabel metal2 35056 14504 35056 14504 0 net63
rlabel metal2 31528 15148 31528 15148 0 net64
rlabel metal2 30520 10808 30520 10808 0 net65
rlabel metal2 19880 14448 19880 14448 0 net66
rlabel metal2 1736 33208 1736 33208 0 net67
rlabel metal2 2856 33208 2856 33208 0 net68
rlabel metal2 3976 33208 3976 33208 0 net69
rlabel metal2 34216 16800 34216 16800 0 net7
rlabel metal2 4984 34706 4984 34706 0 net70
rlabel metal2 5992 33208 5992 33208 0 net71
rlabel metal2 7448 32760 7448 32760 0 net72
rlabel metal3 8960 32760 8960 32760 0 net73
rlabel metal2 9520 33208 9520 33208 0 net74
rlabel metal2 22792 13888 22792 13888 0 net75
rlabel metal2 22344 14000 22344 14000 0 net76
rlabel metal2 22568 21392 22568 21392 0 net8
rlabel metal2 34272 26488 34272 26488 0 net9
rlabel metal2 33656 31752 33656 31752 0 rst_latency\[0\]
rlabel metal2 34440 29960 34440 29960 0 rst_latency\[1\]
rlabel metal3 35224 5040 35224 5040 0 rst_n
rlabel metal2 25816 22232 25816 22232 0 scratch\[0\]
rlabel metal2 24360 23688 24360 23688 0 scratch\[1\]
rlabel metal2 28168 23072 28168 23072 0 scratch\[2\]
rlabel metal2 27888 25704 27888 25704 0 scratch\[3\]
rlabel metal2 34888 26040 34888 26040 0 scratch\[4\]
rlabel metal2 35224 23632 35224 23632 0 scratch\[5\]
rlabel metal2 1848 2982 1848 2982 0 sram_addr[0]
rlabel metal2 3416 2478 3416 2478 0 sram_addr[1]
rlabel metal3 4480 3416 4480 3416 0 sram_addr[2]
rlabel metal2 6664 4200 6664 4200 0 sram_addr[3]
rlabel metal2 8120 2030 8120 2030 0 sram_addr[4]
rlabel metal2 9688 2058 9688 2058 0 sram_addr[5]
rlabel metal3 35616 22568 35616 22568 0 sram_gwe
rlabel metal2 11256 3654 11256 3654 0 sram_in[0]
rlabel metal2 12824 2058 12824 2058 0 sram_in[1]
rlabel metal2 14392 1302 14392 1302 0 sram_in[2]
rlabel metal2 15960 2198 15960 2198 0 sram_in[3]
rlabel metal3 18088 3640 18088 3640 0 sram_in[4]
rlabel metal3 20496 3640 20496 3640 0 sram_in[5]
rlabel metal3 21280 5656 21280 5656 0 sram_in[6]
rlabel metal3 23912 3640 23912 3640 0 sram_in[7]
rlabel metal2 23800 2478 23800 2478 0 sram_out[0]
rlabel metal2 25368 2086 25368 2086 0 sram_out[1]
rlabel metal2 27104 2744 27104 2744 0 sram_out[2]
rlabel metal3 30240 3528 30240 3528 0 sram_out[3]
rlabel metal3 31080 3416 31080 3416 0 sram_out[4]
rlabel metal3 32032 3528 32032 3528 0 sram_out[5]
rlabel metal2 33264 4200 33264 4200 0 sram_out[6]
rlabel metal2 34944 3080 34944 3080 0 sram_out[7]
<< properties >>
string FIXED_BBOX 0 0 37000 37000
<< end >>
