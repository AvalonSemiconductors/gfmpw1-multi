magic
tech gf180mcuD
magscale 1 10
timestamp 1702047371
<< metal1 >>
rect 1344 56474 58576 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 58576 56474
rect 1344 56388 58576 56422
rect 22430 56306 22482 56318
rect 22430 56242 22482 56254
rect 22654 56306 22706 56318
rect 22654 56242 22706 56254
rect 27022 56306 27074 56318
rect 27022 56242 27074 56254
rect 37438 56306 37490 56318
rect 37438 56242 37490 56254
rect 37662 56306 37714 56318
rect 37662 56242 37714 56254
rect 52446 56306 52498 56318
rect 52446 56242 52498 56254
rect 57822 56194 57874 56206
rect 52658 56142 52670 56194
rect 52722 56142 52734 56194
rect 57822 56130 57874 56142
rect 26686 56082 26738 56094
rect 26686 56018 26738 56030
rect 27134 56082 27186 56094
rect 27134 56018 27186 56030
rect 27358 56082 27410 56094
rect 57598 56082 57650 56094
rect 52882 56030 52894 56082
rect 52946 56030 52958 56082
rect 27358 56018 27410 56030
rect 57598 56018 57650 56030
rect 58158 56082 58210 56094
rect 58158 56018 58210 56030
rect 38222 55970 38274 55982
rect 23090 55918 23102 55970
rect 23154 55918 23166 55970
rect 38222 55906 38274 55918
rect 1344 55690 58576 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 58576 55690
rect 1344 55604 58576 55638
rect 57598 55410 57650 55422
rect 20402 55358 20414 55410
rect 20466 55358 20478 55410
rect 25778 55358 25790 55410
rect 25842 55358 25854 55410
rect 29138 55358 29150 55410
rect 29202 55358 29214 55410
rect 36418 55358 36430 55410
rect 36482 55358 36494 55410
rect 40226 55358 40238 55410
rect 40290 55358 40302 55410
rect 42690 55358 42702 55410
rect 42754 55358 42766 55410
rect 48850 55358 48862 55410
rect 48914 55358 48926 55410
rect 52098 55358 52110 55410
rect 52162 55358 52174 55410
rect 55570 55358 55582 55410
rect 55634 55358 55646 55410
rect 57598 55346 57650 55358
rect 21646 55298 21698 55310
rect 17490 55246 17502 55298
rect 17554 55246 17566 55298
rect 21646 55234 21698 55246
rect 21982 55298 22034 55310
rect 40798 55298 40850 55310
rect 22978 55246 22990 55298
rect 23042 55246 23054 55298
rect 27682 55246 27694 55298
rect 27746 55246 27758 55298
rect 32050 55246 32062 55298
rect 32114 55246 32126 55298
rect 33506 55246 33518 55298
rect 33570 55246 33582 55298
rect 37314 55246 37326 55298
rect 37378 55246 37390 55298
rect 21982 55234 22034 55246
rect 40798 55234 40850 55246
rect 41022 55298 41074 55310
rect 42366 55298 42418 55310
rect 41234 55246 41246 55298
rect 41298 55246 41310 55298
rect 46050 55246 46062 55298
rect 46114 55246 46126 55298
rect 49298 55246 49310 55298
rect 49362 55246 49374 55298
rect 52658 55246 52670 55298
rect 52722 55246 52734 55298
rect 41022 55234 41074 55246
rect 42366 55234 42418 55246
rect 21310 55186 21362 55198
rect 27358 55186 27410 55198
rect 18274 55134 18286 55186
rect 18338 55134 18350 55186
rect 23650 55134 23662 55186
rect 23714 55134 23726 55186
rect 21310 55122 21362 55134
rect 27358 55122 27410 55134
rect 27470 55186 27522 55198
rect 40686 55186 40738 55198
rect 31266 55134 31278 55186
rect 31330 55134 31342 55186
rect 34290 55134 34302 55186
rect 34354 55134 34366 55186
rect 38098 55134 38110 55186
rect 38162 55134 38174 55186
rect 46722 55134 46734 55186
rect 46786 55134 46798 55186
rect 49970 55134 49982 55186
rect 50034 55134 50046 55186
rect 53442 55134 53454 55186
rect 53506 55134 53518 55186
rect 27470 55122 27522 55134
rect 40686 55122 40738 55134
rect 21646 55074 21698 55086
rect 42590 55074 42642 55086
rect 26898 55022 26910 55074
rect 26962 55022 26974 55074
rect 21646 55010 21698 55022
rect 42590 55010 42642 55022
rect 57486 55074 57538 55086
rect 57486 55010 57538 55022
rect 1344 54906 58576 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 58576 54906
rect 1344 54820 58576 54854
rect 22766 54738 22818 54750
rect 22766 54674 22818 54686
rect 23774 54738 23826 54750
rect 23774 54674 23826 54686
rect 40238 54738 40290 54750
rect 41806 54738 41858 54750
rect 41458 54686 41470 54738
rect 41522 54686 41534 54738
rect 40238 54674 40290 54686
rect 41806 54674 41858 54686
rect 47406 54738 47458 54750
rect 47406 54674 47458 54686
rect 54462 54738 54514 54750
rect 54462 54674 54514 54686
rect 40126 54626 40178 54638
rect 54574 54626 54626 54638
rect 25442 54574 25454 54626
rect 25506 54574 25518 54626
rect 36866 54574 36878 54626
rect 36930 54574 36942 54626
rect 42130 54574 42142 54626
rect 42194 54574 42206 54626
rect 51986 54574 51998 54626
rect 52050 54574 52062 54626
rect 40126 54562 40178 54574
rect 54574 54562 54626 54574
rect 36542 54514 36594 54526
rect 17490 54462 17502 54514
rect 17554 54462 17566 54514
rect 20626 54462 20638 54514
rect 20690 54462 20702 54514
rect 21858 54462 21870 54514
rect 21922 54462 21934 54514
rect 22978 54462 22990 54514
rect 23042 54462 23054 54514
rect 23538 54462 23550 54514
rect 23602 54462 23614 54514
rect 29026 54462 29038 54514
rect 29090 54462 29102 54514
rect 31378 54462 31390 54514
rect 31442 54462 31454 54514
rect 36542 54450 36594 54462
rect 40910 54514 40962 54526
rect 45490 54462 45502 54514
rect 45554 54462 45566 54514
rect 46498 54462 46510 54514
rect 46562 54462 46574 54514
rect 46722 54462 46734 54514
rect 46786 54462 46798 54514
rect 47618 54462 47630 54514
rect 47682 54462 47694 54514
rect 52882 54462 52894 54514
rect 52946 54462 52958 54514
rect 40910 54450 40962 54462
rect 22318 54402 22370 54414
rect 18162 54350 18174 54402
rect 18226 54350 18238 54402
rect 20290 54350 20302 54402
rect 20354 54350 20366 54402
rect 20962 54350 20974 54402
rect 21026 54350 21038 54402
rect 21522 54350 21534 54402
rect 21586 54350 21598 54402
rect 22318 54338 22370 54350
rect 22654 54402 22706 54414
rect 22654 54338 22706 54350
rect 24782 54402 24834 54414
rect 46958 54402 47010 54414
rect 42578 54350 42590 54402
rect 42642 54350 42654 54402
rect 44706 54350 44718 54402
rect 44770 54350 44782 54402
rect 24782 54338 24834 54350
rect 46958 54338 47010 54350
rect 47294 54402 47346 54414
rect 47294 54338 47346 54350
rect 48302 54402 48354 54414
rect 48302 54338 48354 54350
rect 23886 54290 23938 54302
rect 23886 54226 23938 54238
rect 31614 54290 31666 54302
rect 31614 54226 31666 54238
rect 31838 54290 31890 54302
rect 31838 54226 31890 54238
rect 31950 54290 32002 54302
rect 31950 54226 32002 54238
rect 40350 54290 40402 54302
rect 40350 54226 40402 54238
rect 41134 54290 41186 54302
rect 41134 54226 41186 54238
rect 54350 54290 54402 54302
rect 54350 54226 54402 54238
rect 1344 54122 58576 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 58576 54122
rect 1344 54036 58576 54070
rect 20638 53954 20690 53966
rect 20638 53890 20690 53902
rect 26910 53954 26962 53966
rect 26910 53890 26962 53902
rect 27134 53954 27186 53966
rect 27134 53890 27186 53902
rect 29486 53954 29538 53966
rect 29486 53890 29538 53902
rect 37438 53954 37490 53966
rect 43150 53954 43202 53966
rect 40338 53902 40350 53954
rect 40402 53902 40414 53954
rect 40562 53902 40574 53954
rect 40626 53951 40638 53954
rect 40898 53951 40910 53954
rect 40626 53905 40910 53951
rect 40626 53902 40638 53905
rect 40898 53902 40910 53905
rect 40962 53902 40974 53954
rect 37438 53890 37490 53902
rect 43150 53890 43202 53902
rect 50766 53954 50818 53966
rect 50766 53890 50818 53902
rect 29374 53842 29426 53854
rect 26114 53790 26126 53842
rect 26178 53790 26190 53842
rect 29374 53778 29426 53790
rect 29710 53842 29762 53854
rect 35870 53842 35922 53854
rect 31266 53790 31278 53842
rect 31330 53790 31342 53842
rect 33394 53790 33406 53842
rect 33458 53790 33470 53842
rect 29710 53778 29762 53790
rect 35870 53778 35922 53790
rect 39118 53842 39170 53854
rect 39118 53778 39170 53790
rect 40014 53842 40066 53854
rect 40014 53778 40066 53790
rect 41134 53842 41186 53854
rect 41134 53778 41186 53790
rect 50542 53842 50594 53854
rect 50542 53778 50594 53790
rect 51438 53842 51490 53854
rect 52770 53790 52782 53842
rect 52834 53790 52846 53842
rect 51438 53778 51490 53790
rect 20190 53730 20242 53742
rect 20190 53666 20242 53678
rect 20302 53730 20354 53742
rect 20302 53666 20354 53678
rect 20526 53730 20578 53742
rect 20526 53666 20578 53678
rect 21870 53730 21922 53742
rect 22878 53730 22930 53742
rect 22082 53678 22094 53730
rect 22146 53678 22158 53730
rect 21870 53666 21922 53678
rect 22878 53666 22930 53678
rect 25230 53730 25282 53742
rect 27246 53730 27298 53742
rect 25890 53678 25902 53730
rect 25954 53678 25966 53730
rect 25230 53666 25282 53678
rect 27246 53666 27298 53678
rect 27582 53730 27634 53742
rect 28254 53730 28306 53742
rect 27906 53678 27918 53730
rect 27970 53678 27982 53730
rect 27582 53666 27634 53678
rect 28254 53666 28306 53678
rect 28478 53730 28530 53742
rect 28478 53666 28530 53678
rect 29822 53730 29874 53742
rect 36094 53730 36146 53742
rect 36990 53730 37042 53742
rect 34066 53678 34078 53730
rect 34130 53678 34142 53730
rect 36418 53678 36430 53730
rect 36482 53678 36494 53730
rect 29822 53666 29874 53678
rect 36094 53666 36146 53678
rect 36990 53666 37042 53678
rect 37102 53730 37154 53742
rect 37102 53666 37154 53678
rect 37326 53730 37378 53742
rect 39790 53730 39842 53742
rect 39442 53678 39454 53730
rect 39506 53678 39518 53730
rect 37326 53666 37378 53678
rect 39790 53666 39842 53678
rect 41358 53730 41410 53742
rect 43038 53730 43090 53742
rect 41682 53678 41694 53730
rect 41746 53678 41758 53730
rect 41358 53666 41410 53678
rect 43038 53666 43090 53678
rect 43374 53730 43426 53742
rect 43374 53666 43426 53678
rect 43486 53730 43538 53742
rect 43486 53666 43538 53678
rect 48638 53730 48690 53742
rect 48638 53666 48690 53678
rect 50430 53730 50482 53742
rect 50430 53666 50482 53678
rect 50878 53730 50930 53742
rect 53678 53730 53730 53742
rect 55022 53730 55074 53742
rect 51650 53678 51662 53730
rect 51714 53678 51726 53730
rect 53218 53678 53230 53730
rect 53282 53678 53294 53730
rect 54226 53678 54238 53730
rect 54290 53678 54302 53730
rect 50878 53666 50930 53678
rect 53678 53666 53730 53678
rect 55022 53666 55074 53678
rect 55358 53730 55410 53742
rect 55358 53666 55410 53678
rect 21758 53618 21810 53630
rect 21758 53554 21810 53566
rect 28366 53618 28418 53630
rect 51326 53618 51378 53630
rect 55582 53618 55634 53630
rect 30930 53566 30942 53618
rect 30994 53566 31006 53618
rect 41570 53566 41582 53618
rect 41634 53566 41646 53618
rect 54002 53566 54014 53618
rect 54066 53566 54078 53618
rect 28366 53554 28418 53566
rect 51326 53554 51378 53566
rect 55582 53554 55634 53566
rect 22990 53506 23042 53518
rect 21298 53454 21310 53506
rect 21362 53454 21374 53506
rect 22990 53442 23042 53454
rect 27246 53506 27298 53518
rect 27246 53442 27298 53454
rect 30606 53506 30658 53518
rect 30606 53442 30658 53454
rect 37998 53506 38050 53518
rect 37998 53442 38050 53454
rect 39230 53506 39282 53518
rect 39230 53442 39282 53454
rect 40798 53506 40850 53518
rect 40798 53442 40850 53454
rect 42142 53506 42194 53518
rect 42142 53442 42194 53454
rect 48750 53506 48802 53518
rect 48750 53442 48802 53454
rect 55246 53506 55298 53518
rect 55246 53442 55298 53454
rect 55918 53506 55970 53518
rect 56242 53454 56254 53506
rect 56306 53454 56318 53506
rect 55918 53442 55970 53454
rect 1344 53338 58576 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 58576 53338
rect 1344 53252 58576 53286
rect 26238 53170 26290 53182
rect 26238 53106 26290 53118
rect 28142 53170 28194 53182
rect 28142 53106 28194 53118
rect 31614 53170 31666 53182
rect 46722 53118 46734 53170
rect 46786 53118 46798 53170
rect 50642 53118 50654 53170
rect 50706 53118 50718 53170
rect 31614 53106 31666 53118
rect 26350 53058 26402 53070
rect 26350 52994 26402 53006
rect 28030 53058 28082 53070
rect 28030 52994 28082 53006
rect 31726 53058 31778 53070
rect 49982 53058 50034 53070
rect 35186 53006 35198 53058
rect 35250 53006 35262 53058
rect 31726 52994 31778 53006
rect 49982 52994 50034 53006
rect 54910 53058 54962 53070
rect 54910 52994 54962 53006
rect 55022 53058 55074 53070
rect 55022 52994 55074 53006
rect 19070 52946 19122 52958
rect 41134 52946 41186 52958
rect 24658 52894 24670 52946
rect 24722 52894 24734 52946
rect 28354 52894 28366 52946
rect 28418 52894 28430 52946
rect 40002 52894 40014 52946
rect 40066 52894 40078 52946
rect 40898 52894 40910 52946
rect 40962 52894 40974 52946
rect 19070 52882 19122 52894
rect 41134 52882 41186 52894
rect 41358 52946 41410 52958
rect 50094 52946 50146 52958
rect 46946 52894 46958 52946
rect 47010 52894 47022 52946
rect 41358 52882 41410 52894
rect 50094 52882 50146 52894
rect 50206 52946 50258 52958
rect 50206 52882 50258 52894
rect 54798 52946 54850 52958
rect 56814 52946 56866 52958
rect 55458 52894 55470 52946
rect 55522 52894 55534 52946
rect 56578 52894 56590 52946
rect 56642 52894 56654 52946
rect 54798 52882 54850 52894
rect 56814 52882 56866 52894
rect 22642 52782 22654 52834
rect 22706 52782 22718 52834
rect 31502 52722 31554 52734
rect 31502 52658 31554 52670
rect 41470 52722 41522 52734
rect 41470 52658 41522 52670
rect 57038 52722 57090 52734
rect 57038 52658 57090 52670
rect 57150 52722 57202 52734
rect 57150 52658 57202 52670
rect 1344 52554 58576 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 58576 52554
rect 1344 52468 58576 52502
rect 31390 52386 31442 52398
rect 31390 52322 31442 52334
rect 31614 52386 31666 52398
rect 31614 52322 31666 52334
rect 35870 52386 35922 52398
rect 35870 52322 35922 52334
rect 37326 52386 37378 52398
rect 37326 52322 37378 52334
rect 43710 52386 43762 52398
rect 43710 52322 43762 52334
rect 45054 52386 45106 52398
rect 45054 52322 45106 52334
rect 45278 52386 45330 52398
rect 45278 52322 45330 52334
rect 45950 52386 46002 52398
rect 46274 52334 46286 52386
rect 46338 52334 46350 52386
rect 45950 52322 46002 52334
rect 35534 52274 35586 52286
rect 49646 52274 49698 52286
rect 18050 52222 18062 52274
rect 18114 52222 18126 52274
rect 20066 52222 20078 52274
rect 20130 52222 20142 52274
rect 26450 52222 26462 52274
rect 26514 52222 26526 52274
rect 28578 52222 28590 52274
rect 28642 52222 28654 52274
rect 38770 52222 38782 52274
rect 38834 52222 38846 52274
rect 40898 52222 40910 52274
rect 40962 52222 40974 52274
rect 44034 52222 44046 52274
rect 44098 52222 44110 52274
rect 55234 52222 55246 52274
rect 55298 52222 55310 52274
rect 57362 52222 57374 52274
rect 57426 52222 57438 52274
rect 35534 52210 35586 52222
rect 49646 52210 49698 52222
rect 22766 52162 22818 52174
rect 15250 52110 15262 52162
rect 15314 52110 15326 52162
rect 22766 52098 22818 52110
rect 22990 52162 23042 52174
rect 22990 52098 23042 52110
rect 23998 52162 24050 52174
rect 23998 52098 24050 52110
rect 24558 52162 24610 52174
rect 36094 52162 36146 52174
rect 41582 52162 41634 52174
rect 25666 52110 25678 52162
rect 25730 52110 25742 52162
rect 31826 52110 31838 52162
rect 31890 52110 31902 52162
rect 36306 52110 36318 52162
rect 36370 52110 36382 52162
rect 37314 52110 37326 52162
rect 37378 52110 37390 52162
rect 37986 52110 37998 52162
rect 38050 52110 38062 52162
rect 24558 52098 24610 52110
rect 36094 52098 36146 52110
rect 41582 52098 41634 52110
rect 42254 52162 42306 52174
rect 45726 52162 45778 52174
rect 42690 52110 42702 52162
rect 42754 52110 42766 52162
rect 44818 52110 44830 52162
rect 44882 52110 44894 52162
rect 42254 52098 42306 52110
rect 45726 52098 45778 52110
rect 48078 52162 48130 52174
rect 48078 52098 48130 52110
rect 48414 52162 48466 52174
rect 48414 52098 48466 52110
rect 48526 52162 48578 52174
rect 48526 52098 48578 52110
rect 48862 52162 48914 52174
rect 48862 52098 48914 52110
rect 49198 52162 49250 52174
rect 49198 52098 49250 52110
rect 49534 52162 49586 52174
rect 50206 52162 50258 52174
rect 49858 52110 49870 52162
rect 49922 52110 49934 52162
rect 58034 52110 58046 52162
rect 58098 52110 58110 52162
rect 49534 52098 49586 52110
rect 50206 52098 50258 52110
rect 19742 52050 19794 52062
rect 15922 51998 15934 52050
rect 15986 51998 15998 52050
rect 19742 51986 19794 51998
rect 19966 52050 20018 52062
rect 19966 51986 20018 51998
rect 35758 52050 35810 52062
rect 35758 51986 35810 51998
rect 36990 52050 37042 52062
rect 45390 52050 45442 52062
rect 42466 51998 42478 52050
rect 42530 51998 42542 52050
rect 36990 51986 37042 51998
rect 45390 51986 45442 51998
rect 48190 52050 48242 52062
rect 48190 51986 48242 51998
rect 50318 52050 50370 52062
rect 50318 51986 50370 51998
rect 51214 52050 51266 52062
rect 51214 51986 51266 51998
rect 23662 51938 23714 51950
rect 23314 51886 23326 51938
rect 23378 51886 23390 51938
rect 23662 51874 23714 51886
rect 31726 51938 31778 51950
rect 31726 51874 31778 51886
rect 32398 51938 32450 51950
rect 43934 51938 43986 51950
rect 41234 51886 41246 51938
rect 41298 51886 41310 51938
rect 32398 51874 32450 51886
rect 43934 51874 43986 51886
rect 48862 51938 48914 51950
rect 48862 51874 48914 51886
rect 51102 51938 51154 51950
rect 51102 51874 51154 51886
rect 1344 51770 58576 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 58576 51770
rect 1344 51684 58576 51718
rect 31950 51602 32002 51614
rect 19394 51550 19406 51602
rect 19458 51550 19470 51602
rect 26450 51550 26462 51602
rect 26514 51550 26526 51602
rect 31266 51550 31278 51602
rect 31330 51550 31342 51602
rect 46834 51550 46846 51602
rect 46898 51550 46910 51602
rect 31950 51538 32002 51550
rect 20302 51490 20354 51502
rect 20302 51426 20354 51438
rect 23662 51490 23714 51502
rect 30830 51490 30882 51502
rect 42478 51490 42530 51502
rect 28018 51438 28030 51490
rect 28082 51438 28094 51490
rect 34962 51438 34974 51490
rect 35026 51438 35038 51490
rect 37762 51438 37774 51490
rect 37826 51438 37838 51490
rect 45378 51438 45390 51490
rect 45442 51438 45454 51490
rect 49634 51438 49646 51490
rect 49698 51438 49710 51490
rect 51202 51438 51214 51490
rect 51266 51438 51278 51490
rect 23662 51426 23714 51438
rect 30830 51426 30882 51438
rect 42478 51426 42530 51438
rect 19966 51378 20018 51390
rect 21086 51378 21138 51390
rect 20626 51326 20638 51378
rect 20690 51326 20702 51378
rect 19966 51314 20018 51326
rect 21086 51314 21138 51326
rect 22990 51378 23042 51390
rect 22990 51314 23042 51326
rect 23998 51378 24050 51390
rect 23998 51314 24050 51326
rect 26126 51378 26178 51390
rect 26126 51314 26178 51326
rect 28366 51378 28418 51390
rect 30718 51378 30770 51390
rect 30482 51326 30494 51378
rect 30546 51326 30558 51378
rect 28366 51314 28418 51326
rect 30718 51314 30770 51326
rect 31614 51378 31666 51390
rect 31614 51314 31666 51326
rect 31838 51378 31890 51390
rect 31838 51314 31890 51326
rect 32286 51378 32338 51390
rect 38222 51378 38274 51390
rect 46510 51378 46562 51390
rect 34178 51326 34190 51378
rect 34242 51326 34254 51378
rect 37538 51326 37550 51378
rect 37602 51326 37614 51378
rect 46050 51326 46062 51378
rect 46114 51326 46126 51378
rect 32286 51314 32338 51326
rect 38222 51314 38274 51326
rect 46510 51314 46562 51326
rect 48862 51378 48914 51390
rect 48862 51314 48914 51326
rect 48974 51378 49026 51390
rect 48974 51314 49026 51326
rect 49198 51378 49250 51390
rect 55358 51378 55410 51390
rect 50194 51326 50206 51378
rect 50258 51326 50270 51378
rect 50642 51326 50654 51378
rect 50706 51326 50718 51378
rect 54562 51326 54574 51378
rect 54626 51326 54638 51378
rect 55682 51326 55694 51378
rect 55746 51326 55758 51378
rect 49198 51314 49250 51326
rect 55358 51314 55410 51326
rect 18846 51266 18898 51278
rect 18846 51202 18898 51214
rect 20190 51266 20242 51278
rect 20190 51202 20242 51214
rect 22766 51266 22818 51278
rect 22766 51202 22818 51214
rect 23326 51266 23378 51278
rect 23326 51202 23378 51214
rect 25790 51266 25842 51278
rect 25790 51202 25842 51214
rect 33182 51266 33234 51278
rect 55918 51266 55970 51278
rect 37090 51214 37102 51266
rect 37154 51214 37166 51266
rect 43250 51214 43262 51266
rect 43314 51214 43326 51266
rect 50978 51214 50990 51266
rect 51042 51214 51054 51266
rect 51650 51214 51662 51266
rect 51714 51214 51726 51266
rect 53778 51214 53790 51266
rect 53842 51214 53854 51266
rect 33182 51202 33234 51214
rect 55918 51202 55970 51214
rect 19070 51154 19122 51166
rect 19070 51090 19122 51102
rect 19854 51154 19906 51166
rect 19854 51090 19906 51102
rect 20862 51154 20914 51166
rect 20862 51090 20914 51102
rect 21198 51154 21250 51166
rect 21198 51090 21250 51102
rect 42590 51154 42642 51166
rect 42590 51090 42642 51102
rect 49310 51154 49362 51166
rect 49310 51090 49362 51102
rect 56030 51154 56082 51166
rect 56030 51090 56082 51102
rect 1344 50986 58576 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 58576 50986
rect 1344 50900 58576 50934
rect 19966 50818 20018 50830
rect 19966 50754 20018 50766
rect 49534 50818 49586 50830
rect 49534 50754 49586 50766
rect 49646 50818 49698 50830
rect 49646 50754 49698 50766
rect 50094 50818 50146 50830
rect 50094 50754 50146 50766
rect 50206 50818 50258 50830
rect 50206 50754 50258 50766
rect 50654 50818 50706 50830
rect 50654 50754 50706 50766
rect 21310 50706 21362 50718
rect 29486 50706 29538 50718
rect 35982 50706 36034 50718
rect 23426 50654 23438 50706
rect 23490 50654 23502 50706
rect 25554 50654 25566 50706
rect 25618 50654 25630 50706
rect 30370 50654 30382 50706
rect 30434 50654 30446 50706
rect 31154 50654 31166 50706
rect 31218 50654 31230 50706
rect 33282 50654 33294 50706
rect 33346 50654 33358 50706
rect 21310 50642 21362 50654
rect 29486 50642 29538 50654
rect 35982 50642 36034 50654
rect 46174 50706 46226 50718
rect 46174 50642 46226 50654
rect 19742 50594 19794 50606
rect 35870 50594 35922 50606
rect 19170 50542 19182 50594
rect 19234 50542 19246 50594
rect 22642 50542 22654 50594
rect 22706 50542 22718 50594
rect 26898 50542 26910 50594
rect 26962 50542 26974 50594
rect 29922 50542 29934 50594
rect 29986 50542 29998 50594
rect 34066 50542 34078 50594
rect 34130 50542 34142 50594
rect 19742 50530 19794 50542
rect 35870 50530 35922 50542
rect 36094 50594 36146 50606
rect 36094 50530 36146 50542
rect 36430 50594 36482 50606
rect 36430 50530 36482 50542
rect 37102 50594 37154 50606
rect 37102 50530 37154 50542
rect 45502 50594 45554 50606
rect 45502 50530 45554 50542
rect 49870 50594 49922 50606
rect 51438 50594 51490 50606
rect 51202 50542 51214 50594
rect 51266 50542 51278 50594
rect 51538 50542 51550 50594
rect 51602 50542 51614 50594
rect 52882 50542 52894 50594
rect 52946 50542 52958 50594
rect 49870 50530 49922 50542
rect 51438 50530 51490 50542
rect 21422 50482 21474 50494
rect 14354 50430 14366 50482
rect 14418 50430 14430 50482
rect 20290 50430 20302 50482
rect 20354 50430 20366 50482
rect 21422 50418 21474 50430
rect 27134 50482 27186 50494
rect 27134 50418 27186 50430
rect 28254 50482 28306 50494
rect 50542 50482 50594 50494
rect 28578 50430 28590 50482
rect 28642 50430 28654 50482
rect 45154 50430 45166 50482
rect 45218 50430 45230 50482
rect 28254 50418 28306 50430
rect 50542 50418 50594 50430
rect 50990 50482 51042 50494
rect 57922 50430 57934 50482
rect 57986 50430 57998 50482
rect 50990 50418 51042 50430
rect 21534 50370 21586 50382
rect 21534 50306 21586 50318
rect 51774 50370 51826 50382
rect 51774 50306 51826 50318
rect 1344 50202 58576 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 58576 50202
rect 1344 50116 58576 50150
rect 25902 50034 25954 50046
rect 25902 49970 25954 49982
rect 26798 50034 26850 50046
rect 26798 49970 26850 49982
rect 30158 50034 30210 50046
rect 30158 49970 30210 49982
rect 30382 50034 30434 50046
rect 30382 49970 30434 49982
rect 37102 50034 37154 50046
rect 37102 49970 37154 49982
rect 41806 50034 41858 50046
rect 41806 49970 41858 49982
rect 50542 50034 50594 50046
rect 50542 49970 50594 49982
rect 50990 50034 51042 50046
rect 50990 49970 51042 49982
rect 52558 50034 52610 50046
rect 52558 49970 52610 49982
rect 57374 50034 57426 50046
rect 57374 49970 57426 49982
rect 58158 50034 58210 50046
rect 58158 49970 58210 49982
rect 37662 49922 37714 49934
rect 30930 49870 30942 49922
rect 30994 49870 31006 49922
rect 31266 49870 31278 49922
rect 31330 49870 31342 49922
rect 37662 49858 37714 49870
rect 41358 49922 41410 49934
rect 41358 49858 41410 49870
rect 50206 49922 50258 49934
rect 50206 49858 50258 49870
rect 50318 49922 50370 49934
rect 50318 49858 50370 49870
rect 56030 49922 56082 49934
rect 56030 49858 56082 49870
rect 56590 49922 56642 49934
rect 56590 49858 56642 49870
rect 56702 49922 56754 49934
rect 56702 49858 56754 49870
rect 25678 49810 25730 49822
rect 14242 49758 14254 49810
rect 14306 49758 14318 49810
rect 25678 49746 25730 49758
rect 26686 49810 26738 49822
rect 31390 49810 31442 49822
rect 30706 49758 30718 49810
rect 30770 49758 30782 49810
rect 26686 49746 26738 49758
rect 31390 49746 31442 49758
rect 36542 49810 36594 49822
rect 36542 49746 36594 49758
rect 40910 49810 40962 49822
rect 40910 49746 40962 49758
rect 41134 49810 41186 49822
rect 56926 49810 56978 49822
rect 48962 49758 48974 49810
rect 49026 49758 49038 49810
rect 49186 49758 49198 49810
rect 49250 49758 49262 49810
rect 55570 49758 55582 49810
rect 55634 49758 55646 49810
rect 55794 49758 55806 49810
rect 55858 49758 55870 49810
rect 41134 49746 41186 49758
rect 56926 49746 56978 49758
rect 57598 49810 57650 49822
rect 57598 49746 57650 49758
rect 19630 49698 19682 49710
rect 11330 49646 11342 49698
rect 11394 49646 11406 49698
rect 13458 49646 13470 49698
rect 13522 49646 13534 49698
rect 19630 49634 19682 49646
rect 25790 49698 25842 49710
rect 25790 49634 25842 49646
rect 26126 49698 26178 49710
rect 26126 49634 26178 49646
rect 31950 49698 32002 49710
rect 31950 49634 32002 49646
rect 41022 49698 41074 49710
rect 41022 49634 41074 49646
rect 41918 49698 41970 49710
rect 41918 49634 41970 49646
rect 42366 49698 42418 49710
rect 42366 49634 42418 49646
rect 48750 49698 48802 49710
rect 48750 49634 48802 49646
rect 26350 49586 26402 49598
rect 26350 49522 26402 49534
rect 26798 49586 26850 49598
rect 26798 49522 26850 49534
rect 36654 49586 36706 49598
rect 36654 49522 36706 49534
rect 42254 49586 42306 49598
rect 42254 49522 42306 49534
rect 1344 49418 58576 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 58576 49418
rect 1344 49332 58576 49366
rect 39118 49250 39170 49262
rect 39118 49186 39170 49198
rect 48526 49250 48578 49262
rect 48526 49186 48578 49198
rect 35646 49138 35698 49150
rect 39678 49138 39730 49150
rect 44158 49138 44210 49150
rect 16146 49086 16158 49138
rect 16210 49086 16222 49138
rect 18386 49086 18398 49138
rect 18450 49086 18462 49138
rect 19954 49086 19966 49138
rect 20018 49086 20030 49138
rect 38546 49086 38558 49138
rect 38610 49086 38622 49138
rect 40898 49086 40910 49138
rect 40962 49086 40974 49138
rect 43138 49086 43150 49138
rect 43202 49086 43214 49138
rect 48178 49086 48190 49138
rect 48242 49086 48254 49138
rect 52994 49086 53006 49138
rect 53058 49086 53070 49138
rect 56018 49086 56030 49138
rect 56082 49086 56094 49138
rect 58146 49086 58158 49138
rect 58210 49086 58222 49138
rect 35646 49074 35698 49086
rect 39678 49074 39730 49086
rect 44158 49074 44210 49086
rect 21982 49026 22034 49038
rect 29934 49026 29986 49038
rect 36990 49026 37042 49038
rect 15362 48974 15374 49026
rect 15426 48974 15438 49026
rect 26338 48974 26350 49026
rect 26402 48974 26414 49026
rect 27682 48974 27694 49026
rect 27746 48974 27758 49026
rect 35410 48974 35422 49026
rect 35474 48974 35486 49026
rect 21982 48962 22034 48974
rect 29934 48962 29986 48974
rect 36990 48962 37042 48974
rect 37214 49026 37266 49038
rect 37214 48962 37266 48974
rect 37438 49026 37490 49038
rect 37438 48962 37490 48974
rect 37550 49026 37602 49038
rect 39342 49026 39394 49038
rect 38098 48974 38110 49026
rect 38162 48974 38174 49026
rect 37550 48962 37602 48974
rect 39342 48962 39394 48974
rect 39566 49026 39618 49038
rect 40798 49026 40850 49038
rect 41358 49026 41410 49038
rect 40338 48974 40350 49026
rect 40402 48974 40414 49026
rect 41010 48974 41022 49026
rect 41074 48974 41086 49026
rect 39566 48962 39618 48974
rect 40798 48962 40850 48974
rect 41358 48962 41410 48974
rect 42142 49026 42194 49038
rect 42142 48962 42194 48974
rect 42478 49026 42530 49038
rect 45390 49026 45442 49038
rect 43026 48974 43038 49026
rect 43090 48974 43102 49026
rect 55234 48974 55246 49026
rect 55298 48974 55310 49026
rect 42478 48962 42530 48974
rect 45390 48962 45442 48974
rect 7982 48914 8034 48926
rect 7982 48850 8034 48862
rect 20302 48914 20354 48926
rect 20302 48850 20354 48862
rect 21646 48914 21698 48926
rect 21646 48850 21698 48862
rect 22094 48914 22146 48926
rect 22094 48850 22146 48862
rect 26574 48914 26626 48926
rect 29822 48914 29874 48926
rect 27794 48862 27806 48914
rect 27858 48862 27870 48914
rect 26574 48850 26626 48862
rect 29822 48850 29874 48862
rect 34862 48914 34914 48926
rect 34862 48850 34914 48862
rect 38558 48914 38610 48926
rect 38558 48850 38610 48862
rect 42590 48914 42642 48926
rect 42590 48850 42642 48862
rect 43374 48914 43426 48926
rect 43374 48850 43426 48862
rect 45166 48914 45218 48926
rect 45166 48850 45218 48862
rect 48302 48914 48354 48926
rect 48302 48850 48354 48862
rect 8094 48802 8146 48814
rect 8094 48738 8146 48750
rect 8318 48802 8370 48814
rect 8318 48738 8370 48750
rect 20078 48802 20130 48814
rect 20078 48738 20130 48750
rect 21534 48802 21586 48814
rect 21534 48738 21586 48750
rect 22318 48802 22370 48814
rect 33630 48802 33682 48814
rect 27234 48750 27246 48802
rect 27298 48750 27310 48802
rect 22318 48738 22370 48750
rect 33630 48738 33682 48750
rect 36206 48802 36258 48814
rect 36206 48738 36258 48750
rect 37662 48802 37714 48814
rect 37662 48738 37714 48750
rect 38334 48802 38386 48814
rect 38334 48738 38386 48750
rect 38670 48802 38722 48814
rect 38670 48738 38722 48750
rect 39790 48802 39842 48814
rect 39790 48738 39842 48750
rect 40574 48802 40626 48814
rect 40574 48738 40626 48750
rect 41470 48802 41522 48814
rect 41470 48738 41522 48750
rect 41694 48802 41746 48814
rect 41694 48738 41746 48750
rect 42254 48802 42306 48814
rect 42254 48738 42306 48750
rect 42366 48802 42418 48814
rect 42366 48738 42418 48750
rect 44270 48802 44322 48814
rect 53454 48802 53506 48814
rect 45714 48750 45726 48802
rect 45778 48750 45790 48802
rect 44270 48738 44322 48750
rect 53454 48738 53506 48750
rect 1344 48634 58576 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 58576 48634
rect 1344 48548 58576 48582
rect 24558 48466 24610 48478
rect 24558 48402 24610 48414
rect 25342 48466 25394 48478
rect 25342 48402 25394 48414
rect 26686 48466 26738 48478
rect 26686 48402 26738 48414
rect 34638 48466 34690 48478
rect 34638 48402 34690 48414
rect 37326 48466 37378 48478
rect 37326 48402 37378 48414
rect 40126 48466 40178 48478
rect 40126 48402 40178 48414
rect 43598 48466 43650 48478
rect 43598 48402 43650 48414
rect 43934 48466 43986 48478
rect 43934 48402 43986 48414
rect 44158 48466 44210 48478
rect 44158 48402 44210 48414
rect 46062 48466 46114 48478
rect 46062 48402 46114 48414
rect 9550 48354 9602 48366
rect 9550 48290 9602 48302
rect 9774 48354 9826 48366
rect 32062 48354 32114 48366
rect 18610 48302 18622 48354
rect 18674 48302 18686 48354
rect 9774 48290 9826 48302
rect 32062 48290 32114 48302
rect 36206 48354 36258 48366
rect 36206 48290 36258 48302
rect 37662 48354 37714 48366
rect 45054 48354 45106 48366
rect 42802 48302 42814 48354
rect 42866 48302 42878 48354
rect 37662 48290 37714 48302
rect 45054 48290 45106 48302
rect 45614 48354 45666 48366
rect 45614 48290 45666 48302
rect 46174 48354 46226 48366
rect 46174 48290 46226 48302
rect 48078 48354 48130 48366
rect 56590 48354 56642 48366
rect 51538 48302 51550 48354
rect 51602 48302 51614 48354
rect 48078 48290 48130 48302
rect 56590 48290 56642 48302
rect 57150 48354 57202 48366
rect 57150 48290 57202 48302
rect 26574 48242 26626 48254
rect 31838 48242 31890 48254
rect 6178 48190 6190 48242
rect 6242 48190 6254 48242
rect 14018 48190 14030 48242
rect 14082 48190 14094 48242
rect 17826 48190 17838 48242
rect 17890 48190 17902 48242
rect 21186 48190 21198 48242
rect 21250 48190 21262 48242
rect 27234 48190 27246 48242
rect 27298 48190 27310 48242
rect 27458 48190 27470 48242
rect 27522 48190 27534 48242
rect 29026 48190 29038 48242
rect 29090 48190 29102 48242
rect 30370 48190 30382 48242
rect 30434 48190 30446 48242
rect 26574 48178 26626 48190
rect 31838 48178 31890 48190
rect 32174 48242 32226 48254
rect 34750 48242 34802 48254
rect 39678 48242 39730 48254
rect 34402 48190 34414 48242
rect 34466 48190 34478 48242
rect 35074 48190 35086 48242
rect 35138 48190 35150 48242
rect 37090 48190 37102 48242
rect 37154 48190 37166 48242
rect 32174 48178 32226 48190
rect 34750 48178 34802 48190
rect 39678 48178 39730 48190
rect 39902 48242 39954 48254
rect 39902 48178 39954 48190
rect 40350 48242 40402 48254
rect 40350 48178 40402 48190
rect 41470 48242 41522 48254
rect 41470 48178 41522 48190
rect 41694 48242 41746 48254
rect 41694 48178 41746 48190
rect 42478 48242 42530 48254
rect 42478 48178 42530 48190
rect 43262 48242 43314 48254
rect 43262 48178 43314 48190
rect 43486 48242 43538 48254
rect 43486 48178 43538 48190
rect 43822 48242 43874 48254
rect 43822 48178 43874 48190
rect 44494 48242 44546 48254
rect 44494 48178 44546 48190
rect 44942 48242 44994 48254
rect 44942 48178 44994 48190
rect 45838 48242 45890 48254
rect 45838 48178 45890 48190
rect 46958 48242 47010 48254
rect 46958 48178 47010 48190
rect 47854 48242 47906 48254
rect 56814 48242 56866 48254
rect 50306 48190 50318 48242
rect 50370 48190 50382 48242
rect 50866 48190 50878 48242
rect 50930 48190 50942 48242
rect 47854 48178 47906 48190
rect 56814 48178 56866 48190
rect 9662 48130 9714 48142
rect 24446 48130 24498 48142
rect 6850 48078 6862 48130
rect 6914 48078 6926 48130
rect 8978 48078 8990 48130
rect 9042 48078 9054 48130
rect 14690 48078 14702 48130
rect 14754 48078 14766 48130
rect 16818 48078 16830 48130
rect 16882 48078 16894 48130
rect 20738 48078 20750 48130
rect 20802 48078 20814 48130
rect 21970 48078 21982 48130
rect 22034 48078 22046 48130
rect 24098 48078 24110 48130
rect 24162 48078 24174 48130
rect 9662 48066 9714 48078
rect 24446 48066 24498 48078
rect 25230 48130 25282 48142
rect 33630 48130 33682 48142
rect 30818 48078 30830 48130
rect 30882 48078 30894 48130
rect 33282 48078 33294 48130
rect 33346 48078 33358 48130
rect 25230 48066 25282 48078
rect 33630 48066 33682 48078
rect 39342 48130 39394 48142
rect 39342 48066 39394 48078
rect 44270 48130 44322 48142
rect 44270 48066 44322 48078
rect 45278 48130 45330 48142
rect 45278 48066 45330 48078
rect 45950 48130 46002 48142
rect 45950 48066 46002 48078
rect 47182 48130 47234 48142
rect 47182 48066 47234 48078
rect 47518 48130 47570 48142
rect 57038 48130 57090 48142
rect 49970 48078 49982 48130
rect 50034 48078 50046 48130
rect 53666 48078 53678 48130
rect 53730 48078 53742 48130
rect 47518 48066 47570 48078
rect 57038 48066 57090 48078
rect 26686 48018 26738 48030
rect 39230 48018 39282 48030
rect 30930 47966 30942 48018
rect 30994 47966 31006 48018
rect 26686 47954 26738 47966
rect 39230 47954 39282 47966
rect 40238 48018 40290 48030
rect 40238 47954 40290 47966
rect 40798 48018 40850 48030
rect 40798 47954 40850 47966
rect 41246 48018 41298 48030
rect 41246 47954 41298 47966
rect 43038 48018 43090 48030
rect 46610 47966 46622 48018
rect 46674 47966 46686 48018
rect 43038 47954 43090 47966
rect 1344 47850 58576 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 58576 47850
rect 1344 47764 58576 47798
rect 38334 47682 38386 47694
rect 17602 47630 17614 47682
rect 17666 47630 17678 47682
rect 27458 47630 27470 47682
rect 27522 47630 27534 47682
rect 38334 47618 38386 47630
rect 43486 47682 43538 47694
rect 43486 47618 43538 47630
rect 45054 47682 45106 47694
rect 45054 47618 45106 47630
rect 15934 47570 15986 47582
rect 20526 47570 20578 47582
rect 6178 47518 6190 47570
rect 6242 47518 6254 47570
rect 20066 47518 20078 47570
rect 20130 47518 20142 47570
rect 15934 47506 15986 47518
rect 20526 47506 20578 47518
rect 21870 47570 21922 47582
rect 28590 47570 28642 47582
rect 38670 47570 38722 47582
rect 26674 47518 26686 47570
rect 26738 47518 26750 47570
rect 27794 47518 27806 47570
rect 27858 47518 27870 47570
rect 31826 47518 31838 47570
rect 31890 47518 31902 47570
rect 33954 47518 33966 47570
rect 34018 47518 34030 47570
rect 34962 47518 34974 47570
rect 35026 47518 35038 47570
rect 21870 47506 21922 47518
rect 28590 47506 28642 47518
rect 38670 47506 38722 47518
rect 40686 47570 40738 47582
rect 51102 47570 51154 47582
rect 47058 47518 47070 47570
rect 47122 47518 47134 47570
rect 55234 47518 55246 47570
rect 55298 47518 55310 47570
rect 57362 47518 57374 47570
rect 57426 47518 57438 47570
rect 40686 47506 40738 47518
rect 51102 47506 51154 47518
rect 16046 47458 16098 47470
rect 10434 47406 10446 47458
rect 10498 47406 10510 47458
rect 16046 47394 16098 47406
rect 16494 47458 16546 47470
rect 16494 47394 16546 47406
rect 16718 47458 16770 47470
rect 16718 47394 16770 47406
rect 17054 47458 17106 47470
rect 17054 47394 17106 47406
rect 17950 47458 18002 47470
rect 17950 47394 18002 47406
rect 18174 47458 18226 47470
rect 21422 47458 21474 47470
rect 19954 47406 19966 47458
rect 20018 47406 20030 47458
rect 18174 47394 18226 47406
rect 21422 47394 21474 47406
rect 21758 47458 21810 47470
rect 21758 47394 21810 47406
rect 22094 47458 22146 47470
rect 24222 47458 24274 47470
rect 37214 47458 37266 47470
rect 38558 47458 38610 47470
rect 22306 47406 22318 47458
rect 22370 47406 22382 47458
rect 23314 47406 23326 47458
rect 23378 47406 23390 47458
rect 26898 47406 26910 47458
rect 26962 47406 26974 47458
rect 27682 47406 27694 47458
rect 27746 47406 27758 47458
rect 29698 47406 29710 47458
rect 29762 47406 29774 47458
rect 30258 47406 30270 47458
rect 30322 47406 30334 47458
rect 31154 47406 31166 47458
rect 31218 47406 31230 47458
rect 34514 47406 34526 47458
rect 34578 47406 34590 47458
rect 35522 47406 35534 47458
rect 35586 47406 35598 47458
rect 37874 47406 37886 47458
rect 37938 47406 37950 47458
rect 22094 47394 22146 47406
rect 24222 47394 24274 47406
rect 37214 47394 37266 47406
rect 38558 47394 38610 47406
rect 38782 47458 38834 47470
rect 38782 47394 38834 47406
rect 44942 47458 44994 47470
rect 54126 47458 54178 47470
rect 50642 47406 50654 47458
rect 50706 47406 50718 47458
rect 53330 47406 53342 47458
rect 53394 47406 53406 47458
rect 53666 47406 53678 47458
rect 53730 47406 53742 47458
rect 58034 47406 58046 47458
rect 58098 47406 58110 47458
rect 44942 47394 44994 47406
rect 54126 47394 54178 47406
rect 14926 47346 14978 47358
rect 14926 47282 14978 47294
rect 15262 47346 15314 47358
rect 15262 47282 15314 47294
rect 15822 47346 15874 47358
rect 28478 47346 28530 47358
rect 30382 47346 30434 47358
rect 36318 47346 36370 47358
rect 22530 47294 22542 47346
rect 22594 47294 22606 47346
rect 29250 47294 29262 47346
rect 29314 47294 29326 47346
rect 35634 47294 35646 47346
rect 35698 47294 35710 47346
rect 15822 47282 15874 47294
rect 28478 47282 28530 47294
rect 30382 47282 30434 47294
rect 36318 47282 36370 47294
rect 37438 47346 37490 47358
rect 37438 47282 37490 47294
rect 37550 47346 37602 47358
rect 43598 47346 43650 47358
rect 38098 47294 38110 47346
rect 38162 47294 38174 47346
rect 37550 47282 37602 47294
rect 43598 47282 43650 47294
rect 53902 47346 53954 47358
rect 53902 47282 53954 47294
rect 11342 47234 11394 47246
rect 11342 47170 11394 47182
rect 16942 47234 16994 47246
rect 16942 47170 16994 47182
rect 18622 47234 18674 47246
rect 24110 47234 24162 47246
rect 36430 47234 36482 47246
rect 23426 47182 23438 47234
rect 23490 47182 23502 47234
rect 23650 47182 23662 47234
rect 23714 47182 23726 47234
rect 29698 47182 29710 47234
rect 29762 47182 29774 47234
rect 18622 47170 18674 47182
rect 24110 47170 24162 47182
rect 36430 47170 36482 47182
rect 40798 47234 40850 47246
rect 40798 47170 40850 47182
rect 52782 47234 52834 47246
rect 52782 47170 52834 47182
rect 52894 47234 52946 47246
rect 52894 47170 52946 47182
rect 53006 47234 53058 47246
rect 53006 47170 53058 47182
rect 54014 47234 54066 47246
rect 54014 47170 54066 47182
rect 54238 47234 54290 47246
rect 54238 47170 54290 47182
rect 1344 47066 58576 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 58576 47066
rect 1344 46980 58576 47014
rect 17502 46898 17554 46910
rect 17502 46834 17554 46846
rect 35534 46898 35586 46910
rect 35534 46834 35586 46846
rect 35982 46898 36034 46910
rect 35982 46834 36034 46846
rect 36766 46898 36818 46910
rect 36766 46834 36818 46846
rect 36990 46898 37042 46910
rect 36990 46834 37042 46846
rect 52446 46898 52498 46910
rect 52446 46834 52498 46846
rect 56590 46898 56642 46910
rect 56590 46834 56642 46846
rect 57150 46898 57202 46910
rect 57150 46834 57202 46846
rect 8766 46786 8818 46798
rect 8766 46722 8818 46734
rect 15038 46786 15090 46798
rect 15038 46722 15090 46734
rect 16270 46786 16322 46798
rect 33070 46786 33122 46798
rect 20178 46734 20190 46786
rect 20242 46734 20254 46786
rect 28578 46734 28590 46786
rect 28642 46734 28654 46786
rect 30930 46734 30942 46786
rect 30994 46734 31006 46786
rect 16270 46722 16322 46734
rect 33070 46722 33122 46734
rect 33182 46786 33234 46798
rect 33182 46722 33234 46734
rect 33742 46786 33794 46798
rect 33742 46722 33794 46734
rect 36542 46786 36594 46798
rect 46062 46786 46114 46798
rect 41122 46734 41134 46786
rect 41186 46734 41198 46786
rect 36542 46722 36594 46734
rect 46062 46722 46114 46734
rect 52110 46786 52162 46798
rect 52110 46722 52162 46734
rect 54126 46786 54178 46798
rect 54126 46722 54178 46734
rect 55470 46786 55522 46798
rect 55470 46722 55522 46734
rect 56702 46786 56754 46798
rect 56702 46722 56754 46734
rect 57038 46786 57090 46798
rect 57038 46722 57090 46734
rect 18734 46674 18786 46686
rect 33406 46674 33458 46686
rect 46174 46674 46226 46686
rect 6962 46622 6974 46674
rect 7026 46622 7038 46674
rect 7746 46622 7758 46674
rect 7810 46622 7822 46674
rect 10210 46622 10222 46674
rect 10274 46622 10286 46674
rect 24322 46622 24334 46674
rect 24386 46622 24398 46674
rect 25778 46622 25790 46674
rect 25842 46622 25854 46674
rect 26450 46622 26462 46674
rect 26514 46622 26526 46674
rect 26898 46622 26910 46674
rect 26962 46622 26974 46674
rect 28354 46622 28366 46674
rect 28418 46622 28430 46674
rect 29474 46622 29486 46674
rect 29538 46622 29550 46674
rect 31490 46622 31502 46674
rect 31554 46622 31566 46674
rect 37202 46622 37214 46674
rect 37266 46622 37278 46674
rect 41010 46622 41022 46674
rect 41074 46622 41086 46674
rect 41570 46622 41582 46674
rect 41634 46622 41646 46674
rect 42018 46622 42030 46674
rect 42082 46622 42094 46674
rect 18734 46610 18786 46622
rect 33406 46610 33458 46622
rect 46174 46610 46226 46622
rect 46286 46674 46338 46686
rect 46286 46610 46338 46622
rect 46622 46674 46674 46686
rect 46622 46610 46674 46622
rect 49870 46674 49922 46686
rect 49870 46610 49922 46622
rect 50094 46674 50146 46686
rect 50094 46610 50146 46622
rect 50318 46674 50370 46686
rect 55246 46674 55298 46686
rect 58158 46674 58210 46686
rect 50866 46622 50878 46674
rect 50930 46622 50942 46674
rect 54674 46622 54686 46674
rect 54738 46622 54750 46674
rect 55010 46622 55022 46674
rect 55074 46622 55086 46674
rect 55682 46622 55694 46674
rect 55746 46622 55758 46674
rect 50318 46610 50370 46622
rect 55246 46610 55298 46622
rect 58158 46610 58210 46622
rect 29262 46562 29314 46574
rect 4162 46510 4174 46562
rect 4226 46510 4238 46562
rect 6290 46510 6302 46562
rect 6354 46510 6366 46562
rect 7634 46510 7646 46562
rect 7698 46510 7710 46562
rect 8866 46510 8878 46562
rect 8930 46510 8942 46562
rect 10882 46510 10894 46562
rect 10946 46510 10958 46562
rect 13010 46510 13022 46562
rect 13074 46510 13086 46562
rect 14914 46510 14926 46562
rect 14978 46510 14990 46562
rect 26114 46510 26126 46562
rect 26178 46510 26190 46562
rect 29262 46498 29314 46510
rect 34190 46562 34242 46574
rect 42702 46562 42754 46574
rect 37090 46510 37102 46562
rect 37154 46510 37166 46562
rect 34190 46498 34242 46510
rect 42702 46498 42754 46510
rect 50206 46562 50258 46574
rect 50206 46498 50258 46510
rect 55358 46562 55410 46574
rect 57698 46510 57710 46562
rect 57762 46510 57774 46562
rect 55358 46498 55410 46510
rect 7422 46450 7474 46462
rect 7422 46386 7474 46398
rect 8542 46450 8594 46462
rect 8542 46386 8594 46398
rect 15262 46450 15314 46462
rect 15262 46386 15314 46398
rect 16158 46450 16210 46462
rect 49646 46450 49698 46462
rect 26450 46398 26462 46450
rect 26514 46398 26526 46450
rect 16158 46386 16210 46398
rect 49646 46386 49698 46398
rect 1344 46282 58576 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 58576 46282
rect 1344 46196 58576 46230
rect 11342 46114 11394 46126
rect 11342 46050 11394 46062
rect 14590 46114 14642 46126
rect 14590 46050 14642 46062
rect 29486 46114 29538 46126
rect 29486 46050 29538 46062
rect 29822 46114 29874 46126
rect 29822 46050 29874 46062
rect 37998 46114 38050 46126
rect 37998 46050 38050 46062
rect 40014 46114 40066 46126
rect 40014 46050 40066 46062
rect 7310 46002 7362 46014
rect 29374 46002 29426 46014
rect 37102 46002 37154 46014
rect 21746 45950 21758 46002
rect 21810 45950 21822 46002
rect 31154 45950 31166 46002
rect 31218 45950 31230 46002
rect 7310 45938 7362 45950
rect 29374 45938 29426 45950
rect 37102 45938 37154 45950
rect 40574 46002 40626 46014
rect 47954 45950 47966 46002
rect 48018 45950 48030 46002
rect 50082 45950 50094 46002
rect 50146 45950 50158 46002
rect 40574 45938 40626 45950
rect 7198 45890 7250 45902
rect 6738 45838 6750 45890
rect 6802 45838 6814 45890
rect 7198 45826 7250 45838
rect 8206 45890 8258 45902
rect 8206 45826 8258 45838
rect 8542 45890 8594 45902
rect 12014 45890 12066 45902
rect 11330 45838 11342 45890
rect 11394 45838 11406 45890
rect 8542 45826 8594 45838
rect 12014 45826 12066 45838
rect 12238 45890 12290 45902
rect 18622 45890 18674 45902
rect 26798 45890 26850 45902
rect 14914 45838 14926 45890
rect 14978 45838 14990 45890
rect 21634 45838 21646 45890
rect 21698 45838 21710 45890
rect 22642 45838 22654 45890
rect 22706 45838 22718 45890
rect 24098 45838 24110 45890
rect 24162 45838 24174 45890
rect 26114 45838 26126 45890
rect 26178 45838 26190 45890
rect 29138 45838 29150 45890
rect 29202 45838 29214 45890
rect 36194 45838 36206 45890
rect 36258 45838 36270 45890
rect 47170 45838 47182 45890
rect 47234 45838 47246 45890
rect 50418 45838 50430 45890
rect 50482 45838 50494 45890
rect 51314 45838 51326 45890
rect 51378 45838 51390 45890
rect 52770 45838 52782 45890
rect 52834 45838 52846 45890
rect 53442 45838 53454 45890
rect 53506 45838 53518 45890
rect 54002 45838 54014 45890
rect 54066 45838 54078 45890
rect 54450 45838 54462 45890
rect 54514 45838 54526 45890
rect 55682 45838 55694 45890
rect 55746 45838 55758 45890
rect 56242 45838 56254 45890
rect 56306 45838 56318 45890
rect 57138 45838 57150 45890
rect 57202 45838 57214 45890
rect 12238 45826 12290 45838
rect 18622 45826 18674 45838
rect 26798 45826 26850 45838
rect 11678 45778 11730 45790
rect 11678 45714 11730 45726
rect 12574 45778 12626 45790
rect 12574 45714 12626 45726
rect 14254 45778 14306 45790
rect 14254 45714 14306 45726
rect 21982 45778 22034 45790
rect 26910 45778 26962 45790
rect 23202 45726 23214 45778
rect 23266 45726 23278 45778
rect 24546 45726 24558 45778
rect 24610 45726 24622 45778
rect 25554 45726 25566 45778
rect 25618 45726 25630 45778
rect 21982 45714 22034 45726
rect 26910 45714 26962 45726
rect 29934 45778 29986 45790
rect 29934 45714 29986 45726
rect 37886 45778 37938 45790
rect 37886 45714 37938 45726
rect 39902 45778 39954 45790
rect 39902 45714 39954 45726
rect 44046 45778 44098 45790
rect 51426 45726 51438 45778
rect 51490 45726 51502 45778
rect 53890 45726 53902 45778
rect 53954 45726 53966 45778
rect 54114 45726 54126 45778
rect 54178 45726 54190 45778
rect 55570 45726 55582 45778
rect 55634 45726 55646 45778
rect 57250 45726 57262 45778
rect 57314 45726 57326 45778
rect 44046 45714 44098 45726
rect 8430 45666 8482 45678
rect 8430 45602 8482 45614
rect 12462 45666 12514 45678
rect 12462 45602 12514 45614
rect 12686 45666 12738 45678
rect 14702 45666 14754 45678
rect 20414 45666 20466 45678
rect 13906 45614 13918 45666
rect 13970 45614 13982 45666
rect 18274 45614 18286 45666
rect 18338 45614 18350 45666
rect 12686 45602 12738 45614
rect 14702 45602 14754 45614
rect 20414 45602 20466 45614
rect 27134 45666 27186 45678
rect 27134 45602 27186 45614
rect 44158 45666 44210 45678
rect 58158 45666 58210 45678
rect 50530 45614 50542 45666
rect 50594 45614 50606 45666
rect 51314 45614 51326 45666
rect 51378 45614 51390 45666
rect 54562 45614 54574 45666
rect 54626 45614 54638 45666
rect 54786 45614 54798 45666
rect 54850 45614 54862 45666
rect 56354 45614 56366 45666
rect 56418 45614 56430 45666
rect 56578 45614 56590 45666
rect 56642 45614 56654 45666
rect 44158 45602 44210 45614
rect 58158 45602 58210 45614
rect 1344 45498 58576 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 58576 45498
rect 1344 45412 58576 45446
rect 13246 45330 13298 45342
rect 13246 45266 13298 45278
rect 14366 45330 14418 45342
rect 19506 45278 19518 45330
rect 19570 45278 19582 45330
rect 57474 45278 57486 45330
rect 57538 45278 57550 45330
rect 14366 45266 14418 45278
rect 14590 45218 14642 45230
rect 20638 45218 20690 45230
rect 9650 45166 9662 45218
rect 9714 45166 9726 45218
rect 16034 45166 16046 45218
rect 16098 45166 16110 45218
rect 14590 45154 14642 45166
rect 20638 45154 20690 45166
rect 21198 45218 21250 45230
rect 21198 45154 21250 45166
rect 31502 45218 31554 45230
rect 56814 45218 56866 45230
rect 40114 45166 40126 45218
rect 40178 45166 40190 45218
rect 44930 45166 44942 45218
rect 44994 45166 45006 45218
rect 52770 45166 52782 45218
rect 52834 45166 52846 45218
rect 57586 45166 57598 45218
rect 57650 45166 57662 45218
rect 31502 45154 31554 45166
rect 56814 45154 56866 45166
rect 9550 45106 9602 45118
rect 9550 45042 9602 45054
rect 9886 45106 9938 45118
rect 11230 45106 11282 45118
rect 10210 45054 10222 45106
rect 10274 45054 10286 45106
rect 9886 45042 9938 45054
rect 11230 45042 11282 45054
rect 13022 45106 13074 45118
rect 13022 45042 13074 45054
rect 13358 45106 13410 45118
rect 13358 45042 13410 45054
rect 14702 45106 14754 45118
rect 14702 45042 14754 45054
rect 14814 45106 14866 45118
rect 15822 45106 15874 45118
rect 15362 45054 15374 45106
rect 15426 45054 15438 45106
rect 16594 45054 16606 45106
rect 16658 45054 16670 45106
rect 22866 45054 22878 45106
rect 22930 45054 22942 45106
rect 23538 45054 23550 45106
rect 23602 45054 23614 45106
rect 23762 45054 23774 45106
rect 23826 45054 23838 45106
rect 25330 45054 25342 45106
rect 25394 45054 25406 45106
rect 26338 45054 26350 45106
rect 26402 45054 26414 45106
rect 27122 45054 27134 45106
rect 27186 45054 27198 45106
rect 28578 45054 28590 45106
rect 28642 45054 28654 45106
rect 29586 45054 29598 45106
rect 29650 45054 29662 45106
rect 32162 45054 32174 45106
rect 32226 45054 32238 45106
rect 36194 45054 36206 45106
rect 36258 45054 36270 45106
rect 40898 45054 40910 45106
rect 40962 45054 40974 45106
rect 44258 45054 44270 45106
rect 44322 45054 44334 45106
rect 50082 45054 50094 45106
rect 50146 45054 50158 45106
rect 51090 45054 51102 45106
rect 51154 45054 51166 45106
rect 56690 45054 56702 45106
rect 56754 45054 56766 45106
rect 57474 45054 57486 45106
rect 57538 45054 57550 45106
rect 14814 45042 14866 45054
rect 15822 45042 15874 45054
rect 10558 44994 10610 45006
rect 20078 44994 20130 45006
rect 30158 44994 30210 45006
rect 33070 44994 33122 45006
rect 16482 44942 16494 44994
rect 16546 44942 16558 44994
rect 20738 44942 20750 44994
rect 20802 44942 20814 44994
rect 22978 44942 22990 44994
rect 23042 44942 23054 44994
rect 23426 44942 23438 44994
rect 23490 44942 23502 44994
rect 32386 44942 32398 44994
rect 32450 44942 32462 44994
rect 10558 44930 10610 44942
rect 20078 44930 20130 44942
rect 30158 44930 30210 44942
rect 33070 44930 33122 44942
rect 33742 44994 33794 45006
rect 49086 44994 49138 45006
rect 49758 44994 49810 45006
rect 41682 44942 41694 44994
rect 41746 44942 41758 44994
rect 43810 44942 43822 44994
rect 43874 44942 43886 44994
rect 47058 44942 47070 44994
rect 47122 44942 47134 44994
rect 49410 44942 49422 44994
rect 49474 44942 49486 44994
rect 33742 44930 33794 44942
rect 49086 44930 49138 44942
rect 49758 44930 49810 44942
rect 11118 44882 11170 44894
rect 11118 44818 11170 44830
rect 19854 44882 19906 44894
rect 19854 44818 19906 44830
rect 20414 44882 20466 44894
rect 30046 44882 30098 44894
rect 26114 44830 26126 44882
rect 26178 44830 26190 44882
rect 20414 44818 20466 44830
rect 30046 44818 30098 44830
rect 33182 44882 33234 44894
rect 33182 44818 33234 44830
rect 1344 44714 58576 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 58576 44714
rect 1344 44628 58576 44662
rect 7422 44546 7474 44558
rect 7422 44482 7474 44494
rect 22878 44546 22930 44558
rect 41918 44546 41970 44558
rect 25330 44494 25342 44546
rect 25394 44494 25406 44546
rect 22878 44482 22930 44494
rect 41918 44482 41970 44494
rect 7646 44434 7698 44446
rect 30606 44434 30658 44446
rect 20290 44382 20302 44434
rect 20354 44382 20366 44434
rect 27010 44382 27022 44434
rect 27074 44382 27086 44434
rect 7646 44370 7698 44382
rect 30606 44370 30658 44382
rect 31502 44434 31554 44446
rect 42030 44434 42082 44446
rect 50542 44434 50594 44446
rect 33618 44382 33630 44434
rect 33682 44382 33694 44434
rect 37762 44382 37774 44434
rect 37826 44382 37838 44434
rect 42466 44382 42478 44434
rect 42530 44382 42542 44434
rect 43474 44382 43486 44434
rect 43538 44382 43550 44434
rect 49746 44382 49758 44434
rect 49810 44382 49822 44434
rect 31502 44370 31554 44382
rect 42030 44370 42082 44382
rect 50542 44370 50594 44382
rect 51998 44434 52050 44446
rect 52994 44382 53006 44434
rect 53058 44382 53070 44434
rect 53666 44382 53678 44434
rect 53730 44382 53742 44434
rect 58146 44382 58158 44434
rect 58210 44382 58222 44434
rect 51998 44370 52050 44382
rect 8878 44322 8930 44334
rect 7858 44270 7870 44322
rect 7922 44270 7934 44322
rect 8878 44258 8930 44270
rect 9662 44322 9714 44334
rect 9662 44258 9714 44270
rect 10110 44322 10162 44334
rect 10110 44258 10162 44270
rect 10670 44322 10722 44334
rect 22990 44322 23042 44334
rect 42814 44322 42866 44334
rect 51550 44322 51602 44334
rect 14242 44270 14254 44322
rect 14306 44270 14318 44322
rect 15138 44270 15150 44322
rect 15202 44270 15214 44322
rect 15474 44270 15486 44322
rect 15538 44270 15550 44322
rect 16258 44270 16270 44322
rect 16322 44270 16334 44322
rect 17378 44270 17390 44322
rect 17442 44270 17454 44322
rect 23426 44270 23438 44322
rect 23490 44270 23502 44322
rect 24546 44270 24558 44322
rect 24610 44270 24622 44322
rect 26450 44270 26462 44322
rect 26514 44270 26526 44322
rect 30258 44270 30270 44322
rect 30322 44270 30334 44322
rect 30930 44270 30942 44322
rect 30994 44270 31006 44322
rect 34402 44270 34414 44322
rect 34466 44270 34478 44322
rect 40674 44270 40686 44322
rect 40738 44270 40750 44322
rect 43026 44270 43038 44322
rect 43090 44270 43102 44322
rect 43362 44270 43374 44322
rect 43426 44270 43438 44322
rect 44034 44270 44046 44322
rect 44098 44270 44110 44322
rect 45490 44270 45502 44322
rect 45554 44270 45566 44322
rect 10670 44258 10722 44270
rect 22990 44258 23042 44270
rect 42814 44258 42866 44270
rect 51550 44258 51602 44270
rect 51774 44322 51826 44334
rect 51774 44258 51826 44270
rect 52110 44322 52162 44334
rect 54350 44322 54402 44334
rect 52770 44270 52782 44322
rect 52834 44270 52846 44322
rect 53554 44270 53566 44322
rect 53618 44270 53630 44322
rect 52110 44258 52162 44270
rect 54350 44258 54402 44270
rect 54686 44322 54738 44334
rect 55234 44270 55246 44322
rect 55298 44270 55310 44322
rect 54686 44258 54738 44270
rect 7310 44210 7362 44222
rect 7310 44146 7362 44158
rect 8206 44210 8258 44222
rect 8206 44146 8258 44158
rect 8430 44210 8482 44222
rect 8430 44146 8482 44158
rect 9102 44210 9154 44222
rect 9102 44146 9154 44158
rect 9438 44210 9490 44222
rect 27358 44210 27410 44222
rect 15922 44158 15934 44210
rect 15986 44158 15998 44210
rect 16594 44158 16606 44210
rect 16658 44158 16670 44210
rect 18162 44158 18174 44210
rect 18226 44158 18238 44210
rect 25778 44158 25790 44210
rect 25842 44158 25854 44210
rect 9438 44146 9490 44158
rect 27358 44146 27410 44158
rect 27806 44210 27858 44222
rect 27806 44146 27858 44158
rect 36318 44210 36370 44222
rect 54462 44210 54514 44222
rect 39890 44158 39902 44210
rect 39954 44158 39966 44210
rect 56018 44158 56030 44210
rect 56082 44158 56094 44210
rect 36318 44146 36370 44158
rect 54462 44146 54514 44158
rect 8542 44098 8594 44110
rect 8542 44034 8594 44046
rect 9214 44098 9266 44110
rect 9214 44034 9266 44046
rect 9998 44098 10050 44110
rect 9998 44034 10050 44046
rect 10222 44098 10274 44110
rect 10222 44034 10274 44046
rect 14590 44098 14642 44110
rect 14590 44034 14642 44046
rect 14702 44098 14754 44110
rect 14702 44034 14754 44046
rect 14814 44098 14866 44110
rect 14814 44034 14866 44046
rect 22878 44098 22930 44110
rect 22878 44034 22930 44046
rect 30494 44098 30546 44110
rect 30494 44034 30546 44046
rect 30718 44098 30770 44110
rect 30718 44034 30770 44046
rect 36206 44098 36258 44110
rect 36206 44034 36258 44046
rect 42478 44098 42530 44110
rect 42478 44034 42530 44046
rect 42590 44098 42642 44110
rect 42590 44034 42642 44046
rect 43598 44098 43650 44110
rect 43598 44034 43650 44046
rect 43822 44098 43874 44110
rect 43822 44034 43874 44046
rect 1344 43930 58576 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 58576 43930
rect 1344 43844 58576 43878
rect 17950 43762 18002 43774
rect 17950 43698 18002 43710
rect 31166 43762 31218 43774
rect 31166 43698 31218 43710
rect 32174 43762 32226 43774
rect 32174 43698 32226 43710
rect 39902 43762 39954 43774
rect 39902 43698 39954 43710
rect 15374 43650 15426 43662
rect 6850 43598 6862 43650
rect 6914 43598 6926 43650
rect 10322 43598 10334 43650
rect 10386 43598 10398 43650
rect 15374 43586 15426 43598
rect 16382 43650 16434 43662
rect 31838 43650 31890 43662
rect 38222 43650 38274 43662
rect 29810 43598 29822 43650
rect 29874 43598 29886 43650
rect 35410 43598 35422 43650
rect 35474 43598 35486 43650
rect 16382 43586 16434 43598
rect 31838 43586 31890 43598
rect 38222 43586 38274 43598
rect 39342 43650 39394 43662
rect 39342 43586 39394 43598
rect 39566 43650 39618 43662
rect 39566 43586 39618 43598
rect 44270 43650 44322 43662
rect 44270 43586 44322 43598
rect 54910 43650 54962 43662
rect 54910 43586 54962 43598
rect 55022 43650 55074 43662
rect 55022 43586 55074 43598
rect 57038 43650 57090 43662
rect 57038 43586 57090 43598
rect 15598 43538 15650 43550
rect 7634 43486 7646 43538
rect 7698 43486 7710 43538
rect 13570 43486 13582 43538
rect 13634 43486 13646 43538
rect 15598 43474 15650 43486
rect 16046 43538 16098 43550
rect 16046 43474 16098 43486
rect 18062 43538 18114 43550
rect 30594 43498 30606 43550
rect 30658 43498 30670 43550
rect 32062 43538 32114 43550
rect 18062 43474 18114 43486
rect 32062 43474 32114 43486
rect 32286 43538 32338 43550
rect 32286 43474 32338 43486
rect 32398 43538 32450 43550
rect 37998 43538 38050 43550
rect 34626 43486 34638 43538
rect 34690 43486 34702 43538
rect 32398 43474 32450 43486
rect 37998 43474 38050 43486
rect 38110 43538 38162 43550
rect 38110 43474 38162 43486
rect 38334 43538 38386 43550
rect 39118 43538 39170 43550
rect 54574 43538 54626 43550
rect 38546 43486 38558 43538
rect 38610 43486 38622 43538
rect 38882 43486 38894 43538
rect 38946 43486 38958 43538
rect 45378 43486 45390 43538
rect 45442 43486 45454 43538
rect 50754 43486 50766 43538
rect 50818 43486 50830 43538
rect 51986 43486 51998 43538
rect 52050 43486 52062 43538
rect 52434 43486 52446 43538
rect 52498 43486 52510 43538
rect 53106 43486 53118 43538
rect 53170 43486 53182 43538
rect 38334 43474 38386 43486
rect 39118 43474 39170 43486
rect 54574 43474 54626 43486
rect 15822 43426 15874 43438
rect 4722 43374 4734 43426
rect 4786 43374 4798 43426
rect 15822 43362 15874 43374
rect 25678 43426 25730 43438
rect 33182 43426 33234 43438
rect 39230 43426 39282 43438
rect 27682 43374 27694 43426
rect 27746 43374 27758 43426
rect 37538 43374 37550 43426
rect 37602 43374 37614 43426
rect 25678 43362 25730 43374
rect 33182 43362 33234 43374
rect 39230 43362 39282 43374
rect 40014 43426 40066 43438
rect 40014 43362 40066 43374
rect 43262 43426 43314 43438
rect 43262 43362 43314 43374
rect 44718 43426 44770 43438
rect 46050 43374 46062 43426
rect 46114 43374 46126 43426
rect 48178 43374 48190 43426
rect 48242 43374 48254 43426
rect 50306 43374 50318 43426
rect 50370 43374 50382 43426
rect 53890 43374 53902 43426
rect 53954 43374 53966 43426
rect 44718 43362 44770 43374
rect 25566 43314 25618 43326
rect 25566 43250 25618 43262
rect 54462 43314 54514 43326
rect 54462 43250 54514 43262
rect 56926 43314 56978 43326
rect 56926 43250 56978 43262
rect 1344 43146 58576 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 58576 43146
rect 1344 43060 58576 43094
rect 46286 42978 46338 42990
rect 9538 42926 9550 42978
rect 9602 42926 9614 42978
rect 46286 42914 46338 42926
rect 46734 42978 46786 42990
rect 52782 42978 52834 42990
rect 51538 42926 51550 42978
rect 51602 42926 51614 42978
rect 46734 42914 46786 42926
rect 52782 42914 52834 42926
rect 55918 42978 55970 42990
rect 55918 42914 55970 42926
rect 56926 42978 56978 42990
rect 56926 42914 56978 42926
rect 21422 42866 21474 42878
rect 18722 42814 18734 42866
rect 18786 42814 18798 42866
rect 25106 42814 25118 42866
rect 25170 42814 25182 42866
rect 27234 42814 27246 42866
rect 27298 42814 27310 42866
rect 36418 42814 36430 42866
rect 36482 42814 36494 42866
rect 51314 42814 51326 42866
rect 51378 42814 51390 42866
rect 21422 42802 21474 42814
rect 9998 42754 10050 42766
rect 9998 42690 10050 42702
rect 10222 42754 10274 42766
rect 10222 42690 10274 42702
rect 13806 42754 13858 42766
rect 13806 42690 13858 42702
rect 14366 42754 14418 42766
rect 30830 42754 30882 42766
rect 37550 42754 37602 42766
rect 20738 42702 20750 42754
rect 20802 42702 20814 42754
rect 24322 42702 24334 42754
rect 24386 42702 24398 42754
rect 30594 42702 30606 42754
rect 30658 42702 30670 42754
rect 31266 42702 31278 42754
rect 31330 42702 31342 42754
rect 33618 42702 33630 42754
rect 33682 42702 33694 42754
rect 14366 42690 14418 42702
rect 30830 42690 30882 42702
rect 37550 42690 37602 42702
rect 37998 42754 38050 42766
rect 37998 42690 38050 42702
rect 46286 42754 46338 42766
rect 46286 42690 46338 42702
rect 46958 42754 47010 42766
rect 52894 42754 52946 42766
rect 50754 42702 50766 42754
rect 50818 42702 50830 42754
rect 50978 42702 50990 42754
rect 51042 42702 51054 42754
rect 51762 42702 51774 42754
rect 51826 42702 51838 42754
rect 46958 42690 47010 42702
rect 52894 42690 52946 42702
rect 53230 42754 53282 42766
rect 53230 42690 53282 42702
rect 56142 42754 56194 42766
rect 56142 42690 56194 42702
rect 10110 42642 10162 42654
rect 10110 42578 10162 42590
rect 10670 42642 10722 42654
rect 10670 42578 10722 42590
rect 11006 42642 11058 42654
rect 11006 42578 11058 42590
rect 14142 42642 14194 42654
rect 14142 42578 14194 42590
rect 22094 42642 22146 42654
rect 22094 42578 22146 42590
rect 29262 42642 29314 42654
rect 30942 42642 30994 42654
rect 46174 42642 46226 42654
rect 29922 42590 29934 42642
rect 29986 42590 29998 42642
rect 34290 42590 34302 42642
rect 34354 42590 34366 42642
rect 29262 42578 29314 42590
rect 30942 42578 30994 42590
rect 46174 42578 46226 42590
rect 52782 42642 52834 42654
rect 52782 42578 52834 42590
rect 53342 42642 53394 42654
rect 53342 42578 53394 42590
rect 55358 42642 55410 42654
rect 55358 42578 55410 42590
rect 55582 42642 55634 42654
rect 55582 42578 55634 42590
rect 56814 42642 56866 42654
rect 56814 42578 56866 42590
rect 13918 42530 13970 42542
rect 13918 42466 13970 42478
rect 21982 42530 22034 42542
rect 21982 42466 22034 42478
rect 27806 42530 27858 42542
rect 27806 42466 27858 42478
rect 29150 42530 29202 42542
rect 29150 42466 29202 42478
rect 29598 42530 29650 42542
rect 29598 42466 29650 42478
rect 31054 42530 31106 42542
rect 31054 42466 31106 42478
rect 31838 42530 31890 42542
rect 31838 42466 31890 42478
rect 37662 42530 37714 42542
rect 37662 42466 37714 42478
rect 37774 42530 37826 42542
rect 37774 42466 37826 42478
rect 37886 42530 37938 42542
rect 37886 42466 37938 42478
rect 38670 42530 38722 42542
rect 38670 42466 38722 42478
rect 39006 42530 39058 42542
rect 39006 42466 39058 42478
rect 39790 42530 39842 42542
rect 39790 42466 39842 42478
rect 45950 42530 46002 42542
rect 45950 42466 46002 42478
rect 55134 42530 55186 42542
rect 55134 42466 55186 42478
rect 56254 42530 56306 42542
rect 56254 42466 56306 42478
rect 1344 42362 58576 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 58576 42362
rect 1344 42276 58576 42310
rect 32062 42194 32114 42206
rect 32062 42130 32114 42142
rect 38110 42194 38162 42206
rect 38110 42130 38162 42142
rect 44830 42194 44882 42206
rect 44830 42130 44882 42142
rect 45278 42194 45330 42206
rect 45278 42130 45330 42142
rect 45502 42194 45554 42206
rect 45502 42130 45554 42142
rect 48078 42194 48130 42206
rect 48078 42130 48130 42142
rect 24110 42082 24162 42094
rect 24110 42018 24162 42030
rect 26014 42082 26066 42094
rect 26014 42018 26066 42030
rect 26462 42082 26514 42094
rect 32286 42082 32338 42094
rect 26898 42030 26910 42082
rect 26962 42030 26974 42082
rect 28690 42030 28702 42082
rect 28754 42030 28766 42082
rect 26462 42018 26514 42030
rect 32286 42018 32338 42030
rect 45166 42082 45218 42094
rect 45166 42018 45218 42030
rect 47966 42082 48018 42094
rect 47966 42018 48018 42030
rect 23774 41970 23826 41982
rect 12002 41918 12014 41970
rect 12066 41918 12078 41970
rect 12674 41918 12686 41970
rect 12738 41918 12750 41970
rect 15362 41918 15374 41970
rect 15426 41918 15438 41970
rect 20402 41918 20414 41970
rect 20466 41918 20478 41970
rect 21186 41918 21198 41970
rect 21250 41918 21262 41970
rect 23774 41906 23826 41918
rect 23886 41970 23938 41982
rect 23886 41906 23938 41918
rect 23998 41970 24050 41982
rect 23998 41906 24050 41918
rect 24222 41970 24274 41982
rect 26238 41970 26290 41982
rect 25778 41918 25790 41970
rect 25842 41918 25854 41970
rect 24222 41906 24274 41918
rect 26238 41906 26290 41918
rect 27246 41970 27298 41982
rect 32398 41970 32450 41982
rect 27906 41918 27918 41970
rect 27970 41918 27982 41970
rect 31826 41918 31838 41970
rect 31890 41918 31902 41970
rect 27246 41906 27298 41918
rect 32398 41906 32450 41918
rect 35310 41970 35362 41982
rect 35310 41906 35362 41918
rect 35422 41970 35474 41982
rect 35422 41906 35474 41918
rect 37214 41970 37266 41982
rect 37774 41970 37826 41982
rect 37538 41918 37550 41970
rect 37602 41918 37614 41970
rect 37214 41906 37266 41918
rect 37774 41906 37826 41918
rect 37998 41970 38050 41982
rect 47630 41970 47682 41982
rect 40898 41918 40910 41970
rect 40962 41918 40974 41970
rect 48962 41918 48974 41970
rect 49026 41918 49038 41970
rect 52210 41918 52222 41970
rect 52274 41918 52286 41970
rect 37998 41906 38050 41918
rect 47630 41906 47682 41918
rect 18622 41858 18674 41870
rect 25342 41858 25394 41870
rect 33070 41858 33122 41870
rect 14802 41806 14814 41858
rect 14866 41806 14878 41858
rect 15250 41806 15262 41858
rect 15314 41806 15326 41858
rect 23314 41806 23326 41858
rect 23378 41806 23390 41858
rect 25890 41806 25902 41858
rect 25954 41806 25966 41858
rect 30818 41806 30830 41858
rect 30882 41806 30894 41858
rect 32274 41806 32286 41858
rect 32338 41806 32350 41858
rect 18622 41794 18674 41806
rect 25342 41794 25394 41806
rect 33070 41794 33122 41806
rect 33630 41858 33682 41870
rect 33630 41794 33682 41806
rect 37886 41858 37938 41870
rect 44494 41858 44546 41870
rect 41682 41806 41694 41858
rect 41746 41806 41758 41858
rect 43810 41806 43822 41858
rect 43874 41806 43886 41858
rect 37886 41794 37938 41806
rect 44494 41794 44546 41806
rect 47182 41858 47234 41870
rect 49634 41806 49646 41858
rect 49698 41806 49710 41858
rect 51762 41806 51774 41858
rect 51826 41806 51838 41858
rect 52882 41806 52894 41858
rect 52946 41806 52958 41858
rect 55010 41806 55022 41858
rect 55074 41806 55086 41858
rect 47182 41794 47234 41806
rect 16606 41746 16658 41758
rect 16606 41682 16658 41694
rect 18734 41746 18786 41758
rect 18734 41682 18786 41694
rect 33182 41746 33234 41758
rect 33182 41682 33234 41694
rect 47518 41746 47570 41758
rect 47518 41682 47570 41694
rect 48078 41746 48130 41758
rect 48078 41682 48130 41694
rect 1344 41578 58576 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 58576 41578
rect 1344 41492 58576 41526
rect 49086 41410 49138 41422
rect 49086 41346 49138 41358
rect 49646 41410 49698 41422
rect 49646 41346 49698 41358
rect 16494 41298 16546 41310
rect 29374 41298 29426 41310
rect 37214 41298 37266 41310
rect 9202 41246 9214 41298
rect 9266 41246 9278 41298
rect 11330 41246 11342 41298
rect 11394 41246 11406 41298
rect 17490 41246 17502 41298
rect 17554 41246 17566 41298
rect 19618 41246 19630 41298
rect 19682 41246 19694 41298
rect 31378 41246 31390 41298
rect 31442 41246 31454 41298
rect 33506 41246 33518 41298
rect 33570 41246 33582 41298
rect 40898 41246 40910 41298
rect 40962 41246 40974 41298
rect 48066 41246 48078 41298
rect 48130 41246 48142 41298
rect 49410 41246 49422 41298
rect 49474 41246 49486 41298
rect 16494 41234 16546 41246
rect 29374 41234 29426 41246
rect 37214 41234 37266 41246
rect 16382 41186 16434 41198
rect 25790 41186 25842 41198
rect 8418 41134 8430 41186
rect 8482 41134 8494 41186
rect 15810 41134 15822 41186
rect 15874 41134 15886 41186
rect 20402 41134 20414 41186
rect 20466 41134 20478 41186
rect 16382 41122 16434 41134
rect 25790 41122 25842 41134
rect 26126 41186 26178 41198
rect 43710 41186 43762 41198
rect 34290 41134 34302 41186
rect 34354 41134 34366 41186
rect 43138 41134 43150 41186
rect 43202 41134 43214 41186
rect 43474 41134 43486 41186
rect 43538 41134 43550 41186
rect 26126 41122 26178 41134
rect 43710 41122 43762 41134
rect 44046 41186 44098 41198
rect 49870 41186 49922 41198
rect 45154 41134 45166 41186
rect 45218 41134 45230 41186
rect 44046 41122 44098 41134
rect 49870 41122 49922 41134
rect 51214 41186 51266 41198
rect 51214 41122 51266 41134
rect 51550 41186 51602 41198
rect 52658 41134 52670 41186
rect 52722 41134 52734 41186
rect 51550 41122 51602 41134
rect 12798 41074 12850 41086
rect 12798 41010 12850 41022
rect 26350 41074 26402 41086
rect 29486 41074 29538 41086
rect 27458 41022 27470 41074
rect 27522 41022 27534 41074
rect 26350 41010 26402 41022
rect 29486 41010 29538 41022
rect 30158 41074 30210 41086
rect 37102 41074 37154 41086
rect 49310 41074 49362 41086
rect 30482 41022 30494 41074
rect 30546 41022 30558 41074
rect 45938 41022 45950 41074
rect 46002 41022 46014 41074
rect 30158 41010 30210 41022
rect 37102 41010 37154 41022
rect 49310 41010 49362 41022
rect 51662 41074 51714 41086
rect 55458 41022 55470 41074
rect 55522 41022 55534 41074
rect 51662 41010 51714 41022
rect 12686 40962 12738 40974
rect 12686 40898 12738 40910
rect 25006 40962 25058 40974
rect 25006 40898 25058 40910
rect 25342 40962 25394 40974
rect 25342 40898 25394 40910
rect 25902 40962 25954 40974
rect 25902 40898 25954 40910
rect 26014 40962 26066 40974
rect 26014 40898 26066 40910
rect 26910 40962 26962 40974
rect 26910 40898 26962 40910
rect 27806 40962 27858 40974
rect 27806 40898 27858 40910
rect 28702 40962 28754 40974
rect 28702 40898 28754 40910
rect 29262 40962 29314 40974
rect 29262 40898 29314 40910
rect 43822 40962 43874 40974
rect 43822 40898 43874 40910
rect 43934 40962 43986 40974
rect 43934 40898 43986 40910
rect 48750 40962 48802 40974
rect 48750 40898 48802 40910
rect 51886 40962 51938 40974
rect 51886 40898 51938 40910
rect 1344 40794 58576 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 58576 40794
rect 1344 40708 58576 40742
rect 17502 40626 17554 40638
rect 17502 40562 17554 40574
rect 18846 40626 18898 40638
rect 18846 40562 18898 40574
rect 18958 40626 19010 40638
rect 18958 40562 19010 40574
rect 19630 40626 19682 40638
rect 19630 40562 19682 40574
rect 24222 40626 24274 40638
rect 40350 40626 40402 40638
rect 38882 40574 38894 40626
rect 38946 40574 38958 40626
rect 39554 40574 39566 40626
rect 39618 40574 39630 40626
rect 24222 40562 24274 40574
rect 40350 40562 40402 40574
rect 41022 40626 41074 40638
rect 41022 40562 41074 40574
rect 42254 40626 42306 40638
rect 42254 40562 42306 40574
rect 43374 40626 43426 40638
rect 52334 40626 52386 40638
rect 44258 40574 44270 40626
rect 44322 40574 44334 40626
rect 49746 40574 49758 40626
rect 49810 40574 49822 40626
rect 43374 40562 43426 40574
rect 52334 40562 52386 40574
rect 54238 40626 54290 40638
rect 54238 40562 54290 40574
rect 54910 40626 54962 40638
rect 54910 40562 54962 40574
rect 18510 40514 18562 40526
rect 42366 40514 42418 40526
rect 8306 40462 8318 40514
rect 8370 40462 8382 40514
rect 12114 40462 12126 40514
rect 12178 40462 12190 40514
rect 27906 40462 27918 40514
rect 27970 40462 27982 40514
rect 36418 40462 36430 40514
rect 36482 40462 36494 40514
rect 41906 40462 41918 40514
rect 41970 40462 41982 40514
rect 18510 40450 18562 40462
rect 42366 40450 42418 40462
rect 44830 40514 44882 40526
rect 44830 40450 44882 40462
rect 44942 40514 44994 40526
rect 44942 40450 44994 40462
rect 45838 40514 45890 40526
rect 45838 40450 45890 40462
rect 53006 40514 53058 40526
rect 53006 40450 53058 40462
rect 54686 40514 54738 40526
rect 54686 40450 54738 40462
rect 55806 40514 55858 40526
rect 57810 40462 57822 40514
rect 57874 40462 57886 40514
rect 55806 40450 55858 40462
rect 9662 40402 9714 40414
rect 16382 40402 16434 40414
rect 4946 40350 4958 40402
rect 5010 40350 5022 40402
rect 11442 40350 11454 40402
rect 11506 40350 11518 40402
rect 16146 40350 16158 40402
rect 16210 40350 16222 40402
rect 9662 40338 9714 40350
rect 16382 40338 16434 40350
rect 16606 40402 16658 40414
rect 18734 40402 18786 40414
rect 16818 40350 16830 40402
rect 16882 40350 16894 40402
rect 16606 40338 16658 40350
rect 18734 40338 18786 40350
rect 19070 40402 19122 40414
rect 24110 40402 24162 40414
rect 20850 40350 20862 40402
rect 20914 40350 20926 40402
rect 19070 40338 19122 40350
rect 24110 40338 24162 40350
rect 24446 40402 24498 40414
rect 39902 40402 39954 40414
rect 43934 40402 43986 40414
rect 24658 40350 24670 40402
rect 24722 40350 24734 40402
rect 29026 40350 29038 40402
rect 29090 40350 29102 40402
rect 35746 40350 35758 40402
rect 35810 40350 35822 40402
rect 39106 40350 39118 40402
rect 39170 40350 39182 40402
rect 41682 40350 41694 40402
rect 41746 40350 41758 40402
rect 24446 40338 24498 40350
rect 39902 40338 39954 40350
rect 43934 40338 43986 40350
rect 45166 40402 45218 40414
rect 45166 40338 45218 40350
rect 45502 40402 45554 40414
rect 45502 40338 45554 40350
rect 45614 40402 45666 40414
rect 45614 40338 45666 40350
rect 46062 40402 46114 40414
rect 46062 40338 46114 40350
rect 49422 40402 49474 40414
rect 49422 40338 49474 40350
rect 51886 40402 51938 40414
rect 51886 40338 51938 40350
rect 52782 40402 52834 40414
rect 52782 40338 52834 40350
rect 53230 40402 53282 40414
rect 53230 40338 53282 40350
rect 54574 40402 54626 40414
rect 54574 40338 54626 40350
rect 57598 40402 57650 40414
rect 58034 40350 58046 40402
rect 58098 40350 58110 40402
rect 57598 40338 57650 40350
rect 16494 40290 16546 40302
rect 24334 40290 24386 40302
rect 14242 40238 14254 40290
rect 14306 40238 14318 40290
rect 21522 40238 21534 40290
rect 21586 40238 21598 40290
rect 23650 40238 23662 40290
rect 23714 40238 23726 40290
rect 16494 40226 16546 40238
rect 24334 40226 24386 40238
rect 34526 40290 34578 40302
rect 46286 40290 46338 40302
rect 38546 40238 38558 40290
rect 38610 40238 38622 40290
rect 40898 40238 40910 40290
rect 40962 40238 40974 40290
rect 34526 40226 34578 40238
rect 46286 40226 46338 40238
rect 53454 40290 53506 40302
rect 53454 40226 53506 40238
rect 55246 40290 55298 40302
rect 55246 40226 55298 40238
rect 41246 40178 41298 40190
rect 41246 40114 41298 40126
rect 52670 40178 52722 40190
rect 52670 40114 52722 40126
rect 55470 40178 55522 40190
rect 55470 40114 55522 40126
rect 55918 40178 55970 40190
rect 55918 40114 55970 40126
rect 56030 40178 56082 40190
rect 56030 40114 56082 40126
rect 1344 40010 58576 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 58576 40010
rect 1344 39924 58576 39958
rect 22318 39842 22370 39854
rect 34514 39790 34526 39842
rect 34578 39839 34590 39842
rect 34738 39839 34750 39842
rect 34578 39793 34750 39839
rect 34578 39790 34590 39793
rect 34738 39790 34750 39793
rect 34802 39790 34814 39842
rect 22318 39778 22370 39790
rect 22430 39730 22482 39742
rect 4610 39678 4622 39730
rect 4674 39678 4686 39730
rect 5618 39678 5630 39730
rect 5682 39678 5694 39730
rect 16370 39678 16382 39730
rect 16434 39678 16446 39730
rect 22430 39666 22482 39678
rect 24782 39730 24834 39742
rect 29710 39730 29762 39742
rect 28130 39678 28142 39730
rect 28194 39678 28206 39730
rect 24782 39666 24834 39678
rect 29710 39666 29762 39678
rect 38110 39730 38162 39742
rect 38110 39666 38162 39678
rect 38558 39730 38610 39742
rect 38558 39666 38610 39678
rect 45390 39730 45442 39742
rect 53678 39730 53730 39742
rect 53106 39678 53118 39730
rect 53170 39678 53182 39730
rect 45390 39666 45442 39678
rect 53678 39666 53730 39678
rect 54350 39730 54402 39742
rect 56018 39678 56030 39730
rect 56082 39678 56094 39730
rect 58146 39678 58158 39730
rect 58210 39678 58222 39730
rect 54350 39666 54402 39678
rect 17166 39618 17218 39630
rect 1810 39566 1822 39618
rect 1874 39566 1886 39618
rect 8418 39566 8430 39618
rect 8482 39566 8494 39618
rect 13458 39566 13470 39618
rect 13522 39566 13534 39618
rect 16706 39566 16718 39618
rect 16770 39566 16782 39618
rect 17166 39554 17218 39566
rect 17278 39618 17330 39630
rect 17278 39554 17330 39566
rect 17838 39618 17890 39630
rect 35758 39618 35810 39630
rect 25330 39566 25342 39618
rect 25394 39566 25406 39618
rect 35298 39566 35310 39618
rect 35362 39566 35374 39618
rect 17838 39554 17890 39566
rect 35758 39554 35810 39566
rect 41022 39618 41074 39630
rect 42142 39618 42194 39630
rect 52670 39618 52722 39630
rect 41906 39566 41918 39618
rect 41970 39566 41982 39618
rect 42578 39566 42590 39618
rect 42642 39566 42654 39618
rect 54786 39566 54798 39618
rect 54850 39566 54862 39618
rect 55234 39566 55246 39618
rect 55298 39566 55310 39618
rect 41022 39554 41074 39566
rect 42142 39554 42194 39566
rect 52670 39554 52722 39566
rect 8878 39506 8930 39518
rect 2482 39454 2494 39506
rect 2546 39454 2558 39506
rect 7746 39454 7758 39506
rect 7810 39454 7822 39506
rect 8878 39442 8930 39454
rect 8990 39506 9042 39518
rect 8990 39442 9042 39454
rect 9662 39506 9714 39518
rect 16942 39506 16994 39518
rect 24894 39506 24946 39518
rect 29262 39506 29314 39518
rect 14242 39454 14254 39506
rect 14306 39454 14318 39506
rect 18722 39454 18734 39506
rect 18786 39454 18798 39506
rect 26002 39454 26014 39506
rect 26066 39454 26078 39506
rect 9662 39442 9714 39454
rect 16942 39442 16994 39454
rect 24894 39442 24946 39454
rect 29262 39442 29314 39454
rect 33518 39506 33570 39518
rect 33518 39442 33570 39454
rect 33742 39506 33794 39518
rect 33742 39442 33794 39454
rect 34078 39506 34130 39518
rect 48526 39506 48578 39518
rect 41346 39454 41358 39506
rect 41410 39454 41422 39506
rect 34078 39442 34130 39454
rect 48526 39442 48578 39454
rect 9214 39394 9266 39406
rect 9214 39330 9266 39342
rect 9326 39394 9378 39406
rect 9326 39330 9378 39342
rect 9550 39394 9602 39406
rect 9550 39330 9602 39342
rect 17054 39394 17106 39406
rect 17054 39330 17106 39342
rect 19070 39394 19122 39406
rect 19070 39330 19122 39342
rect 19630 39394 19682 39406
rect 19630 39330 19682 39342
rect 29150 39394 29202 39406
rect 29150 39330 29202 39342
rect 33182 39394 33234 39406
rect 33182 39330 33234 39342
rect 33406 39394 33458 39406
rect 33406 39330 33458 39342
rect 33966 39394 34018 39406
rect 33966 39330 34018 39342
rect 34526 39394 34578 39406
rect 34526 39330 34578 39342
rect 36318 39394 36370 39406
rect 36318 39330 36370 39342
rect 37774 39394 37826 39406
rect 37774 39330 37826 39342
rect 42254 39394 42306 39406
rect 42254 39330 42306 39342
rect 42366 39394 42418 39406
rect 42366 39330 42418 39342
rect 43150 39394 43202 39406
rect 43150 39330 43202 39342
rect 44942 39394 44994 39406
rect 44942 39330 44994 39342
rect 47406 39394 47458 39406
rect 49086 39394 49138 39406
rect 48626 39342 48638 39394
rect 48690 39391 48702 39394
rect 48850 39391 48862 39394
rect 48690 39345 48862 39391
rect 48690 39342 48702 39345
rect 48850 39342 48862 39345
rect 48914 39342 48926 39394
rect 49410 39342 49422 39394
rect 49474 39342 49486 39394
rect 47406 39330 47458 39342
rect 49086 39330 49138 39342
rect 1344 39226 58576 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 58576 39226
rect 1344 39140 58576 39174
rect 5966 39058 6018 39070
rect 5966 38994 6018 39006
rect 7534 39058 7586 39070
rect 7534 38994 7586 39006
rect 14702 39058 14754 39070
rect 14702 38994 14754 39006
rect 19070 39058 19122 39070
rect 19070 38994 19122 39006
rect 19630 39058 19682 39070
rect 19630 38994 19682 39006
rect 36990 39058 37042 39070
rect 36990 38994 37042 39006
rect 37214 39058 37266 39070
rect 37214 38994 37266 39006
rect 37886 39058 37938 39070
rect 37886 38994 37938 39006
rect 38222 39058 38274 39070
rect 38222 38994 38274 39006
rect 45390 39058 45442 39070
rect 55470 39058 55522 39070
rect 46610 39006 46622 39058
rect 46674 39006 46686 39058
rect 45390 38994 45442 39006
rect 55470 38994 55522 39006
rect 55918 39058 55970 39070
rect 55918 38994 55970 39006
rect 56142 39058 56194 39070
rect 56142 38994 56194 39006
rect 5182 38946 5234 38958
rect 5182 38882 5234 38894
rect 5294 38946 5346 38958
rect 5294 38882 5346 38894
rect 5742 38946 5794 38958
rect 5742 38882 5794 38894
rect 7310 38946 7362 38958
rect 7310 38882 7362 38894
rect 14814 38946 14866 38958
rect 14814 38882 14866 38894
rect 18510 38946 18562 38958
rect 18510 38882 18562 38894
rect 30270 38946 30322 38958
rect 30270 38882 30322 38894
rect 32510 38946 32562 38958
rect 49310 38946 49362 38958
rect 34850 38894 34862 38946
rect 34914 38894 34926 38946
rect 35746 38894 35758 38946
rect 35810 38894 35822 38946
rect 32510 38882 32562 38894
rect 49310 38882 49362 38894
rect 55806 38946 55858 38958
rect 55806 38882 55858 38894
rect 5630 38834 5682 38846
rect 1810 38782 1822 38834
rect 1874 38782 1886 38834
rect 5630 38770 5682 38782
rect 6190 38834 6242 38846
rect 6190 38770 6242 38782
rect 6302 38834 6354 38846
rect 6302 38770 6354 38782
rect 6414 38834 6466 38846
rect 6414 38770 6466 38782
rect 6750 38834 6802 38846
rect 6750 38770 6802 38782
rect 7198 38834 7250 38846
rect 7198 38770 7250 38782
rect 7646 38834 7698 38846
rect 7646 38770 7698 38782
rect 8542 38834 8594 38846
rect 8542 38770 8594 38782
rect 8766 38834 8818 38846
rect 8766 38770 8818 38782
rect 9102 38834 9154 38846
rect 18734 38834 18786 38846
rect 12450 38782 12462 38834
rect 12514 38782 12526 38834
rect 9102 38770 9154 38782
rect 18734 38770 18786 38782
rect 18958 38834 19010 38846
rect 30606 38834 30658 38846
rect 37550 38834 37602 38846
rect 20402 38782 20414 38834
rect 20466 38782 20478 38834
rect 26898 38782 26910 38834
rect 26962 38782 26974 38834
rect 34962 38782 34974 38834
rect 35026 38782 35038 38834
rect 36642 38782 36654 38834
rect 36706 38782 36718 38834
rect 18958 38770 19010 38782
rect 30606 38770 30658 38782
rect 37550 38770 37602 38782
rect 39230 38834 39282 38846
rect 45726 38834 45778 38846
rect 43810 38782 43822 38834
rect 43874 38782 43886 38834
rect 39230 38770 39282 38782
rect 45726 38770 45778 38782
rect 45950 38834 46002 38846
rect 45950 38770 46002 38782
rect 46286 38834 46338 38846
rect 47518 38834 47570 38846
rect 46834 38782 46846 38834
rect 46898 38782 46910 38834
rect 46286 38770 46338 38782
rect 47518 38770 47570 38782
rect 47966 38834 48018 38846
rect 47966 38770 48018 38782
rect 48190 38834 48242 38846
rect 48190 38770 48242 38782
rect 48750 38834 48802 38846
rect 48750 38770 48802 38782
rect 48862 38834 48914 38846
rect 48862 38770 48914 38782
rect 48974 38834 49026 38846
rect 54910 38834 54962 38846
rect 52882 38782 52894 38834
rect 52946 38782 52958 38834
rect 48974 38770 49026 38782
rect 54910 38770 54962 38782
rect 57710 38834 57762 38846
rect 57710 38770 57762 38782
rect 8878 38722 8930 38734
rect 18062 38722 18114 38734
rect 2482 38670 2494 38722
rect 2546 38670 2558 38722
rect 4610 38670 4622 38722
rect 4674 38670 4686 38722
rect 9538 38670 9550 38722
rect 9602 38670 9614 38722
rect 11666 38670 11678 38722
rect 11730 38670 11742 38722
rect 8878 38658 8930 38670
rect 18062 38658 18114 38670
rect 18846 38722 18898 38734
rect 18846 38658 18898 38670
rect 20078 38722 20130 38734
rect 45838 38722 45890 38734
rect 21186 38670 21198 38722
rect 21250 38670 21262 38722
rect 23314 38670 23326 38722
rect 23378 38670 23390 38722
rect 27570 38670 27582 38722
rect 27634 38670 27646 38722
rect 29698 38670 29710 38722
rect 29762 38670 29774 38722
rect 30370 38670 30382 38722
rect 30434 38670 30446 38722
rect 35746 38670 35758 38722
rect 35810 38670 35822 38722
rect 38658 38670 38670 38722
rect 38722 38670 38734 38722
rect 40898 38670 40910 38722
rect 40962 38670 40974 38722
rect 43026 38670 43038 38722
rect 43090 38670 43102 38722
rect 20078 38658 20130 38670
rect 45838 38658 45890 38670
rect 47742 38722 47794 38734
rect 57150 38722 57202 38734
rect 49970 38670 49982 38722
rect 50034 38670 50046 38722
rect 52098 38670 52110 38722
rect 52162 38670 52174 38722
rect 47742 38658 47794 38670
rect 57150 38658 57202 38670
rect 5182 38610 5234 38622
rect 5182 38546 5234 38558
rect 17950 38610 18002 38622
rect 17950 38546 18002 38558
rect 30046 38610 30098 38622
rect 30046 38546 30098 38558
rect 30830 38610 30882 38622
rect 30830 38546 30882 38558
rect 36878 38610 36930 38622
rect 36878 38546 36930 38558
rect 1344 38442 58576 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 58576 38442
rect 1344 38356 58576 38390
rect 7646 38274 7698 38286
rect 7646 38210 7698 38222
rect 8766 38274 8818 38286
rect 8766 38210 8818 38222
rect 34190 38274 34242 38286
rect 42030 38274 42082 38286
rect 34402 38222 34414 38274
rect 34466 38271 34478 38274
rect 34962 38271 34974 38274
rect 34466 38225 34974 38271
rect 34466 38222 34478 38225
rect 34962 38222 34974 38225
rect 35026 38222 35038 38274
rect 34190 38210 34242 38222
rect 42030 38210 42082 38222
rect 5854 38162 5906 38174
rect 23662 38162 23714 38174
rect 17042 38110 17054 38162
rect 17106 38110 17118 38162
rect 19170 38110 19182 38162
rect 19234 38110 19246 38162
rect 5854 38098 5906 38110
rect 23662 38098 23714 38110
rect 28030 38162 28082 38174
rect 34078 38162 34130 38174
rect 33506 38110 33518 38162
rect 33570 38110 33582 38162
rect 28030 38098 28082 38110
rect 34078 38098 34130 38110
rect 34750 38162 34802 38174
rect 41918 38162 41970 38174
rect 44270 38162 44322 38174
rect 40002 38110 40014 38162
rect 40066 38110 40078 38162
rect 43698 38110 43710 38162
rect 43762 38110 43774 38162
rect 45042 38110 45054 38162
rect 45106 38110 45118 38162
rect 34750 38098 34802 38110
rect 41918 38098 41970 38110
rect 44270 38098 44322 38110
rect 6078 38050 6130 38062
rect 6078 37986 6130 37998
rect 6526 38050 6578 38062
rect 6526 37986 6578 37998
rect 6862 38050 6914 38062
rect 6862 37986 6914 37998
rect 7534 38050 7586 38062
rect 7534 37986 7586 37998
rect 8878 38050 8930 38062
rect 22990 38050 23042 38062
rect 30046 38050 30098 38062
rect 35646 38050 35698 38062
rect 16370 37998 16382 38050
rect 16434 37998 16446 38050
rect 27570 37998 27582 38050
rect 27634 37998 27646 38050
rect 30594 37998 30606 38050
rect 30658 37998 30670 38050
rect 8878 37986 8930 37998
rect 22990 37986 23042 37998
rect 30046 37986 30098 37998
rect 35646 37986 35698 37998
rect 36318 38050 36370 38062
rect 50542 38050 50594 38062
rect 37202 37998 37214 38050
rect 37266 37998 37278 38050
rect 43586 37998 43598 38050
rect 43650 37998 43662 38050
rect 48738 37998 48750 38050
rect 48802 37998 48814 38050
rect 55906 37998 55918 38050
rect 55970 37998 55982 38050
rect 58146 37998 58158 38050
rect 58210 37998 58222 38050
rect 36318 37986 36370 37998
rect 50542 37986 50594 37998
rect 5742 37938 5794 37950
rect 5742 37874 5794 37886
rect 6302 37938 6354 37950
rect 6302 37874 6354 37886
rect 11006 37938 11058 37950
rect 11006 37874 11058 37886
rect 11342 37938 11394 37950
rect 11342 37874 11394 37886
rect 28702 37938 28754 37950
rect 28702 37874 28754 37886
rect 29262 37938 29314 37950
rect 29262 37874 29314 37886
rect 29374 37938 29426 37950
rect 29374 37874 29426 37886
rect 29710 37938 29762 37950
rect 54910 37938 54962 37950
rect 31378 37886 31390 37938
rect 31442 37886 31454 37938
rect 37874 37886 37886 37938
rect 37938 37886 37950 37938
rect 58034 37886 58046 37938
rect 58098 37886 58110 37938
rect 29710 37874 29762 37886
rect 54910 37874 54962 37886
rect 6750 37826 6802 37838
rect 6750 37762 6802 37774
rect 7646 37826 7698 37838
rect 7646 37762 7698 37774
rect 8766 37826 8818 37838
rect 8766 37762 8818 37774
rect 11902 37826 11954 37838
rect 11902 37762 11954 37774
rect 22766 37826 22818 37838
rect 22766 37762 22818 37774
rect 23102 37826 23154 37838
rect 23102 37762 23154 37774
rect 23326 37826 23378 37838
rect 23326 37762 23378 37774
rect 23550 37826 23602 37838
rect 23550 37762 23602 37774
rect 23774 37826 23826 37838
rect 23774 37762 23826 37774
rect 23998 37826 24050 37838
rect 23998 37762 24050 37774
rect 29038 37826 29090 37838
rect 29038 37762 29090 37774
rect 29822 37826 29874 37838
rect 35298 37774 35310 37826
rect 35362 37774 35374 37826
rect 35970 37774 35982 37826
rect 36034 37774 36046 37826
rect 54450 37774 54462 37826
rect 54514 37774 54526 37826
rect 29822 37762 29874 37774
rect 1344 37658 58576 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 58576 37658
rect 1344 37572 58576 37606
rect 5518 37490 5570 37502
rect 5518 37426 5570 37438
rect 5742 37490 5794 37502
rect 32062 37490 32114 37502
rect 7186 37438 7198 37490
rect 7250 37438 7262 37490
rect 5742 37426 5794 37438
rect 29038 37434 29090 37446
rect 4958 37378 5010 37390
rect 4958 37314 5010 37326
rect 15710 37378 15762 37390
rect 15710 37314 15762 37326
rect 18958 37378 19010 37390
rect 18958 37314 19010 37326
rect 20750 37378 20802 37390
rect 20750 37314 20802 37326
rect 22878 37378 22930 37390
rect 22878 37314 22930 37326
rect 22990 37378 23042 37390
rect 22990 37314 23042 37326
rect 28926 37378 28978 37390
rect 32062 37426 32114 37438
rect 35982 37490 36034 37502
rect 35982 37426 36034 37438
rect 36094 37490 36146 37502
rect 36094 37426 36146 37438
rect 36990 37490 37042 37502
rect 36990 37426 37042 37438
rect 37550 37490 37602 37502
rect 37550 37426 37602 37438
rect 48862 37490 48914 37502
rect 48862 37426 48914 37438
rect 29038 37370 29090 37382
rect 36542 37378 36594 37390
rect 48750 37378 48802 37390
rect 28926 37314 28978 37326
rect 45602 37326 45614 37378
rect 45666 37326 45678 37378
rect 36542 37314 36594 37326
rect 48750 37314 48802 37326
rect 49310 37378 49362 37390
rect 49310 37314 49362 37326
rect 4734 37266 4786 37278
rect 4734 37202 4786 37214
rect 5070 37266 5122 37278
rect 5070 37202 5122 37214
rect 5406 37266 5458 37278
rect 5406 37202 5458 37214
rect 7534 37266 7586 37278
rect 7534 37202 7586 37214
rect 8318 37266 8370 37278
rect 8318 37202 8370 37214
rect 8542 37266 8594 37278
rect 16046 37266 16098 37278
rect 19742 37266 19794 37278
rect 11666 37214 11678 37266
rect 11730 37214 11742 37266
rect 12562 37214 12574 37266
rect 12626 37214 12638 37266
rect 19506 37214 19518 37266
rect 19570 37214 19582 37266
rect 8542 37202 8594 37214
rect 16046 37202 16098 37214
rect 19742 37202 19794 37214
rect 22542 37266 22594 37278
rect 22542 37202 22594 37214
rect 23214 37266 23266 37278
rect 23214 37202 23266 37214
rect 23438 37266 23490 37278
rect 23438 37202 23490 37214
rect 23662 37266 23714 37278
rect 23662 37202 23714 37214
rect 24110 37266 24162 37278
rect 24110 37202 24162 37214
rect 28702 37266 28754 37278
rect 28702 37202 28754 37214
rect 29486 37266 29538 37278
rect 29486 37202 29538 37214
rect 31614 37266 31666 37278
rect 31614 37202 31666 37214
rect 31950 37266 32002 37278
rect 31950 37202 32002 37214
rect 32286 37266 32338 37278
rect 32286 37202 32338 37214
rect 35310 37266 35362 37278
rect 35310 37202 35362 37214
rect 35534 37266 35586 37278
rect 35534 37202 35586 37214
rect 36206 37266 36258 37278
rect 36206 37202 36258 37214
rect 36878 37266 36930 37278
rect 36878 37202 36930 37214
rect 37102 37266 37154 37278
rect 37102 37202 37154 37214
rect 42030 37266 42082 37278
rect 42030 37202 42082 37214
rect 42590 37266 42642 37278
rect 48974 37266 49026 37278
rect 44930 37214 44942 37266
rect 44994 37214 45006 37266
rect 56018 37214 56030 37266
rect 56082 37214 56094 37266
rect 42590 37202 42642 37214
rect 48974 37202 49026 37214
rect 12126 37154 12178 37166
rect 20190 37154 20242 37166
rect 13234 37102 13246 37154
rect 13298 37102 13310 37154
rect 15362 37102 15374 37154
rect 15426 37102 15438 37154
rect 12126 37090 12178 37102
rect 20190 37090 20242 37102
rect 23550 37154 23602 37166
rect 23550 37090 23602 37102
rect 28254 37154 28306 37166
rect 28254 37090 28306 37102
rect 30158 37154 30210 37166
rect 30158 37090 30210 37102
rect 31278 37154 31330 37166
rect 31278 37090 31330 37102
rect 33182 37154 33234 37166
rect 38670 37154 38722 37166
rect 38322 37102 38334 37154
rect 38386 37102 38398 37154
rect 33182 37090 33234 37102
rect 38670 37090 38722 37102
rect 43038 37154 43090 37166
rect 48190 37154 48242 37166
rect 47730 37102 47742 37154
rect 47794 37102 47806 37154
rect 43038 37090 43090 37102
rect 48190 37090 48242 37102
rect 49758 37154 49810 37166
rect 56590 37154 56642 37166
rect 53106 37102 53118 37154
rect 53170 37102 53182 37154
rect 55234 37102 55246 37154
rect 55298 37102 55310 37154
rect 49758 37090 49810 37102
rect 56590 37090 56642 37102
rect 56702 37154 56754 37166
rect 56702 37090 56754 37102
rect 58158 37154 58210 37166
rect 58158 37090 58210 37102
rect 7982 37042 8034 37054
rect 7982 36978 8034 36990
rect 8094 37042 8146 37054
rect 8094 36978 8146 36990
rect 8654 37042 8706 37054
rect 8654 36978 8706 36990
rect 49646 37042 49698 37054
rect 57810 36990 57822 37042
rect 57874 37039 57886 37042
rect 58146 37039 58158 37042
rect 57874 36993 58158 37039
rect 57874 36990 57886 36993
rect 58146 36990 58158 36993
rect 58210 36990 58222 37042
rect 49646 36978 49698 36990
rect 1344 36874 58576 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 58576 36874
rect 1344 36788 58576 36822
rect 12350 36594 12402 36606
rect 43374 36594 43426 36606
rect 4610 36542 4622 36594
rect 4674 36542 4686 36594
rect 16370 36542 16382 36594
rect 16434 36542 16446 36594
rect 27122 36542 27134 36594
rect 27186 36542 27198 36594
rect 12350 36530 12402 36542
rect 43374 36530 43426 36542
rect 44830 36594 44882 36606
rect 52110 36594 52162 36606
rect 45938 36542 45950 36594
rect 46002 36542 46014 36594
rect 49410 36542 49422 36594
rect 49474 36542 49486 36594
rect 51538 36542 51550 36594
rect 51602 36542 51614 36594
rect 52770 36542 52782 36594
rect 52834 36542 52846 36594
rect 54338 36542 54350 36594
rect 54402 36542 54414 36594
rect 58146 36542 58158 36594
rect 58210 36542 58222 36594
rect 44830 36530 44882 36542
rect 52110 36530 52162 36542
rect 13582 36482 13634 36494
rect 1810 36430 1822 36482
rect 1874 36430 1886 36482
rect 13582 36418 13634 36430
rect 13694 36482 13746 36494
rect 13694 36418 13746 36430
rect 14142 36482 14194 36494
rect 14142 36418 14194 36430
rect 16606 36482 16658 36494
rect 20526 36482 20578 36494
rect 27358 36482 27410 36494
rect 16706 36430 16718 36482
rect 16770 36430 16782 36482
rect 20066 36430 20078 36482
rect 20130 36430 20142 36482
rect 24210 36430 24222 36482
rect 24274 36430 24286 36482
rect 16606 36418 16658 36430
rect 20526 36418 20578 36430
rect 27358 36418 27410 36430
rect 28030 36482 28082 36494
rect 28030 36418 28082 36430
rect 31950 36482 32002 36494
rect 31950 36418 32002 36430
rect 32398 36482 32450 36494
rect 32398 36418 32450 36430
rect 32622 36482 32674 36494
rect 32622 36418 32674 36430
rect 33518 36482 33570 36494
rect 33518 36418 33570 36430
rect 35198 36482 35250 36494
rect 35198 36418 35250 36430
rect 35870 36482 35922 36494
rect 35870 36418 35922 36430
rect 36318 36482 36370 36494
rect 41582 36482 41634 36494
rect 38322 36430 38334 36482
rect 38386 36430 38398 36482
rect 36318 36418 36370 36430
rect 41582 36418 41634 36430
rect 42478 36482 42530 36494
rect 53902 36482 53954 36494
rect 43810 36430 43822 36482
rect 43874 36430 43886 36482
rect 45266 36430 45278 36482
rect 45330 36430 45342 36482
rect 46274 36430 46286 36482
rect 46338 36430 46350 36482
rect 48738 36430 48750 36482
rect 48802 36430 48814 36482
rect 55346 36430 55358 36482
rect 55410 36430 55422 36482
rect 42478 36418 42530 36430
rect 53902 36418 53954 36430
rect 5742 36370 5794 36382
rect 2482 36318 2494 36370
rect 2546 36318 2558 36370
rect 5742 36306 5794 36318
rect 5854 36370 5906 36382
rect 27806 36370 27858 36382
rect 24994 36318 25006 36370
rect 25058 36318 25070 36370
rect 5854 36306 5906 36318
rect 27806 36306 27858 36318
rect 35646 36370 35698 36382
rect 35646 36306 35698 36318
rect 37998 36370 38050 36382
rect 37998 36306 38050 36318
rect 46846 36370 46898 36382
rect 46846 36306 46898 36318
rect 52782 36370 52834 36382
rect 52782 36306 52834 36318
rect 53342 36370 53394 36382
rect 53342 36306 53394 36318
rect 54910 36370 54962 36382
rect 56018 36318 56030 36370
rect 56082 36318 56094 36370
rect 54910 36306 54962 36318
rect 5518 36258 5570 36270
rect 5518 36194 5570 36206
rect 13806 36258 13858 36270
rect 15710 36258 15762 36270
rect 15362 36206 15374 36258
rect 15426 36206 15438 36258
rect 13806 36194 13858 36206
rect 15710 36194 15762 36206
rect 17502 36258 17554 36270
rect 17502 36194 17554 36206
rect 21422 36258 21474 36270
rect 21422 36194 21474 36206
rect 27582 36258 27634 36270
rect 27582 36194 27634 36206
rect 28478 36258 28530 36270
rect 28478 36194 28530 36206
rect 31838 36258 31890 36270
rect 31838 36194 31890 36206
rect 32510 36258 32562 36270
rect 32510 36194 32562 36206
rect 33070 36258 33122 36270
rect 33070 36194 33122 36206
rect 33294 36258 33346 36270
rect 33294 36194 33346 36206
rect 33406 36258 33458 36270
rect 33406 36194 33458 36206
rect 33966 36258 34018 36270
rect 33966 36194 34018 36206
rect 34974 36258 35026 36270
rect 34974 36194 35026 36206
rect 35758 36258 35810 36270
rect 35758 36194 35810 36206
rect 38110 36258 38162 36270
rect 38110 36194 38162 36206
rect 39230 36258 39282 36270
rect 39230 36194 39282 36206
rect 42142 36258 42194 36270
rect 42142 36194 42194 36206
rect 43038 36258 43090 36270
rect 43038 36194 43090 36206
rect 51998 36258 52050 36270
rect 51998 36194 52050 36206
rect 52894 36258 52946 36270
rect 52894 36194 52946 36206
rect 53118 36258 53170 36270
rect 53118 36194 53170 36206
rect 54014 36258 54066 36270
rect 54014 36194 54066 36206
rect 54238 36258 54290 36270
rect 54238 36194 54290 36206
rect 54350 36258 54402 36270
rect 54350 36194 54402 36206
rect 1344 36090 58576 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 58576 36090
rect 1344 36004 58576 36038
rect 4510 35922 4562 35934
rect 4510 35858 4562 35870
rect 8318 35922 8370 35934
rect 8318 35858 8370 35870
rect 8542 35922 8594 35934
rect 8542 35858 8594 35870
rect 10558 35922 10610 35934
rect 10558 35858 10610 35870
rect 13358 35922 13410 35934
rect 13358 35858 13410 35870
rect 13694 35922 13746 35934
rect 13694 35858 13746 35870
rect 13806 35922 13858 35934
rect 13806 35858 13858 35870
rect 14254 35922 14306 35934
rect 14254 35858 14306 35870
rect 15374 35922 15426 35934
rect 26126 35922 26178 35934
rect 22866 35870 22878 35922
rect 22930 35870 22942 35922
rect 15374 35858 15426 35870
rect 26126 35858 26178 35870
rect 28702 35922 28754 35934
rect 33182 35922 33234 35934
rect 44158 35922 44210 35934
rect 54910 35922 54962 35934
rect 29026 35870 29038 35922
rect 29090 35870 29102 35922
rect 40226 35870 40238 35922
rect 40290 35870 40302 35922
rect 47170 35870 47182 35922
rect 47234 35870 47246 35922
rect 28702 35858 28754 35870
rect 33182 35858 33234 35870
rect 44158 35858 44210 35870
rect 54910 35858 54962 35870
rect 55582 35922 55634 35934
rect 55582 35858 55634 35870
rect 4734 35810 4786 35822
rect 4734 35746 4786 35758
rect 6078 35810 6130 35822
rect 6078 35746 6130 35758
rect 7758 35810 7810 35822
rect 7758 35746 7810 35758
rect 7870 35810 7922 35822
rect 7870 35746 7922 35758
rect 8206 35810 8258 35822
rect 8206 35746 8258 35758
rect 8878 35810 8930 35822
rect 8878 35746 8930 35758
rect 10110 35810 10162 35822
rect 10110 35746 10162 35758
rect 15150 35810 15202 35822
rect 15150 35746 15202 35758
rect 16270 35810 16322 35822
rect 26574 35810 26626 35822
rect 30046 35810 30098 35822
rect 20626 35758 20638 35810
rect 20690 35758 20702 35810
rect 27682 35758 27694 35810
rect 27746 35758 27758 35810
rect 16270 35746 16322 35758
rect 26574 35746 26626 35758
rect 30046 35746 30098 35758
rect 32510 35810 32562 35822
rect 32510 35746 32562 35758
rect 35870 35810 35922 35822
rect 55134 35810 55186 35822
rect 41794 35758 41806 35810
rect 41858 35758 41870 35810
rect 47842 35758 47854 35810
rect 47906 35758 47918 35810
rect 48962 35758 48974 35810
rect 49026 35758 49038 35810
rect 35870 35746 35922 35758
rect 55134 35746 55186 35758
rect 4286 35698 4338 35710
rect 4286 35634 4338 35646
rect 4958 35698 5010 35710
rect 5518 35698 5570 35710
rect 5282 35646 5294 35698
rect 5346 35646 5358 35698
rect 4958 35634 5010 35646
rect 5518 35634 5570 35646
rect 5742 35698 5794 35710
rect 5742 35634 5794 35646
rect 8766 35698 8818 35710
rect 8766 35634 8818 35646
rect 9102 35698 9154 35710
rect 9102 35634 9154 35646
rect 9438 35698 9490 35710
rect 9438 35634 9490 35646
rect 9886 35698 9938 35710
rect 9886 35634 9938 35646
rect 13582 35698 13634 35710
rect 13582 35634 13634 35646
rect 15374 35698 15426 35710
rect 15374 35634 15426 35646
rect 15710 35698 15762 35710
rect 15710 35634 15762 35646
rect 16158 35698 16210 35710
rect 16158 35634 16210 35646
rect 16382 35698 16434 35710
rect 26014 35698 26066 35710
rect 19954 35646 19966 35698
rect 20018 35646 20030 35698
rect 16382 35634 16434 35646
rect 26014 35634 26066 35646
rect 26350 35698 26402 35710
rect 26350 35634 26402 35646
rect 28030 35698 28082 35710
rect 28030 35634 28082 35646
rect 28366 35698 28418 35710
rect 28366 35634 28418 35646
rect 31950 35698 32002 35710
rect 31950 35634 32002 35646
rect 32174 35698 32226 35710
rect 32174 35634 32226 35646
rect 36206 35698 36258 35710
rect 36206 35634 36258 35646
rect 36430 35698 36482 35710
rect 38558 35698 38610 35710
rect 38210 35646 38222 35698
rect 38274 35646 38286 35698
rect 36430 35634 36482 35646
rect 38558 35634 38610 35646
rect 39006 35698 39058 35710
rect 39678 35698 39730 35710
rect 39442 35646 39454 35698
rect 39506 35646 39518 35698
rect 39006 35634 39058 35646
rect 39678 35634 39730 35646
rect 39790 35698 39842 35710
rect 39790 35634 39842 35646
rect 42142 35698 42194 35710
rect 42142 35634 42194 35646
rect 46846 35698 46898 35710
rect 46846 35634 46898 35646
rect 47518 35698 47570 35710
rect 54686 35698 54738 35710
rect 52882 35646 52894 35698
rect 52946 35646 52958 35698
rect 54450 35646 54462 35698
rect 54514 35646 54526 35698
rect 47518 35634 47570 35646
rect 54686 35634 54738 35646
rect 56030 35698 56082 35710
rect 56030 35634 56082 35646
rect 5966 35586 6018 35598
rect 5966 35522 6018 35534
rect 9662 35586 9714 35598
rect 9662 35522 9714 35534
rect 27022 35586 27074 35598
rect 27022 35522 27074 35534
rect 29598 35586 29650 35598
rect 29598 35522 29650 35534
rect 32062 35586 32114 35598
rect 32062 35522 32114 35534
rect 36318 35586 36370 35598
rect 36318 35522 36370 35534
rect 42590 35586 42642 35598
rect 42590 35522 42642 35534
rect 43262 35586 43314 35598
rect 43262 35522 43314 35534
rect 45614 35586 45666 35598
rect 45614 35522 45666 35534
rect 54798 35586 54850 35598
rect 54798 35522 54850 35534
rect 55470 35586 55522 35598
rect 55470 35522 55522 35534
rect 56702 35586 56754 35598
rect 56702 35522 56754 35534
rect 7758 35474 7810 35486
rect 29374 35474 29426 35486
rect 38894 35474 38946 35486
rect 16818 35422 16830 35474
rect 16882 35422 16894 35474
rect 37874 35422 37886 35474
rect 37938 35422 37950 35474
rect 7758 35410 7810 35422
rect 29374 35410 29426 35422
rect 38894 35410 38946 35422
rect 1344 35306 58576 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 58576 35306
rect 1344 35220 58576 35254
rect 28366 35138 28418 35150
rect 28018 35086 28030 35138
rect 28082 35086 28094 35138
rect 28366 35074 28418 35086
rect 41246 35138 41298 35150
rect 41246 35074 41298 35086
rect 41582 35138 41634 35150
rect 41582 35074 41634 35086
rect 40462 35026 40514 35038
rect 8418 34974 8430 35026
rect 8482 34974 8494 35026
rect 10546 34974 10558 35026
rect 10610 34974 10622 35026
rect 16482 34974 16494 35026
rect 16546 34974 16558 35026
rect 30482 34974 30494 35026
rect 30546 34974 30558 35026
rect 37762 34974 37774 35026
rect 37826 34974 37838 35026
rect 39890 34974 39902 35026
rect 39954 34974 39966 35026
rect 49746 34974 49758 35026
rect 49810 34974 49822 35026
rect 40462 34962 40514 34974
rect 5182 34914 5234 34926
rect 5182 34850 5234 34862
rect 5854 34914 5906 34926
rect 5854 34850 5906 34862
rect 6078 34914 6130 34926
rect 19182 34914 19234 34926
rect 11330 34862 11342 34914
rect 11394 34862 11406 34914
rect 17378 34862 17390 34914
rect 17442 34862 17454 34914
rect 6078 34850 6130 34862
rect 19182 34850 19234 34862
rect 25678 34914 25730 34926
rect 25678 34850 25730 34862
rect 26014 34914 26066 34926
rect 26014 34850 26066 34862
rect 28590 34914 28642 34926
rect 33070 34914 33122 34926
rect 29698 34862 29710 34914
rect 29762 34862 29774 34914
rect 28590 34850 28642 34862
rect 33070 34850 33122 34862
rect 33630 34914 33682 34926
rect 33630 34850 33682 34862
rect 34638 34914 34690 34926
rect 34638 34850 34690 34862
rect 34750 34914 34802 34926
rect 42142 34914 42194 34926
rect 37090 34862 37102 34914
rect 37154 34862 37166 34914
rect 41906 34862 41918 34914
rect 41970 34862 41982 34914
rect 34750 34850 34802 34862
rect 42142 34850 42194 34862
rect 43262 34914 43314 34926
rect 43262 34850 43314 34862
rect 49646 34914 49698 34926
rect 49646 34850 49698 34862
rect 49982 34914 50034 34926
rect 52110 34914 52162 34926
rect 50194 34862 50206 34914
rect 50258 34862 50270 34914
rect 52882 34862 52894 34914
rect 52946 34862 52958 34914
rect 49982 34850 50034 34862
rect 52110 34850 52162 34862
rect 4286 34802 4338 34814
rect 4286 34738 4338 34750
rect 4622 34802 4674 34814
rect 4622 34738 4674 34750
rect 4846 34802 4898 34814
rect 4846 34738 4898 34750
rect 4958 34802 5010 34814
rect 4958 34738 5010 34750
rect 5630 34802 5682 34814
rect 5630 34738 5682 34750
rect 33518 34802 33570 34814
rect 33518 34738 33570 34750
rect 42366 34802 42418 34814
rect 42366 34738 42418 34750
rect 42590 34802 42642 34814
rect 42590 34738 42642 34750
rect 43150 34802 43202 34814
rect 55458 34750 55470 34802
rect 55522 34750 55534 34802
rect 43150 34738 43202 34750
rect 4398 34690 4450 34702
rect 4398 34626 4450 34638
rect 5742 34690 5794 34702
rect 5742 34626 5794 34638
rect 25790 34690 25842 34702
rect 25790 34626 25842 34638
rect 26462 34690 26514 34702
rect 26462 34626 26514 34638
rect 27246 34690 27298 34702
rect 33294 34690 33346 34702
rect 32722 34638 32734 34690
rect 32786 34638 32798 34690
rect 27246 34626 27298 34638
rect 33294 34626 33346 34638
rect 35086 34690 35138 34702
rect 35086 34626 35138 34638
rect 40910 34690 40962 34702
rect 40910 34626 40962 34638
rect 41470 34690 41522 34702
rect 41470 34626 41522 34638
rect 42254 34690 42306 34702
rect 42254 34626 42306 34638
rect 48414 34690 48466 34702
rect 48414 34626 48466 34638
rect 49198 34690 49250 34702
rect 49198 34626 49250 34638
rect 49758 34690 49810 34702
rect 49758 34626 49810 34638
rect 1344 34522 58576 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 58576 34522
rect 1344 34436 58576 34470
rect 16382 34354 16434 34366
rect 8530 34302 8542 34354
rect 8594 34302 8606 34354
rect 16382 34290 16434 34302
rect 33630 34354 33682 34366
rect 39342 34354 39394 34366
rect 34626 34302 34638 34354
rect 34690 34302 34702 34354
rect 36082 34302 36094 34354
rect 36146 34302 36158 34354
rect 41794 34302 41806 34354
rect 41858 34302 41870 34354
rect 33630 34290 33682 34302
rect 39342 34290 39394 34302
rect 11342 34242 11394 34254
rect 33182 34242 33234 34254
rect 27906 34190 27918 34242
rect 27970 34190 27982 34242
rect 11342 34178 11394 34190
rect 33182 34178 33234 34190
rect 34078 34242 34130 34254
rect 38222 34242 38274 34254
rect 35186 34190 35198 34242
rect 35250 34190 35262 34242
rect 34078 34178 34130 34190
rect 38222 34178 38274 34190
rect 39566 34242 39618 34254
rect 46398 34242 46450 34254
rect 43922 34190 43934 34242
rect 43986 34190 43998 34242
rect 51986 34190 51998 34242
rect 52050 34190 52062 34242
rect 39566 34178 39618 34190
rect 46398 34178 46450 34190
rect 9662 34130 9714 34142
rect 16270 34130 16322 34142
rect 26686 34130 26738 34142
rect 8194 34078 8206 34130
rect 8258 34078 8270 34130
rect 8754 34078 8766 34130
rect 8818 34078 8830 34130
rect 11106 34078 11118 34130
rect 11170 34078 11182 34130
rect 11778 34078 11790 34130
rect 11842 34078 11854 34130
rect 19506 34078 19518 34130
rect 19570 34078 19582 34130
rect 20290 34078 20302 34130
rect 20354 34078 20366 34130
rect 21858 34078 21870 34130
rect 21922 34078 21934 34130
rect 9662 34066 9714 34078
rect 16270 34066 16322 34078
rect 26686 34066 26738 34078
rect 27582 34130 27634 34142
rect 35074 34078 35086 34130
rect 35138 34078 35150 34130
rect 38882 34078 38894 34130
rect 38946 34078 38958 34130
rect 41570 34078 41582 34130
rect 41634 34078 41646 34130
rect 43250 34078 43262 34130
rect 43314 34078 43326 34130
rect 47618 34078 47630 34130
rect 47682 34078 47694 34130
rect 51202 34078 51214 34130
rect 51266 34078 51278 34130
rect 27582 34066 27634 34078
rect 15710 34018 15762 34030
rect 27246 34018 27298 34030
rect 4946 33966 4958 34018
rect 5010 33966 5022 34018
rect 12450 33966 12462 34018
rect 12514 33966 12526 34018
rect 14578 33966 14590 34018
rect 14642 33966 14654 34018
rect 17378 33966 17390 34018
rect 17442 33966 17454 34018
rect 22530 33966 22542 34018
rect 22594 33966 22606 34018
rect 24658 33966 24670 34018
rect 24722 33966 24734 34018
rect 15710 33954 15762 33966
rect 27246 33954 27298 33966
rect 28366 34018 28418 34030
rect 28366 33954 28418 33966
rect 33742 34018 33794 34030
rect 47294 34018 47346 34030
rect 54574 34018 54626 34030
rect 46050 33966 46062 34018
rect 46114 33966 46126 34018
rect 54114 33966 54126 34018
rect 54178 33966 54190 34018
rect 33742 33954 33794 33966
rect 47294 33954 47346 33966
rect 54574 33954 54626 33966
rect 16046 33906 16098 33918
rect 16046 33842 16098 33854
rect 16382 33906 16434 33918
rect 16382 33842 16434 33854
rect 33294 33906 33346 33918
rect 33294 33842 33346 33854
rect 34302 33906 34354 33918
rect 34302 33842 34354 33854
rect 39230 33906 39282 33918
rect 39230 33842 39282 33854
rect 46510 33906 46562 33918
rect 46510 33842 46562 33854
rect 47630 33906 47682 33918
rect 47630 33842 47682 33854
rect 47966 33906 48018 33918
rect 47966 33842 48018 33854
rect 1344 33738 58576 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 58576 33738
rect 1344 33652 58576 33686
rect 12350 33570 12402 33582
rect 12350 33506 12402 33518
rect 35758 33570 35810 33582
rect 35758 33506 35810 33518
rect 37774 33570 37826 33582
rect 37774 33506 37826 33518
rect 38670 33570 38722 33582
rect 38994 33518 39006 33570
rect 39058 33518 39070 33570
rect 38670 33506 38722 33518
rect 11678 33458 11730 33470
rect 2482 33406 2494 33458
rect 2546 33406 2558 33458
rect 4610 33406 4622 33458
rect 4674 33406 4686 33458
rect 9874 33406 9886 33458
rect 9938 33406 9950 33458
rect 11678 33394 11730 33406
rect 12462 33458 12514 33470
rect 12462 33394 12514 33406
rect 20862 33458 20914 33470
rect 50766 33458 50818 33470
rect 21858 33406 21870 33458
rect 21922 33406 21934 33458
rect 36082 33406 36094 33458
rect 36146 33406 36158 33458
rect 41906 33406 41918 33458
rect 41970 33406 41982 33458
rect 47394 33406 47406 33458
rect 47458 33406 47470 33458
rect 49522 33406 49534 33458
rect 49586 33406 49598 33458
rect 54786 33406 54798 33458
rect 54850 33406 54862 33458
rect 56018 33406 56030 33458
rect 56082 33406 56094 33458
rect 58146 33406 58158 33458
rect 58210 33406 58222 33458
rect 20862 33394 20914 33406
rect 50766 33394 50818 33406
rect 6414 33346 6466 33358
rect 29710 33346 29762 33358
rect 37550 33346 37602 33358
rect 1810 33294 1822 33346
rect 1874 33294 1886 33346
rect 6962 33294 6974 33346
rect 7026 33294 7038 33346
rect 12674 33294 12686 33346
rect 12738 33294 12750 33346
rect 25218 33294 25230 33346
rect 25282 33294 25294 33346
rect 27458 33294 27470 33346
rect 27522 33294 27534 33346
rect 29922 33294 29934 33346
rect 29986 33294 29998 33346
rect 6414 33282 6466 33294
rect 29710 33282 29762 33294
rect 37550 33282 37602 33294
rect 38446 33346 38498 33358
rect 42030 33346 42082 33358
rect 41794 33294 41806 33346
rect 41858 33294 41870 33346
rect 38446 33282 38498 33294
rect 42030 33282 42082 33294
rect 42254 33346 42306 33358
rect 42254 33282 42306 33294
rect 42926 33346 42978 33358
rect 53006 33346 53058 33358
rect 46610 33294 46622 33346
rect 46674 33294 46686 33346
rect 51874 33294 51886 33346
rect 51938 33294 51950 33346
rect 42926 33282 42978 33294
rect 53006 33282 53058 33294
rect 53342 33346 53394 33358
rect 53554 33294 53566 33346
rect 53618 33294 53630 33346
rect 54898 33294 54910 33346
rect 54962 33294 54974 33346
rect 55346 33294 55358 33346
rect 55410 33294 55422 33346
rect 53342 33282 53394 33294
rect 16606 33234 16658 33246
rect 7746 33182 7758 33234
rect 7810 33182 7822 33234
rect 16606 33170 16658 33182
rect 20302 33234 20354 33246
rect 35982 33234 36034 33246
rect 27682 33182 27694 33234
rect 27746 33182 27758 33234
rect 31938 33182 31950 33234
rect 32002 33182 32014 33234
rect 20302 33170 20354 33182
rect 35982 33170 36034 33182
rect 42478 33234 42530 33246
rect 42478 33170 42530 33182
rect 49982 33234 50034 33246
rect 49982 33170 50034 33182
rect 50318 33234 50370 33246
rect 50318 33170 50370 33182
rect 52670 33234 52722 33246
rect 52670 33170 52722 33182
rect 52782 33234 52834 33246
rect 52782 33170 52834 33182
rect 54238 33234 54290 33246
rect 54238 33170 54290 33182
rect 54574 33234 54626 33246
rect 54574 33170 54626 33182
rect 16382 33122 16434 33134
rect 6066 33070 6078 33122
rect 6130 33070 6142 33122
rect 16382 33058 16434 33070
rect 16494 33122 16546 33134
rect 16494 33058 16546 33070
rect 20190 33122 20242 33134
rect 20190 33058 20242 33070
rect 28254 33122 28306 33134
rect 50878 33122 50930 33134
rect 38098 33070 38110 33122
rect 38162 33070 38174 33122
rect 52098 33070 52110 33122
rect 52162 33070 52174 33122
rect 28254 33058 28306 33070
rect 50878 33058 50930 33070
rect 1344 32954 58576 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 58576 32954
rect 1344 32868 58576 32902
rect 5742 32786 5794 32798
rect 5742 32722 5794 32734
rect 5966 32786 6018 32798
rect 22430 32786 22482 32798
rect 17378 32734 17390 32786
rect 17442 32734 17454 32786
rect 5966 32722 6018 32734
rect 22430 32722 22482 32734
rect 22654 32786 22706 32798
rect 22654 32722 22706 32734
rect 23326 32786 23378 32798
rect 23326 32722 23378 32734
rect 23550 32786 23602 32798
rect 23550 32722 23602 32734
rect 25230 32786 25282 32798
rect 25230 32722 25282 32734
rect 31166 32786 31218 32798
rect 31166 32722 31218 32734
rect 31838 32786 31890 32798
rect 31838 32722 31890 32734
rect 34190 32786 34242 32798
rect 34190 32722 34242 32734
rect 50766 32786 50818 32798
rect 50766 32722 50818 32734
rect 50878 32786 50930 32798
rect 50878 32722 50930 32734
rect 51774 32786 51826 32798
rect 51774 32722 51826 32734
rect 54014 32786 54066 32798
rect 54014 32722 54066 32734
rect 54238 32786 54290 32798
rect 54238 32722 54290 32734
rect 57374 32786 57426 32798
rect 57374 32722 57426 32734
rect 58158 32786 58210 32798
rect 58158 32722 58210 32734
rect 5294 32674 5346 32686
rect 22318 32674 22370 32686
rect 14690 32622 14702 32674
rect 14754 32622 14766 32674
rect 19618 32622 19630 32674
rect 19682 32622 19694 32674
rect 5294 32610 5346 32622
rect 22318 32610 22370 32622
rect 24446 32674 24498 32686
rect 24446 32610 24498 32622
rect 25678 32674 25730 32686
rect 25678 32610 25730 32622
rect 30942 32674 30994 32686
rect 30942 32610 30994 32622
rect 34638 32674 34690 32686
rect 34638 32610 34690 32622
rect 41358 32674 41410 32686
rect 41358 32610 41410 32622
rect 48190 32674 48242 32686
rect 48190 32610 48242 32622
rect 49198 32674 49250 32686
rect 49198 32610 49250 32622
rect 50318 32674 50370 32686
rect 50318 32610 50370 32622
rect 51998 32674 52050 32686
rect 51998 32610 52050 32622
rect 52670 32674 52722 32686
rect 52670 32610 52722 32622
rect 4846 32562 4898 32574
rect 1810 32510 1822 32562
rect 1874 32510 1886 32562
rect 4846 32498 4898 32510
rect 5518 32562 5570 32574
rect 5518 32498 5570 32510
rect 6078 32562 6130 32574
rect 17726 32562 17778 32574
rect 22542 32562 22594 32574
rect 13906 32510 13918 32562
rect 13970 32510 13982 32562
rect 18946 32510 18958 32562
rect 19010 32510 19022 32562
rect 22082 32510 22094 32562
rect 22146 32510 22158 32562
rect 6078 32498 6130 32510
rect 17726 32498 17778 32510
rect 22542 32498 22594 32510
rect 24110 32562 24162 32574
rect 24110 32498 24162 32510
rect 24222 32562 24274 32574
rect 25454 32562 25506 32574
rect 31278 32562 31330 32574
rect 24658 32510 24670 32562
rect 24722 32510 24734 32562
rect 27570 32510 27582 32562
rect 27634 32510 27646 32562
rect 30706 32510 30718 32562
rect 30770 32510 30782 32562
rect 24222 32498 24274 32510
rect 25454 32498 25506 32510
rect 31278 32498 31330 32510
rect 33854 32562 33906 32574
rect 49086 32562 49138 32574
rect 34066 32510 34078 32562
rect 34130 32510 34142 32562
rect 41794 32510 41806 32562
rect 41858 32510 41870 32562
rect 47730 32510 47742 32562
rect 47794 32510 47806 32562
rect 33854 32498 33906 32510
rect 49086 32498 49138 32510
rect 49758 32562 49810 32574
rect 49758 32498 49810 32510
rect 50542 32562 50594 32574
rect 50542 32498 50594 32510
rect 51662 32562 51714 32574
rect 52558 32562 52610 32574
rect 52210 32510 52222 32562
rect 52274 32510 52286 32562
rect 51662 32498 51714 32510
rect 52558 32498 52610 32510
rect 53118 32562 53170 32574
rect 54450 32510 54462 32562
rect 54514 32510 54526 32562
rect 53118 32498 53170 32510
rect 5070 32450 5122 32462
rect 17950 32450 18002 32462
rect 23662 32450 23714 32462
rect 2482 32398 2494 32450
rect 2546 32398 2558 32450
rect 4610 32398 4622 32450
rect 4674 32398 4686 32450
rect 16818 32398 16830 32450
rect 16882 32398 16894 32450
rect 21746 32398 21758 32450
rect 21810 32398 21822 32450
rect 5070 32386 5122 32398
rect 17950 32386 18002 32398
rect 23662 32386 23714 32398
rect 24334 32450 24386 32462
rect 24334 32386 24386 32398
rect 25342 32450 25394 32462
rect 25342 32386 25394 32398
rect 26350 32450 26402 32462
rect 31054 32450 31106 32462
rect 28242 32398 28254 32450
rect 28306 32398 28318 32450
rect 30370 32398 30382 32450
rect 30434 32398 30446 32450
rect 26350 32386 26402 32398
rect 31054 32386 31106 32398
rect 41470 32450 41522 32462
rect 49646 32450 49698 32462
rect 51886 32450 51938 32462
rect 42578 32398 42590 32450
rect 42642 32398 42654 32450
rect 44706 32398 44718 32450
rect 44770 32398 44782 32450
rect 47282 32398 47294 32450
rect 47346 32398 47358 32450
rect 50866 32398 50878 32450
rect 50930 32398 50942 32450
rect 57698 32398 57710 32450
rect 57762 32398 57774 32450
rect 41470 32386 41522 32398
rect 49646 32386 49698 32398
rect 51886 32386 51938 32398
rect 53342 32338 53394 32350
rect 53902 32338 53954 32350
rect 53666 32286 53678 32338
rect 53730 32286 53742 32338
rect 53342 32274 53394 32286
rect 53902 32274 53954 32286
rect 1344 32170 58576 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 58576 32170
rect 1344 32084 58576 32118
rect 4846 32002 4898 32014
rect 37214 32002 37266 32014
rect 35186 31950 35198 32002
rect 35250 31950 35262 32002
rect 4846 31938 4898 31950
rect 37214 31938 37266 31950
rect 7758 31890 7810 31902
rect 16830 31890 16882 31902
rect 29150 31890 29202 31902
rect 9986 31838 9998 31890
rect 10050 31838 10062 31890
rect 24098 31838 24110 31890
rect 24162 31838 24174 31890
rect 26226 31838 26238 31890
rect 26290 31838 26302 31890
rect 7758 31826 7810 31838
rect 16830 31826 16882 31838
rect 29150 31826 29202 31838
rect 29262 31890 29314 31902
rect 36990 31890 37042 31902
rect 52670 31890 52722 31902
rect 32274 31838 32286 31890
rect 32338 31838 32350 31890
rect 34402 31838 34414 31890
rect 34466 31838 34478 31890
rect 35410 31838 35422 31890
rect 35474 31838 35486 31890
rect 41794 31838 41806 31890
rect 41858 31838 41870 31890
rect 47730 31838 47742 31890
rect 47794 31838 47806 31890
rect 29262 31826 29314 31838
rect 36990 31826 37042 31838
rect 52670 31826 52722 31838
rect 54462 31890 54514 31902
rect 58146 31838 58158 31890
rect 58210 31838 58222 31890
rect 54462 31826 54514 31838
rect 4174 31778 4226 31790
rect 4174 31714 4226 31726
rect 7310 31778 7362 31790
rect 8542 31778 8594 31790
rect 22206 31778 22258 31790
rect 8194 31726 8206 31778
rect 8258 31726 8270 31778
rect 12898 31726 12910 31778
rect 12962 31726 12974 31778
rect 7310 31714 7362 31726
rect 8542 31714 8594 31726
rect 22206 31714 22258 31726
rect 22430 31778 22482 31790
rect 22430 31714 22482 31726
rect 22542 31778 22594 31790
rect 44382 31778 44434 31790
rect 48638 31778 48690 31790
rect 23314 31726 23326 31778
rect 23378 31726 23390 31778
rect 31490 31726 31502 31778
rect 31554 31726 31566 31778
rect 35074 31726 35086 31778
rect 35138 31726 35150 31778
rect 35298 31726 35310 31778
rect 35362 31726 35374 31778
rect 43810 31726 43822 31778
rect 43874 31726 43886 31778
rect 44930 31726 44942 31778
rect 44994 31726 45006 31778
rect 22542 31714 22594 31726
rect 44382 31714 44434 31726
rect 48638 31714 48690 31726
rect 48750 31778 48802 31790
rect 48750 31714 48802 31726
rect 53006 31778 53058 31790
rect 54686 31778 54738 31790
rect 53218 31726 53230 31778
rect 53282 31726 53294 31778
rect 54226 31726 54238 31778
rect 54290 31726 54302 31778
rect 55346 31726 55358 31778
rect 55410 31726 55422 31778
rect 53006 31714 53058 31726
rect 54686 31714 54738 31726
rect 4846 31666 4898 31678
rect 4734 31610 4786 31622
rect 4286 31554 4338 31566
rect 4286 31490 4338 31502
rect 4510 31554 4562 31566
rect 4846 31602 4898 31614
rect 7870 31666 7922 31678
rect 7870 31602 7922 31614
rect 8654 31666 8706 31678
rect 16718 31666 16770 31678
rect 12114 31614 12126 31666
rect 12178 31614 12190 31666
rect 8654 31602 8706 31614
rect 16718 31602 16770 31614
rect 20414 31666 20466 31678
rect 20414 31602 20466 31614
rect 21982 31666 22034 31678
rect 21982 31602 22034 31614
rect 22318 31666 22370 31678
rect 48190 31666 48242 31678
rect 53678 31666 53730 31678
rect 30818 31614 30830 31666
rect 30882 31614 30894 31666
rect 45602 31614 45614 31666
rect 45666 31614 45678 31666
rect 49522 31614 49534 31666
rect 49586 31614 49598 31666
rect 52770 31614 52782 31666
rect 52834 31614 52846 31666
rect 22318 31602 22370 31614
rect 48190 31602 48242 31614
rect 53678 31602 53730 31614
rect 54798 31666 54850 31678
rect 56018 31614 56030 31666
rect 56082 31614 56094 31666
rect 54798 31602 54850 31614
rect 4734 31546 4786 31558
rect 5966 31554 6018 31566
rect 5618 31502 5630 31554
rect 5682 31502 5694 31554
rect 4510 31490 4562 31502
rect 5966 31490 6018 31502
rect 7646 31554 7698 31566
rect 7646 31490 7698 31502
rect 8766 31554 8818 31566
rect 8766 31490 8818 31502
rect 16942 31554 16994 31566
rect 16942 31490 16994 31502
rect 17166 31554 17218 31566
rect 17166 31490 17218 31502
rect 20302 31554 20354 31566
rect 20302 31490 20354 31502
rect 31166 31554 31218 31566
rect 48414 31554 48466 31566
rect 37538 31502 37550 31554
rect 37602 31502 37614 31554
rect 31166 31490 31218 31502
rect 48414 31490 48466 31502
rect 48526 31554 48578 31566
rect 48526 31490 48578 31502
rect 49198 31554 49250 31566
rect 49198 31490 49250 31502
rect 1344 31386 58576 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 58576 31386
rect 1344 31300 58576 31334
rect 5966 31218 6018 31230
rect 5966 31154 6018 31166
rect 7758 31218 7810 31230
rect 7758 31154 7810 31166
rect 8206 31218 8258 31230
rect 8206 31154 8258 31166
rect 11230 31218 11282 31230
rect 11230 31154 11282 31166
rect 17390 31218 17442 31230
rect 17390 31154 17442 31166
rect 17838 31218 17890 31230
rect 17838 31154 17890 31166
rect 22990 31218 23042 31230
rect 22990 31154 23042 31166
rect 25678 31218 25730 31230
rect 31726 31218 31778 31230
rect 30706 31166 30718 31218
rect 30770 31166 30782 31218
rect 25678 31154 25730 31166
rect 31726 31154 31778 31166
rect 33182 31218 33234 31230
rect 33182 31154 33234 31166
rect 34750 31218 34802 31230
rect 34750 31154 34802 31166
rect 35534 31218 35586 31230
rect 35534 31154 35586 31166
rect 41358 31218 41410 31230
rect 41358 31154 41410 31166
rect 41582 31218 41634 31230
rect 41582 31154 41634 31166
rect 41694 31218 41746 31230
rect 41694 31154 41746 31166
rect 42366 31218 42418 31230
rect 42366 31154 42418 31166
rect 42590 31218 42642 31230
rect 42590 31154 42642 31166
rect 47518 31218 47570 31230
rect 47518 31154 47570 31166
rect 52894 31218 52946 31230
rect 52894 31154 52946 31166
rect 4510 31106 4562 31118
rect 4510 31042 4562 31054
rect 4734 31106 4786 31118
rect 9550 31106 9602 31118
rect 10558 31106 10610 31118
rect 5618 31054 5630 31106
rect 5682 31054 5694 31106
rect 9874 31054 9886 31106
rect 9938 31054 9950 31106
rect 4734 31042 4786 31054
rect 9550 31042 9602 31054
rect 10558 31042 10610 31054
rect 10782 31106 10834 31118
rect 22430 31106 22482 31118
rect 19730 31054 19742 31106
rect 19794 31054 19806 31106
rect 10782 31042 10834 31054
rect 22430 31042 22482 31054
rect 33854 31106 33906 31118
rect 33854 31042 33906 31054
rect 34862 31106 34914 31118
rect 45502 31106 45554 31118
rect 35970 31054 35982 31106
rect 36034 31054 36046 31106
rect 34862 31042 34914 31054
rect 45502 31042 45554 31054
rect 47406 31106 47458 31118
rect 47406 31042 47458 31054
rect 48750 31106 48802 31118
rect 48750 31042 48802 31054
rect 53342 31106 53394 31118
rect 53342 31042 53394 31054
rect 5182 30994 5234 31006
rect 8542 30994 8594 31006
rect 7522 30942 7534 30994
rect 7586 30942 7598 30994
rect 5182 30930 5234 30942
rect 8542 30930 8594 30942
rect 10446 30994 10498 31006
rect 10446 30930 10498 30942
rect 10894 30994 10946 31006
rect 10894 30930 10946 30942
rect 11230 30994 11282 31006
rect 11230 30930 11282 30942
rect 11454 30994 11506 31006
rect 17614 30994 17666 31006
rect 25342 30994 25394 31006
rect 13010 30942 13022 30994
rect 13074 30942 13086 30994
rect 18946 30942 18958 30994
rect 19010 30942 19022 30994
rect 11454 30930 11506 30942
rect 17614 30930 17666 30942
rect 25342 30930 25394 30942
rect 25790 30994 25842 31006
rect 25790 30930 25842 30942
rect 26014 30994 26066 31006
rect 31054 30994 31106 31006
rect 31950 30994 32002 31006
rect 33742 30994 33794 31006
rect 34526 30994 34578 31006
rect 29474 30942 29486 30994
rect 29538 30942 29550 30994
rect 31490 30942 31502 30994
rect 31554 30942 31566 30994
rect 32162 30942 32174 30994
rect 32226 30942 32238 30994
rect 33506 30942 33518 30994
rect 33570 30942 33582 30994
rect 34290 30942 34302 30994
rect 34354 30942 34366 30994
rect 26014 30930 26066 30942
rect 31054 30930 31106 30942
rect 31950 30930 32002 30942
rect 33742 30930 33794 30942
rect 34526 30930 34578 30942
rect 36318 30994 36370 31006
rect 36318 30930 36370 30942
rect 36542 30994 36594 31006
rect 45838 30994 45890 31006
rect 37426 30942 37438 30994
rect 37490 30942 37502 30994
rect 41122 30942 41134 30994
rect 41186 30942 41198 30994
rect 42130 30942 42142 30994
rect 42194 30942 42206 30994
rect 42802 30942 42814 30994
rect 42866 30942 42878 30994
rect 36542 30930 36594 30942
rect 45838 30930 45890 30942
rect 48974 30994 49026 31006
rect 48974 30930 49026 30942
rect 53006 30994 53058 31006
rect 53006 30930 53058 30942
rect 4958 30882 5010 30894
rect 17502 30882 17554 30894
rect 31838 30882 31890 30894
rect 36990 30882 37042 30894
rect 41470 30882 41522 30894
rect 13794 30830 13806 30882
rect 13858 30830 13870 30882
rect 15922 30830 15934 30882
rect 15986 30830 15998 30882
rect 21858 30830 21870 30882
rect 21922 30830 21934 30882
rect 26562 30830 26574 30882
rect 26626 30830 26638 30882
rect 28690 30830 28702 30882
rect 28754 30830 28766 30882
rect 34850 30830 34862 30882
rect 34914 30830 34926 30882
rect 38210 30830 38222 30882
rect 38274 30830 38286 30882
rect 40338 30830 40350 30882
rect 40402 30830 40414 30882
rect 4958 30818 5010 30830
rect 17502 30818 17554 30830
rect 31838 30818 31890 30830
rect 36990 30818 37042 30830
rect 41470 30818 41522 30830
rect 42478 30882 42530 30894
rect 42478 30818 42530 30830
rect 45614 30882 45666 30894
rect 45614 30818 45666 30830
rect 7870 30770 7922 30782
rect 7870 30706 7922 30718
rect 22542 30770 22594 30782
rect 22542 30706 22594 30718
rect 45950 30770 46002 30782
rect 45950 30706 46002 30718
rect 49310 30770 49362 30782
rect 49310 30706 49362 30718
rect 53454 30770 53506 30782
rect 53454 30706 53506 30718
rect 1344 30602 58576 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 58576 30602
rect 1344 30516 58576 30550
rect 16158 30434 16210 30446
rect 16158 30370 16210 30382
rect 25118 30434 25170 30446
rect 45726 30434 45778 30446
rect 41906 30382 41918 30434
rect 41970 30431 41982 30434
rect 42354 30431 42366 30434
rect 41970 30385 42366 30431
rect 41970 30382 41982 30385
rect 42354 30382 42366 30385
rect 42418 30382 42430 30434
rect 25118 30370 25170 30382
rect 45726 30370 45778 30382
rect 24894 30322 24946 30334
rect 4610 30270 4622 30322
rect 4674 30270 4686 30322
rect 24894 30258 24946 30270
rect 26238 30322 26290 30334
rect 26238 30258 26290 30270
rect 53678 30322 53730 30334
rect 53678 30258 53730 30270
rect 54462 30322 54514 30334
rect 54462 30258 54514 30270
rect 5518 30210 5570 30222
rect 1810 30158 1822 30210
rect 1874 30158 1886 30210
rect 2482 30158 2494 30210
rect 2546 30158 2558 30210
rect 5518 30146 5570 30158
rect 5854 30210 5906 30222
rect 5854 30146 5906 30158
rect 11006 30210 11058 30222
rect 11006 30146 11058 30158
rect 16382 30210 16434 30222
rect 24558 30210 24610 30222
rect 16706 30158 16718 30210
rect 16770 30158 16782 30210
rect 18722 30158 18734 30210
rect 18786 30158 18798 30210
rect 16382 30146 16434 30158
rect 24558 30146 24610 30158
rect 29934 30210 29986 30222
rect 29934 30146 29986 30158
rect 30158 30210 30210 30222
rect 36318 30210 36370 30222
rect 30594 30158 30606 30210
rect 30658 30158 30670 30210
rect 30158 30146 30210 30158
rect 36318 30146 36370 30158
rect 37550 30210 37602 30222
rect 37550 30146 37602 30158
rect 39342 30210 39394 30222
rect 39342 30146 39394 30158
rect 39454 30210 39506 30222
rect 39454 30146 39506 30158
rect 40910 30210 40962 30222
rect 40910 30146 40962 30158
rect 41918 30210 41970 30222
rect 41918 30146 41970 30158
rect 50990 30210 51042 30222
rect 53566 30210 53618 30222
rect 54350 30210 54402 30222
rect 53330 30158 53342 30210
rect 53394 30158 53406 30210
rect 54002 30158 54014 30210
rect 54066 30158 54078 30210
rect 50990 30146 51042 30158
rect 53566 30146 53618 30158
rect 54350 30146 54402 30158
rect 55246 30210 55298 30222
rect 55246 30146 55298 30158
rect 6190 30098 6242 30110
rect 6190 30034 6242 30046
rect 6526 30098 6578 30110
rect 6526 30034 6578 30046
rect 10670 30098 10722 30110
rect 19294 30098 19346 30110
rect 16818 30046 16830 30098
rect 16882 30046 16894 30098
rect 10670 30034 10722 30046
rect 19294 30034 19346 30046
rect 24670 30098 24722 30110
rect 42366 30098 42418 30110
rect 34962 30046 34974 30098
rect 35026 30046 35038 30098
rect 24670 30034 24722 30046
rect 42366 30034 42418 30046
rect 45390 30098 45442 30110
rect 45390 30034 45442 30046
rect 45614 30098 45666 30110
rect 45614 30034 45666 30046
rect 5742 29986 5794 29998
rect 5742 29922 5794 29934
rect 7086 29986 7138 29998
rect 7086 29922 7138 29934
rect 10782 29986 10834 29998
rect 24446 29986 24498 29998
rect 15810 29934 15822 29986
rect 15874 29934 15886 29986
rect 20402 29934 20414 29986
rect 20466 29934 20478 29986
rect 10782 29922 10834 29934
rect 24446 29922 24498 29934
rect 30270 29986 30322 29998
rect 30270 29922 30322 29934
rect 36206 29986 36258 29998
rect 36206 29922 36258 29934
rect 36990 29986 37042 29998
rect 36990 29922 37042 29934
rect 40798 29986 40850 29998
rect 40798 29922 40850 29934
rect 51102 29986 51154 29998
rect 51102 29922 51154 29934
rect 53790 29986 53842 29998
rect 53790 29922 53842 29934
rect 1344 29818 58576 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 58576 29818
rect 1344 29732 58576 29766
rect 11566 29650 11618 29662
rect 5842 29598 5854 29650
rect 5906 29598 5918 29650
rect 8978 29598 8990 29650
rect 9042 29598 9054 29650
rect 11566 29586 11618 29598
rect 16270 29650 16322 29662
rect 19406 29650 19458 29662
rect 19058 29598 19070 29650
rect 19122 29598 19134 29650
rect 16270 29586 16322 29598
rect 19406 29586 19458 29598
rect 19854 29650 19906 29662
rect 19854 29586 19906 29598
rect 27470 29650 27522 29662
rect 27470 29586 27522 29598
rect 33182 29650 33234 29662
rect 33182 29586 33234 29598
rect 37438 29650 37490 29662
rect 37438 29586 37490 29598
rect 37886 29650 37938 29662
rect 37886 29586 37938 29598
rect 47966 29650 48018 29662
rect 47966 29586 48018 29598
rect 49646 29650 49698 29662
rect 49646 29586 49698 29598
rect 51550 29650 51602 29662
rect 51550 29586 51602 29598
rect 51774 29650 51826 29662
rect 51774 29586 51826 29598
rect 55806 29650 55858 29662
rect 55806 29586 55858 29598
rect 11678 29538 11730 29550
rect 4498 29486 4510 29538
rect 4562 29486 4574 29538
rect 5954 29486 5966 29538
rect 6018 29486 6030 29538
rect 11678 29474 11730 29486
rect 16382 29538 16434 29550
rect 16382 29474 16434 29486
rect 26462 29538 26514 29550
rect 44046 29538 44098 29550
rect 50990 29538 51042 29550
rect 30370 29486 30382 29538
rect 30434 29486 30446 29538
rect 35970 29486 35982 29538
rect 36034 29486 36046 29538
rect 47394 29486 47406 29538
rect 47458 29486 47470 29538
rect 50754 29486 50766 29538
rect 50818 29486 50830 29538
rect 26462 29474 26514 29486
rect 44046 29474 44098 29486
rect 50990 29474 51042 29486
rect 4958 29426 5010 29438
rect 8654 29426 8706 29438
rect 5394 29374 5406 29426
rect 5458 29374 5470 29426
rect 4958 29362 5010 29374
rect 8654 29362 8706 29374
rect 11342 29426 11394 29438
rect 27358 29426 27410 29438
rect 16034 29374 16046 29426
rect 16098 29374 16110 29426
rect 21298 29374 21310 29426
rect 21362 29374 21374 29426
rect 27234 29374 27246 29426
rect 27298 29374 27310 29426
rect 11342 29362 11394 29374
rect 27358 29362 27410 29374
rect 27582 29426 27634 29438
rect 37774 29426 37826 29438
rect 46958 29426 47010 29438
rect 29586 29374 29598 29426
rect 29650 29374 29662 29426
rect 36642 29374 36654 29426
rect 36706 29374 36718 29426
rect 37986 29374 37998 29426
rect 38050 29374 38062 29426
rect 43810 29374 43822 29426
rect 43874 29374 43886 29426
rect 27582 29362 27634 29374
rect 37774 29362 37826 29374
rect 46958 29362 47010 29374
rect 47182 29426 47234 29438
rect 49310 29426 49362 29438
rect 47506 29374 47518 29426
rect 47570 29374 47582 29426
rect 47182 29362 47234 29374
rect 49310 29362 49362 29374
rect 49646 29426 49698 29438
rect 49646 29362 49698 29374
rect 49982 29426 50034 29438
rect 51102 29426 51154 29438
rect 50642 29374 50654 29426
rect 50706 29374 50718 29426
rect 49982 29362 50034 29374
rect 51102 29362 51154 29374
rect 52222 29426 52274 29438
rect 54786 29374 54798 29426
rect 54850 29374 54862 29426
rect 55010 29374 55022 29426
rect 55074 29374 55086 29426
rect 52222 29362 52274 29374
rect 11118 29314 11170 29326
rect 25230 29314 25282 29326
rect 22082 29262 22094 29314
rect 22146 29262 22158 29314
rect 24210 29262 24222 29314
rect 24274 29262 24286 29314
rect 11118 29250 11170 29262
rect 25230 29250 25282 29262
rect 28142 29314 28194 29326
rect 44494 29314 44546 29326
rect 32498 29262 32510 29314
rect 32562 29262 32574 29314
rect 33842 29262 33854 29314
rect 33906 29262 33918 29314
rect 28142 29250 28194 29262
rect 44494 29250 44546 29262
rect 45054 29314 45106 29326
rect 45054 29250 45106 29262
rect 46622 29314 46674 29326
rect 46622 29250 46674 29262
rect 51662 29314 51714 29326
rect 51662 29250 51714 29262
rect 55246 29314 55298 29326
rect 55246 29250 55298 29262
rect 55582 29314 55634 29326
rect 55582 29250 55634 29262
rect 25342 29202 25394 29214
rect 25342 29138 25394 29150
rect 26574 29202 26626 29214
rect 26574 29138 26626 29150
rect 26910 29202 26962 29214
rect 26910 29138 26962 29150
rect 44606 29202 44658 29214
rect 44606 29138 44658 29150
rect 50206 29202 50258 29214
rect 50206 29138 50258 29150
rect 55918 29202 55970 29214
rect 55918 29138 55970 29150
rect 1344 29034 58576 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 58576 29034
rect 1344 28948 58576 28982
rect 15934 28866 15986 28878
rect 8866 28814 8878 28866
rect 8930 28814 8942 28866
rect 15934 28802 15986 28814
rect 26014 28866 26066 28878
rect 26014 28802 26066 28814
rect 27246 28866 27298 28878
rect 46062 28866 46114 28878
rect 45602 28814 45614 28866
rect 45666 28814 45678 28866
rect 27246 28802 27298 28814
rect 46062 28802 46114 28814
rect 50318 28866 50370 28878
rect 50318 28802 50370 28814
rect 54798 28866 54850 28878
rect 54798 28802 54850 28814
rect 12126 28754 12178 28766
rect 22318 28754 22370 28766
rect 18386 28702 18398 28754
rect 18450 28702 18462 28754
rect 12126 28690 12178 28702
rect 22318 28690 22370 28702
rect 26574 28754 26626 28766
rect 26574 28690 26626 28702
rect 29822 28754 29874 28766
rect 29822 28690 29874 28702
rect 31054 28754 31106 28766
rect 48526 28754 48578 28766
rect 39890 28702 39902 28754
rect 39954 28702 39966 28754
rect 42018 28702 42030 28754
rect 42082 28702 42094 28754
rect 43474 28702 43486 28754
rect 43538 28702 43550 28754
rect 31054 28690 31106 28702
rect 48526 28690 48578 28702
rect 50430 28754 50482 28766
rect 50430 28690 50482 28702
rect 52782 28754 52834 28766
rect 53890 28702 53902 28754
rect 53954 28702 53966 28754
rect 56018 28702 56030 28754
rect 56082 28702 56094 28754
rect 58146 28702 58158 28754
rect 58210 28702 58222 28754
rect 52782 28690 52834 28702
rect 6862 28642 6914 28654
rect 6862 28578 6914 28590
rect 8654 28642 8706 28654
rect 9662 28642 9714 28654
rect 8866 28590 8878 28642
rect 8930 28590 8942 28642
rect 8654 28578 8706 28590
rect 9662 28578 9714 28590
rect 9886 28642 9938 28654
rect 9886 28578 9938 28590
rect 10110 28642 10162 28654
rect 10110 28578 10162 28590
rect 10894 28642 10946 28654
rect 10894 28578 10946 28590
rect 11342 28642 11394 28654
rect 11342 28578 11394 28590
rect 11566 28642 11618 28654
rect 11566 28578 11618 28590
rect 12014 28642 12066 28654
rect 12014 28578 12066 28590
rect 12238 28642 12290 28654
rect 12238 28578 12290 28590
rect 12462 28642 12514 28654
rect 12462 28578 12514 28590
rect 16158 28642 16210 28654
rect 16158 28578 16210 28590
rect 16494 28642 16546 28654
rect 16494 28578 16546 28590
rect 17166 28642 17218 28654
rect 27358 28642 27410 28654
rect 17714 28590 17726 28642
rect 17778 28590 17790 28642
rect 23090 28590 23102 28642
rect 23154 28590 23166 28642
rect 23538 28590 23550 28642
rect 23602 28590 23614 28642
rect 24434 28590 24446 28642
rect 24498 28590 24510 28642
rect 26338 28590 26350 28642
rect 26402 28590 26414 28642
rect 17166 28578 17218 28590
rect 27358 28578 27410 28590
rect 29038 28642 29090 28654
rect 29038 28578 29090 28590
rect 38222 28642 38274 28654
rect 44270 28642 44322 28654
rect 39218 28590 39230 28642
rect 39282 28590 39294 28642
rect 43810 28590 43822 28642
rect 43874 28590 43886 28642
rect 38222 28578 38274 28590
rect 44270 28578 44322 28590
rect 44942 28642 44994 28654
rect 44942 28578 44994 28590
rect 45166 28642 45218 28654
rect 47182 28642 47234 28654
rect 46386 28590 46398 28642
rect 46450 28590 46462 28642
rect 45166 28578 45218 28590
rect 47182 28578 47234 28590
rect 47854 28642 47906 28654
rect 47854 28578 47906 28590
rect 50990 28642 51042 28654
rect 50990 28578 51042 28590
rect 51326 28642 51378 28654
rect 51326 28578 51378 28590
rect 51550 28642 51602 28654
rect 51550 28578 51602 28590
rect 52110 28642 52162 28654
rect 52110 28578 52162 28590
rect 52670 28642 52722 28654
rect 54238 28642 54290 28654
rect 54910 28642 54962 28654
rect 53778 28590 53790 28642
rect 53842 28590 53854 28642
rect 54450 28590 54462 28642
rect 54514 28590 54526 28642
rect 55346 28590 55358 28642
rect 55410 28590 55422 28642
rect 52670 28578 52722 28590
rect 54238 28578 54290 28590
rect 54910 28578 54962 28590
rect 4398 28530 4450 28542
rect 4398 28466 4450 28478
rect 4510 28530 4562 28542
rect 4510 28466 4562 28478
rect 7646 28530 7698 28542
rect 7646 28466 7698 28478
rect 7982 28530 8034 28542
rect 7982 28466 8034 28478
rect 8318 28530 8370 28542
rect 8318 28466 8370 28478
rect 9438 28530 9490 28542
rect 9438 28466 9490 28478
rect 10558 28530 10610 28542
rect 10558 28466 10610 28478
rect 11118 28530 11170 28542
rect 11118 28466 11170 28478
rect 16718 28530 16770 28542
rect 26686 28530 26738 28542
rect 22754 28478 22766 28530
rect 22818 28478 22830 28530
rect 23762 28478 23774 28530
rect 23826 28478 23838 28530
rect 16718 28466 16770 28478
rect 26686 28466 26738 28478
rect 29262 28530 29314 28542
rect 29262 28466 29314 28478
rect 29374 28530 29426 28542
rect 29374 28466 29426 28478
rect 45054 28530 45106 28542
rect 45054 28466 45106 28478
rect 47406 28530 47458 28542
rect 47406 28466 47458 28478
rect 48190 28530 48242 28542
rect 48190 28466 48242 28478
rect 51998 28530 52050 28542
rect 51998 28466 52050 28478
rect 4174 28418 4226 28430
rect 9102 28418 9154 28430
rect 6514 28366 6526 28418
rect 6578 28366 6590 28418
rect 4174 28354 4226 28366
rect 9102 28354 9154 28366
rect 10670 28418 10722 28430
rect 10670 28354 10722 28366
rect 11342 28418 11394 28430
rect 16606 28418 16658 28430
rect 26462 28418 26514 28430
rect 15586 28366 15598 28418
rect 15650 28366 15662 28418
rect 20626 28366 20638 28418
rect 20690 28366 20702 28418
rect 23538 28366 23550 28418
rect 23602 28366 23614 28418
rect 11342 28354 11394 28366
rect 16606 28354 16658 28366
rect 26462 28354 26514 28366
rect 27246 28418 27298 28430
rect 27246 28354 27298 28366
rect 27806 28418 27858 28430
rect 27806 28354 27858 28366
rect 30942 28418 30994 28430
rect 46174 28418 46226 28430
rect 38546 28366 38558 28418
rect 38610 28366 38622 28418
rect 30942 28354 30994 28366
rect 46174 28354 46226 28366
rect 47630 28418 47682 28430
rect 47630 28354 47682 28366
rect 48414 28418 48466 28430
rect 48414 28354 48466 28366
rect 48638 28418 48690 28430
rect 48638 28354 48690 28366
rect 51102 28418 51154 28430
rect 51102 28354 51154 28366
rect 51774 28418 51826 28430
rect 51774 28354 51826 28366
rect 54014 28418 54066 28430
rect 54014 28354 54066 28366
rect 1344 28250 58576 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 58576 28250
rect 1344 28164 58576 28198
rect 5070 28082 5122 28094
rect 5070 28018 5122 28030
rect 7758 28082 7810 28094
rect 7758 28018 7810 28030
rect 8318 28082 8370 28094
rect 8318 28018 8370 28030
rect 11454 28082 11506 28094
rect 11454 28018 11506 28030
rect 12126 28082 12178 28094
rect 12126 28018 12178 28030
rect 25790 28082 25842 28094
rect 25790 28018 25842 28030
rect 27358 28082 27410 28094
rect 27358 28018 27410 28030
rect 31278 28082 31330 28094
rect 31278 28018 31330 28030
rect 32174 28082 32226 28094
rect 32174 28018 32226 28030
rect 34302 28082 34354 28094
rect 34302 28018 34354 28030
rect 47518 28082 47570 28094
rect 47518 28018 47570 28030
rect 54014 28082 54066 28094
rect 54014 28018 54066 28030
rect 11230 27970 11282 27982
rect 11230 27906 11282 27918
rect 11790 27970 11842 27982
rect 11790 27906 11842 27918
rect 11902 27970 11954 27982
rect 11902 27906 11954 27918
rect 23886 27970 23938 27982
rect 23886 27906 23938 27918
rect 28590 27970 28642 27982
rect 28590 27906 28642 27918
rect 28702 27970 28754 27982
rect 28702 27906 28754 27918
rect 33742 27970 33794 27982
rect 33742 27906 33794 27918
rect 34078 27970 34130 27982
rect 34078 27906 34130 27918
rect 34414 27970 34466 27982
rect 34414 27906 34466 27918
rect 4846 27858 4898 27870
rect 1810 27806 1822 27858
rect 1874 27806 1886 27858
rect 4846 27794 4898 27806
rect 5182 27858 5234 27870
rect 5182 27794 5234 27806
rect 8430 27858 8482 27870
rect 8430 27794 8482 27806
rect 8654 27858 8706 27870
rect 8654 27794 8706 27806
rect 8766 27858 8818 27870
rect 8766 27794 8818 27806
rect 11118 27858 11170 27870
rect 26014 27858 26066 27870
rect 13906 27806 13918 27858
rect 13970 27806 13982 27858
rect 20962 27806 20974 27858
rect 21026 27806 21038 27858
rect 11118 27794 11170 27806
rect 26014 27794 26066 27806
rect 28366 27858 28418 27870
rect 31502 27858 31554 27870
rect 31154 27806 31166 27858
rect 31218 27806 31230 27858
rect 28366 27794 28418 27806
rect 31502 27794 31554 27806
rect 33294 27858 33346 27870
rect 33294 27794 33346 27806
rect 33518 27858 33570 27870
rect 33518 27794 33570 27806
rect 36430 27858 36482 27870
rect 36430 27794 36482 27806
rect 36654 27858 36706 27870
rect 36654 27794 36706 27806
rect 37326 27858 37378 27870
rect 37326 27794 37378 27806
rect 38558 27858 38610 27870
rect 38558 27794 38610 27806
rect 38782 27858 38834 27870
rect 44046 27858 44098 27870
rect 41010 27806 41022 27858
rect 41074 27806 41086 27858
rect 38782 27794 38834 27806
rect 44046 27794 44098 27806
rect 44382 27858 44434 27870
rect 44382 27794 44434 27806
rect 44718 27858 44770 27870
rect 45278 27858 45330 27870
rect 45042 27806 45054 27858
rect 45106 27806 45118 27858
rect 44718 27794 44770 27806
rect 45278 27794 45330 27806
rect 45502 27858 45554 27870
rect 45502 27794 45554 27806
rect 47742 27858 47794 27870
rect 47742 27794 47794 27806
rect 48190 27858 48242 27870
rect 48190 27794 48242 27806
rect 9662 27746 9714 27758
rect 2482 27694 2494 27746
rect 2546 27694 2558 27746
rect 4610 27694 4622 27746
rect 4674 27694 4686 27746
rect 9662 27682 9714 27694
rect 10222 27746 10274 27758
rect 24334 27746 24386 27758
rect 14690 27694 14702 27746
rect 14754 27694 14766 27746
rect 16818 27694 16830 27746
rect 16882 27694 16894 27746
rect 21298 27694 21310 27746
rect 21362 27694 21374 27746
rect 10222 27682 10274 27694
rect 24334 27682 24386 27694
rect 25566 27746 25618 27758
rect 25566 27682 25618 27694
rect 25902 27746 25954 27758
rect 25902 27682 25954 27694
rect 26798 27746 26850 27758
rect 26798 27682 26850 27694
rect 31390 27746 31442 27758
rect 31390 27682 31442 27694
rect 33630 27746 33682 27758
rect 44270 27746 44322 27758
rect 41682 27694 41694 27746
rect 41746 27694 41758 27746
rect 43810 27694 43822 27746
rect 43874 27694 43886 27746
rect 33630 27682 33682 27694
rect 44270 27682 44322 27694
rect 45614 27746 45666 27758
rect 45614 27682 45666 27694
rect 47630 27746 47682 27758
rect 47630 27682 47682 27694
rect 54126 27746 54178 27758
rect 54126 27682 54178 27694
rect 8206 27634 8258 27646
rect 8206 27570 8258 27582
rect 23998 27634 24050 27646
rect 23998 27570 24050 27582
rect 24446 27634 24498 27646
rect 24446 27570 24498 27582
rect 25342 27634 25394 27646
rect 25342 27570 25394 27582
rect 30830 27634 30882 27646
rect 30830 27570 30882 27582
rect 33070 27634 33122 27646
rect 37550 27634 37602 27646
rect 36978 27582 36990 27634
rect 37042 27582 37054 27634
rect 37874 27582 37886 27634
rect 37938 27582 37950 27634
rect 39106 27582 39118 27634
rect 39170 27582 39182 27634
rect 33070 27570 33122 27582
rect 37550 27570 37602 27582
rect 1344 27466 58576 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 58576 27466
rect 1344 27380 58576 27414
rect 16270 27298 16322 27310
rect 16270 27234 16322 27246
rect 16606 27298 16658 27310
rect 16606 27234 16658 27246
rect 29934 27298 29986 27310
rect 29934 27234 29986 27246
rect 51214 27298 51266 27310
rect 51214 27234 51266 27246
rect 3950 27186 4002 27198
rect 3950 27122 4002 27134
rect 21646 27186 21698 27198
rect 21646 27122 21698 27134
rect 22094 27186 22146 27198
rect 22094 27122 22146 27134
rect 34750 27186 34802 27198
rect 34750 27122 34802 27134
rect 37550 27186 37602 27198
rect 37550 27122 37602 27134
rect 38334 27186 38386 27198
rect 38334 27122 38386 27134
rect 3838 27074 3890 27086
rect 3838 27010 3890 27022
rect 4174 27074 4226 27086
rect 4174 27010 4226 27022
rect 4958 27074 5010 27086
rect 4958 27010 5010 27022
rect 5630 27074 5682 27086
rect 5630 27010 5682 27022
rect 7534 27074 7586 27086
rect 7534 27010 7586 27022
rect 9102 27074 9154 27086
rect 26798 27074 26850 27086
rect 16258 27022 16270 27074
rect 16322 27022 16334 27074
rect 22754 27022 22766 27074
rect 22818 27022 22830 27074
rect 24098 27022 24110 27074
rect 24162 27022 24174 27074
rect 25890 27022 25902 27074
rect 25954 27022 25966 27074
rect 9102 27010 9154 27022
rect 26798 27010 26850 27022
rect 27134 27074 27186 27086
rect 27134 27010 27186 27022
rect 29822 27074 29874 27086
rect 32958 27074 33010 27086
rect 49758 27074 49810 27086
rect 50990 27074 51042 27086
rect 52110 27074 52162 27086
rect 30258 27022 30270 27074
rect 30322 27022 30334 27074
rect 31938 27022 31950 27074
rect 32002 27022 32014 27074
rect 33730 27022 33742 27074
rect 33794 27022 33806 27074
rect 37090 27022 37102 27074
rect 37154 27022 37166 27074
rect 45378 27022 45390 27074
rect 45442 27022 45454 27074
rect 50194 27022 50206 27074
rect 50258 27022 50270 27074
rect 51426 27022 51438 27074
rect 51490 27022 51502 27074
rect 52882 27022 52894 27074
rect 52946 27022 52958 27074
rect 29822 27010 29874 27022
rect 32958 27010 33010 27022
rect 49758 27010 49810 27022
rect 50990 27010 51042 27022
rect 52110 27010 52162 27022
rect 4398 26962 4450 26974
rect 4398 26898 4450 26910
rect 4846 26962 4898 26974
rect 4846 26898 4898 26910
rect 5742 26962 5794 26974
rect 5742 26898 5794 26910
rect 7198 26962 7250 26974
rect 7198 26898 7250 26910
rect 7982 26962 8034 26974
rect 7982 26898 8034 26910
rect 8206 26962 8258 26974
rect 8206 26898 8258 26910
rect 8542 26962 8594 26974
rect 8542 26898 8594 26910
rect 8766 26962 8818 26974
rect 8766 26898 8818 26910
rect 8990 26962 9042 26974
rect 27022 26962 27074 26974
rect 22418 26910 22430 26962
rect 22482 26910 22494 26962
rect 25666 26910 25678 26962
rect 25730 26910 25742 26962
rect 8990 26898 9042 26910
rect 27022 26898 27074 26910
rect 27582 26962 27634 26974
rect 34862 26962 34914 26974
rect 30930 26910 30942 26962
rect 30994 26910 31006 26962
rect 27582 26898 27634 26910
rect 34862 26898 34914 26910
rect 38782 26962 38834 26974
rect 38782 26898 38834 26910
rect 43822 26962 43874 26974
rect 49870 26962 49922 26974
rect 47170 26910 47182 26962
rect 47234 26910 47246 26962
rect 50082 26910 50094 26962
rect 50146 26910 50158 26962
rect 55346 26910 55358 26962
rect 55410 26910 55422 26962
rect 43822 26898 43874 26910
rect 49870 26898 49922 26910
rect 4622 26850 4674 26862
rect 4622 26786 4674 26798
rect 5966 26850 6018 26862
rect 5966 26786 6018 26798
rect 8430 26850 8482 26862
rect 29710 26850 29762 26862
rect 45614 26850 45666 26862
rect 23426 26798 23438 26850
rect 23490 26798 23502 26850
rect 30258 26798 30270 26850
rect 30322 26798 30334 26850
rect 8430 26786 8482 26798
rect 29710 26786 29762 26798
rect 45614 26786 45666 26798
rect 47518 26850 47570 26862
rect 47518 26786 47570 26798
rect 50654 26850 50706 26862
rect 50654 26786 50706 26798
rect 51326 26850 51378 26862
rect 51326 26786 51378 26798
rect 1344 26682 58576 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 58576 26682
rect 1344 26596 58576 26630
rect 3278 26514 3330 26526
rect 3278 26450 3330 26462
rect 26350 26514 26402 26526
rect 26350 26450 26402 26462
rect 26574 26514 26626 26526
rect 26574 26450 26626 26462
rect 27246 26514 27298 26526
rect 27246 26450 27298 26462
rect 31614 26514 31666 26526
rect 31614 26450 31666 26462
rect 32174 26514 32226 26526
rect 32174 26450 32226 26462
rect 36542 26514 36594 26526
rect 38110 26514 38162 26526
rect 37090 26462 37102 26514
rect 37154 26462 37166 26514
rect 36542 26450 36594 26462
rect 38110 26450 38162 26462
rect 39006 26514 39058 26526
rect 39006 26450 39058 26462
rect 53006 26514 53058 26526
rect 53006 26450 53058 26462
rect 57598 26514 57650 26526
rect 58158 26514 58210 26526
rect 57810 26462 57822 26514
rect 57874 26462 57886 26514
rect 57598 26450 57650 26462
rect 58158 26450 58210 26462
rect 3166 26402 3218 26414
rect 31726 26402 31778 26414
rect 50654 26402 50706 26414
rect 13010 26350 13022 26402
rect 13074 26350 13086 26402
rect 20066 26350 20078 26402
rect 20130 26350 20142 26402
rect 24098 26350 24110 26402
rect 24162 26350 24174 26402
rect 30034 26350 30046 26402
rect 30098 26350 30110 26402
rect 33842 26350 33854 26402
rect 33906 26350 33918 26402
rect 37762 26350 37774 26402
rect 37826 26350 37838 26402
rect 41122 26350 41134 26402
rect 41186 26350 41198 26402
rect 3166 26338 3218 26350
rect 31726 26338 31778 26350
rect 50654 26338 50706 26350
rect 52334 26402 52386 26414
rect 52334 26338 52386 26350
rect 54238 26402 54290 26414
rect 54238 26338 54290 26350
rect 54350 26402 54402 26414
rect 54350 26338 54402 26350
rect 55470 26402 55522 26414
rect 55470 26338 55522 26350
rect 3502 26290 3554 26302
rect 9774 26290 9826 26302
rect 22878 26290 22930 26302
rect 25454 26290 25506 26302
rect 4946 26238 4958 26290
rect 5010 26238 5022 26290
rect 13794 26238 13806 26290
rect 13858 26238 13870 26290
rect 16594 26238 16606 26290
rect 16658 26238 16670 26290
rect 19282 26238 19294 26290
rect 19346 26238 19358 26290
rect 23090 26238 23102 26290
rect 23154 26238 23166 26290
rect 24322 26238 24334 26290
rect 24386 26238 24398 26290
rect 3502 26226 3554 26238
rect 9774 26226 9826 26238
rect 22878 26226 22930 26238
rect 25454 26226 25506 26238
rect 26126 26290 26178 26302
rect 37438 26290 37490 26302
rect 46622 26290 46674 26302
rect 30706 26238 30718 26290
rect 30770 26238 30782 26290
rect 33058 26238 33070 26290
rect 33122 26238 33134 26290
rect 46162 26238 46174 26290
rect 46226 26238 46238 26290
rect 26126 26226 26178 26238
rect 37438 26226 37490 26238
rect 46622 26226 46674 26238
rect 49982 26290 50034 26302
rect 49982 26226 50034 26238
rect 50430 26290 50482 26302
rect 52894 26290 52946 26302
rect 52658 26238 52670 26290
rect 52722 26238 52734 26290
rect 50430 26226 50482 26238
rect 52894 26226 52946 26238
rect 53118 26290 53170 26302
rect 54126 26290 54178 26302
rect 53330 26238 53342 26290
rect 53394 26238 53406 26290
rect 53118 26226 53170 26238
rect 54126 26226 54178 26238
rect 55022 26290 55074 26302
rect 55022 26226 55074 26238
rect 55694 26290 55746 26302
rect 55694 26226 55746 26238
rect 26462 26178 26514 26190
rect 36654 26178 36706 26190
rect 7970 26126 7982 26178
rect 8034 26126 8046 26178
rect 10882 26126 10894 26178
rect 10946 26126 10958 26178
rect 16146 26126 16158 26178
rect 16210 26126 16222 26178
rect 22194 26126 22206 26178
rect 22258 26126 22270 26178
rect 24210 26126 24222 26178
rect 24274 26126 24286 26178
rect 27906 26126 27918 26178
rect 27970 26126 27982 26178
rect 35970 26126 35982 26178
rect 36034 26126 36046 26178
rect 26462 26114 26514 26126
rect 36654 26114 36706 26126
rect 38558 26178 38610 26190
rect 38558 26114 38610 26126
rect 39678 26178 39730 26190
rect 39678 26114 39730 26126
rect 50542 26178 50594 26190
rect 50542 26114 50594 26126
rect 52222 26178 52274 26190
rect 52222 26114 52274 26126
rect 55246 26178 55298 26190
rect 55246 26114 55298 26126
rect 25566 26066 25618 26078
rect 15810 26014 15822 26066
rect 15874 26014 15886 26066
rect 25566 26002 25618 26014
rect 25902 26066 25954 26078
rect 25902 26002 25954 26014
rect 31614 26066 31666 26078
rect 31614 26002 31666 26014
rect 39566 26066 39618 26078
rect 54786 26014 54798 26066
rect 54850 26014 54862 26066
rect 39566 26002 39618 26014
rect 1344 25898 58576 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 58576 25898
rect 1344 25812 58576 25846
rect 6638 25730 6690 25742
rect 6638 25666 6690 25678
rect 49310 25730 49362 25742
rect 49310 25666 49362 25678
rect 53342 25730 53394 25742
rect 53342 25666 53394 25678
rect 22654 25618 22706 25630
rect 36430 25618 36482 25630
rect 8754 25566 8766 25618
rect 8818 25566 8830 25618
rect 10882 25566 10894 25618
rect 10946 25566 10958 25618
rect 23426 25566 23438 25618
rect 23490 25566 23502 25618
rect 25218 25566 25230 25618
rect 25282 25566 25294 25618
rect 27346 25566 27358 25618
rect 27410 25566 27422 25618
rect 31378 25566 31390 25618
rect 31442 25566 31454 25618
rect 22654 25554 22706 25566
rect 36430 25554 36482 25566
rect 37886 25618 37938 25630
rect 53454 25618 53506 25630
rect 39330 25566 39342 25618
rect 39394 25566 39406 25618
rect 41458 25566 41470 25618
rect 41522 25566 41534 25618
rect 45714 25566 45726 25618
rect 45778 25566 45790 25618
rect 47842 25566 47854 25618
rect 47906 25566 47918 25618
rect 49746 25566 49758 25618
rect 49810 25566 49822 25618
rect 51202 25566 51214 25618
rect 51266 25566 51278 25618
rect 58146 25566 58158 25618
rect 58210 25566 58222 25618
rect 37886 25554 37938 25566
rect 53454 25554 53506 25566
rect 3614 25506 3666 25518
rect 3614 25442 3666 25454
rect 4062 25506 4114 25518
rect 4062 25442 4114 25454
rect 4286 25506 4338 25518
rect 4286 25442 4338 25454
rect 5630 25506 5682 25518
rect 5630 25442 5682 25454
rect 5966 25506 6018 25518
rect 5966 25442 6018 25454
rect 6302 25506 6354 25518
rect 6302 25442 6354 25454
rect 6526 25506 6578 25518
rect 6526 25442 6578 25454
rect 7310 25506 7362 25518
rect 7310 25442 7362 25454
rect 7646 25506 7698 25518
rect 28590 25506 28642 25518
rect 37326 25506 37378 25518
rect 43374 25506 43426 25518
rect 49198 25506 49250 25518
rect 54462 25506 54514 25518
rect 7970 25454 7982 25506
rect 8034 25454 8046 25506
rect 18050 25454 18062 25506
rect 18114 25454 18126 25506
rect 22978 25454 22990 25506
rect 23042 25454 23054 25506
rect 28130 25454 28142 25506
rect 28194 25454 28206 25506
rect 29362 25454 29374 25506
rect 29426 25454 29438 25506
rect 38658 25454 38670 25506
rect 38722 25454 38734 25506
rect 43698 25454 43710 25506
rect 43762 25454 43774 25506
rect 45042 25454 45054 25506
rect 45106 25454 45118 25506
rect 49634 25454 49646 25506
rect 49698 25454 49710 25506
rect 50754 25454 50766 25506
rect 50818 25454 50830 25506
rect 7646 25442 7698 25454
rect 28590 25442 28642 25454
rect 37326 25442 37378 25454
rect 43374 25442 43426 25454
rect 49198 25442 49250 25454
rect 54462 25442 54514 25454
rect 54686 25506 54738 25518
rect 54898 25454 54910 25506
rect 54962 25454 54974 25506
rect 55346 25454 55358 25506
rect 55410 25454 55422 25506
rect 54686 25442 54738 25454
rect 6638 25394 6690 25406
rect 6638 25330 6690 25342
rect 7422 25394 7474 25406
rect 42926 25394 42978 25406
rect 13906 25342 13918 25394
rect 13970 25342 13982 25394
rect 23314 25342 23326 25394
rect 23378 25342 23390 25394
rect 7422 25330 7474 25342
rect 42926 25330 42978 25342
rect 44270 25394 44322 25406
rect 51774 25394 51826 25406
rect 50082 25342 50094 25394
rect 50146 25342 50158 25394
rect 44270 25330 44322 25342
rect 51774 25330 51826 25342
rect 52670 25394 52722 25406
rect 52670 25330 52722 25342
rect 52782 25394 52834 25406
rect 56018 25342 56030 25394
rect 56082 25342 56094 25394
rect 52782 25330 52834 25342
rect 3838 25282 3890 25294
rect 3838 25218 3890 25230
rect 5966 25282 6018 25294
rect 5966 25218 6018 25230
rect 19182 25282 19234 25294
rect 19182 25218 19234 25230
rect 51214 25282 51266 25294
rect 51214 25218 51266 25230
rect 51326 25282 51378 25294
rect 51326 25218 51378 25230
rect 51550 25282 51602 25294
rect 51550 25218 51602 25230
rect 54798 25282 54850 25294
rect 54798 25218 54850 25230
rect 1344 25114 58576 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 58576 25114
rect 1344 25028 58576 25062
rect 30382 24946 30434 24958
rect 30382 24882 30434 24894
rect 37438 24946 37490 24958
rect 37438 24882 37490 24894
rect 40014 24946 40066 24958
rect 40014 24882 40066 24894
rect 40126 24946 40178 24958
rect 49198 24946 49250 24958
rect 45266 24894 45278 24946
rect 45330 24894 45342 24946
rect 40126 24882 40178 24894
rect 49198 24882 49250 24894
rect 50990 24946 51042 24958
rect 50990 24882 51042 24894
rect 55918 24946 55970 24958
rect 55918 24882 55970 24894
rect 24110 24834 24162 24846
rect 2482 24782 2494 24834
rect 2546 24782 2558 24834
rect 5730 24782 5742 24834
rect 5794 24782 5806 24834
rect 24110 24770 24162 24782
rect 24222 24834 24274 24846
rect 24222 24770 24274 24782
rect 30270 24834 30322 24846
rect 30270 24770 30322 24782
rect 37998 24834 38050 24846
rect 37998 24770 38050 24782
rect 40350 24834 40402 24846
rect 40350 24770 40402 24782
rect 44718 24834 44770 24846
rect 44718 24770 44770 24782
rect 49310 24834 49362 24846
rect 49310 24770 49362 24782
rect 49422 24834 49474 24846
rect 49422 24770 49474 24782
rect 51102 24834 51154 24846
rect 51102 24770 51154 24782
rect 35534 24722 35586 24734
rect 1810 24670 1822 24722
rect 1874 24670 1886 24722
rect 5058 24670 5070 24722
rect 5122 24670 5134 24722
rect 10770 24670 10782 24722
rect 10834 24670 10846 24722
rect 13906 24670 13918 24722
rect 13970 24670 13982 24722
rect 22194 24670 22206 24722
rect 22258 24670 22270 24722
rect 35534 24658 35586 24670
rect 35982 24722 36034 24734
rect 35982 24658 36034 24670
rect 36206 24722 36258 24734
rect 36206 24658 36258 24670
rect 37550 24722 37602 24734
rect 37550 24658 37602 24670
rect 38222 24722 38274 24734
rect 38222 24658 38274 24670
rect 39342 24722 39394 24734
rect 39902 24722 39954 24734
rect 49086 24722 49138 24734
rect 54574 24722 54626 24734
rect 56702 24722 56754 24734
rect 39666 24670 39678 24722
rect 39730 24670 39742 24722
rect 41122 24670 41134 24722
rect 41186 24670 41198 24722
rect 49858 24670 49870 24722
rect 49922 24670 49934 24722
rect 56018 24670 56030 24722
rect 56082 24670 56094 24722
rect 56914 24670 56926 24722
rect 56978 24670 56990 24722
rect 39342 24658 39394 24670
rect 39902 24658 39954 24670
rect 49086 24658 49138 24670
rect 54574 24658 54626 24670
rect 56702 24658 56754 24670
rect 9774 24610 9826 24622
rect 18062 24610 18114 24622
rect 36094 24610 36146 24622
rect 4610 24558 4622 24610
rect 4674 24558 4686 24610
rect 7858 24558 7870 24610
rect 7922 24558 7934 24610
rect 11442 24558 11454 24610
rect 11506 24558 11518 24610
rect 13570 24558 13582 24610
rect 13634 24558 13646 24610
rect 14690 24558 14702 24610
rect 14754 24558 14766 24610
rect 16818 24558 16830 24610
rect 16882 24558 16894 24610
rect 18610 24558 18622 24610
rect 18674 24558 18686 24610
rect 9774 24546 9826 24558
rect 18062 24546 18114 24558
rect 36094 24546 36146 24558
rect 36766 24610 36818 24622
rect 36766 24546 36818 24558
rect 38110 24610 38162 24622
rect 44942 24610 44994 24622
rect 41794 24558 41806 24610
rect 41858 24558 41870 24610
rect 43922 24558 43934 24610
rect 43986 24558 43998 24610
rect 38110 24546 38162 24558
rect 44942 24546 44994 24558
rect 55582 24610 55634 24622
rect 55582 24546 55634 24558
rect 24110 24498 24162 24510
rect 24110 24434 24162 24446
rect 54798 24498 54850 24510
rect 55806 24498 55858 24510
rect 55122 24446 55134 24498
rect 55186 24446 55198 24498
rect 54798 24434 54850 24446
rect 55806 24434 55858 24446
rect 56590 24498 56642 24510
rect 56590 24434 56642 24446
rect 1344 24330 58576 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 58576 24330
rect 1344 24244 58576 24278
rect 8990 24162 9042 24174
rect 8642 24110 8654 24162
rect 8706 24110 8718 24162
rect 8990 24098 9042 24110
rect 9662 24162 9714 24174
rect 9662 24098 9714 24110
rect 12350 24162 12402 24174
rect 12350 24098 12402 24110
rect 15822 24162 15874 24174
rect 15822 24098 15874 24110
rect 41806 24162 41858 24174
rect 41806 24098 41858 24110
rect 49422 24162 49474 24174
rect 49422 24098 49474 24110
rect 53790 24162 53842 24174
rect 53790 24098 53842 24110
rect 15934 24050 15986 24062
rect 48862 24050 48914 24062
rect 20738 23998 20750 24050
rect 20802 23998 20814 24050
rect 33170 23998 33182 24050
rect 33234 23998 33246 24050
rect 15934 23986 15986 23998
rect 48862 23986 48914 23998
rect 49870 24050 49922 24062
rect 56018 23998 56030 24050
rect 56082 23998 56094 24050
rect 58146 23998 58158 24050
rect 58210 23998 58222 24050
rect 49870 23986 49922 23998
rect 9214 23938 9266 23950
rect 9214 23874 9266 23886
rect 9774 23938 9826 23950
rect 14254 23938 14306 23950
rect 22318 23938 22370 23950
rect 12338 23886 12350 23938
rect 12402 23886 12414 23938
rect 14578 23886 14590 23938
rect 14642 23886 14654 23938
rect 17826 23886 17838 23938
rect 17890 23886 17902 23938
rect 9774 23874 9826 23886
rect 14254 23874 14306 23886
rect 22318 23874 22370 23886
rect 22766 23938 22818 23950
rect 22766 23874 22818 23886
rect 23326 23938 23378 23950
rect 23326 23874 23378 23886
rect 23662 23938 23714 23950
rect 23662 23874 23714 23886
rect 24222 23938 24274 23950
rect 24222 23874 24274 23886
rect 31838 23938 31890 23950
rect 31838 23874 31890 23886
rect 32174 23938 32226 23950
rect 41246 23938 41298 23950
rect 46398 23938 46450 23950
rect 35970 23886 35982 23938
rect 36034 23886 36046 23938
rect 37426 23886 37438 23938
rect 37490 23886 37502 23938
rect 40786 23886 40798 23938
rect 40850 23886 40862 23938
rect 41458 23886 41470 23938
rect 41522 23886 41534 23938
rect 45266 23886 45278 23938
rect 45330 23886 45342 23938
rect 45938 23886 45950 23938
rect 46002 23886 46014 23938
rect 32174 23874 32226 23886
rect 41246 23874 41298 23886
rect 46398 23874 46450 23886
rect 49086 23938 49138 23950
rect 55346 23886 55358 23938
rect 55410 23886 55422 23938
rect 49086 23874 49138 23886
rect 12686 23826 12738 23838
rect 12686 23762 12738 23774
rect 14142 23826 14194 23838
rect 22094 23826 22146 23838
rect 18610 23774 18622 23826
rect 18674 23774 18686 23826
rect 14142 23762 14194 23774
rect 22094 23762 22146 23774
rect 22206 23826 22258 23838
rect 22206 23762 22258 23774
rect 23886 23826 23938 23838
rect 23886 23762 23938 23774
rect 31502 23826 31554 23838
rect 36878 23826 36930 23838
rect 35298 23774 35310 23826
rect 35362 23774 35374 23826
rect 31502 23762 31554 23774
rect 36878 23762 36930 23774
rect 38558 23826 38610 23838
rect 38558 23762 38610 23774
rect 41134 23826 41186 23838
rect 41134 23762 41186 23774
rect 41918 23826 41970 23838
rect 49758 23826 49810 23838
rect 45042 23774 45054 23826
rect 45106 23774 45118 23826
rect 45714 23774 45726 23826
rect 45778 23774 45790 23826
rect 46722 23774 46734 23826
rect 46786 23774 46798 23826
rect 41918 23762 41970 23774
rect 49758 23762 49810 23774
rect 49982 23826 50034 23838
rect 49982 23762 50034 23774
rect 53902 23826 53954 23838
rect 53902 23762 53954 23774
rect 9662 23714 9714 23726
rect 9662 23650 9714 23662
rect 10222 23714 10274 23726
rect 10222 23650 10274 23662
rect 14030 23714 14082 23726
rect 14030 23650 14082 23662
rect 15038 23714 15090 23726
rect 15038 23650 15090 23662
rect 16046 23714 16098 23726
rect 16046 23650 16098 23662
rect 16718 23714 16770 23726
rect 23998 23714 24050 23726
rect 21634 23662 21646 23714
rect 21698 23662 21710 23714
rect 16718 23650 16770 23662
rect 23998 23650 24050 23662
rect 31950 23714 32002 23726
rect 31950 23650 32002 23662
rect 32510 23714 32562 23726
rect 32510 23650 32562 23662
rect 36990 23714 37042 23726
rect 36990 23650 37042 23662
rect 37214 23714 37266 23726
rect 37214 23650 37266 23662
rect 38446 23714 38498 23726
rect 38446 23650 38498 23662
rect 41022 23714 41074 23726
rect 41022 23650 41074 23662
rect 1344 23546 58576 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 58576 23546
rect 1344 23460 58576 23494
rect 9662 23378 9714 23390
rect 9662 23314 9714 23326
rect 17390 23378 17442 23390
rect 17390 23314 17442 23326
rect 21982 23378 22034 23390
rect 21982 23314 22034 23326
rect 33294 23378 33346 23390
rect 33294 23314 33346 23326
rect 47406 23378 47458 23390
rect 47406 23314 47458 23326
rect 49086 23378 49138 23390
rect 49086 23314 49138 23326
rect 49870 23378 49922 23390
rect 49870 23314 49922 23326
rect 53006 23378 53058 23390
rect 53006 23314 53058 23326
rect 19294 23266 19346 23278
rect 47630 23266 47682 23278
rect 21634 23214 21646 23266
rect 21698 23214 21710 23266
rect 35298 23214 35310 23266
rect 35362 23214 35374 23266
rect 19294 23202 19346 23214
rect 47630 23202 47682 23214
rect 49982 23266 50034 23278
rect 49982 23202 50034 23214
rect 55694 23266 55746 23278
rect 55694 23202 55746 23214
rect 55918 23266 55970 23278
rect 55918 23202 55970 23214
rect 14030 23154 14082 23166
rect 1810 23102 1822 23154
rect 1874 23102 1886 23154
rect 14030 23090 14082 23102
rect 17614 23154 17666 23166
rect 19406 23154 19458 23166
rect 17938 23102 17950 23154
rect 18002 23102 18014 23154
rect 17614 23090 17666 23102
rect 19406 23090 19458 23102
rect 19742 23154 19794 23166
rect 23214 23154 23266 23166
rect 25342 23154 25394 23166
rect 22866 23102 22878 23154
rect 22930 23102 22942 23154
rect 23874 23102 23886 23154
rect 23938 23102 23950 23154
rect 19742 23090 19794 23102
rect 23214 23090 23266 23102
rect 25342 23090 25394 23102
rect 26574 23154 26626 23166
rect 26574 23090 26626 23102
rect 27022 23154 27074 23166
rect 27022 23090 27074 23102
rect 27246 23154 27298 23166
rect 27246 23090 27298 23102
rect 28254 23154 28306 23166
rect 28254 23090 28306 23102
rect 28814 23154 28866 23166
rect 33070 23154 33122 23166
rect 32050 23102 32062 23154
rect 32114 23102 32126 23154
rect 28814 23090 28866 23102
rect 33070 23090 33122 23102
rect 33742 23154 33794 23166
rect 47966 23154 48018 23166
rect 39778 23102 39790 23154
rect 39842 23102 39854 23154
rect 33742 23090 33794 23102
rect 47966 23090 48018 23102
rect 48302 23154 48354 23166
rect 48302 23090 48354 23102
rect 48862 23154 48914 23166
rect 48862 23090 48914 23102
rect 48974 23154 49026 23166
rect 48974 23090 49026 23102
rect 49198 23154 49250 23166
rect 52334 23154 52386 23166
rect 49410 23102 49422 23154
rect 49474 23102 49486 23154
rect 51762 23102 51774 23154
rect 51826 23102 51838 23154
rect 49198 23090 49250 23102
rect 52334 23090 52386 23102
rect 55022 23154 55074 23166
rect 55022 23090 55074 23102
rect 55246 23154 55298 23166
rect 55246 23090 55298 23102
rect 9550 23042 9602 23054
rect 2482 22990 2494 23042
rect 2546 22990 2558 23042
rect 4610 22990 4622 23042
rect 4674 22990 4686 23042
rect 9550 22978 9602 22990
rect 17502 23042 17554 23054
rect 17502 22978 17554 22990
rect 20302 23042 20354 23054
rect 26350 23042 26402 23054
rect 24658 22990 24670 23042
rect 24722 22990 24734 23042
rect 20302 22978 20354 22990
rect 26350 22978 26402 22990
rect 26798 23042 26850 23054
rect 26798 22978 26850 22990
rect 27918 23042 27970 23054
rect 32510 23042 32562 23054
rect 29138 22990 29150 23042
rect 29202 22990 29214 23042
rect 31266 22990 31278 23042
rect 31330 22990 31342 23042
rect 27918 22978 27970 22990
rect 32510 22978 32562 22990
rect 33182 23042 33234 23054
rect 33182 22978 33234 22990
rect 40238 23042 40290 23054
rect 40238 22978 40290 22990
rect 41918 23042 41970 23054
rect 41918 22978 41970 22990
rect 48078 23042 48130 23054
rect 48078 22978 48130 22990
rect 52446 23042 52498 23054
rect 52446 22978 52498 22990
rect 52782 23042 52834 23054
rect 52782 22978 52834 22990
rect 13806 22930 13858 22942
rect 13458 22878 13470 22930
rect 13522 22878 13534 22930
rect 13806 22866 13858 22878
rect 19630 22930 19682 22942
rect 19630 22866 19682 22878
rect 42030 22930 42082 22942
rect 42030 22866 42082 22878
rect 49758 22930 49810 22942
rect 49758 22866 49810 22878
rect 53118 22930 53170 22942
rect 55582 22930 55634 22942
rect 54674 22878 54686 22930
rect 54738 22878 54750 22930
rect 53118 22866 53170 22878
rect 55582 22866 55634 22878
rect 1344 22762 58576 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 58576 22762
rect 1344 22676 58576 22710
rect 4734 22594 4786 22606
rect 35982 22594 36034 22606
rect 32050 22542 32062 22594
rect 32114 22542 32126 22594
rect 4734 22530 4786 22542
rect 35982 22530 36034 22542
rect 36430 22594 36482 22606
rect 36430 22530 36482 22542
rect 51998 22594 52050 22606
rect 51998 22530 52050 22542
rect 52782 22594 52834 22606
rect 52782 22530 52834 22542
rect 3390 22482 3442 22494
rect 3390 22418 3442 22430
rect 3950 22482 4002 22494
rect 35534 22482 35586 22494
rect 52110 22482 52162 22494
rect 9538 22430 9550 22482
rect 9602 22430 9614 22482
rect 12898 22430 12910 22482
rect 12962 22430 12974 22482
rect 18162 22430 18174 22482
rect 18226 22430 18238 22482
rect 25666 22430 25678 22482
rect 25730 22430 25742 22482
rect 27794 22430 27806 22482
rect 27858 22430 27870 22482
rect 37986 22430 37998 22482
rect 38050 22430 38062 22482
rect 40114 22430 40126 22482
rect 40178 22430 40190 22482
rect 42130 22430 42142 22482
rect 42194 22430 42206 22482
rect 44258 22430 44270 22482
rect 44322 22430 44334 22482
rect 45378 22430 45390 22482
rect 45442 22430 45454 22482
rect 58146 22430 58158 22482
rect 58210 22430 58222 22482
rect 3950 22418 4002 22430
rect 35534 22418 35586 22430
rect 52110 22418 52162 22430
rect 4174 22370 4226 22382
rect 4174 22306 4226 22318
rect 5630 22370 5682 22382
rect 5630 22306 5682 22318
rect 5854 22370 5906 22382
rect 24782 22370 24834 22382
rect 31390 22370 31442 22382
rect 6738 22318 6750 22370
rect 6802 22318 6814 22370
rect 10098 22318 10110 22370
rect 10162 22318 10174 22370
rect 15250 22318 15262 22370
rect 15314 22318 15326 22370
rect 23090 22318 23102 22370
rect 23154 22318 23166 22370
rect 23986 22318 23998 22370
rect 24050 22318 24062 22370
rect 28578 22318 28590 22370
rect 28642 22318 28654 22370
rect 5854 22306 5906 22318
rect 24782 22306 24834 22318
rect 31390 22306 31442 22318
rect 31614 22370 31666 22382
rect 31614 22306 31666 22318
rect 32734 22370 32786 22382
rect 32734 22306 32786 22318
rect 35758 22370 35810 22382
rect 52894 22370 52946 22382
rect 37202 22318 37214 22370
rect 37266 22318 37278 22370
rect 41346 22318 41358 22370
rect 41410 22318 41422 22370
rect 50418 22318 50430 22370
rect 50482 22318 50494 22370
rect 55234 22318 55246 22370
rect 55298 22318 55310 22370
rect 35758 22306 35810 22318
rect 52894 22306 52946 22318
rect 5070 22258 5122 22270
rect 25342 22258 25394 22270
rect 7410 22206 7422 22258
rect 7474 22206 7486 22258
rect 10770 22206 10782 22258
rect 10834 22206 10846 22258
rect 16034 22206 16046 22258
rect 16098 22206 16110 22258
rect 23762 22206 23774 22258
rect 23826 22206 23838 22258
rect 5070 22194 5122 22206
rect 25342 22194 25394 22206
rect 31502 22258 31554 22270
rect 31502 22194 31554 22206
rect 52782 22258 52834 22270
rect 56018 22206 56030 22258
rect 56082 22206 56094 22258
rect 52782 22194 52834 22206
rect 4846 22146 4898 22158
rect 33182 22146 33234 22158
rect 3602 22094 3614 22146
rect 3666 22094 3678 22146
rect 6178 22094 6190 22146
rect 6242 22094 6254 22146
rect 22642 22094 22654 22146
rect 22706 22094 22718 22146
rect 23426 22094 23438 22146
rect 23490 22094 23502 22146
rect 4846 22082 4898 22094
rect 33182 22082 33234 22094
rect 50878 22146 50930 22158
rect 50878 22082 50930 22094
rect 1344 21978 58576 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 58576 21978
rect 1344 21892 58576 21926
rect 8878 21810 8930 21822
rect 8878 21746 8930 21758
rect 12798 21810 12850 21822
rect 12798 21746 12850 21758
rect 13470 21810 13522 21822
rect 19182 21810 19234 21822
rect 16146 21758 16158 21810
rect 16210 21758 16222 21810
rect 13470 21746 13522 21758
rect 19182 21746 19234 21758
rect 23550 21810 23602 21822
rect 23550 21746 23602 21758
rect 24558 21810 24610 21822
rect 24558 21746 24610 21758
rect 27246 21810 27298 21822
rect 27246 21746 27298 21758
rect 27358 21810 27410 21822
rect 27358 21746 27410 21758
rect 28254 21810 28306 21822
rect 28254 21746 28306 21758
rect 36766 21810 36818 21822
rect 36766 21746 36818 21758
rect 38110 21810 38162 21822
rect 38110 21746 38162 21758
rect 38782 21810 38834 21822
rect 38782 21746 38834 21758
rect 39006 21810 39058 21822
rect 39006 21746 39058 21758
rect 39118 21810 39170 21822
rect 39118 21746 39170 21758
rect 41246 21810 41298 21822
rect 41246 21746 41298 21758
rect 48974 21810 49026 21822
rect 48974 21746 49026 21758
rect 49534 21810 49586 21822
rect 49534 21746 49586 21758
rect 12686 21698 12738 21710
rect 6402 21646 6414 21698
rect 6466 21646 6478 21698
rect 12686 21634 12738 21646
rect 16606 21698 16658 21710
rect 16606 21634 16658 21646
rect 16830 21698 16882 21710
rect 16830 21634 16882 21646
rect 37438 21698 37490 21710
rect 37438 21634 37490 21646
rect 39342 21698 39394 21710
rect 39342 21634 39394 21646
rect 41582 21698 41634 21710
rect 41582 21634 41634 21646
rect 43374 21698 43426 21710
rect 48750 21698 48802 21710
rect 55806 21698 55858 21710
rect 46050 21646 46062 21698
rect 46114 21646 46126 21698
rect 53106 21646 53118 21698
rect 53170 21646 53182 21698
rect 57810 21646 57822 21698
rect 57874 21646 57886 21698
rect 43374 21634 43426 21646
rect 48750 21634 48802 21646
rect 55806 21634 55858 21646
rect 13246 21586 13298 21598
rect 8418 21534 8430 21586
rect 8482 21534 8494 21586
rect 13246 21522 13298 21534
rect 13918 21586 13970 21598
rect 13918 21522 13970 21534
rect 14478 21586 14530 21598
rect 14478 21522 14530 21534
rect 14702 21586 14754 21598
rect 14702 21522 14754 21534
rect 15822 21586 15874 21598
rect 17726 21586 17778 21598
rect 17378 21534 17390 21586
rect 17442 21534 17454 21586
rect 15822 21522 15874 21534
rect 17726 21522 17778 21534
rect 17950 21586 18002 21598
rect 17950 21522 18002 21534
rect 18846 21586 18898 21598
rect 18846 21522 18898 21534
rect 19182 21586 19234 21598
rect 19182 21522 19234 21534
rect 19518 21586 19570 21598
rect 19518 21522 19570 21534
rect 22430 21586 22482 21598
rect 23774 21586 23826 21598
rect 27134 21586 27186 21598
rect 22642 21534 22654 21586
rect 22706 21534 22718 21586
rect 24098 21534 24110 21586
rect 24162 21534 24174 21586
rect 22430 21522 22482 21534
rect 23774 21522 23826 21534
rect 27134 21522 27186 21534
rect 27806 21586 27858 21598
rect 36542 21586 36594 21598
rect 38894 21586 38946 21598
rect 41134 21586 41186 21598
rect 33058 21534 33070 21586
rect 33122 21534 33134 21586
rect 36306 21534 36318 21586
rect 36370 21534 36382 21586
rect 36978 21534 36990 21586
rect 37042 21534 37054 21586
rect 40898 21534 40910 21586
rect 40962 21534 40974 21586
rect 27806 21522 27858 21534
rect 36542 21522 36594 21534
rect 38894 21522 38946 21534
rect 41134 21522 41186 21534
rect 41358 21586 41410 21598
rect 55358 21586 55410 21598
rect 42466 21534 42478 21586
rect 42530 21534 42542 21586
rect 45378 21534 45390 21586
rect 45442 21534 45454 21586
rect 53890 21534 53902 21586
rect 53954 21534 53966 21586
rect 41358 21522 41410 21534
rect 55358 21522 55410 21534
rect 55470 21586 55522 21598
rect 55470 21522 55522 21534
rect 58158 21586 58210 21598
rect 58158 21522 58210 21534
rect 13358 21474 13410 21486
rect 23214 21474 23266 21486
rect 16482 21422 16494 21474
rect 16546 21422 16558 21474
rect 13358 21410 13410 21422
rect 23214 21410 23266 21422
rect 23662 21474 23714 21486
rect 23662 21410 23714 21422
rect 26798 21474 26850 21486
rect 32510 21474 32562 21486
rect 36654 21474 36706 21486
rect 39790 21474 39842 21486
rect 27794 21422 27806 21474
rect 27858 21422 27870 21474
rect 33842 21422 33854 21474
rect 33906 21422 33918 21474
rect 35970 21422 35982 21474
rect 36034 21422 36046 21474
rect 37314 21422 37326 21474
rect 37378 21422 37390 21474
rect 26798 21410 26850 21422
rect 12910 21362 12962 21374
rect 14130 21310 14142 21362
rect 14194 21310 14206 21362
rect 27809 21359 27855 21422
rect 32510 21410 32562 21422
rect 36654 21410 36706 21422
rect 39790 21410 39842 21422
rect 42926 21474 42978 21486
rect 49422 21474 49474 21486
rect 55694 21474 55746 21486
rect 48178 21422 48190 21474
rect 48242 21422 48254 21474
rect 49074 21422 49086 21474
rect 49138 21422 49150 21474
rect 50978 21422 50990 21474
rect 51042 21422 51054 21474
rect 42926 21410 42978 21422
rect 49422 21410 49474 21422
rect 55694 21410 55746 21422
rect 57598 21474 57650 21486
rect 57598 21410 57650 21422
rect 37662 21362 37714 21374
rect 28242 21359 28254 21362
rect 27809 21313 28254 21359
rect 28242 21310 28254 21313
rect 28306 21310 28318 21362
rect 12910 21298 12962 21310
rect 37662 21298 37714 21310
rect 1344 21194 58576 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 58576 21194
rect 1344 21108 58576 21142
rect 22654 21026 22706 21038
rect 22654 20962 22706 20974
rect 23214 21026 23266 21038
rect 23214 20962 23266 20974
rect 23438 21026 23490 21038
rect 23438 20962 23490 20974
rect 34526 21026 34578 21038
rect 34526 20962 34578 20974
rect 5742 20914 5794 20926
rect 22990 20914 23042 20926
rect 4610 20862 4622 20914
rect 4674 20862 4686 20914
rect 17826 20862 17838 20914
rect 17890 20862 17902 20914
rect 19954 20862 19966 20914
rect 20018 20862 20030 20914
rect 5742 20850 5794 20862
rect 22990 20850 23042 20862
rect 26798 20914 26850 20926
rect 26798 20850 26850 20862
rect 27246 20914 27298 20926
rect 34638 20914 34690 20926
rect 32050 20862 32062 20914
rect 32114 20862 32126 20914
rect 27246 20850 27298 20862
rect 34638 20850 34690 20862
rect 39790 20914 39842 20926
rect 39790 20850 39842 20862
rect 5854 20802 5906 20814
rect 1810 20750 1822 20802
rect 1874 20750 1886 20802
rect 5854 20738 5906 20750
rect 6302 20802 6354 20814
rect 6302 20738 6354 20750
rect 13470 20802 13522 20814
rect 13470 20738 13522 20750
rect 13582 20802 13634 20814
rect 24334 20802 24386 20814
rect 37326 20802 37378 20814
rect 20738 20750 20750 20802
rect 20802 20750 20814 20802
rect 24770 20750 24782 20802
rect 24834 20750 24846 20802
rect 29138 20750 29150 20802
rect 29202 20750 29214 20802
rect 13582 20738 13634 20750
rect 24334 20738 24386 20750
rect 37326 20738 37378 20750
rect 37662 20802 37714 20814
rect 37662 20738 37714 20750
rect 39230 20802 39282 20814
rect 52882 20750 52894 20802
rect 52946 20750 52958 20802
rect 39230 20738 39282 20750
rect 7646 20690 7698 20702
rect 2482 20638 2494 20690
rect 2546 20638 2558 20690
rect 7298 20638 7310 20690
rect 7362 20638 7374 20690
rect 7646 20626 7698 20638
rect 7982 20690 8034 20702
rect 7982 20626 8034 20638
rect 13918 20690 13970 20702
rect 13918 20626 13970 20638
rect 22430 20690 22482 20702
rect 22430 20626 22482 20638
rect 23886 20690 23938 20702
rect 23886 20626 23938 20638
rect 24110 20690 24162 20702
rect 29922 20638 29934 20690
rect 29986 20638 29998 20690
rect 36978 20638 36990 20690
rect 37042 20638 37054 20690
rect 55346 20638 55358 20690
rect 55410 20638 55422 20690
rect 24110 20626 24162 20638
rect 5630 20578 5682 20590
rect 5630 20514 5682 20526
rect 6974 20578 7026 20590
rect 6974 20514 7026 20526
rect 13694 20578 13746 20590
rect 13694 20514 13746 20526
rect 22542 20578 22594 20590
rect 22542 20514 22594 20526
rect 24446 20578 24498 20590
rect 24446 20514 24498 20526
rect 24558 20578 24610 20590
rect 24558 20514 24610 20526
rect 27134 20578 27186 20590
rect 27134 20514 27186 20526
rect 35982 20578 36034 20590
rect 39342 20578 39394 20590
rect 42254 20578 42306 20590
rect 37986 20526 37998 20578
rect 38050 20526 38062 20578
rect 41906 20526 41918 20578
rect 41970 20526 41982 20578
rect 35982 20514 36034 20526
rect 39342 20514 39394 20526
rect 42254 20514 42306 20526
rect 42702 20578 42754 20590
rect 42702 20514 42754 20526
rect 52110 20578 52162 20590
rect 52110 20514 52162 20526
rect 1344 20410 58576 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 58576 20410
rect 1344 20324 58576 20358
rect 4062 20242 4114 20254
rect 4062 20178 4114 20190
rect 19518 20242 19570 20254
rect 19518 20178 19570 20190
rect 3278 20130 3330 20142
rect 3278 20066 3330 20078
rect 3838 20130 3890 20142
rect 3838 20066 3890 20078
rect 4958 20130 5010 20142
rect 6638 20130 6690 20142
rect 13806 20130 13858 20142
rect 6290 20078 6302 20130
rect 6354 20078 6366 20130
rect 8418 20078 8430 20130
rect 8482 20078 8494 20130
rect 4958 20066 5010 20078
rect 6638 20066 6690 20078
rect 13806 20066 13858 20078
rect 14030 20130 14082 20142
rect 14030 20066 14082 20078
rect 17614 20130 17666 20142
rect 17614 20066 17666 20078
rect 19406 20130 19458 20142
rect 19406 20066 19458 20078
rect 20526 20130 20578 20142
rect 20526 20066 20578 20078
rect 30494 20130 30546 20142
rect 41918 20130 41970 20142
rect 41570 20078 41582 20130
rect 41634 20078 41646 20130
rect 30494 20066 30546 20078
rect 41918 20066 41970 20078
rect 42366 20130 42418 20142
rect 42366 20066 42418 20078
rect 42814 20130 42866 20142
rect 42814 20066 42866 20078
rect 49086 20130 49138 20142
rect 49086 20066 49138 20078
rect 49758 20130 49810 20142
rect 49758 20066 49810 20078
rect 54798 20130 54850 20142
rect 54798 20066 54850 20078
rect 56142 20130 56194 20142
rect 56142 20066 56194 20078
rect 4510 20018 4562 20030
rect 12910 20018 12962 20030
rect 9650 19966 9662 20018
rect 9714 19966 9726 20018
rect 4510 19954 4562 19966
rect 12910 19954 12962 19966
rect 13134 20018 13186 20030
rect 19630 20018 19682 20030
rect 13458 19966 13470 20018
rect 13522 19966 13534 20018
rect 13134 19954 13186 19966
rect 19630 19954 19682 19966
rect 20078 20018 20130 20030
rect 25902 20018 25954 20030
rect 23538 19966 23550 20018
rect 23602 19966 23614 20018
rect 23762 19966 23774 20018
rect 23826 19966 23838 20018
rect 20078 19954 20130 19966
rect 25902 19954 25954 19966
rect 26462 20018 26514 20030
rect 27358 20018 27410 20030
rect 26898 19966 26910 20018
rect 26962 19966 26974 20018
rect 26462 19954 26514 19966
rect 27358 19954 27410 19966
rect 27694 20018 27746 20030
rect 27694 19954 27746 19966
rect 29822 20018 29874 20030
rect 29822 19954 29874 19966
rect 30830 20018 30882 20030
rect 30830 19954 30882 19966
rect 31502 20018 31554 20030
rect 49422 20018 49474 20030
rect 31938 19966 31950 20018
rect 32002 19966 32014 20018
rect 44594 19966 44606 20018
rect 44658 19966 44670 20018
rect 31502 19954 31554 19966
rect 49422 19954 49474 19966
rect 49534 20018 49586 20030
rect 49534 19954 49586 19966
rect 49870 20018 49922 20030
rect 49870 19954 49922 19966
rect 54462 20018 54514 20030
rect 54462 19954 54514 19966
rect 54574 20018 54626 20030
rect 55010 19966 55022 20018
rect 55074 19966 55086 20018
rect 54574 19954 54626 19966
rect 3950 19906 4002 19918
rect 3154 19854 3166 19906
rect 3218 19854 3230 19906
rect 3950 19842 4002 19854
rect 8990 19906 9042 19918
rect 13918 19906 13970 19918
rect 10322 19854 10334 19906
rect 10386 19854 10398 19906
rect 12450 19854 12462 19906
rect 12514 19854 12526 19906
rect 8990 19842 9042 19854
rect 13918 19842 13970 19854
rect 17502 19906 17554 19918
rect 28254 19906 28306 19918
rect 23202 19854 23214 19906
rect 23266 19854 23278 19906
rect 17502 19842 17554 19854
rect 28254 19842 28306 19854
rect 29598 19906 29650 19918
rect 29598 19842 29650 19854
rect 30158 19906 30210 19918
rect 33182 19906 33234 19918
rect 49646 19906 49698 19918
rect 32274 19854 32286 19906
rect 32338 19854 32350 19906
rect 45378 19854 45390 19906
rect 45442 19854 45454 19906
rect 47506 19854 47518 19906
rect 47570 19854 47582 19906
rect 30158 19842 30210 19854
rect 33182 19842 33234 19854
rect 49646 19842 49698 19854
rect 50318 19906 50370 19918
rect 50318 19842 50370 19854
rect 54686 19906 54738 19918
rect 54686 19842 54738 19854
rect 55470 19906 55522 19918
rect 55470 19842 55522 19854
rect 3502 19794 3554 19806
rect 3502 19730 3554 19742
rect 8766 19794 8818 19806
rect 8766 19730 8818 19742
rect 17390 19794 17442 19806
rect 50430 19794 50482 19806
rect 23986 19742 23998 19794
rect 24050 19742 24062 19794
rect 17390 19730 17442 19742
rect 50430 19730 50482 19742
rect 55582 19794 55634 19806
rect 55582 19730 55634 19742
rect 1344 19626 58576 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 58576 19626
rect 1344 19540 58576 19574
rect 40686 19346 40738 19358
rect 14914 19294 14926 19346
rect 14978 19294 14990 19346
rect 17042 19294 17054 19346
rect 17106 19294 17118 19346
rect 40686 19282 40738 19294
rect 42142 19346 42194 19358
rect 42142 19282 42194 19294
rect 42590 19346 42642 19358
rect 42590 19282 42642 19294
rect 46958 19346 47010 19358
rect 53790 19346 53842 19358
rect 48626 19294 48638 19346
rect 48690 19294 48702 19346
rect 50754 19294 50766 19346
rect 50818 19294 50830 19346
rect 52770 19294 52782 19346
rect 52834 19294 52846 19346
rect 54786 19294 54798 19346
rect 54850 19294 54862 19346
rect 56018 19294 56030 19346
rect 56082 19294 56094 19346
rect 58146 19294 58158 19346
rect 58210 19294 58222 19346
rect 46958 19282 47010 19294
rect 53790 19282 53842 19294
rect 13470 19234 13522 19246
rect 13470 19170 13522 19182
rect 14142 19234 14194 19246
rect 27694 19234 27746 19246
rect 17714 19182 17726 19234
rect 17778 19182 17790 19234
rect 27346 19182 27358 19234
rect 27410 19182 27422 19234
rect 14142 19170 14194 19182
rect 27694 19170 27746 19182
rect 28254 19234 28306 19246
rect 28254 19170 28306 19182
rect 43038 19234 43090 19246
rect 43038 19170 43090 19182
rect 43262 19234 43314 19246
rect 43262 19170 43314 19182
rect 44942 19234 44994 19246
rect 52110 19234 52162 19246
rect 45490 19182 45502 19234
rect 45554 19182 45566 19234
rect 46610 19182 46622 19234
rect 46674 19182 46686 19234
rect 51426 19182 51438 19234
rect 51490 19182 51502 19234
rect 44942 19170 44994 19182
rect 52110 19170 52162 19182
rect 52894 19234 52946 19246
rect 52894 19170 52946 19182
rect 53230 19234 53282 19246
rect 53230 19170 53282 19182
rect 54686 19234 54738 19246
rect 55346 19182 55358 19234
rect 55410 19182 55422 19234
rect 54686 19170 54738 19182
rect 6638 19122 6690 19134
rect 31614 19122 31666 19134
rect 22530 19070 22542 19122
rect 22594 19070 22606 19122
rect 6638 19058 6690 19070
rect 31614 19058 31666 19070
rect 31950 19122 32002 19134
rect 31950 19058 32002 19070
rect 32174 19122 32226 19134
rect 32174 19058 32226 19070
rect 34750 19122 34802 19134
rect 34750 19058 34802 19070
rect 37998 19122 38050 19134
rect 37998 19058 38050 19070
rect 43598 19122 43650 19134
rect 43598 19058 43650 19070
rect 44830 19122 44882 19134
rect 52782 19122 52834 19134
rect 48290 19070 48302 19122
rect 48354 19070 48366 19122
rect 44830 19058 44882 19070
rect 52782 19058 52834 19070
rect 53118 19122 53170 19134
rect 53118 19058 53170 19070
rect 54238 19122 54290 19134
rect 54238 19058 54290 19070
rect 54462 19122 54514 19134
rect 54462 19058 54514 19070
rect 6414 19010 6466 19022
rect 6414 18946 6466 18958
rect 6526 19010 6578 19022
rect 6526 18946 6578 18958
rect 9214 19010 9266 19022
rect 9214 18946 9266 18958
rect 13582 19010 13634 19022
rect 13582 18946 13634 18958
rect 13694 19010 13746 19022
rect 13694 18946 13746 18958
rect 21758 19010 21810 19022
rect 21758 18946 21810 18958
rect 31726 19010 31778 19022
rect 31726 18946 31778 18958
rect 32622 19010 32674 19022
rect 32622 18946 32674 18958
rect 34638 19010 34690 19022
rect 34638 18946 34690 18958
rect 38222 19010 38274 19022
rect 38222 18946 38274 18958
rect 38334 19010 38386 19022
rect 38334 18946 38386 18958
rect 38446 19010 38498 19022
rect 38446 18946 38498 18958
rect 38558 19010 38610 19022
rect 38558 18946 38610 18958
rect 41246 19010 41298 19022
rect 41246 18946 41298 18958
rect 41582 19010 41634 19022
rect 41582 18946 41634 18958
rect 43486 19010 43538 19022
rect 43486 18946 43538 18958
rect 43934 19010 43986 19022
rect 47966 19010 48018 19022
rect 44258 18958 44270 19010
rect 44322 18958 44334 19010
rect 43934 18946 43986 18958
rect 47966 18946 48018 18958
rect 51998 19010 52050 19022
rect 51998 18946 52050 18958
rect 54798 19010 54850 19022
rect 54798 18946 54850 18958
rect 1344 18842 58576 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 58576 18842
rect 1344 18756 58576 18790
rect 3502 18674 3554 18686
rect 3502 18610 3554 18622
rect 16494 18674 16546 18686
rect 16494 18610 16546 18622
rect 19070 18674 19122 18686
rect 19070 18610 19122 18622
rect 26350 18674 26402 18686
rect 26350 18610 26402 18622
rect 26574 18674 26626 18686
rect 26574 18610 26626 18622
rect 45166 18674 45218 18686
rect 45166 18610 45218 18622
rect 45390 18674 45442 18686
rect 49074 18622 49086 18674
rect 49138 18622 49150 18674
rect 45390 18610 45442 18622
rect 14366 18562 14418 18574
rect 6626 18510 6638 18562
rect 6690 18510 6702 18562
rect 14366 18498 14418 18510
rect 16718 18562 16770 18574
rect 16718 18498 16770 18510
rect 18622 18562 18674 18574
rect 18622 18498 18674 18510
rect 18958 18562 19010 18574
rect 18958 18498 19010 18510
rect 32174 18562 32226 18574
rect 32174 18498 32226 18510
rect 33630 18562 33682 18574
rect 33630 18498 33682 18510
rect 38558 18562 38610 18574
rect 54462 18562 54514 18574
rect 42690 18510 42702 18562
rect 42754 18510 42766 18562
rect 44146 18510 44158 18562
rect 44210 18510 44222 18562
rect 51874 18510 51886 18562
rect 51938 18510 51950 18562
rect 38558 18498 38610 18510
rect 54462 18498 54514 18510
rect 55358 18562 55410 18574
rect 55358 18498 55410 18510
rect 3726 18450 3778 18462
rect 2818 18398 2830 18450
rect 2882 18398 2894 18450
rect 3726 18386 3778 18398
rect 4174 18450 4226 18462
rect 13470 18450 13522 18462
rect 16046 18450 16098 18462
rect 7410 18398 7422 18450
rect 7474 18398 7486 18450
rect 10210 18398 10222 18450
rect 10274 18398 10286 18450
rect 14018 18398 14030 18450
rect 14082 18398 14094 18450
rect 14690 18398 14702 18450
rect 14754 18398 14766 18450
rect 4174 18386 4226 18398
rect 13470 18386 13522 18398
rect 16046 18386 16098 18398
rect 16606 18450 16658 18462
rect 16606 18386 16658 18398
rect 17390 18450 17442 18462
rect 17390 18386 17442 18398
rect 17614 18450 17666 18462
rect 19294 18450 19346 18462
rect 17938 18398 17950 18450
rect 18002 18398 18014 18450
rect 18386 18398 18398 18450
rect 18450 18398 18462 18450
rect 17614 18386 17666 18398
rect 19294 18386 19346 18398
rect 22990 18450 23042 18462
rect 24110 18450 24162 18462
rect 23202 18398 23214 18450
rect 23266 18398 23278 18450
rect 23874 18398 23886 18450
rect 23938 18398 23950 18450
rect 22990 18386 23042 18398
rect 24110 18386 24162 18398
rect 24222 18450 24274 18462
rect 24222 18386 24274 18398
rect 24446 18450 24498 18462
rect 24446 18386 24498 18398
rect 25230 18450 25282 18462
rect 25230 18386 25282 18398
rect 32062 18450 32114 18462
rect 32062 18386 32114 18398
rect 32286 18450 32338 18462
rect 33854 18450 33906 18462
rect 37774 18450 37826 18462
rect 33506 18398 33518 18450
rect 33570 18398 33582 18450
rect 34290 18398 34302 18450
rect 34354 18398 34366 18450
rect 37538 18398 37550 18450
rect 37602 18398 37614 18450
rect 32286 18386 32338 18398
rect 33854 18386 33906 18398
rect 37774 18386 37826 18398
rect 37998 18450 38050 18462
rect 37998 18386 38050 18398
rect 38110 18450 38162 18462
rect 38110 18386 38162 18398
rect 40462 18450 40514 18462
rect 41694 18450 41746 18462
rect 42254 18450 42306 18462
rect 41234 18398 41246 18450
rect 41298 18398 41310 18450
rect 42018 18398 42030 18450
rect 42082 18398 42094 18450
rect 40462 18386 40514 18398
rect 41694 18386 41746 18398
rect 42254 18386 42306 18398
rect 42366 18450 42418 18462
rect 42366 18386 42418 18398
rect 43038 18450 43090 18462
rect 44718 18450 44770 18462
rect 43922 18398 43934 18450
rect 43986 18398 43998 18450
rect 43038 18386 43090 18398
rect 44718 18386 44770 18398
rect 45054 18450 45106 18462
rect 45054 18386 45106 18398
rect 48750 18450 48802 18462
rect 56030 18450 56082 18462
rect 51202 18398 51214 18450
rect 51266 18398 51278 18450
rect 48750 18386 48802 18398
rect 56030 18386 56082 18398
rect 3166 18338 3218 18350
rect 3166 18274 3218 18286
rect 3614 18338 3666 18350
rect 7758 18338 7810 18350
rect 14478 18338 14530 18350
rect 4498 18286 4510 18338
rect 4562 18286 4574 18338
rect 10994 18286 11006 18338
rect 11058 18286 11070 18338
rect 13122 18286 13134 18338
rect 13186 18286 13198 18338
rect 3614 18274 3666 18286
rect 7758 18274 7810 18286
rect 14478 18274 14530 18286
rect 22318 18338 22370 18350
rect 22318 18274 22370 18286
rect 22766 18338 22818 18350
rect 22766 18274 22818 18286
rect 25342 18338 25394 18350
rect 33742 18338 33794 18350
rect 37886 18338 37938 18350
rect 27010 18286 27022 18338
rect 27074 18286 27086 18338
rect 35074 18286 35086 18338
rect 35138 18286 35150 18338
rect 37202 18286 37214 18338
rect 37266 18286 37278 18338
rect 25342 18274 25394 18286
rect 33742 18274 33794 18286
rect 37886 18274 37938 18286
rect 39118 18338 39170 18350
rect 39118 18274 39170 18286
rect 45726 18338 45778 18350
rect 45726 18274 45778 18286
rect 48190 18338 48242 18350
rect 54002 18286 54014 18338
rect 54066 18286 54078 18338
rect 48190 18274 48242 18286
rect 2830 18226 2882 18238
rect 2830 18162 2882 18174
rect 7982 18226 8034 18238
rect 13694 18226 13746 18238
rect 8306 18174 8318 18226
rect 8370 18174 8382 18226
rect 7982 18162 8034 18174
rect 13694 18162 13746 18174
rect 22654 18226 22706 18238
rect 22654 18162 22706 18174
rect 23438 18226 23490 18238
rect 33182 18226 33234 18238
rect 31602 18174 31614 18226
rect 31666 18174 31678 18226
rect 23438 18162 23490 18174
rect 33182 18162 33234 18174
rect 38670 18226 38722 18238
rect 38670 18162 38722 18174
rect 54350 18226 54402 18238
rect 54350 18162 54402 18174
rect 55470 18226 55522 18238
rect 55470 18162 55522 18174
rect 1344 18058 58576 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 58576 18058
rect 1344 17972 58576 18006
rect 35422 17890 35474 17902
rect 35422 17826 35474 17838
rect 36094 17890 36146 17902
rect 36094 17826 36146 17838
rect 6750 17778 6802 17790
rect 28590 17778 28642 17790
rect 32734 17778 32786 17790
rect 2482 17726 2494 17778
rect 2546 17726 2558 17778
rect 4610 17726 4622 17778
rect 4674 17726 4686 17778
rect 19282 17726 19294 17778
rect 19346 17726 19358 17778
rect 20402 17726 20414 17778
rect 20466 17726 20478 17778
rect 23426 17726 23438 17778
rect 23490 17726 23502 17778
rect 25554 17726 25566 17778
rect 25618 17726 25630 17778
rect 32162 17726 32174 17778
rect 32226 17726 32238 17778
rect 6750 17714 6802 17726
rect 28590 17714 28642 17726
rect 32734 17714 32786 17726
rect 35534 17778 35586 17790
rect 35534 17714 35586 17726
rect 36206 17778 36258 17790
rect 42478 17778 42530 17790
rect 37314 17726 37326 17778
rect 37378 17726 37390 17778
rect 39442 17726 39454 17778
rect 39506 17726 39518 17778
rect 41906 17726 41918 17778
rect 41970 17726 41982 17778
rect 36206 17714 36258 17726
rect 42478 17714 42530 17726
rect 46958 17778 47010 17790
rect 46958 17714 47010 17726
rect 6638 17666 6690 17678
rect 1810 17614 1822 17666
rect 1874 17614 1886 17666
rect 6290 17614 6302 17666
rect 6354 17614 6366 17666
rect 6638 17602 6690 17614
rect 6862 17666 6914 17678
rect 6862 17602 6914 17614
rect 7758 17666 7810 17678
rect 18398 17666 18450 17678
rect 33630 17666 33682 17678
rect 14354 17614 14366 17666
rect 14418 17614 14430 17666
rect 17826 17614 17838 17666
rect 17890 17614 17902 17666
rect 19170 17614 19182 17666
rect 19234 17614 19246 17666
rect 22642 17614 22654 17666
rect 22706 17614 22718 17666
rect 29250 17614 29262 17666
rect 29314 17614 29326 17666
rect 7758 17602 7810 17614
rect 18398 17602 18450 17614
rect 33630 17602 33682 17614
rect 34190 17666 34242 17678
rect 41470 17666 41522 17678
rect 40226 17614 40238 17666
rect 40290 17614 40302 17666
rect 40898 17614 40910 17666
rect 40962 17614 40974 17666
rect 52882 17614 52894 17666
rect 52946 17614 52958 17666
rect 34190 17602 34242 17614
rect 41470 17602 41522 17614
rect 15038 17554 15090 17566
rect 7410 17502 7422 17554
rect 7474 17502 7486 17554
rect 14130 17502 14142 17554
rect 14194 17502 14206 17554
rect 15038 17490 15090 17502
rect 15374 17554 15426 17566
rect 15374 17490 15426 17502
rect 18062 17554 18114 17566
rect 19742 17554 19794 17566
rect 18274 17502 18286 17554
rect 18338 17502 18350 17554
rect 18062 17490 18114 17502
rect 19742 17490 19794 17502
rect 20078 17554 20130 17566
rect 20078 17490 20130 17502
rect 20302 17554 20354 17566
rect 20302 17490 20354 17502
rect 27582 17554 27634 17566
rect 27582 17490 27634 17502
rect 27806 17554 27858 17566
rect 27806 17490 27858 17502
rect 27918 17554 27970 17566
rect 41134 17554 41186 17566
rect 30034 17502 30046 17554
rect 30098 17502 30110 17554
rect 55346 17502 55358 17554
rect 55410 17502 55422 17554
rect 27918 17490 27970 17502
rect 41134 17490 41186 17502
rect 17390 17442 17442 17454
rect 17390 17378 17442 17390
rect 21422 17442 21474 17454
rect 21422 17378 21474 17390
rect 28142 17442 28194 17454
rect 28142 17378 28194 17390
rect 33742 17442 33794 17454
rect 33742 17378 33794 17390
rect 33966 17442 34018 17454
rect 33966 17378 34018 17390
rect 34302 17442 34354 17454
rect 34302 17378 34354 17390
rect 34526 17442 34578 17454
rect 34526 17378 34578 17390
rect 52110 17442 52162 17454
rect 52110 17378 52162 17390
rect 1344 17274 58576 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 58576 17274
rect 1344 17188 58576 17222
rect 15710 17106 15762 17118
rect 3266 17054 3278 17106
rect 3330 17054 3342 17106
rect 15710 17042 15762 17054
rect 23886 17106 23938 17118
rect 23886 17042 23938 17054
rect 25342 17106 25394 17118
rect 25342 17042 25394 17054
rect 41022 17106 41074 17118
rect 41022 17042 41074 17054
rect 44270 17106 44322 17118
rect 44270 17042 44322 17054
rect 44494 17106 44546 17118
rect 44494 17042 44546 17054
rect 45278 17106 45330 17118
rect 45278 17042 45330 17054
rect 46510 17106 46562 17118
rect 46510 17042 46562 17054
rect 51438 17106 51490 17118
rect 51438 17042 51490 17054
rect 51774 17106 51826 17118
rect 51774 17042 51826 17054
rect 52782 17106 52834 17118
rect 52782 17042 52834 17054
rect 22990 16994 23042 17006
rect 10210 16942 10222 16994
rect 10274 16942 10286 16994
rect 16034 16942 16046 16994
rect 16098 16942 16110 16994
rect 21522 16942 21534 16994
rect 21586 16942 21598 16994
rect 22990 16930 23042 16942
rect 23326 16994 23378 17006
rect 23326 16930 23378 16942
rect 24670 16994 24722 17006
rect 30718 16994 30770 17006
rect 46734 16994 46786 17006
rect 27906 16942 27918 16994
rect 27970 16942 27982 16994
rect 42242 16942 42254 16994
rect 42306 16942 42318 16994
rect 24670 16930 24722 16942
rect 30718 16930 30770 16942
rect 46734 16930 46786 16942
rect 47630 16994 47682 17006
rect 47630 16930 47682 16942
rect 49646 16994 49698 17006
rect 49646 16930 49698 16942
rect 3838 16882 3890 16894
rect 15262 16882 15314 16894
rect 24110 16882 24162 16894
rect 31054 16882 31106 16894
rect 41918 16882 41970 16894
rect 44942 16882 44994 16894
rect 13794 16830 13806 16882
rect 13858 16830 13870 16882
rect 22306 16830 22318 16882
rect 22370 16830 22382 16882
rect 28690 16830 28702 16882
rect 28754 16830 28766 16882
rect 31266 16830 31278 16882
rect 31330 16830 31342 16882
rect 41458 16830 41470 16882
rect 41522 16830 41534 16882
rect 42466 16830 42478 16882
rect 42530 16830 42542 16882
rect 3838 16818 3890 16830
rect 15262 16818 15314 16830
rect 24110 16818 24162 16830
rect 31054 16818 31106 16830
rect 41918 16818 41970 16830
rect 44942 16818 44994 16830
rect 46174 16882 46226 16894
rect 46174 16818 46226 16830
rect 47518 16882 47570 16894
rect 49310 16882 49362 16894
rect 47842 16830 47854 16882
rect 47906 16830 47918 16882
rect 47518 16818 47570 16830
rect 49310 16818 49362 16830
rect 52334 16882 52386 16894
rect 52334 16818 52386 16830
rect 54014 16882 54066 16894
rect 54014 16818 54066 16830
rect 3614 16770 3666 16782
rect 30830 16770 30882 16782
rect 19394 16718 19406 16770
rect 19458 16718 19470 16770
rect 25778 16718 25790 16770
rect 25842 16718 25854 16770
rect 3614 16706 3666 16718
rect 30830 16706 30882 16718
rect 44382 16770 44434 16782
rect 44382 16706 44434 16718
rect 47294 16770 47346 16782
rect 47294 16706 47346 16718
rect 46846 16658 46898 16670
rect 46846 16594 46898 16606
rect 48302 16658 48354 16670
rect 48302 16594 48354 16606
rect 53902 16658 53954 16670
rect 53902 16594 53954 16606
rect 1344 16490 58576 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 58576 16490
rect 1344 16404 58576 16438
rect 30830 16322 30882 16334
rect 30830 16258 30882 16270
rect 14702 16210 14754 16222
rect 25566 16210 25618 16222
rect 8866 16158 8878 16210
rect 8930 16158 8942 16210
rect 15474 16158 15486 16210
rect 15538 16158 15550 16210
rect 14702 16146 14754 16158
rect 25566 16146 25618 16158
rect 27022 16210 27074 16222
rect 27022 16146 27074 16158
rect 27358 16210 27410 16222
rect 31726 16210 31778 16222
rect 42030 16210 42082 16222
rect 48190 16210 48242 16222
rect 28130 16158 28142 16210
rect 28194 16158 28206 16210
rect 35970 16158 35982 16210
rect 36034 16158 36046 16210
rect 47730 16158 47742 16210
rect 47794 16158 47806 16210
rect 48850 16158 48862 16210
rect 48914 16158 48926 16210
rect 50978 16158 50990 16210
rect 51042 16158 51054 16210
rect 56018 16158 56030 16210
rect 56082 16158 56094 16210
rect 58146 16158 58158 16210
rect 58210 16158 58222 16210
rect 27358 16146 27410 16158
rect 31726 16146 31778 16158
rect 42030 16146 42082 16158
rect 48190 16146 48242 16158
rect 6750 16098 6802 16110
rect 6750 16034 6802 16046
rect 7198 16098 7250 16110
rect 7982 16098 8034 16110
rect 7746 16046 7758 16098
rect 7810 16046 7822 16098
rect 7198 16034 7250 16046
rect 7982 16034 8034 16046
rect 8094 16098 8146 16110
rect 13806 16098 13858 16110
rect 15038 16098 15090 16110
rect 11666 16046 11678 16098
rect 11730 16046 11742 16098
rect 14242 16046 14254 16098
rect 14306 16046 14318 16098
rect 8094 16034 8146 16046
rect 13806 16034 13858 16046
rect 15038 16034 15090 16046
rect 17838 16098 17890 16110
rect 17838 16034 17890 16046
rect 23886 16098 23938 16110
rect 25006 16098 25058 16110
rect 31054 16098 31106 16110
rect 38334 16098 38386 16110
rect 24322 16046 24334 16098
rect 24386 16046 24398 16098
rect 27794 16046 27806 16098
rect 27858 16046 27870 16098
rect 31266 16046 31278 16098
rect 31330 16046 31342 16098
rect 31938 16046 31950 16098
rect 32002 16046 32014 16098
rect 23886 16034 23938 16046
rect 25006 16034 25058 16046
rect 31054 16034 31106 16046
rect 38334 16034 38386 16046
rect 43934 16098 43986 16110
rect 44258 16046 44270 16098
rect 44322 16046 44334 16098
rect 44930 16046 44942 16098
rect 44994 16046 45006 16098
rect 51650 16046 51662 16098
rect 51714 16046 51726 16098
rect 52994 16046 53006 16098
rect 53058 16046 53070 16098
rect 55234 16046 55246 16098
rect 55298 16046 55310 16098
rect 43934 16034 43986 16046
rect 7422 15986 7474 15998
rect 30718 15986 30770 15998
rect 10994 15934 11006 15986
rect 11058 15934 11070 15986
rect 7422 15922 7474 15934
rect 30718 15922 30770 15934
rect 31614 15986 31666 15998
rect 31614 15922 31666 15934
rect 36430 15986 36482 15998
rect 36430 15922 36482 15934
rect 37886 15986 37938 15998
rect 37886 15922 37938 15934
rect 44046 15986 44098 15998
rect 53230 15986 53282 15998
rect 45602 15934 45614 15986
rect 45666 15934 45678 15986
rect 44046 15922 44098 15934
rect 53230 15922 53282 15934
rect 53342 15986 53394 15998
rect 54574 15986 54626 15998
rect 53778 15934 53790 15986
rect 53842 15934 53854 15986
rect 53342 15922 53394 15934
rect 54574 15922 54626 15934
rect 6974 15874 7026 15886
rect 18174 15874 18226 15886
rect 8530 15822 8542 15874
rect 8594 15822 8606 15874
rect 13458 15822 13470 15874
rect 13522 15822 13534 15874
rect 6974 15810 7026 15822
rect 18174 15810 18226 15822
rect 38110 15874 38162 15886
rect 38110 15810 38162 15822
rect 38222 15874 38274 15886
rect 38222 15810 38274 15822
rect 38446 15874 38498 15886
rect 48078 15874 48130 15886
rect 43474 15822 43486 15874
rect 43538 15822 43550 15874
rect 38446 15810 38498 15822
rect 48078 15810 48130 15822
rect 54910 15874 54962 15886
rect 54910 15810 54962 15822
rect 1344 15706 58576 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 58576 15706
rect 1344 15620 58576 15654
rect 14478 15538 14530 15550
rect 14478 15474 14530 15486
rect 29262 15538 29314 15550
rect 29262 15474 29314 15486
rect 46510 15538 46562 15550
rect 53678 15538 53730 15550
rect 49298 15486 49310 15538
rect 49362 15486 49374 15538
rect 52994 15486 53006 15538
rect 53058 15486 53070 15538
rect 46510 15474 46562 15486
rect 53678 15474 53730 15486
rect 10110 15426 10162 15438
rect 5506 15374 5518 15426
rect 5570 15374 5582 15426
rect 10110 15362 10162 15374
rect 10558 15426 10610 15438
rect 10558 15362 10610 15374
rect 14814 15426 14866 15438
rect 23662 15426 23714 15438
rect 18162 15374 18174 15426
rect 18226 15374 18238 15426
rect 14814 15362 14866 15374
rect 23662 15362 23714 15374
rect 28926 15426 28978 15438
rect 28926 15362 28978 15374
rect 29038 15426 29090 15438
rect 33630 15426 33682 15438
rect 30370 15374 30382 15426
rect 30434 15374 30446 15426
rect 29038 15362 29090 15374
rect 33630 15362 33682 15374
rect 33742 15426 33794 15438
rect 33742 15362 33794 15374
rect 34414 15426 34466 15438
rect 34414 15362 34466 15374
rect 38446 15426 38498 15438
rect 38446 15362 38498 15374
rect 52110 15426 52162 15438
rect 52110 15362 52162 15374
rect 53454 15426 53506 15438
rect 57810 15374 57822 15426
rect 57874 15374 57886 15426
rect 53454 15362 53506 15374
rect 3838 15314 3890 15326
rect 7982 15314 8034 15326
rect 4834 15262 4846 15314
rect 4898 15262 4910 15314
rect 3838 15250 3890 15262
rect 7982 15250 8034 15262
rect 8318 15314 8370 15326
rect 8318 15250 8370 15262
rect 8542 15314 8594 15326
rect 8542 15250 8594 15262
rect 9662 15314 9714 15326
rect 9662 15250 9714 15262
rect 9998 15314 10050 15326
rect 9998 15250 10050 15262
rect 13246 15314 13298 15326
rect 13246 15250 13298 15262
rect 13582 15314 13634 15326
rect 13582 15250 13634 15262
rect 13806 15314 13858 15326
rect 23774 15314 23826 15326
rect 36430 15314 36482 15326
rect 17490 15262 17502 15314
rect 17554 15262 17566 15314
rect 29586 15262 29598 15314
rect 29650 15262 29662 15314
rect 34066 15262 34078 15314
rect 34130 15262 34142 15314
rect 35970 15262 35982 15314
rect 36034 15262 36046 15314
rect 13806 15250 13858 15262
rect 23774 15250 23826 15262
rect 36430 15250 36482 15262
rect 36654 15314 36706 15326
rect 47294 15314 47346 15326
rect 48750 15314 48802 15326
rect 52670 15314 52722 15326
rect 37650 15262 37662 15314
rect 37714 15262 37726 15314
rect 46162 15262 46174 15314
rect 46226 15262 46238 15314
rect 46722 15262 46734 15314
rect 46786 15262 46798 15314
rect 47730 15262 47742 15314
rect 47794 15262 47806 15314
rect 51874 15262 51886 15314
rect 51938 15262 51950 15314
rect 36654 15250 36706 15262
rect 47294 15250 47346 15262
rect 48750 15250 48802 15262
rect 52670 15250 52722 15262
rect 53342 15314 53394 15326
rect 53342 15250 53394 15262
rect 57598 15314 57650 15326
rect 57598 15250 57650 15262
rect 58158 15314 58210 15326
rect 58158 15250 58210 15262
rect 4062 15202 4114 15214
rect 8206 15202 8258 15214
rect 7634 15150 7646 15202
rect 7698 15150 7710 15202
rect 4062 15138 4114 15150
rect 8206 15138 8258 15150
rect 9774 15202 9826 15214
rect 9774 15138 9826 15150
rect 13358 15202 13410 15214
rect 28590 15202 28642 15214
rect 34302 15202 34354 15214
rect 48190 15202 48242 15214
rect 20290 15150 20302 15202
rect 20354 15150 20366 15202
rect 32498 15150 32510 15202
rect 32562 15150 32574 15202
rect 41122 15150 41134 15202
rect 41186 15150 41198 15202
rect 13358 15138 13410 15150
rect 28590 15138 28642 15150
rect 34302 15138 34354 15150
rect 48190 15138 48242 15150
rect 48974 15202 49026 15214
rect 48974 15138 49026 15150
rect 49758 15202 49810 15214
rect 49758 15138 49810 15150
rect 52446 15202 52498 15214
rect 52446 15138 52498 15150
rect 23662 15090 23714 15102
rect 3490 15038 3502 15090
rect 3554 15038 3566 15090
rect 23662 15026 23714 15038
rect 33630 15090 33682 15102
rect 38558 15090 38610 15102
rect 35298 15038 35310 15090
rect 35362 15038 35374 15090
rect 33630 15026 33682 15038
rect 38558 15026 38610 15038
rect 1344 14922 58576 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 58576 14922
rect 1344 14836 58576 14870
rect 31278 14754 31330 14766
rect 30930 14702 30942 14754
rect 30994 14702 31006 14754
rect 31278 14690 31330 14702
rect 7646 14642 7698 14654
rect 4610 14590 4622 14642
rect 4674 14590 4686 14642
rect 7646 14578 7698 14590
rect 13918 14642 13970 14654
rect 13918 14578 13970 14590
rect 17054 14642 17106 14654
rect 31502 14642 31554 14654
rect 54338 14646 54350 14698
rect 54402 14646 54414 14698
rect 22978 14590 22990 14642
rect 23042 14590 23054 14642
rect 36978 14590 36990 14642
rect 37042 14590 37054 14642
rect 39106 14590 39118 14642
rect 39170 14590 39182 14642
rect 43810 14590 43822 14642
rect 43874 14590 43886 14642
rect 45042 14590 45054 14642
rect 45106 14590 45118 14642
rect 53666 14590 53678 14642
rect 53730 14590 53742 14642
rect 56018 14590 56030 14642
rect 56082 14590 56094 14642
rect 58146 14590 58158 14642
rect 58210 14590 58222 14642
rect 17054 14578 17106 14590
rect 31502 14578 31554 14590
rect 7534 14530 7586 14542
rect 1810 14478 1822 14530
rect 1874 14478 1886 14530
rect 7534 14466 7586 14478
rect 7758 14530 7810 14542
rect 7758 14466 7810 14478
rect 8206 14530 8258 14542
rect 14030 14530 14082 14542
rect 13458 14478 13470 14530
rect 13522 14478 13534 14530
rect 8206 14466 8258 14478
rect 14030 14466 14082 14478
rect 20526 14530 20578 14542
rect 20526 14466 20578 14478
rect 20750 14530 20802 14542
rect 35534 14530 35586 14542
rect 22866 14478 22878 14530
rect 22930 14478 22942 14530
rect 24098 14478 24110 14530
rect 24162 14478 24174 14530
rect 24994 14478 25006 14530
rect 25058 14478 25070 14530
rect 20750 14466 20802 14478
rect 35534 14466 35586 14478
rect 35982 14530 36034 14542
rect 35982 14466 36034 14478
rect 36318 14530 36370 14542
rect 50542 14530 50594 14542
rect 54574 14530 54626 14542
rect 39890 14478 39902 14530
rect 39954 14478 39966 14530
rect 40898 14478 40910 14530
rect 40962 14478 40974 14530
rect 48626 14478 48638 14530
rect 48690 14478 48702 14530
rect 53330 14478 53342 14530
rect 53394 14478 53406 14530
rect 55346 14478 55358 14530
rect 55410 14478 55422 14530
rect 36318 14466 36370 14478
rect 50542 14466 50594 14478
rect 54574 14466 54626 14478
rect 16158 14418 16210 14430
rect 2482 14366 2494 14418
rect 2546 14366 2558 14418
rect 16158 14354 16210 14366
rect 17390 14418 17442 14430
rect 17390 14354 17442 14366
rect 17502 14418 17554 14430
rect 17502 14354 17554 14366
rect 17726 14418 17778 14430
rect 17726 14354 17778 14366
rect 20190 14418 20242 14430
rect 20190 14354 20242 14366
rect 23326 14418 23378 14430
rect 23326 14354 23378 14366
rect 24334 14418 24386 14430
rect 24334 14354 24386 14366
rect 24670 14418 24722 14430
rect 24670 14354 24722 14366
rect 35198 14418 35250 14430
rect 35198 14354 35250 14366
rect 35758 14418 35810 14430
rect 35758 14354 35810 14366
rect 40462 14418 40514 14430
rect 54014 14418 54066 14430
rect 41682 14366 41694 14418
rect 41746 14366 41758 14418
rect 40462 14354 40514 14366
rect 54014 14354 54066 14366
rect 13806 14306 13858 14318
rect 13806 14242 13858 14254
rect 16270 14306 16322 14318
rect 16270 14242 16322 14254
rect 16494 14306 16546 14318
rect 16494 14242 16546 14254
rect 20526 14306 20578 14318
rect 20526 14242 20578 14254
rect 24782 14306 24834 14318
rect 24782 14242 24834 14254
rect 34974 14306 35026 14318
rect 34974 14242 35026 14254
rect 35310 14306 35362 14318
rect 35310 14242 35362 14254
rect 36094 14306 36146 14318
rect 36094 14242 36146 14254
rect 36206 14306 36258 14318
rect 36206 14242 36258 14254
rect 40574 14306 40626 14318
rect 54898 14254 54910 14306
rect 54962 14254 54974 14306
rect 40574 14242 40626 14254
rect 1344 14138 58576 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 58576 14138
rect 1344 14052 58576 14086
rect 3054 13970 3106 13982
rect 3054 13906 3106 13918
rect 3614 13970 3666 13982
rect 3614 13906 3666 13918
rect 3838 13970 3890 13982
rect 3838 13906 3890 13918
rect 4622 13970 4674 13982
rect 4622 13906 4674 13918
rect 15486 13970 15538 13982
rect 15486 13906 15538 13918
rect 15598 13970 15650 13982
rect 16718 13970 16770 13982
rect 25342 13970 25394 13982
rect 16370 13918 16382 13970
rect 16434 13918 16446 13970
rect 24658 13918 24670 13970
rect 24722 13918 24734 13970
rect 15598 13906 15650 13918
rect 16718 13906 16770 13918
rect 25342 13906 25394 13918
rect 35758 13970 35810 13982
rect 35758 13906 35810 13918
rect 41582 13970 41634 13982
rect 41582 13906 41634 13918
rect 41694 13970 41746 13982
rect 41694 13906 41746 13918
rect 51998 13970 52050 13982
rect 51998 13906 52050 13918
rect 15934 13858 15986 13870
rect 11106 13806 11118 13858
rect 11170 13806 11182 13858
rect 15934 13794 15986 13806
rect 24110 13858 24162 13870
rect 24110 13794 24162 13806
rect 25230 13858 25282 13870
rect 25230 13794 25282 13806
rect 25454 13858 25506 13870
rect 41918 13858 41970 13870
rect 29586 13806 29598 13858
rect 29650 13806 29662 13858
rect 33842 13806 33854 13858
rect 33906 13806 33918 13858
rect 34290 13806 34302 13858
rect 34354 13806 34366 13858
rect 37762 13806 37774 13858
rect 37826 13806 37838 13858
rect 25454 13794 25506 13806
rect 41918 13794 41970 13806
rect 47518 13858 47570 13870
rect 47518 13794 47570 13806
rect 50654 13858 50706 13870
rect 50654 13794 50706 13806
rect 52894 13858 52946 13870
rect 52894 13794 52946 13806
rect 55694 13858 55746 13870
rect 55694 13794 55746 13806
rect 56030 13858 56082 13870
rect 56030 13794 56082 13806
rect 13582 13746 13634 13758
rect 4162 13694 4174 13746
rect 4226 13694 4238 13746
rect 10322 13694 10334 13746
rect 10386 13694 10398 13746
rect 13582 13682 13634 13694
rect 13694 13746 13746 13758
rect 13694 13682 13746 13694
rect 15710 13746 15762 13758
rect 15710 13682 15762 13694
rect 18174 13746 18226 13758
rect 24334 13746 24386 13758
rect 23426 13694 23438 13746
rect 23490 13694 23502 13746
rect 18174 13682 18226 13694
rect 24334 13682 24386 13694
rect 26910 13746 26962 13758
rect 41358 13746 41410 13758
rect 28466 13694 28478 13746
rect 28530 13694 28542 13746
rect 34850 13694 34862 13746
rect 34914 13694 34926 13746
rect 35970 13694 35982 13746
rect 36034 13694 36046 13746
rect 37986 13694 37998 13746
rect 38050 13694 38062 13746
rect 26910 13682 26962 13694
rect 41358 13682 41410 13694
rect 41470 13746 41522 13758
rect 41470 13682 41522 13694
rect 46286 13746 46338 13758
rect 46286 13682 46338 13694
rect 46510 13746 46562 13758
rect 46510 13682 46562 13694
rect 46734 13746 46786 13758
rect 46734 13682 46786 13694
rect 48078 13746 48130 13758
rect 48078 13682 48130 13694
rect 49198 13746 49250 13758
rect 49198 13682 49250 13694
rect 49310 13746 49362 13758
rect 49310 13682 49362 13694
rect 49534 13746 49586 13758
rect 50542 13746 50594 13758
rect 49746 13694 49758 13746
rect 49810 13694 49822 13746
rect 52434 13694 52446 13746
rect 52498 13694 52510 13746
rect 52658 13694 52670 13746
rect 52722 13694 52734 13746
rect 49534 13682 49586 13694
rect 50542 13682 50594 13694
rect 3278 13634 3330 13646
rect 2930 13582 2942 13634
rect 2994 13582 3006 13634
rect 3278 13570 3330 13582
rect 3726 13634 3778 13646
rect 33518 13634 33570 13646
rect 13234 13582 13246 13634
rect 13298 13582 13310 13634
rect 19170 13582 19182 13634
rect 19234 13582 19246 13634
rect 3726 13570 3778 13582
rect 33518 13570 33570 13582
rect 42590 13634 42642 13646
rect 42590 13570 42642 13582
rect 45950 13634 46002 13646
rect 45950 13570 46002 13582
rect 46398 13634 46450 13646
rect 49422 13634 49474 13646
rect 47170 13582 47182 13634
rect 47234 13582 47246 13634
rect 46398 13570 46450 13582
rect 49422 13570 49474 13582
rect 50206 13634 50258 13646
rect 50206 13570 50258 13582
rect 51886 13634 51938 13646
rect 51886 13570 51938 13582
rect 54014 13634 54066 13646
rect 54014 13570 54066 13582
rect 42702 13522 42754 13534
rect 42702 13458 42754 13470
rect 48190 13522 48242 13534
rect 48190 13458 48242 13470
rect 50094 13522 50146 13534
rect 50094 13458 50146 13470
rect 53006 13522 53058 13534
rect 53006 13458 53058 13470
rect 1344 13354 58576 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 58576 13354
rect 1344 13268 58576 13302
rect 21310 13186 21362 13198
rect 21310 13122 21362 13134
rect 30830 13186 30882 13198
rect 30830 13122 30882 13134
rect 37886 13186 37938 13198
rect 37886 13122 37938 13134
rect 21422 13074 21474 13086
rect 29822 13074 29874 13086
rect 37102 13074 37154 13086
rect 9202 13022 9214 13074
rect 9266 13022 9278 13074
rect 18162 13022 18174 13074
rect 18226 13022 18238 13074
rect 23650 13022 23662 13074
rect 23714 13022 23726 13074
rect 25778 13022 25790 13074
rect 25842 13022 25854 13074
rect 35858 13022 35870 13074
rect 35922 13022 35934 13074
rect 21422 13010 21474 13022
rect 29822 13010 29874 13022
rect 37102 13010 37154 13022
rect 37662 13074 37714 13086
rect 37662 13010 37714 13022
rect 38670 13074 38722 13086
rect 38670 13010 38722 13022
rect 39118 13074 39170 13086
rect 39118 13010 39170 13022
rect 39902 13074 39954 13086
rect 41346 13022 41358 13074
rect 41410 13022 41422 13074
rect 56018 13022 56030 13074
rect 56082 13022 56094 13074
rect 58146 13022 58158 13074
rect 58210 13022 58222 13074
rect 39902 13010 39954 13022
rect 9998 12962 10050 12974
rect 22654 12962 22706 12974
rect 6290 12910 6302 12962
rect 6354 12910 6366 12962
rect 10322 12910 10334 12962
rect 10386 12910 10398 12962
rect 20066 12910 20078 12962
rect 20130 12910 20142 12962
rect 9998 12898 10050 12910
rect 22654 12898 22706 12910
rect 22990 12962 23042 12974
rect 27582 12962 27634 12974
rect 28254 12962 28306 12974
rect 26562 12910 26574 12962
rect 26626 12910 26638 12962
rect 27122 12910 27134 12962
rect 27186 12910 27198 12962
rect 28018 12910 28030 12962
rect 28082 12910 28094 12962
rect 22990 12898 23042 12910
rect 27582 12898 27634 12910
rect 28254 12898 28306 12910
rect 28366 12962 28418 12974
rect 28366 12898 28418 12910
rect 28590 12962 28642 12974
rect 28590 12898 28642 12910
rect 30158 12962 30210 12974
rect 30158 12898 30210 12910
rect 30718 12962 30770 12974
rect 30718 12898 30770 12910
rect 31278 12962 31330 12974
rect 31278 12898 31330 12910
rect 31614 12962 31666 12974
rect 31614 12898 31666 12910
rect 31838 12962 31890 12974
rect 31838 12898 31890 12910
rect 33854 12962 33906 12974
rect 33854 12898 33906 12910
rect 34638 12962 34690 12974
rect 50990 12962 51042 12974
rect 35074 12910 35086 12962
rect 35138 12910 35150 12962
rect 35746 12910 35758 12962
rect 35810 12910 35822 12962
rect 43474 12910 43486 12962
rect 43538 12910 43550 12962
rect 44258 12910 44270 12962
rect 44322 12910 44334 12962
rect 45266 12910 45278 12962
rect 45330 12910 45342 12962
rect 34638 12898 34690 12910
rect 50990 12898 51042 12910
rect 52670 12962 52722 12974
rect 52670 12898 52722 12910
rect 53006 12962 53058 12974
rect 53218 12910 53230 12962
rect 53282 12910 53294 12962
rect 55234 12910 55246 12962
rect 55298 12910 55310 12962
rect 53006 12898 53058 12910
rect 4510 12850 4562 12862
rect 10110 12850 10162 12862
rect 7074 12798 7086 12850
rect 7138 12798 7150 12850
rect 4510 12786 4562 12798
rect 10110 12786 10162 12798
rect 30382 12850 30434 12862
rect 30382 12786 30434 12798
rect 30830 12850 30882 12862
rect 30830 12786 30882 12798
rect 33966 12850 34018 12862
rect 52894 12850 52946 12862
rect 36082 12798 36094 12850
rect 36146 12798 36158 12850
rect 47282 12798 47294 12850
rect 47346 12798 47358 12850
rect 33966 12786 34018 12798
rect 52894 12786 52946 12798
rect 54014 12850 54066 12862
rect 54014 12786 54066 12798
rect 4286 12738 4338 12750
rect 4286 12674 4338 12686
rect 4398 12738 4450 12750
rect 21982 12738 22034 12750
rect 9538 12686 9550 12738
rect 9602 12686 9614 12738
rect 4398 12674 4450 12686
rect 21982 12674 22034 12686
rect 22766 12738 22818 12750
rect 22766 12674 22818 12686
rect 27358 12738 27410 12750
rect 27358 12674 27410 12686
rect 31726 12738 31778 12750
rect 31726 12674 31778 12686
rect 36990 12738 37042 12750
rect 40574 12738 40626 12750
rect 38210 12686 38222 12738
rect 38274 12686 38286 12738
rect 36990 12674 37042 12686
rect 40574 12674 40626 12686
rect 45054 12738 45106 12750
rect 45054 12674 45106 12686
rect 50878 12738 50930 12750
rect 50878 12674 50930 12686
rect 53678 12738 53730 12750
rect 53678 12674 53730 12686
rect 53902 12738 53954 12750
rect 53902 12674 53954 12686
rect 54462 12738 54514 12750
rect 54462 12674 54514 12686
rect 1344 12570 58576 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 58576 12570
rect 1344 12484 58576 12518
rect 9550 12402 9602 12414
rect 9550 12338 9602 12350
rect 17502 12402 17554 12414
rect 17502 12338 17554 12350
rect 41022 12402 41074 12414
rect 41022 12338 41074 12350
rect 41358 12402 41410 12414
rect 41358 12338 41410 12350
rect 42142 12402 42194 12414
rect 42142 12338 42194 12350
rect 42254 12402 42306 12414
rect 42254 12338 42306 12350
rect 42366 12402 42418 12414
rect 42366 12338 42418 12350
rect 42478 12402 42530 12414
rect 42478 12338 42530 12350
rect 43038 12402 43090 12414
rect 43038 12338 43090 12350
rect 45278 12402 45330 12414
rect 45278 12338 45330 12350
rect 45502 12402 45554 12414
rect 45502 12338 45554 12350
rect 48078 12402 48130 12414
rect 48078 12338 48130 12350
rect 48974 12402 49026 12414
rect 48974 12338 49026 12350
rect 49086 12402 49138 12414
rect 49086 12338 49138 12350
rect 49198 12402 49250 12414
rect 49198 12338 49250 12350
rect 49758 12402 49810 12414
rect 49758 12338 49810 12350
rect 49982 12402 50034 12414
rect 55022 12402 55074 12414
rect 50754 12350 50766 12402
rect 50818 12350 50830 12402
rect 50978 12350 50990 12402
rect 51042 12350 51054 12402
rect 49982 12338 50034 12350
rect 55022 12338 55074 12350
rect 12574 12290 12626 12302
rect 6290 12238 6302 12290
rect 6354 12238 6366 12290
rect 12574 12226 12626 12238
rect 14254 12290 14306 12302
rect 14254 12226 14306 12238
rect 15262 12290 15314 12302
rect 41918 12290 41970 12302
rect 19954 12238 19966 12290
rect 20018 12238 20030 12290
rect 27570 12238 27582 12290
rect 27634 12238 27646 12290
rect 15262 12226 15314 12238
rect 41918 12226 41970 12238
rect 45166 12290 45218 12302
rect 50206 12290 50258 12302
rect 55694 12290 55746 12302
rect 45826 12238 45838 12290
rect 45890 12238 45902 12290
rect 46722 12238 46734 12290
rect 46786 12238 46798 12290
rect 52098 12238 52110 12290
rect 52162 12238 52174 12290
rect 45166 12226 45218 12238
rect 50206 12226 50258 12238
rect 55694 12226 55746 12238
rect 9774 12178 9826 12190
rect 8754 12126 8766 12178
rect 8818 12126 8830 12178
rect 9774 12114 9826 12126
rect 10222 12178 10274 12190
rect 10222 12114 10274 12126
rect 12238 12178 12290 12190
rect 12238 12114 12290 12126
rect 12798 12178 12850 12190
rect 12798 12114 12850 12126
rect 14590 12178 14642 12190
rect 15598 12178 15650 12190
rect 14914 12126 14926 12178
rect 14978 12126 14990 12178
rect 14590 12114 14642 12126
rect 15598 12114 15650 12126
rect 15710 12178 15762 12190
rect 15710 12114 15762 12126
rect 15934 12178 15986 12190
rect 41134 12178 41186 12190
rect 49310 12178 49362 12190
rect 52782 12178 52834 12190
rect 16146 12126 16158 12178
rect 16210 12126 16222 12178
rect 19170 12126 19182 12178
rect 19234 12126 19246 12178
rect 26786 12126 26798 12178
rect 26850 12126 26862 12178
rect 39666 12126 39678 12178
rect 39730 12126 39742 12178
rect 41570 12126 41582 12178
rect 41634 12126 41646 12178
rect 45938 12126 45950 12178
rect 46002 12126 46014 12178
rect 46610 12126 46622 12178
rect 46674 12126 46686 12178
rect 47506 12126 47518 12178
rect 47570 12126 47582 12178
rect 48738 12126 48750 12178
rect 48802 12126 48814 12178
rect 51202 12126 51214 12178
rect 51266 12126 51278 12178
rect 51762 12126 51774 12178
rect 51826 12126 51838 12178
rect 15934 12114 15986 12126
rect 41134 12114 41186 12126
rect 49310 12114 49362 12126
rect 52782 12114 52834 12126
rect 53006 12178 53058 12190
rect 53006 12114 53058 12126
rect 54462 12178 54514 12190
rect 54462 12114 54514 12126
rect 54574 12178 54626 12190
rect 54574 12114 54626 12126
rect 55358 12178 55410 12190
rect 55358 12114 55410 12126
rect 9662 12066 9714 12078
rect 9662 12002 9714 12014
rect 12350 12066 12402 12078
rect 12350 12002 12402 12014
rect 17614 12066 17666 12078
rect 40014 12066 40066 12078
rect 22082 12014 22094 12066
rect 22146 12014 22158 12066
rect 29698 12014 29710 12066
rect 29762 12014 29774 12066
rect 34626 12014 34638 12066
rect 34690 12014 34702 12066
rect 17614 12002 17666 12014
rect 40014 12002 40066 12014
rect 41246 12066 41298 12078
rect 41246 12002 41298 12014
rect 49870 12066 49922 12078
rect 49870 12002 49922 12014
rect 14926 11954 14978 11966
rect 14926 11890 14978 11902
rect 40126 11954 40178 11966
rect 53902 11954 53954 11966
rect 53330 11902 53342 11954
rect 53394 11902 53406 11954
rect 40126 11890 40178 11902
rect 53902 11890 53954 11902
rect 54014 11954 54066 11966
rect 54014 11890 54066 11902
rect 54238 11954 54290 11966
rect 54238 11890 54290 11902
rect 1344 11786 58576 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 58576 11786
rect 1344 11700 58576 11734
rect 45502 11618 45554 11630
rect 8978 11566 8990 11618
rect 9042 11615 9054 11618
rect 9650 11615 9662 11618
rect 9042 11569 9662 11615
rect 9042 11566 9054 11569
rect 9650 11566 9662 11569
rect 9714 11566 9726 11618
rect 45502 11554 45554 11566
rect 46958 11618 47010 11630
rect 46958 11554 47010 11566
rect 5742 11506 5794 11518
rect 2482 11454 2494 11506
rect 2546 11454 2558 11506
rect 4610 11454 4622 11506
rect 4674 11454 4686 11506
rect 5742 11442 5794 11454
rect 6638 11506 6690 11518
rect 6638 11442 6690 11454
rect 8430 11506 8482 11518
rect 13582 11506 13634 11518
rect 42814 11506 42866 11518
rect 10770 11454 10782 11506
rect 10834 11454 10846 11506
rect 12898 11454 12910 11506
rect 12962 11454 12974 11506
rect 16146 11454 16158 11506
rect 16210 11454 16222 11506
rect 18274 11454 18286 11506
rect 18338 11454 18350 11506
rect 24210 11454 24222 11506
rect 24274 11454 24286 11506
rect 25106 11454 25118 11506
rect 25170 11454 25182 11506
rect 31826 11454 31838 11506
rect 31890 11454 31902 11506
rect 33954 11454 33966 11506
rect 34018 11454 34030 11506
rect 37986 11454 37998 11506
rect 38050 11454 38062 11506
rect 40114 11454 40126 11506
rect 40178 11454 40190 11506
rect 8430 11442 8482 11454
rect 13582 11442 13634 11454
rect 42814 11442 42866 11454
rect 45726 11506 45778 11518
rect 45726 11442 45778 11454
rect 46062 11506 46114 11518
rect 46062 11442 46114 11454
rect 47070 11506 47122 11518
rect 47070 11442 47122 11454
rect 51998 11506 52050 11518
rect 55234 11454 55246 11506
rect 55298 11454 55310 11506
rect 57362 11454 57374 11506
rect 57426 11454 57438 11506
rect 51998 11442 52050 11454
rect 5854 11394 5906 11406
rect 1810 11342 1822 11394
rect 1874 11342 1886 11394
rect 5854 11330 5906 11342
rect 6302 11394 6354 11406
rect 6302 11330 6354 11342
rect 8318 11394 8370 11406
rect 8318 11330 8370 11342
rect 8654 11394 8706 11406
rect 8654 11330 8706 11342
rect 8878 11394 8930 11406
rect 13470 11394 13522 11406
rect 10098 11342 10110 11394
rect 10162 11342 10174 11394
rect 8878 11330 8930 11342
rect 13470 11330 13522 11342
rect 13694 11394 13746 11406
rect 13694 11330 13746 11342
rect 14590 11394 14642 11406
rect 41918 11394 41970 11406
rect 15474 11342 15486 11394
rect 15538 11342 15550 11394
rect 21298 11342 21310 11394
rect 21362 11342 21374 11394
rect 24770 11342 24782 11394
rect 24834 11342 24846 11394
rect 31154 11342 31166 11394
rect 31218 11342 31230 11394
rect 40898 11342 40910 11394
rect 40962 11342 40974 11394
rect 14590 11330 14642 11342
rect 41918 11330 41970 11342
rect 45950 11394 46002 11406
rect 48190 11394 48242 11406
rect 47282 11342 47294 11394
rect 47346 11342 47358 11394
rect 49634 11342 49646 11394
rect 49698 11342 49710 11394
rect 50194 11342 50206 11394
rect 50258 11342 50270 11394
rect 50978 11342 50990 11394
rect 51042 11342 51054 11394
rect 53106 11342 53118 11394
rect 53170 11342 53182 11394
rect 53554 11342 53566 11394
rect 53618 11342 53630 11394
rect 58034 11342 58046 11394
rect 58098 11342 58110 11394
rect 45950 11330 46002 11342
rect 48190 11330 48242 11342
rect 5630 11282 5682 11294
rect 5630 11218 5682 11230
rect 13918 11282 13970 11294
rect 13918 11218 13970 11230
rect 14478 11282 14530 11294
rect 26462 11282 26514 11294
rect 22082 11230 22094 11282
rect 22146 11230 22158 11282
rect 14478 11218 14530 11230
rect 26462 11218 26514 11230
rect 42254 11282 42306 11294
rect 42254 11218 42306 11230
rect 42478 11282 42530 11294
rect 42478 11218 42530 11230
rect 48078 11282 48130 11294
rect 48078 11218 48130 11230
rect 49422 11282 49474 11294
rect 51438 11282 51490 11294
rect 50866 11230 50878 11282
rect 50930 11230 50942 11282
rect 53666 11230 53678 11282
rect 53730 11230 53742 11282
rect 49422 11218 49474 11230
rect 51438 11218 51490 11230
rect 9326 11170 9378 11182
rect 9326 11106 9378 11118
rect 14254 11170 14306 11182
rect 14254 11106 14306 11118
rect 25678 11170 25730 11182
rect 25678 11106 25730 11118
rect 26574 11170 26626 11182
rect 26574 11106 26626 11118
rect 42030 11170 42082 11182
rect 42030 11106 42082 11118
rect 42142 11170 42194 11182
rect 42142 11106 42194 11118
rect 42926 11170 42978 11182
rect 42926 11106 42978 11118
rect 46174 11170 46226 11182
rect 46174 11106 46226 11118
rect 47854 11170 47906 11182
rect 47854 11106 47906 11118
rect 51326 11170 51378 11182
rect 51326 11106 51378 11118
rect 52110 11170 52162 11182
rect 52770 11118 52782 11170
rect 52834 11118 52846 11170
rect 52994 11118 53006 11170
rect 53058 11118 53070 11170
rect 52110 11106 52162 11118
rect 1344 11002 58576 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 58576 11002
rect 1344 10916 58576 10950
rect 5518 10834 5570 10846
rect 4162 10782 4174 10834
rect 4226 10782 4238 10834
rect 5518 10770 5570 10782
rect 6638 10834 6690 10846
rect 6638 10770 6690 10782
rect 23662 10834 23714 10846
rect 38222 10834 38274 10846
rect 37426 10782 37438 10834
rect 37490 10782 37502 10834
rect 23662 10770 23714 10782
rect 38222 10770 38274 10782
rect 53566 10834 53618 10846
rect 53566 10770 53618 10782
rect 14254 10722 14306 10734
rect 14254 10658 14306 10670
rect 15598 10722 15650 10734
rect 15598 10658 15650 10670
rect 23102 10722 23154 10734
rect 23102 10658 23154 10670
rect 24110 10722 24162 10734
rect 49758 10722 49810 10734
rect 35186 10670 35198 10722
rect 35250 10670 35262 10722
rect 41570 10670 41582 10722
rect 41634 10670 41646 10722
rect 24110 10658 24162 10670
rect 49758 10658 49810 10670
rect 50094 10722 50146 10734
rect 50094 10658 50146 10670
rect 50318 10722 50370 10734
rect 50318 10658 50370 10670
rect 4510 10610 4562 10622
rect 4510 10546 4562 10558
rect 4734 10610 4786 10622
rect 4734 10546 4786 10558
rect 5630 10610 5682 10622
rect 5630 10546 5682 10558
rect 5742 10610 5794 10622
rect 5742 10546 5794 10558
rect 6190 10610 6242 10622
rect 6190 10546 6242 10558
rect 14030 10610 14082 10622
rect 14030 10546 14082 10558
rect 14366 10610 14418 10622
rect 14366 10546 14418 10558
rect 14814 10610 14866 10622
rect 14814 10546 14866 10558
rect 15038 10610 15090 10622
rect 15038 10546 15090 10558
rect 15262 10610 15314 10622
rect 22542 10610 22594 10622
rect 18946 10558 18958 10610
rect 19010 10558 19022 10610
rect 15262 10546 15314 10558
rect 22542 10546 22594 10558
rect 22654 10610 22706 10622
rect 22654 10546 22706 10558
rect 22878 10610 22930 10622
rect 23886 10610 23938 10622
rect 39342 10610 39394 10622
rect 23426 10558 23438 10610
rect 23490 10558 23502 10610
rect 28130 10558 28142 10610
rect 28194 10558 28206 10610
rect 29362 10558 29374 10610
rect 29426 10558 29438 10610
rect 34514 10558 34526 10610
rect 34578 10558 34590 10610
rect 38994 10558 39006 10610
rect 39058 10558 39070 10610
rect 22878 10546 22930 10558
rect 23886 10546 23938 10558
rect 39342 10546 39394 10558
rect 40014 10610 40066 10622
rect 46846 10610 46898 10622
rect 45602 10558 45614 10610
rect 45666 10558 45678 10610
rect 40014 10546 40066 10558
rect 46846 10546 46898 10558
rect 47182 10610 47234 10622
rect 47182 10546 47234 10558
rect 47630 10610 47682 10622
rect 47630 10546 47682 10558
rect 18510 10498 18562 10510
rect 22766 10498 22818 10510
rect 19618 10446 19630 10498
rect 19682 10446 19694 10498
rect 21746 10446 21758 10498
rect 21810 10446 21822 10498
rect 18510 10434 18562 10446
rect 22766 10434 22818 10446
rect 23774 10498 23826 10510
rect 48862 10498 48914 10510
rect 25330 10446 25342 10498
rect 25394 10446 25406 10498
rect 27458 10446 27470 10498
rect 27522 10446 27534 10498
rect 30146 10446 30158 10498
rect 30210 10446 30222 10498
rect 32274 10446 32286 10498
rect 32338 10446 32350 10498
rect 23774 10434 23826 10446
rect 48862 10434 48914 10446
rect 49870 10498 49922 10510
rect 49870 10434 49922 10446
rect 53678 10498 53730 10510
rect 53678 10434 53730 10446
rect 47406 10386 47458 10398
rect 39442 10334 39454 10386
rect 39506 10334 39518 10386
rect 47406 10322 47458 10334
rect 48078 10386 48130 10398
rect 48078 10322 48130 10334
rect 48750 10386 48802 10398
rect 48750 10322 48802 10334
rect 53790 10386 53842 10398
rect 53790 10322 53842 10334
rect 1344 10218 58576 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 58576 10218
rect 1344 10132 58576 10166
rect 19966 10050 20018 10062
rect 19966 9986 20018 9998
rect 20302 10050 20354 10062
rect 20302 9986 20354 9998
rect 22206 10050 22258 10062
rect 27806 10050 27858 10062
rect 26786 9998 26798 10050
rect 26850 9998 26862 10050
rect 47730 9998 47742 10050
rect 47794 9998 47806 10050
rect 22206 9986 22258 9998
rect 27806 9986 27858 9998
rect 5630 9938 5682 9950
rect 20750 9938 20802 9950
rect 5058 9886 5070 9938
rect 5122 9886 5134 9938
rect 7298 9886 7310 9938
rect 7362 9886 7374 9938
rect 5630 9874 5682 9886
rect 20750 9874 20802 9886
rect 22094 9938 22146 9950
rect 22094 9874 22146 9886
rect 30158 9938 30210 9950
rect 30158 9874 30210 9886
rect 37998 9938 38050 9950
rect 49410 9886 49422 9938
rect 49474 9886 49486 9938
rect 55458 9886 55470 9938
rect 55522 9886 55534 9938
rect 37998 9874 38050 9886
rect 5854 9826 5906 9838
rect 19070 9826 19122 9838
rect 26238 9826 26290 9838
rect 2146 9774 2158 9826
rect 2210 9774 2222 9826
rect 6850 9774 6862 9826
rect 6914 9774 6926 9826
rect 10098 9774 10110 9826
rect 10162 9774 10174 9826
rect 14914 9774 14926 9826
rect 14978 9774 14990 9826
rect 21858 9774 21870 9826
rect 21922 9774 21934 9826
rect 5854 9762 5906 9774
rect 19070 9762 19122 9774
rect 26238 9762 26290 9774
rect 26574 9826 26626 9838
rect 29822 9826 29874 9838
rect 27010 9774 27022 9826
rect 27074 9774 27086 9826
rect 26574 9762 26626 9774
rect 29822 9762 29874 9774
rect 30046 9826 30098 9838
rect 30046 9762 30098 9774
rect 30382 9826 30434 9838
rect 30382 9762 30434 9774
rect 30606 9826 30658 9838
rect 37662 9826 37714 9838
rect 31378 9774 31390 9826
rect 31442 9774 31454 9826
rect 30606 9762 30658 9774
rect 37662 9762 37714 9774
rect 38334 9826 38386 9838
rect 38334 9762 38386 9774
rect 39230 9826 39282 9838
rect 39230 9762 39282 9774
rect 39454 9826 39506 9838
rect 39454 9762 39506 9774
rect 39566 9826 39618 9838
rect 39566 9762 39618 9774
rect 41022 9826 41074 9838
rect 41022 9762 41074 9774
rect 42590 9826 42642 9838
rect 42590 9762 42642 9774
rect 47406 9826 47458 9838
rect 49870 9826 49922 9838
rect 47954 9774 47966 9826
rect 48018 9774 48030 9826
rect 48514 9774 48526 9826
rect 48578 9774 48590 9826
rect 48850 9774 48862 9826
rect 48914 9774 48926 9826
rect 47406 9762 47458 9774
rect 49870 9762 49922 9774
rect 50542 9826 50594 9838
rect 50542 9762 50594 9774
rect 52110 9826 52162 9838
rect 52882 9774 52894 9826
rect 52946 9774 52958 9826
rect 52110 9762 52162 9774
rect 28142 9714 28194 9726
rect 2930 9662 2942 9714
rect 2994 9662 3006 9714
rect 6178 9662 6190 9714
rect 6242 9662 6254 9714
rect 9426 9662 9438 9714
rect 9490 9662 9502 9714
rect 17378 9662 17390 9714
rect 17442 9662 17454 9714
rect 28142 9650 28194 9662
rect 30718 9714 30770 9726
rect 30718 9650 30770 9662
rect 30830 9714 30882 9726
rect 30830 9650 30882 9662
rect 30942 9714 30994 9726
rect 30942 9650 30994 9662
rect 33966 9714 34018 9726
rect 33966 9650 34018 9662
rect 34302 9714 34354 9726
rect 34302 9650 34354 9662
rect 41470 9714 41522 9726
rect 42242 9662 42254 9714
rect 42306 9662 42318 9714
rect 41470 9650 41522 9662
rect 6638 9602 6690 9614
rect 20078 9602 20130 9614
rect 27918 9602 27970 9614
rect 19394 9550 19406 9602
rect 19458 9550 19470 9602
rect 26674 9550 26686 9602
rect 26738 9550 26750 9602
rect 6638 9538 6690 9550
rect 20078 9538 20130 9550
rect 27918 9538 27970 9550
rect 28590 9602 28642 9614
rect 28590 9538 28642 9550
rect 34190 9602 34242 9614
rect 39118 9602 39170 9614
rect 38658 9550 38670 9602
rect 38722 9550 38734 9602
rect 34190 9538 34242 9550
rect 39118 9538 39170 9550
rect 39342 9602 39394 9614
rect 39342 9538 39394 9550
rect 40910 9602 40962 9614
rect 40910 9538 40962 9550
rect 41134 9602 41186 9614
rect 41134 9538 41186 9550
rect 41246 9602 41298 9614
rect 41246 9538 41298 9550
rect 49982 9602 50034 9614
rect 49982 9538 50034 9550
rect 50094 9602 50146 9614
rect 50094 9538 50146 9550
rect 1344 9434 58576 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 58576 9434
rect 1344 9348 58576 9382
rect 6078 9266 6130 9278
rect 6078 9202 6130 9214
rect 7310 9266 7362 9278
rect 7310 9202 7362 9214
rect 8654 9266 8706 9278
rect 8654 9202 8706 9214
rect 9662 9266 9714 9278
rect 9662 9202 9714 9214
rect 10670 9266 10722 9278
rect 10670 9202 10722 9214
rect 12238 9266 12290 9278
rect 16270 9266 16322 9278
rect 14802 9214 14814 9266
rect 14866 9214 14878 9266
rect 12238 9202 12290 9214
rect 16270 9202 16322 9214
rect 25454 9266 25506 9278
rect 25454 9202 25506 9214
rect 28814 9266 28866 9278
rect 28814 9202 28866 9214
rect 29262 9266 29314 9278
rect 29262 9202 29314 9214
rect 30382 9266 30434 9278
rect 30382 9202 30434 9214
rect 49086 9266 49138 9278
rect 49086 9202 49138 9214
rect 49758 9266 49810 9278
rect 49758 9202 49810 9214
rect 49870 9266 49922 9278
rect 49870 9202 49922 9214
rect 51326 9266 51378 9278
rect 51326 9202 51378 9214
rect 52782 9266 52834 9278
rect 52782 9202 52834 9214
rect 57598 9266 57650 9278
rect 58158 9266 58210 9278
rect 57810 9214 57822 9266
rect 57874 9214 57886 9266
rect 57598 9202 57650 9214
rect 58158 9202 58210 9214
rect 5966 9154 6018 9166
rect 5966 9090 6018 9102
rect 7198 9154 7250 9166
rect 7198 9090 7250 9102
rect 8766 9154 8818 9166
rect 8766 9090 8818 9102
rect 8990 9154 9042 9166
rect 8990 9090 9042 9102
rect 9774 9154 9826 9166
rect 29150 9154 29202 9166
rect 16482 9102 16494 9154
rect 16546 9102 16558 9154
rect 18162 9102 18174 9154
rect 18226 9102 18238 9154
rect 9774 9090 9826 9102
rect 29150 9090 29202 9102
rect 40126 9154 40178 9166
rect 40126 9090 40178 9102
rect 41246 9154 41298 9166
rect 48078 9154 48130 9166
rect 43698 9102 43710 9154
rect 43762 9102 43774 9154
rect 41246 9090 41298 9102
rect 48078 9090 48130 9102
rect 49982 9154 50034 9166
rect 49982 9090 50034 9102
rect 52894 9154 52946 9166
rect 52894 9090 52946 9102
rect 56926 9154 56978 9166
rect 56926 9090 56978 9102
rect 8430 9042 8482 9054
rect 6290 8990 6302 9042
rect 6354 8990 6366 9042
rect 8430 8978 8482 8990
rect 9550 9042 9602 9054
rect 9550 8978 9602 8990
rect 10222 9042 10274 9054
rect 15150 9042 15202 9054
rect 29486 9042 29538 9054
rect 46174 9042 46226 9054
rect 12562 8990 12574 9042
rect 12626 8990 12638 9042
rect 14018 8990 14030 9042
rect 14082 8990 14094 9042
rect 16706 8990 16718 9042
rect 16770 8990 16782 9042
rect 17378 8990 17390 9042
rect 17442 8990 17454 9042
rect 20962 8990 20974 9042
rect 21026 8990 21038 9042
rect 36194 8990 36206 9042
rect 36258 8990 36270 9042
rect 36530 8990 36542 9042
rect 36594 8990 36606 9042
rect 42914 8990 42926 9042
rect 42978 8990 42990 9042
rect 10222 8978 10274 8990
rect 15150 8978 15202 8990
rect 29486 8978 29538 8990
rect 46174 8978 46226 8990
rect 48190 9042 48242 9054
rect 48190 8978 48242 8990
rect 48750 9042 48802 9054
rect 48750 8978 48802 8990
rect 48974 9042 49026 9054
rect 48974 8978 49026 8990
rect 49422 9042 49474 9054
rect 51214 9042 51266 9054
rect 50978 8990 50990 9042
rect 51042 8990 51054 9042
rect 49422 8978 49474 8990
rect 51214 8978 51266 8990
rect 51438 9042 51490 9054
rect 53006 9042 53058 9054
rect 51650 8990 51662 9042
rect 51714 8990 51726 9042
rect 51438 8978 51490 8990
rect 53006 8978 53058 8990
rect 53230 9042 53282 9054
rect 53230 8978 53282 8990
rect 53454 9042 53506 9054
rect 54238 9042 54290 9054
rect 53778 8990 53790 9042
rect 53842 8990 53854 9042
rect 53454 8978 53506 8990
rect 54238 8978 54290 8990
rect 54574 9042 54626 9054
rect 54574 8978 54626 8990
rect 55246 9042 55298 9054
rect 55246 8978 55298 8990
rect 55470 9042 55522 9054
rect 55470 8978 55522 8990
rect 56590 9042 56642 9054
rect 56590 8978 56642 8990
rect 12910 8930 12962 8942
rect 12910 8866 12962 8878
rect 13470 8930 13522 8942
rect 15598 8930 15650 8942
rect 20750 8930 20802 8942
rect 52334 8930 52386 8942
rect 14242 8878 14254 8930
rect 14306 8878 14318 8930
rect 20290 8878 20302 8930
rect 20354 8878 20366 8930
rect 33282 8878 33294 8930
rect 33346 8878 33358 8930
rect 35410 8878 35422 8930
rect 35474 8878 35486 8930
rect 37314 8878 37326 8930
rect 37378 8878 37390 8930
rect 39442 8878 39454 8930
rect 39506 8878 39518 8930
rect 45826 8878 45838 8930
rect 45890 8878 45902 8930
rect 13470 8866 13522 8878
rect 15598 8866 15650 8878
rect 20750 8866 20802 8878
rect 52334 8866 52386 8878
rect 7310 8818 7362 8830
rect 7310 8754 7362 8766
rect 12574 8818 12626 8830
rect 12574 8754 12626 8766
rect 20638 8818 20690 8830
rect 20638 8754 20690 8766
rect 40238 8818 40290 8830
rect 40238 8754 40290 8766
rect 41358 8818 41410 8830
rect 41358 8754 41410 8766
rect 46286 8818 46338 8830
rect 46286 8754 46338 8766
rect 54014 8818 54066 8830
rect 54014 8754 54066 8766
rect 54462 8818 54514 8830
rect 54898 8766 54910 8818
rect 54962 8766 54974 8818
rect 54462 8754 54514 8766
rect 1344 8650 58576 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 58576 8650
rect 1344 8564 58576 8598
rect 37998 8482 38050 8494
rect 37998 8418 38050 8430
rect 47182 8482 47234 8494
rect 47182 8418 47234 8430
rect 47630 8482 47682 8494
rect 47630 8418 47682 8430
rect 8654 8370 8706 8382
rect 26462 8370 26514 8382
rect 38110 8370 38162 8382
rect 17266 8318 17278 8370
rect 17330 8318 17342 8370
rect 19394 8318 19406 8370
rect 19458 8318 19470 8370
rect 24210 8318 24222 8370
rect 24274 8318 24286 8370
rect 35074 8318 35086 8370
rect 35138 8318 35150 8370
rect 8654 8306 8706 8318
rect 26462 8306 26514 8318
rect 38110 8306 38162 8318
rect 40462 8370 40514 8382
rect 49758 8370 49810 8382
rect 42130 8318 42142 8370
rect 42194 8318 42206 8370
rect 44258 8318 44270 8370
rect 44322 8318 44334 8370
rect 40462 8306 40514 8318
rect 49758 8306 49810 8318
rect 50318 8370 50370 8382
rect 54002 8318 54014 8370
rect 54066 8318 54078 8370
rect 55234 8318 55246 8370
rect 55298 8318 55310 8370
rect 57362 8318 57374 8370
rect 57426 8318 57438 8370
rect 50318 8306 50370 8318
rect 25790 8258 25842 8270
rect 9202 8206 9214 8258
rect 9266 8206 9278 8258
rect 20178 8206 20190 8258
rect 20242 8206 20254 8258
rect 21298 8206 21310 8258
rect 21362 8206 21374 8258
rect 24770 8206 24782 8258
rect 24834 8206 24846 8258
rect 25554 8206 25566 8258
rect 25618 8206 25630 8258
rect 25790 8194 25842 8206
rect 33966 8258 34018 8270
rect 33966 8194 34018 8206
rect 34750 8258 34802 8270
rect 41458 8206 41470 8258
rect 41522 8206 41534 8258
rect 49970 8206 49982 8258
rect 50034 8206 50046 8258
rect 52882 8206 52894 8258
rect 52946 8206 52958 8258
rect 53890 8206 53902 8258
rect 53954 8206 53966 8258
rect 58034 8206 58046 8258
rect 58098 8206 58110 8258
rect 34750 8194 34802 8206
rect 8990 8146 9042 8158
rect 25902 8146 25954 8158
rect 8754 8094 8766 8146
rect 8818 8094 8830 8146
rect 22082 8094 22094 8146
rect 22146 8094 22158 8146
rect 8990 8082 9042 8094
rect 25902 8082 25954 8094
rect 33854 8146 33906 8158
rect 33854 8082 33906 8094
rect 34190 8146 34242 8158
rect 34190 8082 34242 8094
rect 34414 8146 34466 8158
rect 34414 8082 34466 8094
rect 46846 8146 46898 8158
rect 46846 8082 46898 8094
rect 47518 8146 47570 8158
rect 54462 8146 54514 8158
rect 53106 8094 53118 8146
rect 53170 8094 53182 8146
rect 47518 8082 47570 8094
rect 54462 8082 54514 8094
rect 54910 8146 54962 8158
rect 54910 8082 54962 8094
rect 9662 8034 9714 8046
rect 30270 8034 30322 8046
rect 34974 8034 35026 8046
rect 24546 7982 24558 8034
rect 24610 7982 24622 8034
rect 30594 7982 30606 8034
rect 30658 7982 30670 8034
rect 9662 7970 9714 7982
rect 30270 7970 30322 7982
rect 34974 7970 35026 7982
rect 47070 8034 47122 8046
rect 47070 7970 47122 7982
rect 47630 8034 47682 8046
rect 47630 7970 47682 7982
rect 49646 8034 49698 8046
rect 49646 7970 49698 7982
rect 49870 8034 49922 8046
rect 49870 7970 49922 7982
rect 1344 7866 58576 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 58576 7866
rect 1344 7780 58576 7814
rect 25454 7698 25506 7710
rect 25454 7634 25506 7646
rect 26014 7698 26066 7710
rect 26014 7634 26066 7646
rect 26126 7698 26178 7710
rect 26126 7634 26178 7646
rect 29822 7698 29874 7710
rect 29822 7634 29874 7646
rect 35646 7698 35698 7710
rect 35646 7634 35698 7646
rect 39902 7698 39954 7710
rect 39902 7634 39954 7646
rect 40014 7698 40066 7710
rect 40014 7634 40066 7646
rect 41358 7698 41410 7710
rect 41358 7634 41410 7646
rect 42702 7698 42754 7710
rect 42702 7634 42754 7646
rect 43598 7698 43650 7710
rect 43598 7634 43650 7646
rect 46062 7698 46114 7710
rect 49982 7698 50034 7710
rect 46946 7646 46958 7698
rect 47010 7646 47022 7698
rect 46062 7634 46114 7646
rect 49982 7634 50034 7646
rect 9998 7586 10050 7598
rect 9998 7522 10050 7534
rect 10334 7586 10386 7598
rect 27134 7586 27186 7598
rect 12002 7534 12014 7586
rect 12066 7534 12078 7586
rect 20178 7534 20190 7586
rect 20242 7534 20254 7586
rect 10334 7522 10386 7534
rect 27134 7522 27186 7534
rect 30270 7586 30322 7598
rect 30270 7522 30322 7534
rect 30606 7586 30658 7598
rect 30606 7522 30658 7534
rect 31726 7586 31778 7598
rect 31726 7522 31778 7534
rect 39230 7586 39282 7598
rect 39230 7522 39282 7534
rect 41134 7586 41186 7598
rect 53118 7586 53170 7598
rect 47058 7534 47070 7586
rect 47122 7534 47134 7586
rect 41134 7522 41186 7534
rect 53118 7522 53170 7534
rect 53230 7586 53282 7598
rect 53230 7522 53282 7534
rect 53342 7586 53394 7598
rect 53342 7522 53394 7534
rect 53790 7586 53842 7598
rect 53790 7522 53842 7534
rect 54014 7586 54066 7598
rect 54014 7522 54066 7534
rect 54350 7586 54402 7598
rect 54350 7522 54402 7534
rect 56926 7586 56978 7598
rect 56926 7522 56978 7534
rect 7310 7474 7362 7486
rect 25902 7474 25954 7486
rect 7746 7422 7758 7474
rect 7810 7422 7822 7474
rect 11218 7422 11230 7474
rect 11282 7422 11294 7474
rect 24658 7422 24670 7474
rect 24722 7422 24734 7474
rect 7310 7410 7362 7422
rect 25902 7410 25954 7422
rect 26238 7474 26290 7486
rect 26910 7474 26962 7486
rect 26450 7422 26462 7474
rect 26514 7422 26526 7474
rect 26238 7410 26290 7422
rect 26910 7410 26962 7422
rect 29486 7474 29538 7486
rect 29486 7410 29538 7422
rect 30830 7474 30882 7486
rect 30830 7410 30882 7422
rect 31614 7474 31666 7486
rect 34862 7474 34914 7486
rect 31938 7422 31950 7474
rect 32002 7422 32014 7474
rect 31614 7410 31666 7422
rect 34862 7410 34914 7422
rect 39678 7474 39730 7486
rect 39678 7410 39730 7422
rect 39790 7474 39842 7486
rect 45950 7474 46002 7486
rect 40226 7422 40238 7474
rect 40290 7422 40302 7474
rect 40898 7422 40910 7474
rect 40962 7422 40974 7474
rect 41570 7422 41582 7474
rect 41634 7422 41646 7474
rect 39790 7410 39842 7422
rect 45950 7410 46002 7422
rect 46398 7474 46450 7486
rect 46398 7410 46450 7422
rect 46622 7474 46674 7486
rect 46622 7410 46674 7422
rect 46846 7474 46898 7486
rect 46846 7410 46898 7422
rect 47406 7474 47458 7486
rect 47406 7410 47458 7422
rect 50094 7474 50146 7486
rect 50094 7410 50146 7422
rect 55022 7474 55074 7486
rect 56590 7474 56642 7486
rect 55346 7422 55358 7474
rect 55410 7422 55422 7474
rect 55022 7410 55074 7422
rect 56590 7410 56642 7422
rect 8206 7362 8258 7374
rect 19070 7362 19122 7374
rect 14130 7310 14142 7362
rect 14194 7310 14206 7362
rect 8206 7298 8258 7310
rect 19070 7298 19122 7310
rect 29710 7362 29762 7374
rect 29710 7298 29762 7310
rect 30382 7362 30434 7374
rect 34638 7362 34690 7374
rect 42254 7362 42306 7374
rect 31154 7310 31166 7362
rect 31218 7310 31230 7362
rect 41122 7310 41134 7362
rect 41186 7310 41198 7362
rect 30382 7298 30434 7310
rect 34638 7298 34690 7310
rect 42254 7298 42306 7310
rect 43150 7362 43202 7374
rect 43150 7298 43202 7310
rect 54238 7362 54290 7374
rect 54238 7298 54290 7310
rect 54798 7362 54850 7374
rect 54798 7298 54850 7310
rect 26798 7250 26850 7262
rect 26798 7186 26850 7198
rect 27358 7250 27410 7262
rect 27358 7186 27410 7198
rect 27582 7250 27634 7262
rect 27582 7186 27634 7198
rect 29822 7250 29874 7262
rect 39118 7250 39170 7262
rect 49982 7250 50034 7262
rect 35186 7198 35198 7250
rect 35250 7198 35262 7250
rect 43026 7198 43038 7250
rect 43090 7247 43102 7250
rect 43586 7247 43598 7250
rect 43090 7201 43598 7247
rect 43090 7198 43102 7201
rect 43586 7198 43598 7201
rect 43650 7198 43662 7250
rect 52658 7198 52670 7250
rect 52722 7198 52734 7250
rect 29822 7186 29874 7198
rect 39118 7186 39170 7198
rect 49982 7186 50034 7198
rect 1344 7082 58576 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 58576 7082
rect 1344 6996 58576 7030
rect 43486 6914 43538 6926
rect 43486 6850 43538 6862
rect 48974 6914 49026 6926
rect 48974 6850 49026 6862
rect 50094 6914 50146 6926
rect 50094 6850 50146 6862
rect 53342 6914 53394 6926
rect 53342 6850 53394 6862
rect 53790 6914 53842 6926
rect 53790 6850 53842 6862
rect 19630 6802 19682 6814
rect 5954 6750 5966 6802
rect 6018 6750 6030 6802
rect 16370 6750 16382 6802
rect 16434 6750 16446 6802
rect 16818 6750 16830 6802
rect 16882 6750 16894 6802
rect 19630 6738 19682 6750
rect 21870 6802 21922 6814
rect 21870 6738 21922 6750
rect 21982 6802 22034 6814
rect 21982 6738 22034 6750
rect 22878 6802 22930 6814
rect 43262 6802 43314 6814
rect 27010 6750 27022 6802
rect 27074 6750 27086 6802
rect 29922 6750 29934 6802
rect 29986 6750 29998 6802
rect 32050 6750 32062 6802
rect 32114 6750 32126 6802
rect 33842 6750 33854 6802
rect 33906 6750 33918 6802
rect 22878 6738 22930 6750
rect 43262 6738 43314 6750
rect 45726 6802 45778 6814
rect 52222 6802 52274 6814
rect 46610 6750 46622 6802
rect 46674 6750 46686 6802
rect 45726 6738 45778 6750
rect 52222 6738 52274 6750
rect 53230 6802 53282 6814
rect 53230 6738 53282 6750
rect 54574 6802 54626 6814
rect 55234 6750 55246 6802
rect 55298 6750 55310 6802
rect 54574 6738 54626 6750
rect 19518 6690 19570 6702
rect 22990 6690 23042 6702
rect 35982 6690 36034 6702
rect 42702 6690 42754 6702
rect 8866 6638 8878 6690
rect 8930 6638 8942 6690
rect 13570 6638 13582 6690
rect 13634 6638 13646 6690
rect 17378 6638 17390 6690
rect 17442 6638 17454 6690
rect 19282 6638 19294 6690
rect 19346 6638 19358 6690
rect 19954 6638 19966 6690
rect 20018 6638 20030 6690
rect 21634 6638 21646 6690
rect 21698 6638 21710 6690
rect 23202 6638 23214 6690
rect 23266 6638 23278 6690
rect 24210 6638 24222 6690
rect 24274 6638 24286 6690
rect 24882 6638 24894 6690
rect 24946 6638 24958 6690
rect 29138 6638 29150 6690
rect 29202 6638 29214 6690
rect 33506 6638 33518 6690
rect 33570 6638 33582 6690
rect 35074 6638 35086 6690
rect 35138 6638 35150 6690
rect 42242 6638 42254 6690
rect 42306 6638 42318 6690
rect 19518 6626 19570 6638
rect 22990 6626 23042 6638
rect 35982 6626 36034 6638
rect 42702 6626 42754 6638
rect 43038 6690 43090 6702
rect 44046 6690 44098 6702
rect 43698 6638 43710 6690
rect 43762 6638 43774 6690
rect 43038 6626 43090 6638
rect 44046 6626 44098 6638
rect 45054 6690 45106 6702
rect 45838 6690 45890 6702
rect 45378 6638 45390 6690
rect 45442 6638 45454 6690
rect 45054 6626 45106 6638
rect 45838 6626 45890 6638
rect 47182 6690 47234 6702
rect 49646 6690 49698 6702
rect 49298 6638 49310 6690
rect 49362 6638 49374 6690
rect 47182 6626 47234 6638
rect 49646 6626 49698 6638
rect 53566 6690 53618 6702
rect 57362 6638 57374 6690
rect 57426 6638 57438 6690
rect 58034 6638 58046 6690
rect 58098 6638 58110 6690
rect 53566 6626 53618 6638
rect 22542 6578 22594 6590
rect 8082 6526 8094 6578
rect 8146 6526 8158 6578
rect 14242 6526 14254 6578
rect 14306 6526 14318 6578
rect 22542 6514 22594 6526
rect 22766 6578 22818 6590
rect 22766 6514 22818 6526
rect 34302 6578 34354 6590
rect 36094 6578 36146 6590
rect 46062 6578 46114 6590
rect 35298 6526 35310 6578
rect 35362 6526 35374 6578
rect 37202 6526 37214 6578
rect 37266 6526 37278 6578
rect 34302 6514 34354 6526
rect 36094 6514 36146 6526
rect 46062 6514 46114 6526
rect 46398 6578 46450 6590
rect 46398 6514 46450 6526
rect 49870 6578 49922 6590
rect 49870 6514 49922 6526
rect 50766 6578 50818 6590
rect 50766 6514 50818 6526
rect 51102 6578 51154 6590
rect 51102 6514 51154 6526
rect 52894 6578 52946 6590
rect 52894 6514 52946 6526
rect 16830 6466 16882 6478
rect 16830 6402 16882 6414
rect 16942 6466 16994 6478
rect 16942 6402 16994 6414
rect 17166 6466 17218 6478
rect 17166 6402 17218 6414
rect 19742 6466 19794 6478
rect 19742 6402 19794 6414
rect 36318 6466 36370 6478
rect 36318 6402 36370 6414
rect 42590 6466 42642 6478
rect 42590 6402 42642 6414
rect 43486 6466 43538 6478
rect 43486 6402 43538 6414
rect 45614 6466 45666 6478
rect 45614 6402 45666 6414
rect 46622 6466 46674 6478
rect 46622 6402 46674 6414
rect 49086 6466 49138 6478
rect 53678 6466 53730 6478
rect 50418 6414 50430 6466
rect 50482 6414 50494 6466
rect 49086 6402 49138 6414
rect 53678 6402 53730 6414
rect 1344 6298 58576 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 58576 6298
rect 1344 6212 58576 6246
rect 7982 6130 8034 6142
rect 7982 6066 8034 6078
rect 16270 6130 16322 6142
rect 16270 6066 16322 6078
rect 16830 6130 16882 6142
rect 16830 6066 16882 6078
rect 17950 6130 18002 6142
rect 26014 6130 26066 6142
rect 21298 6078 21310 6130
rect 21362 6078 21374 6130
rect 23538 6078 23550 6130
rect 23602 6078 23614 6130
rect 17950 6066 18002 6078
rect 26014 6066 26066 6078
rect 26686 6130 26738 6142
rect 26686 6066 26738 6078
rect 49646 6130 49698 6142
rect 49646 6066 49698 6078
rect 7870 6018 7922 6030
rect 7870 5954 7922 5966
rect 8094 6018 8146 6030
rect 8094 5954 8146 5966
rect 8542 6018 8594 6030
rect 8542 5954 8594 5966
rect 16382 6018 16434 6030
rect 16382 5954 16434 5966
rect 17390 6018 17442 6030
rect 17390 5954 17442 5966
rect 25230 6018 25282 6030
rect 25230 5954 25282 5966
rect 26462 6018 26514 6030
rect 33854 6018 33906 6030
rect 29138 5966 29150 6018
rect 29202 5966 29214 6018
rect 26462 5954 26514 5966
rect 33854 5954 33906 5966
rect 34974 6018 35026 6030
rect 47854 6018 47906 6030
rect 38210 5966 38222 6018
rect 38274 5966 38286 6018
rect 34974 5954 35026 5966
rect 47854 5954 47906 5966
rect 50094 6018 50146 6030
rect 50094 5954 50146 5966
rect 50206 6018 50258 6030
rect 50206 5954 50258 5966
rect 17614 5906 17666 5918
rect 15698 5854 15710 5906
rect 15762 5854 15774 5906
rect 16034 5854 16046 5906
rect 16098 5854 16110 5906
rect 17614 5842 17666 5854
rect 17838 5906 17890 5918
rect 17838 5842 17890 5854
rect 21646 5906 21698 5918
rect 24446 5906 24498 5918
rect 34638 5906 34690 5918
rect 47406 5906 47458 5918
rect 23762 5854 23774 5906
rect 23826 5854 23838 5906
rect 25442 5854 25454 5906
rect 25506 5854 25518 5906
rect 25778 5854 25790 5906
rect 25842 5854 25854 5906
rect 27122 5854 27134 5906
rect 27186 5854 27198 5906
rect 34402 5854 34414 5906
rect 34466 5854 34478 5906
rect 35298 5854 35310 5906
rect 35362 5854 35374 5906
rect 37538 5854 37550 5906
rect 37602 5854 37614 5906
rect 46162 5854 46174 5906
rect 46226 5854 46238 5906
rect 46946 5854 46958 5906
rect 47010 5854 47022 5906
rect 21646 5842 21698 5854
rect 24446 5842 24498 5854
rect 34638 5842 34690 5854
rect 47406 5842 47458 5854
rect 50318 5906 50370 5918
rect 56018 5854 56030 5906
rect 56082 5854 56094 5906
rect 50318 5842 50370 5854
rect 17726 5794 17778 5806
rect 13346 5742 13358 5794
rect 13410 5742 13422 5794
rect 17726 5730 17778 5742
rect 24334 5794 24386 5806
rect 24334 5730 24386 5742
rect 26574 5794 26626 5806
rect 46510 5794 46562 5806
rect 40338 5742 40350 5794
rect 40402 5742 40414 5794
rect 41122 5742 41134 5794
rect 41186 5742 41198 5794
rect 26574 5730 26626 5742
rect 46510 5730 46562 5742
rect 47966 5794 48018 5806
rect 53106 5742 53118 5794
rect 53170 5742 53182 5794
rect 55234 5742 55246 5794
rect 55298 5742 55310 5794
rect 47966 5730 48018 5742
rect 35310 5682 35362 5694
rect 25778 5630 25790 5682
rect 25842 5630 25854 5682
rect 50754 5630 50766 5682
rect 50818 5630 50830 5682
rect 35310 5618 35362 5630
rect 1344 5514 58576 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 58576 5514
rect 1344 5428 58576 5462
rect 16270 5346 16322 5358
rect 16270 5282 16322 5294
rect 30046 5346 30098 5358
rect 30046 5282 30098 5294
rect 44830 5346 44882 5358
rect 44830 5282 44882 5294
rect 45726 5346 45778 5358
rect 45726 5282 45778 5294
rect 19182 5234 19234 5246
rect 24110 5234 24162 5246
rect 10658 5182 10670 5234
rect 10722 5182 10734 5234
rect 12786 5182 12798 5234
rect 12850 5182 12862 5234
rect 15922 5182 15934 5234
rect 15986 5182 15998 5234
rect 18722 5182 18734 5234
rect 18786 5182 18798 5234
rect 19506 5182 19518 5234
rect 19570 5182 19582 5234
rect 19182 5170 19234 5182
rect 24110 5170 24162 5182
rect 26238 5234 26290 5246
rect 26238 5170 26290 5182
rect 26686 5234 26738 5246
rect 26686 5170 26738 5182
rect 27470 5234 27522 5246
rect 42702 5234 42754 5246
rect 33506 5182 33518 5234
rect 33570 5182 33582 5234
rect 35634 5182 35646 5234
rect 35698 5182 35710 5234
rect 41346 5182 41358 5234
rect 41410 5182 41422 5234
rect 27470 5170 27522 5182
rect 42702 5170 42754 5182
rect 45502 5234 45554 5246
rect 52222 5234 52274 5246
rect 46386 5182 46398 5234
rect 46450 5182 46462 5234
rect 54674 5182 54686 5234
rect 54738 5182 54750 5234
rect 45502 5170 45554 5182
rect 52222 5170 52274 5182
rect 18398 5122 18450 5134
rect 9314 5070 9326 5122
rect 9378 5070 9390 5122
rect 9986 5070 9998 5122
rect 10050 5070 10062 5122
rect 18162 5070 18174 5122
rect 18226 5070 18238 5122
rect 18398 5058 18450 5070
rect 20750 5122 20802 5134
rect 20750 5058 20802 5070
rect 21646 5122 21698 5134
rect 21646 5058 21698 5070
rect 22430 5122 22482 5134
rect 26574 5122 26626 5134
rect 30718 5122 30770 5134
rect 50990 5122 51042 5134
rect 22754 5070 22766 5122
rect 22818 5070 22830 5122
rect 23090 5070 23102 5122
rect 23154 5070 23166 5122
rect 26898 5070 26910 5122
rect 26962 5070 26974 5122
rect 29698 5070 29710 5122
rect 29762 5070 29774 5122
rect 36306 5070 36318 5122
rect 36370 5070 36382 5122
rect 38546 5070 38558 5122
rect 38610 5070 38622 5122
rect 41682 5070 41694 5122
rect 41746 5070 41758 5122
rect 49298 5070 49310 5122
rect 49362 5070 49374 5122
rect 52658 5070 52670 5122
rect 52722 5070 52734 5122
rect 22430 5058 22482 5070
rect 26574 5058 26626 5070
rect 30718 5058 30770 5070
rect 50990 5058 51042 5070
rect 16046 5010 16098 5022
rect 16046 4946 16098 4958
rect 18734 5010 18786 5022
rect 18734 4946 18786 4958
rect 19406 5010 19458 5022
rect 21422 5010 21474 5022
rect 20402 4958 20414 5010
rect 20466 4958 20478 5010
rect 19406 4946 19458 4958
rect 21422 4946 21474 4958
rect 21982 5010 22034 5022
rect 31502 5010 31554 5022
rect 30370 4958 30382 5010
rect 30434 4958 30446 5010
rect 21982 4946 22034 4958
rect 31502 4946 31554 4958
rect 31838 5010 31890 5022
rect 44942 5010 44994 5022
rect 39218 4958 39230 5010
rect 39282 4958 39294 5010
rect 48514 4958 48526 5010
rect 48578 4958 48590 5010
rect 31838 4946 31890 4958
rect 44942 4946 44994 4958
rect 9550 4898 9602 4910
rect 9550 4834 9602 4846
rect 18622 4898 18674 4910
rect 18622 4834 18674 4846
rect 21758 4898 21810 4910
rect 21758 4834 21810 4846
rect 21870 4898 21922 4910
rect 21870 4834 21922 4846
rect 22542 4898 22594 4910
rect 22542 4834 22594 4846
rect 29934 4898 29986 4910
rect 51326 4898 51378 4910
rect 46050 4846 46062 4898
rect 46114 4846 46126 4898
rect 29934 4834 29986 4846
rect 51326 4834 51378 4846
rect 1344 4730 58576 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 58576 4730
rect 1344 4644 58576 4678
rect 33294 4562 33346 4574
rect 33294 4498 33346 4510
rect 34414 4562 34466 4574
rect 34414 4498 34466 4510
rect 34526 4562 34578 4574
rect 34526 4498 34578 4510
rect 47742 4562 47794 4574
rect 47742 4498 47794 4510
rect 54126 4562 54178 4574
rect 54126 4498 54178 4510
rect 33182 4450 33234 4462
rect 10882 4398 10894 4450
rect 10946 4398 10958 4450
rect 14578 4398 14590 4450
rect 14642 4398 14654 4450
rect 19954 4398 19966 4450
rect 20018 4398 20030 4450
rect 22082 4398 22094 4450
rect 22146 4398 22158 4450
rect 26002 4398 26014 4450
rect 26066 4398 26078 4450
rect 30034 4398 30046 4450
rect 30098 4398 30110 4450
rect 33182 4386 33234 4398
rect 34638 4450 34690 4462
rect 47406 4450 47458 4462
rect 36866 4398 36878 4450
rect 36930 4398 36942 4450
rect 41906 4398 41918 4450
rect 41970 4398 41982 4450
rect 34638 4386 34690 4398
rect 47406 4386 47458 4398
rect 48078 4450 48130 4462
rect 53790 4450 53842 4462
rect 52658 4398 52670 4450
rect 52722 4398 52734 4450
rect 57810 4398 57822 4450
rect 57874 4398 57886 4450
rect 48078 4386 48130 4398
rect 53790 4386 53842 4398
rect 58158 4338 58210 4350
rect 10210 4286 10222 4338
rect 10274 4286 10286 4338
rect 13794 4286 13806 4338
rect 13858 4286 13870 4338
rect 20626 4286 20638 4338
rect 20690 4286 20702 4338
rect 21298 4286 21310 4338
rect 21362 4286 21374 4338
rect 25218 4286 25230 4338
rect 25282 4286 25294 4338
rect 29250 4286 29262 4338
rect 29314 4286 29326 4338
rect 36194 4286 36206 4338
rect 36258 4286 36270 4338
rect 41122 4286 41134 4338
rect 41186 4286 41198 4338
rect 44482 4286 44494 4338
rect 44546 4286 44558 4338
rect 53442 4286 53454 4338
rect 53506 4286 53518 4338
rect 58158 4274 58210 4286
rect 48862 4226 48914 4238
rect 57598 4226 57650 4238
rect 13010 4174 13022 4226
rect 13074 4174 13086 4226
rect 16706 4174 16718 4226
rect 16770 4174 16782 4226
rect 17826 4174 17838 4226
rect 17890 4174 17902 4226
rect 24210 4174 24222 4226
rect 24274 4174 24286 4226
rect 28130 4174 28142 4226
rect 28194 4174 28206 4226
rect 32162 4174 32174 4226
rect 32226 4174 32238 4226
rect 38994 4174 39006 4226
rect 39058 4174 39070 4226
rect 44034 4174 44046 4226
rect 44098 4174 44110 4226
rect 50530 4174 50542 4226
rect 50594 4174 50606 4226
rect 48862 4162 48914 4174
rect 57598 4162 57650 4174
rect 45390 4114 45442 4126
rect 45390 4050 45442 4062
rect 1344 3946 58576 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 58576 3946
rect 1344 3860 58576 3894
rect 22094 3666 22146 3678
rect 18834 3614 18846 3666
rect 18898 3614 18910 3666
rect 22094 3602 22146 3614
rect 26126 3666 26178 3678
rect 26126 3602 26178 3614
rect 40798 3666 40850 3678
rect 40798 3602 40850 3614
rect 43150 3666 43202 3678
rect 44370 3614 44382 3666
rect 44434 3614 44446 3666
rect 46498 3614 46510 3666
rect 46562 3614 46574 3666
rect 43150 3602 43202 3614
rect 20066 3502 20078 3554
rect 20130 3502 20142 3554
rect 21074 3502 21086 3554
rect 21138 3502 21150 3554
rect 25218 3502 25230 3554
rect 25282 3502 25294 3554
rect 36642 3502 36654 3554
rect 36706 3502 36718 3554
rect 39778 3502 39790 3554
rect 39842 3502 39854 3554
rect 43698 3502 43710 3554
rect 43762 3502 43774 3554
rect 47394 3502 47406 3554
rect 47458 3502 47470 3554
rect 48962 3390 48974 3442
rect 49026 3390 49038 3442
rect 2942 3330 2994 3342
rect 2942 3266 2994 3278
rect 5518 3330 5570 3342
rect 5518 3266 5570 3278
rect 6974 3330 7026 3342
rect 6974 3266 7026 3278
rect 9326 3330 9378 3342
rect 9326 3266 9378 3278
rect 11006 3330 11058 3342
rect 11006 3266 11058 3278
rect 13134 3330 13186 3342
rect 13134 3266 13186 3278
rect 15038 3330 15090 3342
rect 15038 3266 15090 3278
rect 17054 3330 17106 3342
rect 17054 3266 17106 3278
rect 28366 3330 28418 3342
rect 28366 3266 28418 3278
rect 29150 3330 29202 3342
rect 29150 3266 29202 3278
rect 31166 3330 31218 3342
rect 31166 3266 31218 3278
rect 33182 3330 33234 3342
rect 33182 3266 33234 3278
rect 35198 3330 35250 3342
rect 35198 3266 35250 3278
rect 37662 3330 37714 3342
rect 37662 3266 37714 3278
rect 50318 3330 50370 3342
rect 50318 3266 50370 3278
rect 51326 3330 51378 3342
rect 51326 3266 51378 3278
rect 53342 3330 53394 3342
rect 53342 3266 53394 3278
rect 55358 3330 55410 3342
rect 55358 3266 55410 3278
rect 57374 3330 57426 3342
rect 57374 3266 57426 3278
rect 1344 3162 58576 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 58576 3162
rect 1344 3076 58576 3110
rect 26898 1710 26910 1762
rect 26962 1759 26974 1762
rect 28354 1759 28366 1762
rect 26962 1713 28366 1759
rect 26962 1710 26974 1713
rect 28354 1710 28366 1713
rect 28418 1710 28430 1762
rect 49074 1710 49086 1762
rect 49138 1759 49150 1762
rect 50306 1759 50318 1762
rect 49138 1713 50318 1759
rect 49138 1710 49150 1713
rect 50306 1710 50318 1713
rect 50370 1710 50382 1762
<< via1 >>
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 22430 56254 22482 56306
rect 22654 56254 22706 56306
rect 27022 56254 27074 56306
rect 37438 56254 37490 56306
rect 37662 56254 37714 56306
rect 52446 56254 52498 56306
rect 52670 56142 52722 56194
rect 57822 56142 57874 56194
rect 26686 56030 26738 56082
rect 27134 56030 27186 56082
rect 27358 56030 27410 56082
rect 52894 56030 52946 56082
rect 57598 56030 57650 56082
rect 58158 56030 58210 56082
rect 23102 55918 23154 55970
rect 38222 55918 38274 55970
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 20414 55358 20466 55410
rect 25790 55358 25842 55410
rect 29150 55358 29202 55410
rect 36430 55358 36482 55410
rect 40238 55358 40290 55410
rect 42702 55358 42754 55410
rect 48862 55358 48914 55410
rect 52110 55358 52162 55410
rect 55582 55358 55634 55410
rect 57598 55358 57650 55410
rect 17502 55246 17554 55298
rect 21646 55246 21698 55298
rect 21982 55246 22034 55298
rect 22990 55246 23042 55298
rect 27694 55246 27746 55298
rect 32062 55246 32114 55298
rect 33518 55246 33570 55298
rect 37326 55246 37378 55298
rect 40798 55246 40850 55298
rect 41022 55246 41074 55298
rect 41246 55246 41298 55298
rect 42366 55246 42418 55298
rect 46062 55246 46114 55298
rect 49310 55246 49362 55298
rect 52670 55246 52722 55298
rect 18286 55134 18338 55186
rect 21310 55134 21362 55186
rect 23662 55134 23714 55186
rect 27358 55134 27410 55186
rect 27470 55134 27522 55186
rect 31278 55134 31330 55186
rect 34302 55134 34354 55186
rect 38110 55134 38162 55186
rect 40686 55134 40738 55186
rect 46734 55134 46786 55186
rect 49982 55134 50034 55186
rect 53454 55134 53506 55186
rect 21646 55022 21698 55074
rect 26910 55022 26962 55074
rect 42590 55022 42642 55074
rect 57486 55022 57538 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 22766 54686 22818 54738
rect 23774 54686 23826 54738
rect 40238 54686 40290 54738
rect 41470 54686 41522 54738
rect 41806 54686 41858 54738
rect 47406 54686 47458 54738
rect 54462 54686 54514 54738
rect 25454 54574 25506 54626
rect 36878 54574 36930 54626
rect 40126 54574 40178 54626
rect 42142 54574 42194 54626
rect 51998 54574 52050 54626
rect 54574 54574 54626 54626
rect 17502 54462 17554 54514
rect 20638 54462 20690 54514
rect 21870 54462 21922 54514
rect 22990 54462 23042 54514
rect 23550 54462 23602 54514
rect 29038 54462 29090 54514
rect 31390 54462 31442 54514
rect 36542 54462 36594 54514
rect 40910 54462 40962 54514
rect 45502 54462 45554 54514
rect 46510 54462 46562 54514
rect 46734 54462 46786 54514
rect 47630 54462 47682 54514
rect 52894 54462 52946 54514
rect 18174 54350 18226 54402
rect 20302 54350 20354 54402
rect 20974 54350 21026 54402
rect 21534 54350 21586 54402
rect 22318 54350 22370 54402
rect 22654 54350 22706 54402
rect 24782 54350 24834 54402
rect 42590 54350 42642 54402
rect 44718 54350 44770 54402
rect 46958 54350 47010 54402
rect 47294 54350 47346 54402
rect 48302 54350 48354 54402
rect 23886 54238 23938 54290
rect 31614 54238 31666 54290
rect 31838 54238 31890 54290
rect 31950 54238 32002 54290
rect 40350 54238 40402 54290
rect 41134 54238 41186 54290
rect 54350 54238 54402 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 20638 53902 20690 53954
rect 26910 53902 26962 53954
rect 27134 53902 27186 53954
rect 29486 53902 29538 53954
rect 37438 53902 37490 53954
rect 40350 53902 40402 53954
rect 40574 53902 40626 53954
rect 40910 53902 40962 53954
rect 43150 53902 43202 53954
rect 50766 53902 50818 53954
rect 26126 53790 26178 53842
rect 29374 53790 29426 53842
rect 29710 53790 29762 53842
rect 31278 53790 31330 53842
rect 33406 53790 33458 53842
rect 35870 53790 35922 53842
rect 39118 53790 39170 53842
rect 40014 53790 40066 53842
rect 41134 53790 41186 53842
rect 50542 53790 50594 53842
rect 51438 53790 51490 53842
rect 52782 53790 52834 53842
rect 20190 53678 20242 53730
rect 20302 53678 20354 53730
rect 20526 53678 20578 53730
rect 21870 53678 21922 53730
rect 22094 53678 22146 53730
rect 22878 53678 22930 53730
rect 25230 53678 25282 53730
rect 25902 53678 25954 53730
rect 27246 53678 27298 53730
rect 27582 53678 27634 53730
rect 27918 53678 27970 53730
rect 28254 53678 28306 53730
rect 28478 53678 28530 53730
rect 29822 53678 29874 53730
rect 34078 53678 34130 53730
rect 36094 53678 36146 53730
rect 36430 53678 36482 53730
rect 36990 53678 37042 53730
rect 37102 53678 37154 53730
rect 37326 53678 37378 53730
rect 39454 53678 39506 53730
rect 39790 53678 39842 53730
rect 41358 53678 41410 53730
rect 41694 53678 41746 53730
rect 43038 53678 43090 53730
rect 43374 53678 43426 53730
rect 43486 53678 43538 53730
rect 48638 53678 48690 53730
rect 50430 53678 50482 53730
rect 50878 53678 50930 53730
rect 51662 53678 51714 53730
rect 53230 53678 53282 53730
rect 53678 53678 53730 53730
rect 54238 53678 54290 53730
rect 55022 53678 55074 53730
rect 55358 53678 55410 53730
rect 21758 53566 21810 53618
rect 28366 53566 28418 53618
rect 30942 53566 30994 53618
rect 41582 53566 41634 53618
rect 51326 53566 51378 53618
rect 54014 53566 54066 53618
rect 55582 53566 55634 53618
rect 21310 53454 21362 53506
rect 22990 53454 23042 53506
rect 27246 53454 27298 53506
rect 30606 53454 30658 53506
rect 37998 53454 38050 53506
rect 39230 53454 39282 53506
rect 40798 53454 40850 53506
rect 42142 53454 42194 53506
rect 48750 53454 48802 53506
rect 55246 53454 55298 53506
rect 55918 53454 55970 53506
rect 56254 53454 56306 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 26238 53118 26290 53170
rect 28142 53118 28194 53170
rect 31614 53118 31666 53170
rect 46734 53118 46786 53170
rect 50654 53118 50706 53170
rect 26350 53006 26402 53058
rect 28030 53006 28082 53058
rect 31726 53006 31778 53058
rect 35198 53006 35250 53058
rect 49982 53006 50034 53058
rect 54910 53006 54962 53058
rect 55022 53006 55074 53058
rect 19070 52894 19122 52946
rect 24670 52894 24722 52946
rect 28366 52894 28418 52946
rect 40014 52894 40066 52946
rect 40910 52894 40962 52946
rect 41134 52894 41186 52946
rect 41358 52894 41410 52946
rect 46958 52894 47010 52946
rect 50094 52894 50146 52946
rect 50206 52894 50258 52946
rect 54798 52894 54850 52946
rect 55470 52894 55522 52946
rect 56590 52894 56642 52946
rect 56814 52894 56866 52946
rect 22654 52782 22706 52834
rect 31502 52670 31554 52722
rect 41470 52670 41522 52722
rect 57038 52670 57090 52722
rect 57150 52670 57202 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 31390 52334 31442 52386
rect 31614 52334 31666 52386
rect 35870 52334 35922 52386
rect 37326 52334 37378 52386
rect 43710 52334 43762 52386
rect 45054 52334 45106 52386
rect 45278 52334 45330 52386
rect 45950 52334 46002 52386
rect 46286 52334 46338 52386
rect 18062 52222 18114 52274
rect 20078 52222 20130 52274
rect 26462 52222 26514 52274
rect 28590 52222 28642 52274
rect 35534 52222 35586 52274
rect 38782 52222 38834 52274
rect 40910 52222 40962 52274
rect 44046 52222 44098 52274
rect 49646 52222 49698 52274
rect 55246 52222 55298 52274
rect 57374 52222 57426 52274
rect 15262 52110 15314 52162
rect 22766 52110 22818 52162
rect 22990 52110 23042 52162
rect 23998 52110 24050 52162
rect 24558 52110 24610 52162
rect 25678 52110 25730 52162
rect 31838 52110 31890 52162
rect 36094 52110 36146 52162
rect 36318 52110 36370 52162
rect 37326 52110 37378 52162
rect 37998 52110 38050 52162
rect 41582 52110 41634 52162
rect 42254 52110 42306 52162
rect 42702 52110 42754 52162
rect 44830 52110 44882 52162
rect 45726 52110 45778 52162
rect 48078 52110 48130 52162
rect 48414 52110 48466 52162
rect 48526 52110 48578 52162
rect 48862 52110 48914 52162
rect 49198 52110 49250 52162
rect 49534 52110 49586 52162
rect 49870 52110 49922 52162
rect 50206 52110 50258 52162
rect 58046 52110 58098 52162
rect 15934 51998 15986 52050
rect 19742 51998 19794 52050
rect 19966 51998 20018 52050
rect 35758 51998 35810 52050
rect 36990 51998 37042 52050
rect 42478 51998 42530 52050
rect 45390 51998 45442 52050
rect 48190 51998 48242 52050
rect 50318 51998 50370 52050
rect 51214 51998 51266 52050
rect 23326 51886 23378 51938
rect 23662 51886 23714 51938
rect 31726 51886 31778 51938
rect 32398 51886 32450 51938
rect 41246 51886 41298 51938
rect 43934 51886 43986 51938
rect 48862 51886 48914 51938
rect 51102 51886 51154 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 19406 51550 19458 51602
rect 26462 51550 26514 51602
rect 31278 51550 31330 51602
rect 31950 51550 32002 51602
rect 46846 51550 46898 51602
rect 20302 51438 20354 51490
rect 23662 51438 23714 51490
rect 28030 51438 28082 51490
rect 30830 51438 30882 51490
rect 34974 51438 35026 51490
rect 37774 51438 37826 51490
rect 42478 51438 42530 51490
rect 45390 51438 45442 51490
rect 49646 51438 49698 51490
rect 51214 51438 51266 51490
rect 19966 51326 20018 51378
rect 20638 51326 20690 51378
rect 21086 51326 21138 51378
rect 22990 51326 23042 51378
rect 23998 51326 24050 51378
rect 26126 51326 26178 51378
rect 28366 51326 28418 51378
rect 30494 51326 30546 51378
rect 30718 51326 30770 51378
rect 31614 51326 31666 51378
rect 31838 51326 31890 51378
rect 32286 51326 32338 51378
rect 34190 51326 34242 51378
rect 37550 51326 37602 51378
rect 38222 51326 38274 51378
rect 46062 51326 46114 51378
rect 46510 51326 46562 51378
rect 48862 51326 48914 51378
rect 48974 51326 49026 51378
rect 49198 51326 49250 51378
rect 50206 51326 50258 51378
rect 50654 51326 50706 51378
rect 54574 51326 54626 51378
rect 55358 51326 55410 51378
rect 55694 51326 55746 51378
rect 18846 51214 18898 51266
rect 20190 51214 20242 51266
rect 22766 51214 22818 51266
rect 23326 51214 23378 51266
rect 25790 51214 25842 51266
rect 33182 51214 33234 51266
rect 37102 51214 37154 51266
rect 43262 51214 43314 51266
rect 50990 51214 51042 51266
rect 51662 51214 51714 51266
rect 53790 51214 53842 51266
rect 55918 51214 55970 51266
rect 19070 51102 19122 51154
rect 19854 51102 19906 51154
rect 20862 51102 20914 51154
rect 21198 51102 21250 51154
rect 42590 51102 42642 51154
rect 49310 51102 49362 51154
rect 56030 51102 56082 51154
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 19966 50766 20018 50818
rect 49534 50766 49586 50818
rect 49646 50766 49698 50818
rect 50094 50766 50146 50818
rect 50206 50766 50258 50818
rect 50654 50766 50706 50818
rect 21310 50654 21362 50706
rect 23438 50654 23490 50706
rect 25566 50654 25618 50706
rect 29486 50654 29538 50706
rect 30382 50654 30434 50706
rect 31166 50654 31218 50706
rect 33294 50654 33346 50706
rect 35982 50654 36034 50706
rect 46174 50654 46226 50706
rect 19182 50542 19234 50594
rect 19742 50542 19794 50594
rect 22654 50542 22706 50594
rect 26910 50542 26962 50594
rect 29934 50542 29986 50594
rect 34078 50542 34130 50594
rect 35870 50542 35922 50594
rect 36094 50542 36146 50594
rect 36430 50542 36482 50594
rect 37102 50542 37154 50594
rect 45502 50542 45554 50594
rect 49870 50542 49922 50594
rect 51214 50542 51266 50594
rect 51438 50542 51490 50594
rect 51550 50542 51602 50594
rect 52894 50542 52946 50594
rect 14366 50430 14418 50482
rect 20302 50430 20354 50482
rect 21422 50430 21474 50482
rect 27134 50430 27186 50482
rect 28254 50430 28306 50482
rect 28590 50430 28642 50482
rect 45166 50430 45218 50482
rect 50542 50430 50594 50482
rect 50990 50430 51042 50482
rect 57934 50430 57986 50482
rect 21534 50318 21586 50370
rect 51774 50318 51826 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 25902 49982 25954 50034
rect 26798 49982 26850 50034
rect 30158 49982 30210 50034
rect 30382 49982 30434 50034
rect 37102 49982 37154 50034
rect 41806 49982 41858 50034
rect 50542 49982 50594 50034
rect 50990 49982 51042 50034
rect 52558 49982 52610 50034
rect 57374 49982 57426 50034
rect 58158 49982 58210 50034
rect 30942 49870 30994 49922
rect 31278 49870 31330 49922
rect 37662 49870 37714 49922
rect 41358 49870 41410 49922
rect 50206 49870 50258 49922
rect 50318 49870 50370 49922
rect 56030 49870 56082 49922
rect 56590 49870 56642 49922
rect 56702 49870 56754 49922
rect 14254 49758 14306 49810
rect 25678 49758 25730 49810
rect 26686 49758 26738 49810
rect 30718 49758 30770 49810
rect 31390 49758 31442 49810
rect 36542 49758 36594 49810
rect 40910 49758 40962 49810
rect 41134 49758 41186 49810
rect 48974 49758 49026 49810
rect 49198 49758 49250 49810
rect 55582 49758 55634 49810
rect 55806 49758 55858 49810
rect 56926 49758 56978 49810
rect 57598 49758 57650 49810
rect 11342 49646 11394 49698
rect 13470 49646 13522 49698
rect 19630 49646 19682 49698
rect 25790 49646 25842 49698
rect 26126 49646 26178 49698
rect 31950 49646 32002 49698
rect 41022 49646 41074 49698
rect 41918 49646 41970 49698
rect 42366 49646 42418 49698
rect 48750 49646 48802 49698
rect 26350 49534 26402 49586
rect 26798 49534 26850 49586
rect 36654 49534 36706 49586
rect 42254 49534 42306 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 39118 49198 39170 49250
rect 48526 49198 48578 49250
rect 16158 49086 16210 49138
rect 18398 49086 18450 49138
rect 19966 49086 20018 49138
rect 35646 49086 35698 49138
rect 38558 49086 38610 49138
rect 39678 49086 39730 49138
rect 40910 49086 40962 49138
rect 43150 49086 43202 49138
rect 44158 49086 44210 49138
rect 48190 49086 48242 49138
rect 53006 49086 53058 49138
rect 56030 49086 56082 49138
rect 58158 49086 58210 49138
rect 15374 48974 15426 49026
rect 21982 48974 22034 49026
rect 26350 48974 26402 49026
rect 27694 48974 27746 49026
rect 29934 48974 29986 49026
rect 35422 48974 35474 49026
rect 36990 48974 37042 49026
rect 37214 48974 37266 49026
rect 37438 48974 37490 49026
rect 37550 48974 37602 49026
rect 38110 48974 38162 49026
rect 39342 48974 39394 49026
rect 39566 48974 39618 49026
rect 40350 48974 40402 49026
rect 40798 48974 40850 49026
rect 41022 48974 41074 49026
rect 41358 48974 41410 49026
rect 42142 48974 42194 49026
rect 42478 48974 42530 49026
rect 43038 48974 43090 49026
rect 45390 48974 45442 49026
rect 55246 48974 55298 49026
rect 7982 48862 8034 48914
rect 20302 48862 20354 48914
rect 21646 48862 21698 48914
rect 22094 48862 22146 48914
rect 26574 48862 26626 48914
rect 27806 48862 27858 48914
rect 29822 48862 29874 48914
rect 34862 48862 34914 48914
rect 38558 48862 38610 48914
rect 42590 48862 42642 48914
rect 43374 48862 43426 48914
rect 45166 48862 45218 48914
rect 48302 48862 48354 48914
rect 8094 48750 8146 48802
rect 8318 48750 8370 48802
rect 20078 48750 20130 48802
rect 21534 48750 21586 48802
rect 22318 48750 22370 48802
rect 27246 48750 27298 48802
rect 33630 48750 33682 48802
rect 36206 48750 36258 48802
rect 37662 48750 37714 48802
rect 38334 48750 38386 48802
rect 38670 48750 38722 48802
rect 39790 48750 39842 48802
rect 40574 48750 40626 48802
rect 41470 48750 41522 48802
rect 41694 48750 41746 48802
rect 42254 48750 42306 48802
rect 42366 48750 42418 48802
rect 44270 48750 44322 48802
rect 45726 48750 45778 48802
rect 53454 48750 53506 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 24558 48414 24610 48466
rect 25342 48414 25394 48466
rect 26686 48414 26738 48466
rect 34638 48414 34690 48466
rect 37326 48414 37378 48466
rect 40126 48414 40178 48466
rect 43598 48414 43650 48466
rect 43934 48414 43986 48466
rect 44158 48414 44210 48466
rect 46062 48414 46114 48466
rect 9550 48302 9602 48354
rect 9774 48302 9826 48354
rect 18622 48302 18674 48354
rect 32062 48302 32114 48354
rect 36206 48302 36258 48354
rect 37662 48302 37714 48354
rect 42814 48302 42866 48354
rect 45054 48302 45106 48354
rect 45614 48302 45666 48354
rect 46174 48302 46226 48354
rect 48078 48302 48130 48354
rect 51550 48302 51602 48354
rect 56590 48302 56642 48354
rect 57150 48302 57202 48354
rect 6190 48190 6242 48242
rect 14030 48190 14082 48242
rect 17838 48190 17890 48242
rect 21198 48190 21250 48242
rect 26574 48190 26626 48242
rect 27246 48190 27298 48242
rect 27470 48190 27522 48242
rect 29038 48190 29090 48242
rect 30382 48190 30434 48242
rect 31838 48190 31890 48242
rect 32174 48190 32226 48242
rect 34414 48190 34466 48242
rect 34750 48190 34802 48242
rect 35086 48190 35138 48242
rect 37102 48190 37154 48242
rect 39678 48190 39730 48242
rect 39902 48190 39954 48242
rect 40350 48190 40402 48242
rect 41470 48190 41522 48242
rect 41694 48190 41746 48242
rect 42478 48190 42530 48242
rect 43262 48190 43314 48242
rect 43486 48190 43538 48242
rect 43822 48190 43874 48242
rect 44494 48190 44546 48242
rect 44942 48190 44994 48242
rect 45838 48190 45890 48242
rect 46958 48190 47010 48242
rect 47854 48190 47906 48242
rect 50318 48190 50370 48242
rect 50878 48190 50930 48242
rect 56814 48190 56866 48242
rect 6862 48078 6914 48130
rect 8990 48078 9042 48130
rect 9662 48078 9714 48130
rect 14702 48078 14754 48130
rect 16830 48078 16882 48130
rect 20750 48078 20802 48130
rect 21982 48078 22034 48130
rect 24110 48078 24162 48130
rect 24446 48078 24498 48130
rect 25230 48078 25282 48130
rect 30830 48078 30882 48130
rect 33294 48078 33346 48130
rect 33630 48078 33682 48130
rect 39342 48078 39394 48130
rect 44270 48078 44322 48130
rect 45278 48078 45330 48130
rect 45950 48078 46002 48130
rect 47182 48078 47234 48130
rect 47518 48078 47570 48130
rect 49982 48078 50034 48130
rect 53678 48078 53730 48130
rect 57038 48078 57090 48130
rect 26686 47966 26738 48018
rect 30942 47966 30994 48018
rect 39230 47966 39282 48018
rect 40238 47966 40290 48018
rect 40798 47966 40850 48018
rect 41246 47966 41298 48018
rect 43038 47966 43090 48018
rect 46622 47966 46674 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 17614 47630 17666 47682
rect 27470 47630 27522 47682
rect 38334 47630 38386 47682
rect 43486 47630 43538 47682
rect 45054 47630 45106 47682
rect 6190 47518 6242 47570
rect 15934 47518 15986 47570
rect 20078 47518 20130 47570
rect 20526 47518 20578 47570
rect 21870 47518 21922 47570
rect 26686 47518 26738 47570
rect 27806 47518 27858 47570
rect 28590 47518 28642 47570
rect 31838 47518 31890 47570
rect 33966 47518 34018 47570
rect 34974 47518 35026 47570
rect 38670 47518 38722 47570
rect 40686 47518 40738 47570
rect 47070 47518 47122 47570
rect 51102 47518 51154 47570
rect 55246 47518 55298 47570
rect 57374 47518 57426 47570
rect 10446 47406 10498 47458
rect 16046 47406 16098 47458
rect 16494 47406 16546 47458
rect 16718 47406 16770 47458
rect 17054 47406 17106 47458
rect 17950 47406 18002 47458
rect 18174 47406 18226 47458
rect 19966 47406 20018 47458
rect 21422 47406 21474 47458
rect 21758 47406 21810 47458
rect 22094 47406 22146 47458
rect 22318 47406 22370 47458
rect 23326 47406 23378 47458
rect 24222 47406 24274 47458
rect 26910 47406 26962 47458
rect 27694 47406 27746 47458
rect 29710 47406 29762 47458
rect 30270 47406 30322 47458
rect 31166 47406 31218 47458
rect 34526 47406 34578 47458
rect 35534 47406 35586 47458
rect 37214 47406 37266 47458
rect 37886 47406 37938 47458
rect 38558 47406 38610 47458
rect 38782 47406 38834 47458
rect 44942 47406 44994 47458
rect 50654 47406 50706 47458
rect 53342 47406 53394 47458
rect 53678 47406 53730 47458
rect 54126 47406 54178 47458
rect 58046 47406 58098 47458
rect 14926 47294 14978 47346
rect 15262 47294 15314 47346
rect 15822 47294 15874 47346
rect 22542 47294 22594 47346
rect 28478 47294 28530 47346
rect 29262 47294 29314 47346
rect 30382 47294 30434 47346
rect 35646 47294 35698 47346
rect 36318 47294 36370 47346
rect 37438 47294 37490 47346
rect 37550 47294 37602 47346
rect 38110 47294 38162 47346
rect 43598 47294 43650 47346
rect 53902 47294 53954 47346
rect 11342 47182 11394 47234
rect 16942 47182 16994 47234
rect 18622 47182 18674 47234
rect 23438 47182 23490 47234
rect 23662 47182 23714 47234
rect 24110 47182 24162 47234
rect 29710 47182 29762 47234
rect 36430 47182 36482 47234
rect 40798 47182 40850 47234
rect 52782 47182 52834 47234
rect 52894 47182 52946 47234
rect 53006 47182 53058 47234
rect 54014 47182 54066 47234
rect 54238 47182 54290 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 17502 46846 17554 46898
rect 35534 46846 35586 46898
rect 35982 46846 36034 46898
rect 36766 46846 36818 46898
rect 36990 46846 37042 46898
rect 52446 46846 52498 46898
rect 56590 46846 56642 46898
rect 57150 46846 57202 46898
rect 8766 46734 8818 46786
rect 15038 46734 15090 46786
rect 16270 46734 16322 46786
rect 20190 46734 20242 46786
rect 28590 46734 28642 46786
rect 30942 46734 30994 46786
rect 33070 46734 33122 46786
rect 33182 46734 33234 46786
rect 33742 46734 33794 46786
rect 36542 46734 36594 46786
rect 41134 46734 41186 46786
rect 46062 46734 46114 46786
rect 52110 46734 52162 46786
rect 54126 46734 54178 46786
rect 55470 46734 55522 46786
rect 56702 46734 56754 46786
rect 57038 46734 57090 46786
rect 6974 46622 7026 46674
rect 7758 46622 7810 46674
rect 10222 46622 10274 46674
rect 18734 46622 18786 46674
rect 24334 46622 24386 46674
rect 25790 46622 25842 46674
rect 26462 46622 26514 46674
rect 26910 46622 26962 46674
rect 28366 46622 28418 46674
rect 29486 46622 29538 46674
rect 31502 46622 31554 46674
rect 33406 46622 33458 46674
rect 37214 46622 37266 46674
rect 41022 46622 41074 46674
rect 41582 46622 41634 46674
rect 42030 46622 42082 46674
rect 46174 46622 46226 46674
rect 46286 46622 46338 46674
rect 46622 46622 46674 46674
rect 49870 46622 49922 46674
rect 50094 46622 50146 46674
rect 50318 46622 50370 46674
rect 50878 46622 50930 46674
rect 54686 46622 54738 46674
rect 55022 46622 55074 46674
rect 55246 46622 55298 46674
rect 55694 46622 55746 46674
rect 58158 46622 58210 46674
rect 4174 46510 4226 46562
rect 6302 46510 6354 46562
rect 7646 46510 7698 46562
rect 8878 46510 8930 46562
rect 10894 46510 10946 46562
rect 13022 46510 13074 46562
rect 14926 46510 14978 46562
rect 26126 46510 26178 46562
rect 29262 46510 29314 46562
rect 34190 46510 34242 46562
rect 37102 46510 37154 46562
rect 42702 46510 42754 46562
rect 50206 46510 50258 46562
rect 55358 46510 55410 46562
rect 57710 46510 57762 46562
rect 7422 46398 7474 46450
rect 8542 46398 8594 46450
rect 15262 46398 15314 46450
rect 16158 46398 16210 46450
rect 26462 46398 26514 46450
rect 49646 46398 49698 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 11342 46062 11394 46114
rect 14590 46062 14642 46114
rect 29486 46062 29538 46114
rect 29822 46062 29874 46114
rect 37998 46062 38050 46114
rect 40014 46062 40066 46114
rect 7310 45950 7362 46002
rect 21758 45950 21810 46002
rect 29374 45950 29426 46002
rect 31166 45950 31218 46002
rect 37102 45950 37154 46002
rect 40574 45950 40626 46002
rect 47966 45950 48018 46002
rect 50094 45950 50146 46002
rect 6750 45838 6802 45890
rect 7198 45838 7250 45890
rect 8206 45838 8258 45890
rect 8542 45838 8594 45890
rect 11342 45838 11394 45890
rect 12014 45838 12066 45890
rect 12238 45838 12290 45890
rect 14926 45838 14978 45890
rect 18622 45838 18674 45890
rect 21646 45838 21698 45890
rect 22654 45838 22706 45890
rect 24110 45838 24162 45890
rect 26126 45838 26178 45890
rect 26798 45838 26850 45890
rect 29150 45838 29202 45890
rect 36206 45838 36258 45890
rect 47182 45838 47234 45890
rect 50430 45838 50482 45890
rect 51326 45838 51378 45890
rect 52782 45838 52834 45890
rect 53454 45838 53506 45890
rect 54014 45838 54066 45890
rect 54462 45838 54514 45890
rect 55694 45838 55746 45890
rect 56254 45838 56306 45890
rect 57150 45838 57202 45890
rect 11678 45726 11730 45778
rect 12574 45726 12626 45778
rect 14254 45726 14306 45778
rect 21982 45726 22034 45778
rect 23214 45726 23266 45778
rect 24558 45726 24610 45778
rect 25566 45726 25618 45778
rect 26910 45726 26962 45778
rect 29934 45726 29986 45778
rect 37886 45726 37938 45778
rect 39902 45726 39954 45778
rect 44046 45726 44098 45778
rect 51438 45726 51490 45778
rect 53902 45726 53954 45778
rect 54126 45726 54178 45778
rect 55582 45726 55634 45778
rect 57262 45726 57314 45778
rect 8430 45614 8482 45666
rect 12462 45614 12514 45666
rect 12686 45614 12738 45666
rect 13918 45614 13970 45666
rect 14702 45614 14754 45666
rect 18286 45614 18338 45666
rect 20414 45614 20466 45666
rect 27134 45614 27186 45666
rect 44158 45614 44210 45666
rect 50542 45614 50594 45666
rect 51326 45614 51378 45666
rect 54574 45614 54626 45666
rect 54798 45614 54850 45666
rect 56366 45614 56418 45666
rect 56590 45614 56642 45666
rect 58158 45614 58210 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 13246 45278 13298 45330
rect 14366 45278 14418 45330
rect 19518 45278 19570 45330
rect 57486 45278 57538 45330
rect 9662 45166 9714 45218
rect 14590 45166 14642 45218
rect 16046 45166 16098 45218
rect 20638 45166 20690 45218
rect 21198 45166 21250 45218
rect 31502 45166 31554 45218
rect 40126 45166 40178 45218
rect 44942 45166 44994 45218
rect 52782 45166 52834 45218
rect 56814 45166 56866 45218
rect 57598 45166 57650 45218
rect 9550 45054 9602 45106
rect 9886 45054 9938 45106
rect 10222 45054 10274 45106
rect 11230 45054 11282 45106
rect 13022 45054 13074 45106
rect 13358 45054 13410 45106
rect 14702 45054 14754 45106
rect 14814 45054 14866 45106
rect 15374 45054 15426 45106
rect 15822 45054 15874 45106
rect 16606 45054 16658 45106
rect 22878 45054 22930 45106
rect 23550 45054 23602 45106
rect 23774 45054 23826 45106
rect 25342 45054 25394 45106
rect 26350 45054 26402 45106
rect 27134 45054 27186 45106
rect 28590 45054 28642 45106
rect 29598 45054 29650 45106
rect 32174 45054 32226 45106
rect 36206 45054 36258 45106
rect 40910 45054 40962 45106
rect 44270 45054 44322 45106
rect 50094 45054 50146 45106
rect 51102 45054 51154 45106
rect 56702 45054 56754 45106
rect 57486 45054 57538 45106
rect 10558 44942 10610 44994
rect 16494 44942 16546 44994
rect 20078 44942 20130 44994
rect 20750 44942 20802 44994
rect 22990 44942 23042 44994
rect 23438 44942 23490 44994
rect 30158 44942 30210 44994
rect 32398 44942 32450 44994
rect 33070 44942 33122 44994
rect 33742 44942 33794 44994
rect 41694 44942 41746 44994
rect 43822 44942 43874 44994
rect 47070 44942 47122 44994
rect 49086 44942 49138 44994
rect 49422 44942 49474 44994
rect 49758 44942 49810 44994
rect 11118 44830 11170 44882
rect 19854 44830 19906 44882
rect 20414 44830 20466 44882
rect 26126 44830 26178 44882
rect 30046 44830 30098 44882
rect 33182 44830 33234 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 7422 44494 7474 44546
rect 22878 44494 22930 44546
rect 25342 44494 25394 44546
rect 41918 44494 41970 44546
rect 7646 44382 7698 44434
rect 20302 44382 20354 44434
rect 27022 44382 27074 44434
rect 30606 44382 30658 44434
rect 31502 44382 31554 44434
rect 33630 44382 33682 44434
rect 37774 44382 37826 44434
rect 42030 44382 42082 44434
rect 42478 44382 42530 44434
rect 43486 44382 43538 44434
rect 49758 44382 49810 44434
rect 50542 44382 50594 44434
rect 51998 44382 52050 44434
rect 53006 44382 53058 44434
rect 53678 44382 53730 44434
rect 58158 44382 58210 44434
rect 7870 44270 7922 44322
rect 8878 44270 8930 44322
rect 9662 44270 9714 44322
rect 10110 44270 10162 44322
rect 10670 44270 10722 44322
rect 14254 44270 14306 44322
rect 15150 44270 15202 44322
rect 15486 44270 15538 44322
rect 16270 44270 16322 44322
rect 17390 44270 17442 44322
rect 22990 44270 23042 44322
rect 23438 44270 23490 44322
rect 24558 44270 24610 44322
rect 26462 44270 26514 44322
rect 30270 44270 30322 44322
rect 30942 44270 30994 44322
rect 34414 44270 34466 44322
rect 40686 44270 40738 44322
rect 42814 44270 42866 44322
rect 43038 44270 43090 44322
rect 43374 44270 43426 44322
rect 44046 44270 44098 44322
rect 45502 44270 45554 44322
rect 51550 44270 51602 44322
rect 51774 44270 51826 44322
rect 52110 44270 52162 44322
rect 52782 44270 52834 44322
rect 53566 44270 53618 44322
rect 54350 44270 54402 44322
rect 54686 44270 54738 44322
rect 55246 44270 55298 44322
rect 7310 44158 7362 44210
rect 8206 44158 8258 44210
rect 8430 44158 8482 44210
rect 9102 44158 9154 44210
rect 9438 44158 9490 44210
rect 15934 44158 15986 44210
rect 16606 44158 16658 44210
rect 18174 44158 18226 44210
rect 25790 44158 25842 44210
rect 27358 44158 27410 44210
rect 27806 44158 27858 44210
rect 36318 44158 36370 44210
rect 39902 44158 39954 44210
rect 54462 44158 54514 44210
rect 56030 44158 56082 44210
rect 8542 44046 8594 44098
rect 9214 44046 9266 44098
rect 9998 44046 10050 44098
rect 10222 44046 10274 44098
rect 14590 44046 14642 44098
rect 14702 44046 14754 44098
rect 14814 44046 14866 44098
rect 22878 44046 22930 44098
rect 30494 44046 30546 44098
rect 30718 44046 30770 44098
rect 36206 44046 36258 44098
rect 42478 44046 42530 44098
rect 42590 44046 42642 44098
rect 43598 44046 43650 44098
rect 43822 44046 43874 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 17950 43710 18002 43762
rect 31166 43710 31218 43762
rect 32174 43710 32226 43762
rect 39902 43710 39954 43762
rect 6862 43598 6914 43650
rect 10334 43598 10386 43650
rect 15374 43598 15426 43650
rect 16382 43598 16434 43650
rect 29822 43598 29874 43650
rect 31838 43598 31890 43650
rect 35422 43598 35474 43650
rect 38222 43598 38274 43650
rect 39342 43598 39394 43650
rect 39566 43598 39618 43650
rect 44270 43598 44322 43650
rect 54910 43598 54962 43650
rect 55022 43598 55074 43650
rect 57038 43598 57090 43650
rect 7646 43486 7698 43538
rect 13582 43486 13634 43538
rect 15598 43486 15650 43538
rect 16046 43486 16098 43538
rect 18062 43486 18114 43538
rect 30606 43498 30658 43550
rect 32062 43486 32114 43538
rect 32286 43486 32338 43538
rect 32398 43486 32450 43538
rect 34638 43486 34690 43538
rect 37998 43486 38050 43538
rect 38110 43486 38162 43538
rect 38334 43486 38386 43538
rect 38558 43486 38610 43538
rect 38894 43486 38946 43538
rect 39118 43486 39170 43538
rect 45390 43486 45442 43538
rect 50766 43486 50818 43538
rect 51998 43486 52050 43538
rect 52446 43486 52498 43538
rect 53118 43486 53170 43538
rect 54574 43486 54626 43538
rect 4734 43374 4786 43426
rect 15822 43374 15874 43426
rect 25678 43374 25730 43426
rect 27694 43374 27746 43426
rect 33182 43374 33234 43426
rect 37550 43374 37602 43426
rect 39230 43374 39282 43426
rect 40014 43374 40066 43426
rect 43262 43374 43314 43426
rect 44718 43374 44770 43426
rect 46062 43374 46114 43426
rect 48190 43374 48242 43426
rect 50318 43374 50370 43426
rect 53902 43374 53954 43426
rect 25566 43262 25618 43314
rect 54462 43262 54514 43314
rect 56926 43262 56978 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 9550 42926 9602 42978
rect 46286 42926 46338 42978
rect 46734 42926 46786 42978
rect 51550 42926 51602 42978
rect 52782 42926 52834 42978
rect 55918 42926 55970 42978
rect 56926 42926 56978 42978
rect 18734 42814 18786 42866
rect 21422 42814 21474 42866
rect 25118 42814 25170 42866
rect 27246 42814 27298 42866
rect 36430 42814 36482 42866
rect 51326 42814 51378 42866
rect 9998 42702 10050 42754
rect 10222 42702 10274 42754
rect 13806 42702 13858 42754
rect 14366 42702 14418 42754
rect 20750 42702 20802 42754
rect 24334 42702 24386 42754
rect 30606 42702 30658 42754
rect 30830 42702 30882 42754
rect 31278 42702 31330 42754
rect 33630 42702 33682 42754
rect 37550 42702 37602 42754
rect 37998 42702 38050 42754
rect 46286 42702 46338 42754
rect 46958 42702 47010 42754
rect 50766 42702 50818 42754
rect 50990 42702 51042 42754
rect 51774 42702 51826 42754
rect 52894 42702 52946 42754
rect 53230 42702 53282 42754
rect 56142 42702 56194 42754
rect 10110 42590 10162 42642
rect 10670 42590 10722 42642
rect 11006 42590 11058 42642
rect 14142 42590 14194 42642
rect 22094 42590 22146 42642
rect 29262 42590 29314 42642
rect 29934 42590 29986 42642
rect 30942 42590 30994 42642
rect 34302 42590 34354 42642
rect 46174 42590 46226 42642
rect 52782 42590 52834 42642
rect 53342 42590 53394 42642
rect 55358 42590 55410 42642
rect 55582 42590 55634 42642
rect 56814 42590 56866 42642
rect 13918 42478 13970 42530
rect 21982 42478 22034 42530
rect 27806 42478 27858 42530
rect 29150 42478 29202 42530
rect 29598 42478 29650 42530
rect 31054 42478 31106 42530
rect 31838 42478 31890 42530
rect 37662 42478 37714 42530
rect 37774 42478 37826 42530
rect 37886 42478 37938 42530
rect 38670 42478 38722 42530
rect 39006 42478 39058 42530
rect 39790 42478 39842 42530
rect 45950 42478 46002 42530
rect 55134 42478 55186 42530
rect 56254 42478 56306 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 32062 42142 32114 42194
rect 38110 42142 38162 42194
rect 44830 42142 44882 42194
rect 45278 42142 45330 42194
rect 45502 42142 45554 42194
rect 48078 42142 48130 42194
rect 24110 42030 24162 42082
rect 26014 42030 26066 42082
rect 26462 42030 26514 42082
rect 26910 42030 26962 42082
rect 28702 42030 28754 42082
rect 32286 42030 32338 42082
rect 45166 42030 45218 42082
rect 47966 42030 48018 42082
rect 12014 41918 12066 41970
rect 12686 41918 12738 41970
rect 15374 41918 15426 41970
rect 20414 41918 20466 41970
rect 21198 41918 21250 41970
rect 23774 41918 23826 41970
rect 23886 41918 23938 41970
rect 23998 41918 24050 41970
rect 24222 41918 24274 41970
rect 25790 41918 25842 41970
rect 26238 41918 26290 41970
rect 27246 41918 27298 41970
rect 27918 41918 27970 41970
rect 31838 41918 31890 41970
rect 32398 41918 32450 41970
rect 35310 41918 35362 41970
rect 35422 41918 35474 41970
rect 37214 41918 37266 41970
rect 37550 41918 37602 41970
rect 37774 41918 37826 41970
rect 37998 41918 38050 41970
rect 40910 41918 40962 41970
rect 47630 41918 47682 41970
rect 48974 41918 49026 41970
rect 52222 41918 52274 41970
rect 14814 41806 14866 41858
rect 15262 41806 15314 41858
rect 18622 41806 18674 41858
rect 23326 41806 23378 41858
rect 25342 41806 25394 41858
rect 25902 41806 25954 41858
rect 30830 41806 30882 41858
rect 32286 41806 32338 41858
rect 33070 41806 33122 41858
rect 33630 41806 33682 41858
rect 37886 41806 37938 41858
rect 41694 41806 41746 41858
rect 43822 41806 43874 41858
rect 44494 41806 44546 41858
rect 47182 41806 47234 41858
rect 49646 41806 49698 41858
rect 51774 41806 51826 41858
rect 52894 41806 52946 41858
rect 55022 41806 55074 41858
rect 16606 41694 16658 41746
rect 18734 41694 18786 41746
rect 33182 41694 33234 41746
rect 47518 41694 47570 41746
rect 48078 41694 48130 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 49086 41358 49138 41410
rect 49646 41358 49698 41410
rect 9214 41246 9266 41298
rect 11342 41246 11394 41298
rect 16494 41246 16546 41298
rect 17502 41246 17554 41298
rect 19630 41246 19682 41298
rect 29374 41246 29426 41298
rect 31390 41246 31442 41298
rect 33518 41246 33570 41298
rect 37214 41246 37266 41298
rect 40910 41246 40962 41298
rect 48078 41246 48130 41298
rect 49422 41246 49474 41298
rect 8430 41134 8482 41186
rect 15822 41134 15874 41186
rect 16382 41134 16434 41186
rect 20414 41134 20466 41186
rect 25790 41134 25842 41186
rect 26126 41134 26178 41186
rect 34302 41134 34354 41186
rect 43150 41134 43202 41186
rect 43486 41134 43538 41186
rect 43710 41134 43762 41186
rect 44046 41134 44098 41186
rect 45166 41134 45218 41186
rect 49870 41134 49922 41186
rect 51214 41134 51266 41186
rect 51550 41134 51602 41186
rect 52670 41134 52722 41186
rect 12798 41022 12850 41074
rect 26350 41022 26402 41074
rect 27470 41022 27522 41074
rect 29486 41022 29538 41074
rect 30158 41022 30210 41074
rect 30494 41022 30546 41074
rect 37102 41022 37154 41074
rect 45950 41022 46002 41074
rect 49310 41022 49362 41074
rect 51662 41022 51714 41074
rect 55470 41022 55522 41074
rect 12686 40910 12738 40962
rect 25006 40910 25058 40962
rect 25342 40910 25394 40962
rect 25902 40910 25954 40962
rect 26014 40910 26066 40962
rect 26910 40910 26962 40962
rect 27806 40910 27858 40962
rect 28702 40910 28754 40962
rect 29262 40910 29314 40962
rect 43822 40910 43874 40962
rect 43934 40910 43986 40962
rect 48750 40910 48802 40962
rect 51886 40910 51938 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 17502 40574 17554 40626
rect 18846 40574 18898 40626
rect 18958 40574 19010 40626
rect 19630 40574 19682 40626
rect 24222 40574 24274 40626
rect 38894 40574 38946 40626
rect 39566 40574 39618 40626
rect 40350 40574 40402 40626
rect 41022 40574 41074 40626
rect 42254 40574 42306 40626
rect 43374 40574 43426 40626
rect 44270 40574 44322 40626
rect 49758 40574 49810 40626
rect 52334 40574 52386 40626
rect 54238 40574 54290 40626
rect 54910 40574 54962 40626
rect 8318 40462 8370 40514
rect 12126 40462 12178 40514
rect 18510 40462 18562 40514
rect 27918 40462 27970 40514
rect 36430 40462 36482 40514
rect 41918 40462 41970 40514
rect 42366 40462 42418 40514
rect 44830 40462 44882 40514
rect 44942 40462 44994 40514
rect 45838 40462 45890 40514
rect 53006 40462 53058 40514
rect 54686 40462 54738 40514
rect 55806 40462 55858 40514
rect 57822 40462 57874 40514
rect 4958 40350 5010 40402
rect 9662 40350 9714 40402
rect 11454 40350 11506 40402
rect 16158 40350 16210 40402
rect 16382 40350 16434 40402
rect 16606 40350 16658 40402
rect 16830 40350 16882 40402
rect 18734 40350 18786 40402
rect 19070 40350 19122 40402
rect 20862 40350 20914 40402
rect 24110 40350 24162 40402
rect 24446 40350 24498 40402
rect 24670 40350 24722 40402
rect 29038 40350 29090 40402
rect 35758 40350 35810 40402
rect 39118 40350 39170 40402
rect 39902 40350 39954 40402
rect 41694 40350 41746 40402
rect 43934 40350 43986 40402
rect 45166 40350 45218 40402
rect 45502 40350 45554 40402
rect 45614 40350 45666 40402
rect 46062 40350 46114 40402
rect 49422 40350 49474 40402
rect 51886 40350 51938 40402
rect 52782 40350 52834 40402
rect 53230 40350 53282 40402
rect 54574 40350 54626 40402
rect 57598 40350 57650 40402
rect 58046 40350 58098 40402
rect 14254 40238 14306 40290
rect 16494 40238 16546 40290
rect 21534 40238 21586 40290
rect 23662 40238 23714 40290
rect 24334 40238 24386 40290
rect 34526 40238 34578 40290
rect 38558 40238 38610 40290
rect 40910 40238 40962 40290
rect 46286 40238 46338 40290
rect 53454 40238 53506 40290
rect 55246 40238 55298 40290
rect 41246 40126 41298 40178
rect 52670 40126 52722 40178
rect 55470 40126 55522 40178
rect 55918 40126 55970 40178
rect 56030 40126 56082 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 22318 39790 22370 39842
rect 34526 39790 34578 39842
rect 34750 39790 34802 39842
rect 4622 39678 4674 39730
rect 5630 39678 5682 39730
rect 16382 39678 16434 39730
rect 22430 39678 22482 39730
rect 24782 39678 24834 39730
rect 28142 39678 28194 39730
rect 29710 39678 29762 39730
rect 38110 39678 38162 39730
rect 38558 39678 38610 39730
rect 45390 39678 45442 39730
rect 53118 39678 53170 39730
rect 53678 39678 53730 39730
rect 54350 39678 54402 39730
rect 56030 39678 56082 39730
rect 58158 39678 58210 39730
rect 1822 39566 1874 39618
rect 8430 39566 8482 39618
rect 13470 39566 13522 39618
rect 16718 39566 16770 39618
rect 17166 39566 17218 39618
rect 17278 39566 17330 39618
rect 17838 39566 17890 39618
rect 25342 39566 25394 39618
rect 35310 39566 35362 39618
rect 35758 39566 35810 39618
rect 41022 39566 41074 39618
rect 41918 39566 41970 39618
rect 42142 39566 42194 39618
rect 42590 39566 42642 39618
rect 52670 39566 52722 39618
rect 54798 39566 54850 39618
rect 55246 39566 55298 39618
rect 2494 39454 2546 39506
rect 7758 39454 7810 39506
rect 8878 39454 8930 39506
rect 8990 39454 9042 39506
rect 9662 39454 9714 39506
rect 14254 39454 14306 39506
rect 16942 39454 16994 39506
rect 18734 39454 18786 39506
rect 24894 39454 24946 39506
rect 26014 39454 26066 39506
rect 29262 39454 29314 39506
rect 33518 39454 33570 39506
rect 33742 39454 33794 39506
rect 34078 39454 34130 39506
rect 41358 39454 41410 39506
rect 48526 39454 48578 39506
rect 9214 39342 9266 39394
rect 9326 39342 9378 39394
rect 9550 39342 9602 39394
rect 17054 39342 17106 39394
rect 19070 39342 19122 39394
rect 19630 39342 19682 39394
rect 29150 39342 29202 39394
rect 33182 39342 33234 39394
rect 33406 39342 33458 39394
rect 33966 39342 34018 39394
rect 34526 39342 34578 39394
rect 36318 39342 36370 39394
rect 37774 39342 37826 39394
rect 42254 39342 42306 39394
rect 42366 39342 42418 39394
rect 43150 39342 43202 39394
rect 44942 39342 44994 39394
rect 47406 39342 47458 39394
rect 48638 39342 48690 39394
rect 48862 39342 48914 39394
rect 49086 39342 49138 39394
rect 49422 39342 49474 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 5966 39006 6018 39058
rect 7534 39006 7586 39058
rect 14702 39006 14754 39058
rect 19070 39006 19122 39058
rect 19630 39006 19682 39058
rect 36990 39006 37042 39058
rect 37214 39006 37266 39058
rect 37886 39006 37938 39058
rect 38222 39006 38274 39058
rect 45390 39006 45442 39058
rect 46622 39006 46674 39058
rect 55470 39006 55522 39058
rect 55918 39006 55970 39058
rect 56142 39006 56194 39058
rect 5182 38894 5234 38946
rect 5294 38894 5346 38946
rect 5742 38894 5794 38946
rect 7310 38894 7362 38946
rect 14814 38894 14866 38946
rect 18510 38894 18562 38946
rect 30270 38894 30322 38946
rect 32510 38894 32562 38946
rect 34862 38894 34914 38946
rect 35758 38894 35810 38946
rect 49310 38894 49362 38946
rect 55806 38894 55858 38946
rect 1822 38782 1874 38834
rect 5630 38782 5682 38834
rect 6190 38782 6242 38834
rect 6302 38782 6354 38834
rect 6414 38782 6466 38834
rect 6750 38782 6802 38834
rect 7198 38782 7250 38834
rect 7646 38782 7698 38834
rect 8542 38782 8594 38834
rect 8766 38782 8818 38834
rect 9102 38782 9154 38834
rect 12462 38782 12514 38834
rect 18734 38782 18786 38834
rect 18958 38782 19010 38834
rect 20414 38782 20466 38834
rect 26910 38782 26962 38834
rect 30606 38782 30658 38834
rect 34974 38782 35026 38834
rect 36654 38782 36706 38834
rect 37550 38782 37602 38834
rect 39230 38782 39282 38834
rect 43822 38782 43874 38834
rect 45726 38782 45778 38834
rect 45950 38782 46002 38834
rect 46286 38782 46338 38834
rect 46846 38782 46898 38834
rect 47518 38782 47570 38834
rect 47966 38782 48018 38834
rect 48190 38782 48242 38834
rect 48750 38782 48802 38834
rect 48862 38782 48914 38834
rect 48974 38782 49026 38834
rect 52894 38782 52946 38834
rect 54910 38782 54962 38834
rect 57710 38782 57762 38834
rect 2494 38670 2546 38722
rect 4622 38670 4674 38722
rect 8878 38670 8930 38722
rect 9550 38670 9602 38722
rect 11678 38670 11730 38722
rect 18062 38670 18114 38722
rect 18846 38670 18898 38722
rect 20078 38670 20130 38722
rect 21198 38670 21250 38722
rect 23326 38670 23378 38722
rect 27582 38670 27634 38722
rect 29710 38670 29762 38722
rect 30382 38670 30434 38722
rect 35758 38670 35810 38722
rect 38670 38670 38722 38722
rect 40910 38670 40962 38722
rect 43038 38670 43090 38722
rect 45838 38670 45890 38722
rect 47742 38670 47794 38722
rect 49982 38670 50034 38722
rect 52110 38670 52162 38722
rect 57150 38670 57202 38722
rect 5182 38558 5234 38610
rect 17950 38558 18002 38610
rect 30046 38558 30098 38610
rect 30830 38558 30882 38610
rect 36878 38558 36930 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 7646 38222 7698 38274
rect 8766 38222 8818 38274
rect 34190 38222 34242 38274
rect 34414 38222 34466 38274
rect 34974 38222 35026 38274
rect 42030 38222 42082 38274
rect 5854 38110 5906 38162
rect 17054 38110 17106 38162
rect 19182 38110 19234 38162
rect 23662 38110 23714 38162
rect 28030 38110 28082 38162
rect 33518 38110 33570 38162
rect 34078 38110 34130 38162
rect 34750 38110 34802 38162
rect 40014 38110 40066 38162
rect 41918 38110 41970 38162
rect 43710 38110 43762 38162
rect 44270 38110 44322 38162
rect 45054 38110 45106 38162
rect 6078 37998 6130 38050
rect 6526 37998 6578 38050
rect 6862 37998 6914 38050
rect 7534 37998 7586 38050
rect 8878 37998 8930 38050
rect 16382 37998 16434 38050
rect 22990 37998 23042 38050
rect 27582 37998 27634 38050
rect 30046 37998 30098 38050
rect 30606 37998 30658 38050
rect 35646 37998 35698 38050
rect 36318 37998 36370 38050
rect 37214 37998 37266 38050
rect 43598 37998 43650 38050
rect 48750 37998 48802 38050
rect 50542 37998 50594 38050
rect 55918 37998 55970 38050
rect 58158 37998 58210 38050
rect 5742 37886 5794 37938
rect 6302 37886 6354 37938
rect 11006 37886 11058 37938
rect 11342 37886 11394 37938
rect 28702 37886 28754 37938
rect 29262 37886 29314 37938
rect 29374 37886 29426 37938
rect 29710 37886 29762 37938
rect 31390 37886 31442 37938
rect 37886 37886 37938 37938
rect 54910 37886 54962 37938
rect 58046 37886 58098 37938
rect 6750 37774 6802 37826
rect 7646 37774 7698 37826
rect 8766 37774 8818 37826
rect 11902 37774 11954 37826
rect 22766 37774 22818 37826
rect 23102 37774 23154 37826
rect 23326 37774 23378 37826
rect 23550 37774 23602 37826
rect 23774 37774 23826 37826
rect 23998 37774 24050 37826
rect 29038 37774 29090 37826
rect 29822 37774 29874 37826
rect 35310 37774 35362 37826
rect 35982 37774 36034 37826
rect 54462 37774 54514 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 5518 37438 5570 37490
rect 5742 37438 5794 37490
rect 7198 37438 7250 37490
rect 4958 37326 5010 37378
rect 15710 37326 15762 37378
rect 18958 37326 19010 37378
rect 20750 37326 20802 37378
rect 22878 37326 22930 37378
rect 22990 37326 23042 37378
rect 28926 37326 28978 37378
rect 29038 37382 29090 37434
rect 32062 37438 32114 37490
rect 35982 37438 36034 37490
rect 36094 37438 36146 37490
rect 36990 37438 37042 37490
rect 37550 37438 37602 37490
rect 48862 37438 48914 37490
rect 36542 37326 36594 37378
rect 45614 37326 45666 37378
rect 48750 37326 48802 37378
rect 49310 37326 49362 37378
rect 4734 37214 4786 37266
rect 5070 37214 5122 37266
rect 5406 37214 5458 37266
rect 7534 37214 7586 37266
rect 8318 37214 8370 37266
rect 8542 37214 8594 37266
rect 11678 37214 11730 37266
rect 12574 37214 12626 37266
rect 16046 37214 16098 37266
rect 19518 37214 19570 37266
rect 19742 37214 19794 37266
rect 22542 37214 22594 37266
rect 23214 37214 23266 37266
rect 23438 37214 23490 37266
rect 23662 37214 23714 37266
rect 24110 37214 24162 37266
rect 28702 37214 28754 37266
rect 29486 37214 29538 37266
rect 31614 37214 31666 37266
rect 31950 37214 32002 37266
rect 32286 37214 32338 37266
rect 35310 37214 35362 37266
rect 35534 37214 35586 37266
rect 36206 37214 36258 37266
rect 36878 37214 36930 37266
rect 37102 37214 37154 37266
rect 42030 37214 42082 37266
rect 42590 37214 42642 37266
rect 44942 37214 44994 37266
rect 48974 37214 49026 37266
rect 56030 37214 56082 37266
rect 12126 37102 12178 37154
rect 13246 37102 13298 37154
rect 15374 37102 15426 37154
rect 20190 37102 20242 37154
rect 23550 37102 23602 37154
rect 28254 37102 28306 37154
rect 30158 37102 30210 37154
rect 31278 37102 31330 37154
rect 33182 37102 33234 37154
rect 38334 37102 38386 37154
rect 38670 37102 38722 37154
rect 43038 37102 43090 37154
rect 47742 37102 47794 37154
rect 48190 37102 48242 37154
rect 49758 37102 49810 37154
rect 53118 37102 53170 37154
rect 55246 37102 55298 37154
rect 56590 37102 56642 37154
rect 56702 37102 56754 37154
rect 58158 37102 58210 37154
rect 7982 36990 8034 37042
rect 8094 36990 8146 37042
rect 8654 36990 8706 37042
rect 49646 36990 49698 37042
rect 57822 36990 57874 37042
rect 58158 36990 58210 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 4622 36542 4674 36594
rect 12350 36542 12402 36594
rect 16382 36542 16434 36594
rect 27134 36542 27186 36594
rect 43374 36542 43426 36594
rect 44830 36542 44882 36594
rect 45950 36542 46002 36594
rect 49422 36542 49474 36594
rect 51550 36542 51602 36594
rect 52110 36542 52162 36594
rect 52782 36542 52834 36594
rect 54350 36542 54402 36594
rect 58158 36542 58210 36594
rect 1822 36430 1874 36482
rect 13582 36430 13634 36482
rect 13694 36430 13746 36482
rect 14142 36430 14194 36482
rect 16606 36430 16658 36482
rect 16718 36430 16770 36482
rect 20078 36430 20130 36482
rect 20526 36430 20578 36482
rect 24222 36430 24274 36482
rect 27358 36430 27410 36482
rect 28030 36430 28082 36482
rect 31950 36430 32002 36482
rect 32398 36430 32450 36482
rect 32622 36430 32674 36482
rect 33518 36430 33570 36482
rect 35198 36430 35250 36482
rect 35870 36430 35922 36482
rect 36318 36430 36370 36482
rect 38334 36430 38386 36482
rect 41582 36430 41634 36482
rect 42478 36430 42530 36482
rect 43822 36430 43874 36482
rect 45278 36430 45330 36482
rect 46286 36430 46338 36482
rect 48750 36430 48802 36482
rect 53902 36430 53954 36482
rect 55358 36430 55410 36482
rect 2494 36318 2546 36370
rect 5742 36318 5794 36370
rect 5854 36318 5906 36370
rect 25006 36318 25058 36370
rect 27806 36318 27858 36370
rect 35646 36318 35698 36370
rect 37998 36318 38050 36370
rect 46846 36318 46898 36370
rect 52782 36318 52834 36370
rect 53342 36318 53394 36370
rect 54910 36318 54962 36370
rect 56030 36318 56082 36370
rect 5518 36206 5570 36258
rect 13806 36206 13858 36258
rect 15374 36206 15426 36258
rect 15710 36206 15762 36258
rect 17502 36206 17554 36258
rect 21422 36206 21474 36258
rect 27582 36206 27634 36258
rect 28478 36206 28530 36258
rect 31838 36206 31890 36258
rect 32510 36206 32562 36258
rect 33070 36206 33122 36258
rect 33294 36206 33346 36258
rect 33406 36206 33458 36258
rect 33966 36206 34018 36258
rect 34974 36206 35026 36258
rect 35758 36206 35810 36258
rect 38110 36206 38162 36258
rect 39230 36206 39282 36258
rect 42142 36206 42194 36258
rect 43038 36206 43090 36258
rect 51998 36206 52050 36258
rect 52894 36206 52946 36258
rect 53118 36206 53170 36258
rect 54014 36206 54066 36258
rect 54238 36206 54290 36258
rect 54350 36206 54402 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 4510 35870 4562 35922
rect 8318 35870 8370 35922
rect 8542 35870 8594 35922
rect 10558 35870 10610 35922
rect 13358 35870 13410 35922
rect 13694 35870 13746 35922
rect 13806 35870 13858 35922
rect 14254 35870 14306 35922
rect 15374 35870 15426 35922
rect 22878 35870 22930 35922
rect 26126 35870 26178 35922
rect 28702 35870 28754 35922
rect 29038 35870 29090 35922
rect 33182 35870 33234 35922
rect 40238 35870 40290 35922
rect 44158 35870 44210 35922
rect 47182 35870 47234 35922
rect 54910 35870 54962 35922
rect 55582 35870 55634 35922
rect 4734 35758 4786 35810
rect 6078 35758 6130 35810
rect 7758 35758 7810 35810
rect 7870 35758 7922 35810
rect 8206 35758 8258 35810
rect 8878 35758 8930 35810
rect 10110 35758 10162 35810
rect 15150 35758 15202 35810
rect 16270 35758 16322 35810
rect 20638 35758 20690 35810
rect 26574 35758 26626 35810
rect 27694 35758 27746 35810
rect 30046 35758 30098 35810
rect 32510 35758 32562 35810
rect 35870 35758 35922 35810
rect 41806 35758 41858 35810
rect 47854 35758 47906 35810
rect 48974 35758 49026 35810
rect 55134 35758 55186 35810
rect 4286 35646 4338 35698
rect 4958 35646 5010 35698
rect 5294 35646 5346 35698
rect 5518 35646 5570 35698
rect 5742 35646 5794 35698
rect 8766 35646 8818 35698
rect 9102 35646 9154 35698
rect 9438 35646 9490 35698
rect 9886 35646 9938 35698
rect 13582 35646 13634 35698
rect 15374 35646 15426 35698
rect 15710 35646 15762 35698
rect 16158 35646 16210 35698
rect 16382 35646 16434 35698
rect 19966 35646 20018 35698
rect 26014 35646 26066 35698
rect 26350 35646 26402 35698
rect 28030 35646 28082 35698
rect 28366 35646 28418 35698
rect 31950 35646 32002 35698
rect 32174 35646 32226 35698
rect 36206 35646 36258 35698
rect 36430 35646 36482 35698
rect 38222 35646 38274 35698
rect 38558 35646 38610 35698
rect 39006 35646 39058 35698
rect 39454 35646 39506 35698
rect 39678 35646 39730 35698
rect 39790 35646 39842 35698
rect 42142 35646 42194 35698
rect 46846 35646 46898 35698
rect 47518 35646 47570 35698
rect 52894 35646 52946 35698
rect 54462 35646 54514 35698
rect 54686 35646 54738 35698
rect 56030 35646 56082 35698
rect 5966 35534 6018 35586
rect 9662 35534 9714 35586
rect 27022 35534 27074 35586
rect 29598 35534 29650 35586
rect 32062 35534 32114 35586
rect 36318 35534 36370 35586
rect 42590 35534 42642 35586
rect 43262 35534 43314 35586
rect 45614 35534 45666 35586
rect 54798 35534 54850 35586
rect 55470 35534 55522 35586
rect 56702 35534 56754 35586
rect 7758 35422 7810 35474
rect 16830 35422 16882 35474
rect 29374 35422 29426 35474
rect 37886 35422 37938 35474
rect 38894 35422 38946 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 28030 35086 28082 35138
rect 28366 35086 28418 35138
rect 41246 35086 41298 35138
rect 41582 35086 41634 35138
rect 8430 34974 8482 35026
rect 10558 34974 10610 35026
rect 16494 34974 16546 35026
rect 30494 34974 30546 35026
rect 37774 34974 37826 35026
rect 39902 34974 39954 35026
rect 40462 34974 40514 35026
rect 49758 34974 49810 35026
rect 5182 34862 5234 34914
rect 5854 34862 5906 34914
rect 6078 34862 6130 34914
rect 11342 34862 11394 34914
rect 17390 34862 17442 34914
rect 19182 34862 19234 34914
rect 25678 34862 25730 34914
rect 26014 34862 26066 34914
rect 28590 34862 28642 34914
rect 29710 34862 29762 34914
rect 33070 34862 33122 34914
rect 33630 34862 33682 34914
rect 34638 34862 34690 34914
rect 34750 34862 34802 34914
rect 37102 34862 37154 34914
rect 41918 34862 41970 34914
rect 42142 34862 42194 34914
rect 43262 34862 43314 34914
rect 49646 34862 49698 34914
rect 49982 34862 50034 34914
rect 50206 34862 50258 34914
rect 52110 34862 52162 34914
rect 52894 34862 52946 34914
rect 4286 34750 4338 34802
rect 4622 34750 4674 34802
rect 4846 34750 4898 34802
rect 4958 34750 5010 34802
rect 5630 34750 5682 34802
rect 33518 34750 33570 34802
rect 42366 34750 42418 34802
rect 42590 34750 42642 34802
rect 43150 34750 43202 34802
rect 55470 34750 55522 34802
rect 4398 34638 4450 34690
rect 5742 34638 5794 34690
rect 25790 34638 25842 34690
rect 26462 34638 26514 34690
rect 27246 34638 27298 34690
rect 32734 34638 32786 34690
rect 33294 34638 33346 34690
rect 35086 34638 35138 34690
rect 40910 34638 40962 34690
rect 41470 34638 41522 34690
rect 42254 34638 42306 34690
rect 48414 34638 48466 34690
rect 49198 34638 49250 34690
rect 49758 34638 49810 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 8542 34302 8594 34354
rect 16382 34302 16434 34354
rect 33630 34302 33682 34354
rect 34638 34302 34690 34354
rect 36094 34302 36146 34354
rect 39342 34302 39394 34354
rect 41806 34302 41858 34354
rect 11342 34190 11394 34242
rect 27918 34190 27970 34242
rect 33182 34190 33234 34242
rect 34078 34190 34130 34242
rect 35198 34190 35250 34242
rect 38222 34190 38274 34242
rect 39566 34190 39618 34242
rect 43934 34190 43986 34242
rect 46398 34190 46450 34242
rect 51998 34190 52050 34242
rect 8206 34078 8258 34130
rect 8766 34078 8818 34130
rect 9662 34078 9714 34130
rect 11118 34078 11170 34130
rect 11790 34078 11842 34130
rect 16270 34078 16322 34130
rect 19518 34078 19570 34130
rect 20302 34078 20354 34130
rect 21870 34078 21922 34130
rect 26686 34078 26738 34130
rect 27582 34078 27634 34130
rect 35086 34078 35138 34130
rect 38894 34078 38946 34130
rect 41582 34078 41634 34130
rect 43262 34078 43314 34130
rect 47630 34078 47682 34130
rect 51214 34078 51266 34130
rect 4958 33966 5010 34018
rect 12462 33966 12514 34018
rect 14590 33966 14642 34018
rect 15710 33966 15762 34018
rect 17390 33966 17442 34018
rect 22542 33966 22594 34018
rect 24670 33966 24722 34018
rect 27246 33966 27298 34018
rect 28366 33966 28418 34018
rect 33742 33966 33794 34018
rect 46062 33966 46114 34018
rect 47294 33966 47346 34018
rect 54126 33966 54178 34018
rect 54574 33966 54626 34018
rect 16046 33854 16098 33906
rect 16382 33854 16434 33906
rect 33294 33854 33346 33906
rect 34302 33854 34354 33906
rect 39230 33854 39282 33906
rect 46510 33854 46562 33906
rect 47630 33854 47682 33906
rect 47966 33854 48018 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 12350 33518 12402 33570
rect 35758 33518 35810 33570
rect 37774 33518 37826 33570
rect 38670 33518 38722 33570
rect 39006 33518 39058 33570
rect 2494 33406 2546 33458
rect 4622 33406 4674 33458
rect 9886 33406 9938 33458
rect 11678 33406 11730 33458
rect 12462 33406 12514 33458
rect 20862 33406 20914 33458
rect 21870 33406 21922 33458
rect 36094 33406 36146 33458
rect 41918 33406 41970 33458
rect 47406 33406 47458 33458
rect 49534 33406 49586 33458
rect 50766 33406 50818 33458
rect 54798 33406 54850 33458
rect 56030 33406 56082 33458
rect 58158 33406 58210 33458
rect 1822 33294 1874 33346
rect 6414 33294 6466 33346
rect 6974 33294 7026 33346
rect 12686 33294 12738 33346
rect 25230 33294 25282 33346
rect 27470 33294 27522 33346
rect 29710 33294 29762 33346
rect 29934 33294 29986 33346
rect 37550 33294 37602 33346
rect 38446 33294 38498 33346
rect 41806 33294 41858 33346
rect 42030 33294 42082 33346
rect 42254 33294 42306 33346
rect 42926 33294 42978 33346
rect 46622 33294 46674 33346
rect 51886 33294 51938 33346
rect 53006 33294 53058 33346
rect 53342 33294 53394 33346
rect 53566 33294 53618 33346
rect 54910 33294 54962 33346
rect 55358 33294 55410 33346
rect 7758 33182 7810 33234
rect 16606 33182 16658 33234
rect 20302 33182 20354 33234
rect 27694 33182 27746 33234
rect 31950 33182 32002 33234
rect 35982 33182 36034 33234
rect 42478 33182 42530 33234
rect 49982 33182 50034 33234
rect 50318 33182 50370 33234
rect 52670 33182 52722 33234
rect 52782 33182 52834 33234
rect 54238 33182 54290 33234
rect 54574 33182 54626 33234
rect 6078 33070 6130 33122
rect 16382 33070 16434 33122
rect 16494 33070 16546 33122
rect 20190 33070 20242 33122
rect 28254 33070 28306 33122
rect 38110 33070 38162 33122
rect 50878 33070 50930 33122
rect 52110 33070 52162 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 5742 32734 5794 32786
rect 5966 32734 6018 32786
rect 17390 32734 17442 32786
rect 22430 32734 22482 32786
rect 22654 32734 22706 32786
rect 23326 32734 23378 32786
rect 23550 32734 23602 32786
rect 25230 32734 25282 32786
rect 31166 32734 31218 32786
rect 31838 32734 31890 32786
rect 34190 32734 34242 32786
rect 50766 32734 50818 32786
rect 50878 32734 50930 32786
rect 51774 32734 51826 32786
rect 54014 32734 54066 32786
rect 54238 32734 54290 32786
rect 57374 32734 57426 32786
rect 58158 32734 58210 32786
rect 5294 32622 5346 32674
rect 14702 32622 14754 32674
rect 19630 32622 19682 32674
rect 22318 32622 22370 32674
rect 24446 32622 24498 32674
rect 25678 32622 25730 32674
rect 30942 32622 30994 32674
rect 34638 32622 34690 32674
rect 41358 32622 41410 32674
rect 48190 32622 48242 32674
rect 49198 32622 49250 32674
rect 50318 32622 50370 32674
rect 51998 32622 52050 32674
rect 52670 32622 52722 32674
rect 1822 32510 1874 32562
rect 4846 32510 4898 32562
rect 5518 32510 5570 32562
rect 6078 32510 6130 32562
rect 13918 32510 13970 32562
rect 17726 32510 17778 32562
rect 18958 32510 19010 32562
rect 22094 32510 22146 32562
rect 22542 32510 22594 32562
rect 24110 32510 24162 32562
rect 24222 32510 24274 32562
rect 24670 32510 24722 32562
rect 25454 32510 25506 32562
rect 27582 32510 27634 32562
rect 30718 32510 30770 32562
rect 31278 32510 31330 32562
rect 33854 32510 33906 32562
rect 34078 32510 34130 32562
rect 41806 32510 41858 32562
rect 47742 32510 47794 32562
rect 49086 32510 49138 32562
rect 49758 32510 49810 32562
rect 50542 32510 50594 32562
rect 51662 32510 51714 32562
rect 52222 32510 52274 32562
rect 52558 32510 52610 32562
rect 53118 32510 53170 32562
rect 54462 32510 54514 32562
rect 2494 32398 2546 32450
rect 4622 32398 4674 32450
rect 5070 32398 5122 32450
rect 16830 32398 16882 32450
rect 17950 32398 18002 32450
rect 21758 32398 21810 32450
rect 23662 32398 23714 32450
rect 24334 32398 24386 32450
rect 25342 32398 25394 32450
rect 26350 32398 26402 32450
rect 28254 32398 28306 32450
rect 30382 32398 30434 32450
rect 31054 32398 31106 32450
rect 41470 32398 41522 32450
rect 42590 32398 42642 32450
rect 44718 32398 44770 32450
rect 47294 32398 47346 32450
rect 49646 32398 49698 32450
rect 50878 32398 50930 32450
rect 51886 32398 51938 32450
rect 57710 32398 57762 32450
rect 53342 32286 53394 32338
rect 53678 32286 53730 32338
rect 53902 32286 53954 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 4846 31950 4898 32002
rect 35198 31950 35250 32002
rect 37214 31950 37266 32002
rect 7758 31838 7810 31890
rect 9998 31838 10050 31890
rect 16830 31838 16882 31890
rect 24110 31838 24162 31890
rect 26238 31838 26290 31890
rect 29150 31838 29202 31890
rect 29262 31838 29314 31890
rect 32286 31838 32338 31890
rect 34414 31838 34466 31890
rect 35422 31838 35474 31890
rect 36990 31838 37042 31890
rect 41806 31838 41858 31890
rect 47742 31838 47794 31890
rect 52670 31838 52722 31890
rect 54462 31838 54514 31890
rect 58158 31838 58210 31890
rect 4174 31726 4226 31778
rect 7310 31726 7362 31778
rect 8206 31726 8258 31778
rect 8542 31726 8594 31778
rect 12910 31726 12962 31778
rect 22206 31726 22258 31778
rect 22430 31726 22482 31778
rect 22542 31726 22594 31778
rect 23326 31726 23378 31778
rect 31502 31726 31554 31778
rect 35086 31726 35138 31778
rect 35310 31726 35362 31778
rect 43822 31726 43874 31778
rect 44382 31726 44434 31778
rect 44942 31726 44994 31778
rect 48638 31726 48690 31778
rect 48750 31726 48802 31778
rect 53006 31726 53058 31778
rect 53230 31726 53282 31778
rect 54238 31726 54290 31778
rect 54686 31726 54738 31778
rect 55358 31726 55410 31778
rect 4286 31502 4338 31554
rect 4510 31502 4562 31554
rect 4734 31558 4786 31610
rect 4846 31614 4898 31666
rect 7870 31614 7922 31666
rect 8654 31614 8706 31666
rect 12126 31614 12178 31666
rect 16718 31614 16770 31666
rect 20414 31614 20466 31666
rect 21982 31614 22034 31666
rect 22318 31614 22370 31666
rect 30830 31614 30882 31666
rect 45614 31614 45666 31666
rect 48190 31614 48242 31666
rect 49534 31614 49586 31666
rect 52782 31614 52834 31666
rect 53678 31614 53730 31666
rect 54798 31614 54850 31666
rect 56030 31614 56082 31666
rect 5630 31502 5682 31554
rect 5966 31502 6018 31554
rect 7646 31502 7698 31554
rect 8766 31502 8818 31554
rect 16942 31502 16994 31554
rect 17166 31502 17218 31554
rect 20302 31502 20354 31554
rect 31166 31502 31218 31554
rect 37550 31502 37602 31554
rect 48414 31502 48466 31554
rect 48526 31502 48578 31554
rect 49198 31502 49250 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 5966 31166 6018 31218
rect 7758 31166 7810 31218
rect 8206 31166 8258 31218
rect 11230 31166 11282 31218
rect 17390 31166 17442 31218
rect 17838 31166 17890 31218
rect 22990 31166 23042 31218
rect 25678 31166 25730 31218
rect 30718 31166 30770 31218
rect 31726 31166 31778 31218
rect 33182 31166 33234 31218
rect 34750 31166 34802 31218
rect 35534 31166 35586 31218
rect 41358 31166 41410 31218
rect 41582 31166 41634 31218
rect 41694 31166 41746 31218
rect 42366 31166 42418 31218
rect 42590 31166 42642 31218
rect 47518 31166 47570 31218
rect 52894 31166 52946 31218
rect 4510 31054 4562 31106
rect 4734 31054 4786 31106
rect 5630 31054 5682 31106
rect 9550 31054 9602 31106
rect 9886 31054 9938 31106
rect 10558 31054 10610 31106
rect 10782 31054 10834 31106
rect 19742 31054 19794 31106
rect 22430 31054 22482 31106
rect 33854 31054 33906 31106
rect 34862 31054 34914 31106
rect 35982 31054 36034 31106
rect 45502 31054 45554 31106
rect 47406 31054 47458 31106
rect 48750 31054 48802 31106
rect 53342 31054 53394 31106
rect 5182 30942 5234 30994
rect 7534 30942 7586 30994
rect 8542 30942 8594 30994
rect 10446 30942 10498 30994
rect 10894 30942 10946 30994
rect 11230 30942 11282 30994
rect 11454 30942 11506 30994
rect 13022 30942 13074 30994
rect 17614 30942 17666 30994
rect 18958 30942 19010 30994
rect 25342 30942 25394 30994
rect 25790 30942 25842 30994
rect 26014 30942 26066 30994
rect 29486 30942 29538 30994
rect 31054 30942 31106 30994
rect 31502 30942 31554 30994
rect 31950 30942 32002 30994
rect 32174 30942 32226 30994
rect 33518 30942 33570 30994
rect 33742 30942 33794 30994
rect 34302 30942 34354 30994
rect 34526 30942 34578 30994
rect 36318 30942 36370 30994
rect 36542 30942 36594 30994
rect 37438 30942 37490 30994
rect 41134 30942 41186 30994
rect 42142 30942 42194 30994
rect 42814 30942 42866 30994
rect 45838 30942 45890 30994
rect 48974 30942 49026 30994
rect 53006 30942 53058 30994
rect 4958 30830 5010 30882
rect 13806 30830 13858 30882
rect 15934 30830 15986 30882
rect 17502 30830 17554 30882
rect 21870 30830 21922 30882
rect 26574 30830 26626 30882
rect 28702 30830 28754 30882
rect 31838 30830 31890 30882
rect 34862 30830 34914 30882
rect 36990 30830 37042 30882
rect 38222 30830 38274 30882
rect 40350 30830 40402 30882
rect 41470 30830 41522 30882
rect 42478 30830 42530 30882
rect 45614 30830 45666 30882
rect 7870 30718 7922 30770
rect 22542 30718 22594 30770
rect 45950 30718 46002 30770
rect 49310 30718 49362 30770
rect 53454 30718 53506 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 16158 30382 16210 30434
rect 25118 30382 25170 30434
rect 41918 30382 41970 30434
rect 42366 30382 42418 30434
rect 45726 30382 45778 30434
rect 4622 30270 4674 30322
rect 24894 30270 24946 30322
rect 26238 30270 26290 30322
rect 53678 30270 53730 30322
rect 54462 30270 54514 30322
rect 1822 30158 1874 30210
rect 2494 30158 2546 30210
rect 5518 30158 5570 30210
rect 5854 30158 5906 30210
rect 11006 30158 11058 30210
rect 16382 30158 16434 30210
rect 16718 30158 16770 30210
rect 18734 30158 18786 30210
rect 24558 30158 24610 30210
rect 29934 30158 29986 30210
rect 30158 30158 30210 30210
rect 30606 30158 30658 30210
rect 36318 30158 36370 30210
rect 37550 30158 37602 30210
rect 39342 30158 39394 30210
rect 39454 30158 39506 30210
rect 40910 30158 40962 30210
rect 41918 30158 41970 30210
rect 50990 30158 51042 30210
rect 53342 30158 53394 30210
rect 53566 30158 53618 30210
rect 54014 30158 54066 30210
rect 54350 30158 54402 30210
rect 55246 30158 55298 30210
rect 6190 30046 6242 30098
rect 6526 30046 6578 30098
rect 10670 30046 10722 30098
rect 16830 30046 16882 30098
rect 19294 30046 19346 30098
rect 24670 30046 24722 30098
rect 34974 30046 35026 30098
rect 42366 30046 42418 30098
rect 45390 30046 45442 30098
rect 45614 30046 45666 30098
rect 5742 29934 5794 29986
rect 7086 29934 7138 29986
rect 10782 29934 10834 29986
rect 15822 29934 15874 29986
rect 20414 29934 20466 29986
rect 24446 29934 24498 29986
rect 30270 29934 30322 29986
rect 36206 29934 36258 29986
rect 36990 29934 37042 29986
rect 40798 29934 40850 29986
rect 51102 29934 51154 29986
rect 53790 29934 53842 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 5854 29598 5906 29650
rect 8990 29598 9042 29650
rect 11566 29598 11618 29650
rect 16270 29598 16322 29650
rect 19070 29598 19122 29650
rect 19406 29598 19458 29650
rect 19854 29598 19906 29650
rect 27470 29598 27522 29650
rect 33182 29598 33234 29650
rect 37438 29598 37490 29650
rect 37886 29598 37938 29650
rect 47966 29598 48018 29650
rect 49646 29598 49698 29650
rect 51550 29598 51602 29650
rect 51774 29598 51826 29650
rect 55806 29598 55858 29650
rect 4510 29486 4562 29538
rect 5966 29486 6018 29538
rect 11678 29486 11730 29538
rect 16382 29486 16434 29538
rect 26462 29486 26514 29538
rect 30382 29486 30434 29538
rect 35982 29486 36034 29538
rect 44046 29486 44098 29538
rect 47406 29486 47458 29538
rect 50766 29486 50818 29538
rect 50990 29486 51042 29538
rect 4958 29374 5010 29426
rect 5406 29374 5458 29426
rect 8654 29374 8706 29426
rect 11342 29374 11394 29426
rect 16046 29374 16098 29426
rect 21310 29374 21362 29426
rect 27246 29374 27298 29426
rect 27358 29374 27410 29426
rect 27582 29374 27634 29426
rect 29598 29374 29650 29426
rect 36654 29374 36706 29426
rect 37774 29374 37826 29426
rect 37998 29374 38050 29426
rect 43822 29374 43874 29426
rect 46958 29374 47010 29426
rect 47182 29374 47234 29426
rect 47518 29374 47570 29426
rect 49310 29374 49362 29426
rect 49646 29374 49698 29426
rect 49982 29374 50034 29426
rect 50654 29374 50706 29426
rect 51102 29374 51154 29426
rect 52222 29374 52274 29426
rect 54798 29374 54850 29426
rect 55022 29374 55074 29426
rect 11118 29262 11170 29314
rect 22094 29262 22146 29314
rect 24222 29262 24274 29314
rect 25230 29262 25282 29314
rect 28142 29262 28194 29314
rect 32510 29262 32562 29314
rect 33854 29262 33906 29314
rect 44494 29262 44546 29314
rect 45054 29262 45106 29314
rect 46622 29262 46674 29314
rect 51662 29262 51714 29314
rect 55246 29262 55298 29314
rect 55582 29262 55634 29314
rect 25342 29150 25394 29202
rect 26574 29150 26626 29202
rect 26910 29150 26962 29202
rect 44606 29150 44658 29202
rect 50206 29150 50258 29202
rect 55918 29150 55970 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 8878 28814 8930 28866
rect 15934 28814 15986 28866
rect 26014 28814 26066 28866
rect 27246 28814 27298 28866
rect 45614 28814 45666 28866
rect 46062 28814 46114 28866
rect 50318 28814 50370 28866
rect 54798 28814 54850 28866
rect 12126 28702 12178 28754
rect 18398 28702 18450 28754
rect 22318 28702 22370 28754
rect 26574 28702 26626 28754
rect 29822 28702 29874 28754
rect 31054 28702 31106 28754
rect 39902 28702 39954 28754
rect 42030 28702 42082 28754
rect 43486 28702 43538 28754
rect 48526 28702 48578 28754
rect 50430 28702 50482 28754
rect 52782 28702 52834 28754
rect 53902 28702 53954 28754
rect 56030 28702 56082 28754
rect 58158 28702 58210 28754
rect 6862 28590 6914 28642
rect 8654 28590 8706 28642
rect 8878 28590 8930 28642
rect 9662 28590 9714 28642
rect 9886 28590 9938 28642
rect 10110 28590 10162 28642
rect 10894 28590 10946 28642
rect 11342 28590 11394 28642
rect 11566 28590 11618 28642
rect 12014 28590 12066 28642
rect 12238 28590 12290 28642
rect 12462 28590 12514 28642
rect 16158 28590 16210 28642
rect 16494 28590 16546 28642
rect 17166 28590 17218 28642
rect 17726 28590 17778 28642
rect 23102 28590 23154 28642
rect 23550 28590 23602 28642
rect 24446 28590 24498 28642
rect 26350 28590 26402 28642
rect 27358 28590 27410 28642
rect 29038 28590 29090 28642
rect 38222 28590 38274 28642
rect 39230 28590 39282 28642
rect 43822 28590 43874 28642
rect 44270 28590 44322 28642
rect 44942 28590 44994 28642
rect 45166 28590 45218 28642
rect 46398 28590 46450 28642
rect 47182 28590 47234 28642
rect 47854 28590 47906 28642
rect 50990 28590 51042 28642
rect 51326 28590 51378 28642
rect 51550 28590 51602 28642
rect 52110 28590 52162 28642
rect 52670 28590 52722 28642
rect 53790 28590 53842 28642
rect 54238 28590 54290 28642
rect 54462 28590 54514 28642
rect 54910 28590 54962 28642
rect 55358 28590 55410 28642
rect 4398 28478 4450 28530
rect 4510 28478 4562 28530
rect 7646 28478 7698 28530
rect 7982 28478 8034 28530
rect 8318 28478 8370 28530
rect 9438 28478 9490 28530
rect 10558 28478 10610 28530
rect 11118 28478 11170 28530
rect 16718 28478 16770 28530
rect 22766 28478 22818 28530
rect 23774 28478 23826 28530
rect 26686 28478 26738 28530
rect 29262 28478 29314 28530
rect 29374 28478 29426 28530
rect 45054 28478 45106 28530
rect 47406 28478 47458 28530
rect 48190 28478 48242 28530
rect 51998 28478 52050 28530
rect 4174 28366 4226 28418
rect 6526 28366 6578 28418
rect 9102 28366 9154 28418
rect 10670 28366 10722 28418
rect 11342 28366 11394 28418
rect 15598 28366 15650 28418
rect 16606 28366 16658 28418
rect 20638 28366 20690 28418
rect 23550 28366 23602 28418
rect 26462 28366 26514 28418
rect 27246 28366 27298 28418
rect 27806 28366 27858 28418
rect 30942 28366 30994 28418
rect 38558 28366 38610 28418
rect 46174 28366 46226 28418
rect 47630 28366 47682 28418
rect 48414 28366 48466 28418
rect 48638 28366 48690 28418
rect 51102 28366 51154 28418
rect 51774 28366 51826 28418
rect 54014 28366 54066 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 5070 28030 5122 28082
rect 7758 28030 7810 28082
rect 8318 28030 8370 28082
rect 11454 28030 11506 28082
rect 12126 28030 12178 28082
rect 25790 28030 25842 28082
rect 27358 28030 27410 28082
rect 31278 28030 31330 28082
rect 32174 28030 32226 28082
rect 34302 28030 34354 28082
rect 47518 28030 47570 28082
rect 54014 28030 54066 28082
rect 11230 27918 11282 27970
rect 11790 27918 11842 27970
rect 11902 27918 11954 27970
rect 23886 27918 23938 27970
rect 28590 27918 28642 27970
rect 28702 27918 28754 27970
rect 33742 27918 33794 27970
rect 34078 27918 34130 27970
rect 34414 27918 34466 27970
rect 1822 27806 1874 27858
rect 4846 27806 4898 27858
rect 5182 27806 5234 27858
rect 8430 27806 8482 27858
rect 8654 27806 8706 27858
rect 8766 27806 8818 27858
rect 11118 27806 11170 27858
rect 13918 27806 13970 27858
rect 20974 27806 21026 27858
rect 26014 27806 26066 27858
rect 28366 27806 28418 27858
rect 31166 27806 31218 27858
rect 31502 27806 31554 27858
rect 33294 27806 33346 27858
rect 33518 27806 33570 27858
rect 36430 27806 36482 27858
rect 36654 27806 36706 27858
rect 37326 27806 37378 27858
rect 38558 27806 38610 27858
rect 38782 27806 38834 27858
rect 41022 27806 41074 27858
rect 44046 27806 44098 27858
rect 44382 27806 44434 27858
rect 44718 27806 44770 27858
rect 45054 27806 45106 27858
rect 45278 27806 45330 27858
rect 45502 27806 45554 27858
rect 47742 27806 47794 27858
rect 48190 27806 48242 27858
rect 2494 27694 2546 27746
rect 4622 27694 4674 27746
rect 9662 27694 9714 27746
rect 10222 27694 10274 27746
rect 14702 27694 14754 27746
rect 16830 27694 16882 27746
rect 21310 27694 21362 27746
rect 24334 27694 24386 27746
rect 25566 27694 25618 27746
rect 25902 27694 25954 27746
rect 26798 27694 26850 27746
rect 31390 27694 31442 27746
rect 33630 27694 33682 27746
rect 41694 27694 41746 27746
rect 43822 27694 43874 27746
rect 44270 27694 44322 27746
rect 45614 27694 45666 27746
rect 47630 27694 47682 27746
rect 54126 27694 54178 27746
rect 8206 27582 8258 27634
rect 23998 27582 24050 27634
rect 24446 27582 24498 27634
rect 25342 27582 25394 27634
rect 30830 27582 30882 27634
rect 33070 27582 33122 27634
rect 36990 27582 37042 27634
rect 37550 27582 37602 27634
rect 37886 27582 37938 27634
rect 39118 27582 39170 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 16270 27246 16322 27298
rect 16606 27246 16658 27298
rect 29934 27246 29986 27298
rect 51214 27246 51266 27298
rect 3950 27134 4002 27186
rect 21646 27134 21698 27186
rect 22094 27134 22146 27186
rect 34750 27134 34802 27186
rect 37550 27134 37602 27186
rect 38334 27134 38386 27186
rect 3838 27022 3890 27074
rect 4174 27022 4226 27074
rect 4958 27022 5010 27074
rect 5630 27022 5682 27074
rect 7534 27022 7586 27074
rect 9102 27022 9154 27074
rect 16270 27022 16322 27074
rect 22766 27022 22818 27074
rect 24110 27022 24162 27074
rect 25902 27022 25954 27074
rect 26798 27022 26850 27074
rect 27134 27022 27186 27074
rect 29822 27022 29874 27074
rect 30270 27022 30322 27074
rect 31950 27022 32002 27074
rect 32958 27022 33010 27074
rect 33742 27022 33794 27074
rect 37102 27022 37154 27074
rect 45390 27022 45442 27074
rect 49758 27022 49810 27074
rect 50206 27022 50258 27074
rect 50990 27022 51042 27074
rect 51438 27022 51490 27074
rect 52110 27022 52162 27074
rect 52894 27022 52946 27074
rect 4398 26910 4450 26962
rect 4846 26910 4898 26962
rect 5742 26910 5794 26962
rect 7198 26910 7250 26962
rect 7982 26910 8034 26962
rect 8206 26910 8258 26962
rect 8542 26910 8594 26962
rect 8766 26910 8818 26962
rect 8990 26910 9042 26962
rect 22430 26910 22482 26962
rect 25678 26910 25730 26962
rect 27022 26910 27074 26962
rect 27582 26910 27634 26962
rect 30942 26910 30994 26962
rect 34862 26910 34914 26962
rect 38782 26910 38834 26962
rect 43822 26910 43874 26962
rect 47182 26910 47234 26962
rect 49870 26910 49922 26962
rect 50094 26910 50146 26962
rect 55358 26910 55410 26962
rect 4622 26798 4674 26850
rect 5966 26798 6018 26850
rect 8430 26798 8482 26850
rect 23438 26798 23490 26850
rect 29710 26798 29762 26850
rect 30270 26798 30322 26850
rect 45614 26798 45666 26850
rect 47518 26798 47570 26850
rect 50654 26798 50706 26850
rect 51326 26798 51378 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 3278 26462 3330 26514
rect 26350 26462 26402 26514
rect 26574 26462 26626 26514
rect 27246 26462 27298 26514
rect 31614 26462 31666 26514
rect 32174 26462 32226 26514
rect 36542 26462 36594 26514
rect 37102 26462 37154 26514
rect 38110 26462 38162 26514
rect 39006 26462 39058 26514
rect 53006 26462 53058 26514
rect 57598 26462 57650 26514
rect 57822 26462 57874 26514
rect 58158 26462 58210 26514
rect 3166 26350 3218 26402
rect 13022 26350 13074 26402
rect 20078 26350 20130 26402
rect 24110 26350 24162 26402
rect 30046 26350 30098 26402
rect 31726 26350 31778 26402
rect 33854 26350 33906 26402
rect 37774 26350 37826 26402
rect 41134 26350 41186 26402
rect 50654 26350 50706 26402
rect 52334 26350 52386 26402
rect 54238 26350 54290 26402
rect 54350 26350 54402 26402
rect 55470 26350 55522 26402
rect 3502 26238 3554 26290
rect 4958 26238 5010 26290
rect 9774 26238 9826 26290
rect 13806 26238 13858 26290
rect 16606 26238 16658 26290
rect 19294 26238 19346 26290
rect 22878 26238 22930 26290
rect 23102 26238 23154 26290
rect 24334 26238 24386 26290
rect 25454 26238 25506 26290
rect 26126 26238 26178 26290
rect 30718 26238 30770 26290
rect 33070 26238 33122 26290
rect 37438 26238 37490 26290
rect 46174 26238 46226 26290
rect 46622 26238 46674 26290
rect 49982 26238 50034 26290
rect 50430 26238 50482 26290
rect 52670 26238 52722 26290
rect 52894 26238 52946 26290
rect 53118 26238 53170 26290
rect 53342 26238 53394 26290
rect 54126 26238 54178 26290
rect 55022 26238 55074 26290
rect 55694 26238 55746 26290
rect 7982 26126 8034 26178
rect 10894 26126 10946 26178
rect 16158 26126 16210 26178
rect 22206 26126 22258 26178
rect 24222 26126 24274 26178
rect 26462 26126 26514 26178
rect 27918 26126 27970 26178
rect 35982 26126 36034 26178
rect 36654 26126 36706 26178
rect 38558 26126 38610 26178
rect 39678 26126 39730 26178
rect 50542 26126 50594 26178
rect 52222 26126 52274 26178
rect 55246 26126 55298 26178
rect 15822 26014 15874 26066
rect 25566 26014 25618 26066
rect 25902 26014 25954 26066
rect 31614 26014 31666 26066
rect 39566 26014 39618 26066
rect 54798 26014 54850 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 6638 25678 6690 25730
rect 49310 25678 49362 25730
rect 53342 25678 53394 25730
rect 8766 25566 8818 25618
rect 10894 25566 10946 25618
rect 22654 25566 22706 25618
rect 23438 25566 23490 25618
rect 25230 25566 25282 25618
rect 27358 25566 27410 25618
rect 31390 25566 31442 25618
rect 36430 25566 36482 25618
rect 37886 25566 37938 25618
rect 39342 25566 39394 25618
rect 41470 25566 41522 25618
rect 45726 25566 45778 25618
rect 47854 25566 47906 25618
rect 49758 25566 49810 25618
rect 51214 25566 51266 25618
rect 53454 25566 53506 25618
rect 58158 25566 58210 25618
rect 3614 25454 3666 25506
rect 4062 25454 4114 25506
rect 4286 25454 4338 25506
rect 5630 25454 5682 25506
rect 5966 25454 6018 25506
rect 6302 25454 6354 25506
rect 6526 25454 6578 25506
rect 7310 25454 7362 25506
rect 7646 25454 7698 25506
rect 7982 25454 8034 25506
rect 18062 25454 18114 25506
rect 22990 25454 23042 25506
rect 28142 25454 28194 25506
rect 28590 25454 28642 25506
rect 29374 25454 29426 25506
rect 37326 25454 37378 25506
rect 38670 25454 38722 25506
rect 43374 25454 43426 25506
rect 43710 25454 43762 25506
rect 45054 25454 45106 25506
rect 49198 25454 49250 25506
rect 49646 25454 49698 25506
rect 50766 25454 50818 25506
rect 54462 25454 54514 25506
rect 54686 25454 54738 25506
rect 54910 25454 54962 25506
rect 55358 25454 55410 25506
rect 6638 25342 6690 25394
rect 7422 25342 7474 25394
rect 13918 25342 13970 25394
rect 23326 25342 23378 25394
rect 42926 25342 42978 25394
rect 44270 25342 44322 25394
rect 50094 25342 50146 25394
rect 51774 25342 51826 25394
rect 52670 25342 52722 25394
rect 52782 25342 52834 25394
rect 56030 25342 56082 25394
rect 3838 25230 3890 25282
rect 5966 25230 6018 25282
rect 19182 25230 19234 25282
rect 51214 25230 51266 25282
rect 51326 25230 51378 25282
rect 51550 25230 51602 25282
rect 54798 25230 54850 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 30382 24894 30434 24946
rect 37438 24894 37490 24946
rect 40014 24894 40066 24946
rect 40126 24894 40178 24946
rect 45278 24894 45330 24946
rect 49198 24894 49250 24946
rect 50990 24894 51042 24946
rect 55918 24894 55970 24946
rect 2494 24782 2546 24834
rect 5742 24782 5794 24834
rect 24110 24782 24162 24834
rect 24222 24782 24274 24834
rect 30270 24782 30322 24834
rect 37998 24782 38050 24834
rect 40350 24782 40402 24834
rect 44718 24782 44770 24834
rect 49310 24782 49362 24834
rect 49422 24782 49474 24834
rect 51102 24782 51154 24834
rect 1822 24670 1874 24722
rect 5070 24670 5122 24722
rect 10782 24670 10834 24722
rect 13918 24670 13970 24722
rect 22206 24670 22258 24722
rect 35534 24670 35586 24722
rect 35982 24670 36034 24722
rect 36206 24670 36258 24722
rect 37550 24670 37602 24722
rect 38222 24670 38274 24722
rect 39342 24670 39394 24722
rect 39678 24670 39730 24722
rect 39902 24670 39954 24722
rect 41134 24670 41186 24722
rect 49086 24670 49138 24722
rect 49870 24670 49922 24722
rect 54574 24670 54626 24722
rect 56030 24670 56082 24722
rect 56702 24670 56754 24722
rect 56926 24670 56978 24722
rect 4622 24558 4674 24610
rect 7870 24558 7922 24610
rect 9774 24558 9826 24610
rect 11454 24558 11506 24610
rect 13582 24558 13634 24610
rect 14702 24558 14754 24610
rect 16830 24558 16882 24610
rect 18062 24558 18114 24610
rect 18622 24558 18674 24610
rect 36094 24558 36146 24610
rect 36766 24558 36818 24610
rect 38110 24558 38162 24610
rect 41806 24558 41858 24610
rect 43934 24558 43986 24610
rect 44942 24558 44994 24610
rect 55582 24558 55634 24610
rect 24110 24446 24162 24498
rect 54798 24446 54850 24498
rect 55134 24446 55186 24498
rect 55806 24446 55858 24498
rect 56590 24446 56642 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 8654 24110 8706 24162
rect 8990 24110 9042 24162
rect 9662 24110 9714 24162
rect 12350 24110 12402 24162
rect 15822 24110 15874 24162
rect 41806 24110 41858 24162
rect 49422 24110 49474 24162
rect 53790 24110 53842 24162
rect 15934 23998 15986 24050
rect 20750 23998 20802 24050
rect 33182 23998 33234 24050
rect 48862 23998 48914 24050
rect 49870 23998 49922 24050
rect 56030 23998 56082 24050
rect 58158 23998 58210 24050
rect 9214 23886 9266 23938
rect 9774 23886 9826 23938
rect 12350 23886 12402 23938
rect 14254 23886 14306 23938
rect 14590 23886 14642 23938
rect 17838 23886 17890 23938
rect 22318 23886 22370 23938
rect 22766 23886 22818 23938
rect 23326 23886 23378 23938
rect 23662 23886 23714 23938
rect 24222 23886 24274 23938
rect 31838 23886 31890 23938
rect 32174 23886 32226 23938
rect 35982 23886 36034 23938
rect 37438 23886 37490 23938
rect 40798 23886 40850 23938
rect 41246 23886 41298 23938
rect 41470 23886 41522 23938
rect 45278 23886 45330 23938
rect 45950 23886 46002 23938
rect 46398 23886 46450 23938
rect 49086 23886 49138 23938
rect 55358 23886 55410 23938
rect 12686 23774 12738 23826
rect 14142 23774 14194 23826
rect 18622 23774 18674 23826
rect 22094 23774 22146 23826
rect 22206 23774 22258 23826
rect 23886 23774 23938 23826
rect 31502 23774 31554 23826
rect 35310 23774 35362 23826
rect 36878 23774 36930 23826
rect 38558 23774 38610 23826
rect 41134 23774 41186 23826
rect 41918 23774 41970 23826
rect 45054 23774 45106 23826
rect 45726 23774 45778 23826
rect 46734 23774 46786 23826
rect 49758 23774 49810 23826
rect 49982 23774 50034 23826
rect 53902 23774 53954 23826
rect 9662 23662 9714 23714
rect 10222 23662 10274 23714
rect 14030 23662 14082 23714
rect 15038 23662 15090 23714
rect 16046 23662 16098 23714
rect 16718 23662 16770 23714
rect 21646 23662 21698 23714
rect 23998 23662 24050 23714
rect 31950 23662 32002 23714
rect 32510 23662 32562 23714
rect 36990 23662 37042 23714
rect 37214 23662 37266 23714
rect 38446 23662 38498 23714
rect 41022 23662 41074 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 9662 23326 9714 23378
rect 17390 23326 17442 23378
rect 21982 23326 22034 23378
rect 33294 23326 33346 23378
rect 47406 23326 47458 23378
rect 49086 23326 49138 23378
rect 49870 23326 49922 23378
rect 53006 23326 53058 23378
rect 19294 23214 19346 23266
rect 21646 23214 21698 23266
rect 35310 23214 35362 23266
rect 47630 23214 47682 23266
rect 49982 23214 50034 23266
rect 55694 23214 55746 23266
rect 55918 23214 55970 23266
rect 1822 23102 1874 23154
rect 14030 23102 14082 23154
rect 17614 23102 17666 23154
rect 17950 23102 18002 23154
rect 19406 23102 19458 23154
rect 19742 23102 19794 23154
rect 22878 23102 22930 23154
rect 23214 23102 23266 23154
rect 23886 23102 23938 23154
rect 25342 23102 25394 23154
rect 26574 23102 26626 23154
rect 27022 23102 27074 23154
rect 27246 23102 27298 23154
rect 28254 23102 28306 23154
rect 28814 23102 28866 23154
rect 32062 23102 32114 23154
rect 33070 23102 33122 23154
rect 33742 23102 33794 23154
rect 39790 23102 39842 23154
rect 47966 23102 48018 23154
rect 48302 23102 48354 23154
rect 48862 23102 48914 23154
rect 48974 23102 49026 23154
rect 49198 23102 49250 23154
rect 49422 23102 49474 23154
rect 51774 23102 51826 23154
rect 52334 23102 52386 23154
rect 55022 23102 55074 23154
rect 55246 23102 55298 23154
rect 2494 22990 2546 23042
rect 4622 22990 4674 23042
rect 9550 22990 9602 23042
rect 17502 22990 17554 23042
rect 20302 22990 20354 23042
rect 24670 22990 24722 23042
rect 26350 22990 26402 23042
rect 26798 22990 26850 23042
rect 27918 22990 27970 23042
rect 29150 22990 29202 23042
rect 31278 22990 31330 23042
rect 32510 22990 32562 23042
rect 33182 22990 33234 23042
rect 40238 22990 40290 23042
rect 41918 22990 41970 23042
rect 48078 22990 48130 23042
rect 52446 22990 52498 23042
rect 52782 22990 52834 23042
rect 13470 22878 13522 22930
rect 13806 22878 13858 22930
rect 19630 22878 19682 22930
rect 42030 22878 42082 22930
rect 49758 22878 49810 22930
rect 53118 22878 53170 22930
rect 54686 22878 54738 22930
rect 55582 22878 55634 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 4734 22542 4786 22594
rect 32062 22542 32114 22594
rect 35982 22542 36034 22594
rect 36430 22542 36482 22594
rect 51998 22542 52050 22594
rect 52782 22542 52834 22594
rect 3390 22430 3442 22482
rect 3950 22430 4002 22482
rect 9550 22430 9602 22482
rect 12910 22430 12962 22482
rect 18174 22430 18226 22482
rect 25678 22430 25730 22482
rect 27806 22430 27858 22482
rect 35534 22430 35586 22482
rect 37998 22430 38050 22482
rect 40126 22430 40178 22482
rect 42142 22430 42194 22482
rect 44270 22430 44322 22482
rect 45390 22430 45442 22482
rect 52110 22430 52162 22482
rect 58158 22430 58210 22482
rect 4174 22318 4226 22370
rect 5630 22318 5682 22370
rect 5854 22318 5906 22370
rect 6750 22318 6802 22370
rect 10110 22318 10162 22370
rect 15262 22318 15314 22370
rect 23102 22318 23154 22370
rect 23998 22318 24050 22370
rect 24782 22318 24834 22370
rect 28590 22318 28642 22370
rect 31390 22318 31442 22370
rect 31614 22318 31666 22370
rect 32734 22318 32786 22370
rect 35758 22318 35810 22370
rect 37214 22318 37266 22370
rect 41358 22318 41410 22370
rect 50430 22318 50482 22370
rect 52894 22318 52946 22370
rect 55246 22318 55298 22370
rect 5070 22206 5122 22258
rect 7422 22206 7474 22258
rect 10782 22206 10834 22258
rect 16046 22206 16098 22258
rect 23774 22206 23826 22258
rect 25342 22206 25394 22258
rect 31502 22206 31554 22258
rect 52782 22206 52834 22258
rect 56030 22206 56082 22258
rect 3614 22094 3666 22146
rect 4846 22094 4898 22146
rect 6190 22094 6242 22146
rect 22654 22094 22706 22146
rect 23438 22094 23490 22146
rect 33182 22094 33234 22146
rect 50878 22094 50930 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 8878 21758 8930 21810
rect 12798 21758 12850 21810
rect 13470 21758 13522 21810
rect 16158 21758 16210 21810
rect 19182 21758 19234 21810
rect 23550 21758 23602 21810
rect 24558 21758 24610 21810
rect 27246 21758 27298 21810
rect 27358 21758 27410 21810
rect 28254 21758 28306 21810
rect 36766 21758 36818 21810
rect 38110 21758 38162 21810
rect 38782 21758 38834 21810
rect 39006 21758 39058 21810
rect 39118 21758 39170 21810
rect 41246 21758 41298 21810
rect 48974 21758 49026 21810
rect 49534 21758 49586 21810
rect 6414 21646 6466 21698
rect 12686 21646 12738 21698
rect 16606 21646 16658 21698
rect 16830 21646 16882 21698
rect 37438 21646 37490 21698
rect 39342 21646 39394 21698
rect 41582 21646 41634 21698
rect 43374 21646 43426 21698
rect 46062 21646 46114 21698
rect 48750 21646 48802 21698
rect 53118 21646 53170 21698
rect 55806 21646 55858 21698
rect 57822 21646 57874 21698
rect 8430 21534 8482 21586
rect 13246 21534 13298 21586
rect 13918 21534 13970 21586
rect 14478 21534 14530 21586
rect 14702 21534 14754 21586
rect 15822 21534 15874 21586
rect 17390 21534 17442 21586
rect 17726 21534 17778 21586
rect 17950 21534 18002 21586
rect 18846 21534 18898 21586
rect 19182 21534 19234 21586
rect 19518 21534 19570 21586
rect 22430 21534 22482 21586
rect 22654 21534 22706 21586
rect 23774 21534 23826 21586
rect 24110 21534 24162 21586
rect 27134 21534 27186 21586
rect 27806 21534 27858 21586
rect 33070 21534 33122 21586
rect 36318 21534 36370 21586
rect 36542 21534 36594 21586
rect 36990 21534 37042 21586
rect 38894 21534 38946 21586
rect 40910 21534 40962 21586
rect 41134 21534 41186 21586
rect 41358 21534 41410 21586
rect 42478 21534 42530 21586
rect 45390 21534 45442 21586
rect 53902 21534 53954 21586
rect 55358 21534 55410 21586
rect 55470 21534 55522 21586
rect 58158 21534 58210 21586
rect 13358 21422 13410 21474
rect 16494 21422 16546 21474
rect 23214 21422 23266 21474
rect 23662 21422 23714 21474
rect 26798 21422 26850 21474
rect 27806 21422 27858 21474
rect 32510 21422 32562 21474
rect 33854 21422 33906 21474
rect 35982 21422 36034 21474
rect 36654 21422 36706 21474
rect 37326 21422 37378 21474
rect 39790 21422 39842 21474
rect 12910 21310 12962 21362
rect 14142 21310 14194 21362
rect 42926 21422 42978 21474
rect 48190 21422 48242 21474
rect 49086 21422 49138 21474
rect 49422 21422 49474 21474
rect 50990 21422 51042 21474
rect 55694 21422 55746 21474
rect 57598 21422 57650 21474
rect 28254 21310 28306 21362
rect 37662 21310 37714 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 22654 20974 22706 21026
rect 23214 20974 23266 21026
rect 23438 20974 23490 21026
rect 34526 20974 34578 21026
rect 4622 20862 4674 20914
rect 5742 20862 5794 20914
rect 17838 20862 17890 20914
rect 19966 20862 20018 20914
rect 22990 20862 23042 20914
rect 26798 20862 26850 20914
rect 27246 20862 27298 20914
rect 32062 20862 32114 20914
rect 34638 20862 34690 20914
rect 39790 20862 39842 20914
rect 1822 20750 1874 20802
rect 5854 20750 5906 20802
rect 6302 20750 6354 20802
rect 13470 20750 13522 20802
rect 13582 20750 13634 20802
rect 20750 20750 20802 20802
rect 24334 20750 24386 20802
rect 24782 20750 24834 20802
rect 29150 20750 29202 20802
rect 37326 20750 37378 20802
rect 37662 20750 37714 20802
rect 39230 20750 39282 20802
rect 52894 20750 52946 20802
rect 2494 20638 2546 20690
rect 7310 20638 7362 20690
rect 7646 20638 7698 20690
rect 7982 20638 8034 20690
rect 13918 20638 13970 20690
rect 22430 20638 22482 20690
rect 23886 20638 23938 20690
rect 24110 20638 24162 20690
rect 29934 20638 29986 20690
rect 36990 20638 37042 20690
rect 55358 20638 55410 20690
rect 5630 20526 5682 20578
rect 6974 20526 7026 20578
rect 13694 20526 13746 20578
rect 22542 20526 22594 20578
rect 24446 20526 24498 20578
rect 24558 20526 24610 20578
rect 27134 20526 27186 20578
rect 35982 20526 36034 20578
rect 37998 20526 38050 20578
rect 39342 20526 39394 20578
rect 41918 20526 41970 20578
rect 42254 20526 42306 20578
rect 42702 20526 42754 20578
rect 52110 20526 52162 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 4062 20190 4114 20242
rect 19518 20190 19570 20242
rect 3278 20078 3330 20130
rect 3838 20078 3890 20130
rect 4958 20078 5010 20130
rect 6302 20078 6354 20130
rect 6638 20078 6690 20130
rect 8430 20078 8482 20130
rect 13806 20078 13858 20130
rect 14030 20078 14082 20130
rect 17614 20078 17666 20130
rect 19406 20078 19458 20130
rect 20526 20078 20578 20130
rect 30494 20078 30546 20130
rect 41582 20078 41634 20130
rect 41918 20078 41970 20130
rect 42366 20078 42418 20130
rect 42814 20078 42866 20130
rect 49086 20078 49138 20130
rect 49758 20078 49810 20130
rect 54798 20078 54850 20130
rect 56142 20078 56194 20130
rect 4510 19966 4562 20018
rect 9662 19966 9714 20018
rect 12910 19966 12962 20018
rect 13134 19966 13186 20018
rect 13470 19966 13522 20018
rect 19630 19966 19682 20018
rect 20078 19966 20130 20018
rect 23550 19966 23602 20018
rect 23774 19966 23826 20018
rect 25902 19966 25954 20018
rect 26462 19966 26514 20018
rect 26910 19966 26962 20018
rect 27358 19966 27410 20018
rect 27694 19966 27746 20018
rect 29822 19966 29874 20018
rect 30830 19966 30882 20018
rect 31502 19966 31554 20018
rect 31950 19966 32002 20018
rect 44606 19966 44658 20018
rect 49422 19966 49474 20018
rect 49534 19966 49586 20018
rect 49870 19966 49922 20018
rect 54462 19966 54514 20018
rect 54574 19966 54626 20018
rect 55022 19966 55074 20018
rect 3166 19854 3218 19906
rect 3950 19854 4002 19906
rect 8990 19854 9042 19906
rect 10334 19854 10386 19906
rect 12462 19854 12514 19906
rect 13918 19854 13970 19906
rect 17502 19854 17554 19906
rect 23214 19854 23266 19906
rect 28254 19854 28306 19906
rect 29598 19854 29650 19906
rect 30158 19854 30210 19906
rect 32286 19854 32338 19906
rect 33182 19854 33234 19906
rect 45390 19854 45442 19906
rect 47518 19854 47570 19906
rect 49646 19854 49698 19906
rect 50318 19854 50370 19906
rect 54686 19854 54738 19906
rect 55470 19854 55522 19906
rect 3502 19742 3554 19794
rect 8766 19742 8818 19794
rect 17390 19742 17442 19794
rect 23998 19742 24050 19794
rect 50430 19742 50482 19794
rect 55582 19742 55634 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 14926 19294 14978 19346
rect 17054 19294 17106 19346
rect 40686 19294 40738 19346
rect 42142 19294 42194 19346
rect 42590 19294 42642 19346
rect 46958 19294 47010 19346
rect 48638 19294 48690 19346
rect 50766 19294 50818 19346
rect 52782 19294 52834 19346
rect 53790 19294 53842 19346
rect 54798 19294 54850 19346
rect 56030 19294 56082 19346
rect 58158 19294 58210 19346
rect 13470 19182 13522 19234
rect 14142 19182 14194 19234
rect 17726 19182 17778 19234
rect 27358 19182 27410 19234
rect 27694 19182 27746 19234
rect 28254 19182 28306 19234
rect 43038 19182 43090 19234
rect 43262 19182 43314 19234
rect 44942 19182 44994 19234
rect 45502 19182 45554 19234
rect 46622 19182 46674 19234
rect 51438 19182 51490 19234
rect 52110 19182 52162 19234
rect 52894 19182 52946 19234
rect 53230 19182 53282 19234
rect 54686 19182 54738 19234
rect 55358 19182 55410 19234
rect 6638 19070 6690 19122
rect 22542 19070 22594 19122
rect 31614 19070 31666 19122
rect 31950 19070 32002 19122
rect 32174 19070 32226 19122
rect 34750 19070 34802 19122
rect 37998 19070 38050 19122
rect 43598 19070 43650 19122
rect 44830 19070 44882 19122
rect 48302 19070 48354 19122
rect 52782 19070 52834 19122
rect 53118 19070 53170 19122
rect 54238 19070 54290 19122
rect 54462 19070 54514 19122
rect 6414 18958 6466 19010
rect 6526 18958 6578 19010
rect 9214 18958 9266 19010
rect 13582 18958 13634 19010
rect 13694 18958 13746 19010
rect 21758 18958 21810 19010
rect 31726 18958 31778 19010
rect 32622 18958 32674 19010
rect 34638 18958 34690 19010
rect 38222 18958 38274 19010
rect 38334 18958 38386 19010
rect 38446 18958 38498 19010
rect 38558 18958 38610 19010
rect 41246 18958 41298 19010
rect 41582 18958 41634 19010
rect 43486 18958 43538 19010
rect 43934 18958 43986 19010
rect 44270 18958 44322 19010
rect 47966 18958 48018 19010
rect 51998 18958 52050 19010
rect 54798 18958 54850 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 3502 18622 3554 18674
rect 16494 18622 16546 18674
rect 19070 18622 19122 18674
rect 26350 18622 26402 18674
rect 26574 18622 26626 18674
rect 45166 18622 45218 18674
rect 45390 18622 45442 18674
rect 49086 18622 49138 18674
rect 6638 18510 6690 18562
rect 14366 18510 14418 18562
rect 16718 18510 16770 18562
rect 18622 18510 18674 18562
rect 18958 18510 19010 18562
rect 32174 18510 32226 18562
rect 33630 18510 33682 18562
rect 38558 18510 38610 18562
rect 42702 18510 42754 18562
rect 44158 18510 44210 18562
rect 51886 18510 51938 18562
rect 54462 18510 54514 18562
rect 55358 18510 55410 18562
rect 2830 18398 2882 18450
rect 3726 18398 3778 18450
rect 4174 18398 4226 18450
rect 7422 18398 7474 18450
rect 10222 18398 10274 18450
rect 13470 18398 13522 18450
rect 14030 18398 14082 18450
rect 14702 18398 14754 18450
rect 16046 18398 16098 18450
rect 16606 18398 16658 18450
rect 17390 18398 17442 18450
rect 17614 18398 17666 18450
rect 17950 18398 18002 18450
rect 18398 18398 18450 18450
rect 19294 18398 19346 18450
rect 22990 18398 23042 18450
rect 23214 18398 23266 18450
rect 23886 18398 23938 18450
rect 24110 18398 24162 18450
rect 24222 18398 24274 18450
rect 24446 18398 24498 18450
rect 25230 18398 25282 18450
rect 32062 18398 32114 18450
rect 32286 18398 32338 18450
rect 33518 18398 33570 18450
rect 33854 18398 33906 18450
rect 34302 18398 34354 18450
rect 37550 18398 37602 18450
rect 37774 18398 37826 18450
rect 37998 18398 38050 18450
rect 38110 18398 38162 18450
rect 40462 18398 40514 18450
rect 41246 18398 41298 18450
rect 41694 18398 41746 18450
rect 42030 18398 42082 18450
rect 42254 18398 42306 18450
rect 42366 18398 42418 18450
rect 43038 18398 43090 18450
rect 43934 18398 43986 18450
rect 44718 18398 44770 18450
rect 45054 18398 45106 18450
rect 48750 18398 48802 18450
rect 51214 18398 51266 18450
rect 56030 18398 56082 18450
rect 3166 18286 3218 18338
rect 3614 18286 3666 18338
rect 4510 18286 4562 18338
rect 7758 18286 7810 18338
rect 11006 18286 11058 18338
rect 13134 18286 13186 18338
rect 14478 18286 14530 18338
rect 22318 18286 22370 18338
rect 22766 18286 22818 18338
rect 25342 18286 25394 18338
rect 27022 18286 27074 18338
rect 33742 18286 33794 18338
rect 35086 18286 35138 18338
rect 37214 18286 37266 18338
rect 37886 18286 37938 18338
rect 39118 18286 39170 18338
rect 45726 18286 45778 18338
rect 48190 18286 48242 18338
rect 54014 18286 54066 18338
rect 2830 18174 2882 18226
rect 7982 18174 8034 18226
rect 8318 18174 8370 18226
rect 13694 18174 13746 18226
rect 22654 18174 22706 18226
rect 23438 18174 23490 18226
rect 31614 18174 31666 18226
rect 33182 18174 33234 18226
rect 38670 18174 38722 18226
rect 54350 18174 54402 18226
rect 55470 18174 55522 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 35422 17838 35474 17890
rect 36094 17838 36146 17890
rect 2494 17726 2546 17778
rect 4622 17726 4674 17778
rect 6750 17726 6802 17778
rect 19294 17726 19346 17778
rect 20414 17726 20466 17778
rect 23438 17726 23490 17778
rect 25566 17726 25618 17778
rect 28590 17726 28642 17778
rect 32174 17726 32226 17778
rect 32734 17726 32786 17778
rect 35534 17726 35586 17778
rect 36206 17726 36258 17778
rect 37326 17726 37378 17778
rect 39454 17726 39506 17778
rect 41918 17726 41970 17778
rect 42478 17726 42530 17778
rect 46958 17726 47010 17778
rect 1822 17614 1874 17666
rect 6302 17614 6354 17666
rect 6638 17614 6690 17666
rect 6862 17614 6914 17666
rect 7758 17614 7810 17666
rect 14366 17614 14418 17666
rect 17838 17614 17890 17666
rect 18398 17614 18450 17666
rect 19182 17614 19234 17666
rect 22654 17614 22706 17666
rect 29262 17614 29314 17666
rect 33630 17614 33682 17666
rect 34190 17614 34242 17666
rect 40238 17614 40290 17666
rect 40910 17614 40962 17666
rect 41470 17614 41522 17666
rect 52894 17614 52946 17666
rect 7422 17502 7474 17554
rect 14142 17502 14194 17554
rect 15038 17502 15090 17554
rect 15374 17502 15426 17554
rect 18062 17502 18114 17554
rect 18286 17502 18338 17554
rect 19742 17502 19794 17554
rect 20078 17502 20130 17554
rect 20302 17502 20354 17554
rect 27582 17502 27634 17554
rect 27806 17502 27858 17554
rect 27918 17502 27970 17554
rect 30046 17502 30098 17554
rect 41134 17502 41186 17554
rect 55358 17502 55410 17554
rect 17390 17390 17442 17442
rect 21422 17390 21474 17442
rect 28142 17390 28194 17442
rect 33742 17390 33794 17442
rect 33966 17390 34018 17442
rect 34302 17390 34354 17442
rect 34526 17390 34578 17442
rect 52110 17390 52162 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 3278 17054 3330 17106
rect 15710 17054 15762 17106
rect 23886 17054 23938 17106
rect 25342 17054 25394 17106
rect 41022 17054 41074 17106
rect 44270 17054 44322 17106
rect 44494 17054 44546 17106
rect 45278 17054 45330 17106
rect 46510 17054 46562 17106
rect 51438 17054 51490 17106
rect 51774 17054 51826 17106
rect 52782 17054 52834 17106
rect 10222 16942 10274 16994
rect 16046 16942 16098 16994
rect 21534 16942 21586 16994
rect 22990 16942 23042 16994
rect 23326 16942 23378 16994
rect 24670 16942 24722 16994
rect 27918 16942 27970 16994
rect 30718 16942 30770 16994
rect 42254 16942 42306 16994
rect 46734 16942 46786 16994
rect 47630 16942 47682 16994
rect 49646 16942 49698 16994
rect 3838 16830 3890 16882
rect 13806 16830 13858 16882
rect 15262 16830 15314 16882
rect 22318 16830 22370 16882
rect 24110 16830 24162 16882
rect 28702 16830 28754 16882
rect 31054 16830 31106 16882
rect 31278 16830 31330 16882
rect 41470 16830 41522 16882
rect 41918 16830 41970 16882
rect 42478 16830 42530 16882
rect 44942 16830 44994 16882
rect 46174 16830 46226 16882
rect 47518 16830 47570 16882
rect 47854 16830 47906 16882
rect 49310 16830 49362 16882
rect 52334 16830 52386 16882
rect 54014 16830 54066 16882
rect 3614 16718 3666 16770
rect 19406 16718 19458 16770
rect 25790 16718 25842 16770
rect 30830 16718 30882 16770
rect 44382 16718 44434 16770
rect 47294 16718 47346 16770
rect 46846 16606 46898 16658
rect 48302 16606 48354 16658
rect 53902 16606 53954 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 30830 16270 30882 16322
rect 8878 16158 8930 16210
rect 14702 16158 14754 16210
rect 15486 16158 15538 16210
rect 25566 16158 25618 16210
rect 27022 16158 27074 16210
rect 27358 16158 27410 16210
rect 28142 16158 28194 16210
rect 31726 16158 31778 16210
rect 35982 16158 36034 16210
rect 42030 16158 42082 16210
rect 47742 16158 47794 16210
rect 48190 16158 48242 16210
rect 48862 16158 48914 16210
rect 50990 16158 51042 16210
rect 56030 16158 56082 16210
rect 58158 16158 58210 16210
rect 6750 16046 6802 16098
rect 7198 16046 7250 16098
rect 7758 16046 7810 16098
rect 7982 16046 8034 16098
rect 8094 16046 8146 16098
rect 11678 16046 11730 16098
rect 13806 16046 13858 16098
rect 14254 16046 14306 16098
rect 15038 16046 15090 16098
rect 17838 16046 17890 16098
rect 23886 16046 23938 16098
rect 24334 16046 24386 16098
rect 25006 16046 25058 16098
rect 27806 16046 27858 16098
rect 31054 16046 31106 16098
rect 31278 16046 31330 16098
rect 31950 16046 32002 16098
rect 38334 16046 38386 16098
rect 43934 16046 43986 16098
rect 44270 16046 44322 16098
rect 44942 16046 44994 16098
rect 51662 16046 51714 16098
rect 53006 16046 53058 16098
rect 55246 16046 55298 16098
rect 7422 15934 7474 15986
rect 11006 15934 11058 15986
rect 30718 15934 30770 15986
rect 31614 15934 31666 15986
rect 36430 15934 36482 15986
rect 37886 15934 37938 15986
rect 44046 15934 44098 15986
rect 45614 15934 45666 15986
rect 53230 15934 53282 15986
rect 53342 15934 53394 15986
rect 53790 15934 53842 15986
rect 54574 15934 54626 15986
rect 6974 15822 7026 15874
rect 8542 15822 8594 15874
rect 13470 15822 13522 15874
rect 18174 15822 18226 15874
rect 38110 15822 38162 15874
rect 38222 15822 38274 15874
rect 38446 15822 38498 15874
rect 43486 15822 43538 15874
rect 48078 15822 48130 15874
rect 54910 15822 54962 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 14478 15486 14530 15538
rect 29262 15486 29314 15538
rect 46510 15486 46562 15538
rect 49310 15486 49362 15538
rect 53006 15486 53058 15538
rect 53678 15486 53730 15538
rect 5518 15374 5570 15426
rect 10110 15374 10162 15426
rect 10558 15374 10610 15426
rect 14814 15374 14866 15426
rect 18174 15374 18226 15426
rect 23662 15374 23714 15426
rect 28926 15374 28978 15426
rect 29038 15374 29090 15426
rect 30382 15374 30434 15426
rect 33630 15374 33682 15426
rect 33742 15374 33794 15426
rect 34414 15374 34466 15426
rect 38446 15374 38498 15426
rect 52110 15374 52162 15426
rect 53454 15374 53506 15426
rect 57822 15374 57874 15426
rect 3838 15262 3890 15314
rect 4846 15262 4898 15314
rect 7982 15262 8034 15314
rect 8318 15262 8370 15314
rect 8542 15262 8594 15314
rect 9662 15262 9714 15314
rect 9998 15262 10050 15314
rect 13246 15262 13298 15314
rect 13582 15262 13634 15314
rect 13806 15262 13858 15314
rect 17502 15262 17554 15314
rect 23774 15262 23826 15314
rect 29598 15262 29650 15314
rect 34078 15262 34130 15314
rect 35982 15262 36034 15314
rect 36430 15262 36482 15314
rect 36654 15262 36706 15314
rect 37662 15262 37714 15314
rect 46174 15262 46226 15314
rect 46734 15262 46786 15314
rect 47294 15262 47346 15314
rect 47742 15262 47794 15314
rect 48750 15262 48802 15314
rect 51886 15262 51938 15314
rect 52670 15262 52722 15314
rect 53342 15262 53394 15314
rect 57598 15262 57650 15314
rect 58158 15262 58210 15314
rect 4062 15150 4114 15202
rect 7646 15150 7698 15202
rect 8206 15150 8258 15202
rect 9774 15150 9826 15202
rect 13358 15150 13410 15202
rect 20302 15150 20354 15202
rect 28590 15150 28642 15202
rect 32510 15150 32562 15202
rect 34302 15150 34354 15202
rect 41134 15150 41186 15202
rect 48190 15150 48242 15202
rect 48974 15150 49026 15202
rect 49758 15150 49810 15202
rect 52446 15150 52498 15202
rect 3502 15038 3554 15090
rect 23662 15038 23714 15090
rect 33630 15038 33682 15090
rect 35310 15038 35362 15090
rect 38558 15038 38610 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 30942 14702 30994 14754
rect 31278 14702 31330 14754
rect 4622 14590 4674 14642
rect 7646 14590 7698 14642
rect 13918 14590 13970 14642
rect 54350 14646 54402 14698
rect 17054 14590 17106 14642
rect 22990 14590 23042 14642
rect 31502 14590 31554 14642
rect 36990 14590 37042 14642
rect 39118 14590 39170 14642
rect 43822 14590 43874 14642
rect 45054 14590 45106 14642
rect 53678 14590 53730 14642
rect 56030 14590 56082 14642
rect 58158 14590 58210 14642
rect 1822 14478 1874 14530
rect 7534 14478 7586 14530
rect 7758 14478 7810 14530
rect 8206 14478 8258 14530
rect 13470 14478 13522 14530
rect 14030 14478 14082 14530
rect 20526 14478 20578 14530
rect 20750 14478 20802 14530
rect 22878 14478 22930 14530
rect 24110 14478 24162 14530
rect 25006 14478 25058 14530
rect 35534 14478 35586 14530
rect 35982 14478 36034 14530
rect 36318 14478 36370 14530
rect 39902 14478 39954 14530
rect 40910 14478 40962 14530
rect 48638 14478 48690 14530
rect 50542 14478 50594 14530
rect 53342 14478 53394 14530
rect 54574 14478 54626 14530
rect 55358 14478 55410 14530
rect 2494 14366 2546 14418
rect 16158 14366 16210 14418
rect 17390 14366 17442 14418
rect 17502 14366 17554 14418
rect 17726 14366 17778 14418
rect 20190 14366 20242 14418
rect 23326 14366 23378 14418
rect 24334 14366 24386 14418
rect 24670 14366 24722 14418
rect 35198 14366 35250 14418
rect 35758 14366 35810 14418
rect 40462 14366 40514 14418
rect 41694 14366 41746 14418
rect 54014 14366 54066 14418
rect 13806 14254 13858 14306
rect 16270 14254 16322 14306
rect 16494 14254 16546 14306
rect 20526 14254 20578 14306
rect 24782 14254 24834 14306
rect 34974 14254 35026 14306
rect 35310 14254 35362 14306
rect 36094 14254 36146 14306
rect 36206 14254 36258 14306
rect 40574 14254 40626 14306
rect 54910 14254 54962 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 3054 13918 3106 13970
rect 3614 13918 3666 13970
rect 3838 13918 3890 13970
rect 4622 13918 4674 13970
rect 15486 13918 15538 13970
rect 15598 13918 15650 13970
rect 16382 13918 16434 13970
rect 16718 13918 16770 13970
rect 24670 13918 24722 13970
rect 25342 13918 25394 13970
rect 35758 13918 35810 13970
rect 41582 13918 41634 13970
rect 41694 13918 41746 13970
rect 51998 13918 52050 13970
rect 11118 13806 11170 13858
rect 15934 13806 15986 13858
rect 24110 13806 24162 13858
rect 25230 13806 25282 13858
rect 25454 13806 25506 13858
rect 29598 13806 29650 13858
rect 33854 13806 33906 13858
rect 34302 13806 34354 13858
rect 37774 13806 37826 13858
rect 41918 13806 41970 13858
rect 47518 13806 47570 13858
rect 50654 13806 50706 13858
rect 52894 13806 52946 13858
rect 55694 13806 55746 13858
rect 56030 13806 56082 13858
rect 4174 13694 4226 13746
rect 10334 13694 10386 13746
rect 13582 13694 13634 13746
rect 13694 13694 13746 13746
rect 15710 13694 15762 13746
rect 18174 13694 18226 13746
rect 23438 13694 23490 13746
rect 24334 13694 24386 13746
rect 26910 13694 26962 13746
rect 28478 13694 28530 13746
rect 34862 13694 34914 13746
rect 35982 13694 36034 13746
rect 37998 13694 38050 13746
rect 41358 13694 41410 13746
rect 41470 13694 41522 13746
rect 46286 13694 46338 13746
rect 46510 13694 46562 13746
rect 46734 13694 46786 13746
rect 48078 13694 48130 13746
rect 49198 13694 49250 13746
rect 49310 13694 49362 13746
rect 49534 13694 49586 13746
rect 49758 13694 49810 13746
rect 50542 13694 50594 13746
rect 52446 13694 52498 13746
rect 52670 13694 52722 13746
rect 2942 13582 2994 13634
rect 3278 13582 3330 13634
rect 3726 13582 3778 13634
rect 13246 13582 13298 13634
rect 19182 13582 19234 13634
rect 33518 13582 33570 13634
rect 42590 13582 42642 13634
rect 45950 13582 46002 13634
rect 46398 13582 46450 13634
rect 47182 13582 47234 13634
rect 49422 13582 49474 13634
rect 50206 13582 50258 13634
rect 51886 13582 51938 13634
rect 54014 13582 54066 13634
rect 42702 13470 42754 13522
rect 48190 13470 48242 13522
rect 50094 13470 50146 13522
rect 53006 13470 53058 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 21310 13134 21362 13186
rect 30830 13134 30882 13186
rect 37886 13134 37938 13186
rect 9214 13022 9266 13074
rect 18174 13022 18226 13074
rect 21422 13022 21474 13074
rect 23662 13022 23714 13074
rect 25790 13022 25842 13074
rect 29822 13022 29874 13074
rect 35870 13022 35922 13074
rect 37102 13022 37154 13074
rect 37662 13022 37714 13074
rect 38670 13022 38722 13074
rect 39118 13022 39170 13074
rect 39902 13022 39954 13074
rect 41358 13022 41410 13074
rect 56030 13022 56082 13074
rect 58158 13022 58210 13074
rect 6302 12910 6354 12962
rect 9998 12910 10050 12962
rect 10334 12910 10386 12962
rect 20078 12910 20130 12962
rect 22654 12910 22706 12962
rect 22990 12910 23042 12962
rect 26574 12910 26626 12962
rect 27134 12910 27186 12962
rect 27582 12910 27634 12962
rect 28030 12910 28082 12962
rect 28254 12910 28306 12962
rect 28366 12910 28418 12962
rect 28590 12910 28642 12962
rect 30158 12910 30210 12962
rect 30718 12910 30770 12962
rect 31278 12910 31330 12962
rect 31614 12910 31666 12962
rect 31838 12910 31890 12962
rect 33854 12910 33906 12962
rect 34638 12910 34690 12962
rect 35086 12910 35138 12962
rect 35758 12910 35810 12962
rect 43486 12910 43538 12962
rect 44270 12910 44322 12962
rect 45278 12910 45330 12962
rect 50990 12910 51042 12962
rect 52670 12910 52722 12962
rect 53006 12910 53058 12962
rect 53230 12910 53282 12962
rect 55246 12910 55298 12962
rect 4510 12798 4562 12850
rect 7086 12798 7138 12850
rect 10110 12798 10162 12850
rect 30382 12798 30434 12850
rect 30830 12798 30882 12850
rect 33966 12798 34018 12850
rect 36094 12798 36146 12850
rect 47294 12798 47346 12850
rect 52894 12798 52946 12850
rect 54014 12798 54066 12850
rect 4286 12686 4338 12738
rect 4398 12686 4450 12738
rect 9550 12686 9602 12738
rect 21982 12686 22034 12738
rect 22766 12686 22818 12738
rect 27358 12686 27410 12738
rect 31726 12686 31778 12738
rect 36990 12686 37042 12738
rect 38222 12686 38274 12738
rect 40574 12686 40626 12738
rect 45054 12686 45106 12738
rect 50878 12686 50930 12738
rect 53678 12686 53730 12738
rect 53902 12686 53954 12738
rect 54462 12686 54514 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 9550 12350 9602 12402
rect 17502 12350 17554 12402
rect 41022 12350 41074 12402
rect 41358 12350 41410 12402
rect 42142 12350 42194 12402
rect 42254 12350 42306 12402
rect 42366 12350 42418 12402
rect 42478 12350 42530 12402
rect 43038 12350 43090 12402
rect 45278 12350 45330 12402
rect 45502 12350 45554 12402
rect 48078 12350 48130 12402
rect 48974 12350 49026 12402
rect 49086 12350 49138 12402
rect 49198 12350 49250 12402
rect 49758 12350 49810 12402
rect 49982 12350 50034 12402
rect 50766 12350 50818 12402
rect 50990 12350 51042 12402
rect 55022 12350 55074 12402
rect 6302 12238 6354 12290
rect 12574 12238 12626 12290
rect 14254 12238 14306 12290
rect 15262 12238 15314 12290
rect 19966 12238 20018 12290
rect 27582 12238 27634 12290
rect 41918 12238 41970 12290
rect 45166 12238 45218 12290
rect 45838 12238 45890 12290
rect 46734 12238 46786 12290
rect 50206 12238 50258 12290
rect 52110 12238 52162 12290
rect 55694 12238 55746 12290
rect 8766 12126 8818 12178
rect 9774 12126 9826 12178
rect 10222 12126 10274 12178
rect 12238 12126 12290 12178
rect 12798 12126 12850 12178
rect 14590 12126 14642 12178
rect 14926 12126 14978 12178
rect 15598 12126 15650 12178
rect 15710 12126 15762 12178
rect 15934 12126 15986 12178
rect 16158 12126 16210 12178
rect 19182 12126 19234 12178
rect 26798 12126 26850 12178
rect 39678 12126 39730 12178
rect 41134 12126 41186 12178
rect 41582 12126 41634 12178
rect 45950 12126 46002 12178
rect 46622 12126 46674 12178
rect 47518 12126 47570 12178
rect 48750 12126 48802 12178
rect 49310 12126 49362 12178
rect 51214 12126 51266 12178
rect 51774 12126 51826 12178
rect 52782 12126 52834 12178
rect 53006 12126 53058 12178
rect 54462 12126 54514 12178
rect 54574 12126 54626 12178
rect 55358 12126 55410 12178
rect 9662 12014 9714 12066
rect 12350 12014 12402 12066
rect 17614 12014 17666 12066
rect 22094 12014 22146 12066
rect 29710 12014 29762 12066
rect 34638 12014 34690 12066
rect 40014 12014 40066 12066
rect 41246 12014 41298 12066
rect 49870 12014 49922 12066
rect 14926 11902 14978 11954
rect 40126 11902 40178 11954
rect 53342 11902 53394 11954
rect 53902 11902 53954 11954
rect 54014 11902 54066 11954
rect 54238 11902 54290 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 8990 11566 9042 11618
rect 9662 11566 9714 11618
rect 45502 11566 45554 11618
rect 46958 11566 47010 11618
rect 2494 11454 2546 11506
rect 4622 11454 4674 11506
rect 5742 11454 5794 11506
rect 6638 11454 6690 11506
rect 8430 11454 8482 11506
rect 10782 11454 10834 11506
rect 12910 11454 12962 11506
rect 13582 11454 13634 11506
rect 16158 11454 16210 11506
rect 18286 11454 18338 11506
rect 24222 11454 24274 11506
rect 25118 11454 25170 11506
rect 31838 11454 31890 11506
rect 33966 11454 34018 11506
rect 37998 11454 38050 11506
rect 40126 11454 40178 11506
rect 42814 11454 42866 11506
rect 45726 11454 45778 11506
rect 46062 11454 46114 11506
rect 47070 11454 47122 11506
rect 51998 11454 52050 11506
rect 55246 11454 55298 11506
rect 57374 11454 57426 11506
rect 1822 11342 1874 11394
rect 5854 11342 5906 11394
rect 6302 11342 6354 11394
rect 8318 11342 8370 11394
rect 8654 11342 8706 11394
rect 8878 11342 8930 11394
rect 10110 11342 10162 11394
rect 13470 11342 13522 11394
rect 13694 11342 13746 11394
rect 14590 11342 14642 11394
rect 15486 11342 15538 11394
rect 21310 11342 21362 11394
rect 24782 11342 24834 11394
rect 31166 11342 31218 11394
rect 40910 11342 40962 11394
rect 41918 11342 41970 11394
rect 45950 11342 46002 11394
rect 47294 11342 47346 11394
rect 48190 11342 48242 11394
rect 49646 11342 49698 11394
rect 50206 11342 50258 11394
rect 50990 11342 51042 11394
rect 53118 11342 53170 11394
rect 53566 11342 53618 11394
rect 58046 11342 58098 11394
rect 5630 11230 5682 11282
rect 13918 11230 13970 11282
rect 14478 11230 14530 11282
rect 22094 11230 22146 11282
rect 26462 11230 26514 11282
rect 42254 11230 42306 11282
rect 42478 11230 42530 11282
rect 48078 11230 48130 11282
rect 49422 11230 49474 11282
rect 50878 11230 50930 11282
rect 51438 11230 51490 11282
rect 53678 11230 53730 11282
rect 9326 11118 9378 11170
rect 14254 11118 14306 11170
rect 25678 11118 25730 11170
rect 26574 11118 26626 11170
rect 42030 11118 42082 11170
rect 42142 11118 42194 11170
rect 42926 11118 42978 11170
rect 46174 11118 46226 11170
rect 47854 11118 47906 11170
rect 51326 11118 51378 11170
rect 52110 11118 52162 11170
rect 52782 11118 52834 11170
rect 53006 11118 53058 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 4174 10782 4226 10834
rect 5518 10782 5570 10834
rect 6638 10782 6690 10834
rect 23662 10782 23714 10834
rect 37438 10782 37490 10834
rect 38222 10782 38274 10834
rect 53566 10782 53618 10834
rect 14254 10670 14306 10722
rect 15598 10670 15650 10722
rect 23102 10670 23154 10722
rect 24110 10670 24162 10722
rect 35198 10670 35250 10722
rect 41582 10670 41634 10722
rect 49758 10670 49810 10722
rect 50094 10670 50146 10722
rect 50318 10670 50370 10722
rect 4510 10558 4562 10610
rect 4734 10558 4786 10610
rect 5630 10558 5682 10610
rect 5742 10558 5794 10610
rect 6190 10558 6242 10610
rect 14030 10558 14082 10610
rect 14366 10558 14418 10610
rect 14814 10558 14866 10610
rect 15038 10558 15090 10610
rect 15262 10558 15314 10610
rect 18958 10558 19010 10610
rect 22542 10558 22594 10610
rect 22654 10558 22706 10610
rect 22878 10558 22930 10610
rect 23438 10558 23490 10610
rect 23886 10558 23938 10610
rect 28142 10558 28194 10610
rect 29374 10558 29426 10610
rect 34526 10558 34578 10610
rect 39006 10558 39058 10610
rect 39342 10558 39394 10610
rect 40014 10558 40066 10610
rect 45614 10558 45666 10610
rect 46846 10558 46898 10610
rect 47182 10558 47234 10610
rect 47630 10558 47682 10610
rect 18510 10446 18562 10498
rect 19630 10446 19682 10498
rect 21758 10446 21810 10498
rect 22766 10446 22818 10498
rect 23774 10446 23826 10498
rect 25342 10446 25394 10498
rect 27470 10446 27522 10498
rect 30158 10446 30210 10498
rect 32286 10446 32338 10498
rect 48862 10446 48914 10498
rect 49870 10446 49922 10498
rect 53678 10446 53730 10498
rect 39454 10334 39506 10386
rect 47406 10334 47458 10386
rect 48078 10334 48130 10386
rect 48750 10334 48802 10386
rect 53790 10334 53842 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19966 9998 20018 10050
rect 20302 9998 20354 10050
rect 22206 9998 22258 10050
rect 26798 9998 26850 10050
rect 27806 9998 27858 10050
rect 47742 9998 47794 10050
rect 5070 9886 5122 9938
rect 5630 9886 5682 9938
rect 7310 9886 7362 9938
rect 20750 9886 20802 9938
rect 22094 9886 22146 9938
rect 30158 9886 30210 9938
rect 37998 9886 38050 9938
rect 49422 9886 49474 9938
rect 55470 9886 55522 9938
rect 2158 9774 2210 9826
rect 5854 9774 5906 9826
rect 6862 9774 6914 9826
rect 10110 9774 10162 9826
rect 14926 9774 14978 9826
rect 19070 9774 19122 9826
rect 21870 9774 21922 9826
rect 26238 9774 26290 9826
rect 26574 9774 26626 9826
rect 27022 9774 27074 9826
rect 29822 9774 29874 9826
rect 30046 9774 30098 9826
rect 30382 9774 30434 9826
rect 30606 9774 30658 9826
rect 31390 9774 31442 9826
rect 37662 9774 37714 9826
rect 38334 9774 38386 9826
rect 39230 9774 39282 9826
rect 39454 9774 39506 9826
rect 39566 9774 39618 9826
rect 41022 9774 41074 9826
rect 42590 9774 42642 9826
rect 47406 9774 47458 9826
rect 47966 9774 48018 9826
rect 48526 9774 48578 9826
rect 48862 9774 48914 9826
rect 49870 9774 49922 9826
rect 50542 9774 50594 9826
rect 52110 9774 52162 9826
rect 52894 9774 52946 9826
rect 2942 9662 2994 9714
rect 6190 9662 6242 9714
rect 9438 9662 9490 9714
rect 17390 9662 17442 9714
rect 28142 9662 28194 9714
rect 30718 9662 30770 9714
rect 30830 9662 30882 9714
rect 30942 9662 30994 9714
rect 33966 9662 34018 9714
rect 34302 9662 34354 9714
rect 41470 9662 41522 9714
rect 42254 9662 42306 9714
rect 6638 9550 6690 9602
rect 19406 9550 19458 9602
rect 20078 9550 20130 9602
rect 26686 9550 26738 9602
rect 27918 9550 27970 9602
rect 28590 9550 28642 9602
rect 34190 9550 34242 9602
rect 38670 9550 38722 9602
rect 39118 9550 39170 9602
rect 39342 9550 39394 9602
rect 40910 9550 40962 9602
rect 41134 9550 41186 9602
rect 41246 9550 41298 9602
rect 49982 9550 50034 9602
rect 50094 9550 50146 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 6078 9214 6130 9266
rect 7310 9214 7362 9266
rect 8654 9214 8706 9266
rect 9662 9214 9714 9266
rect 10670 9214 10722 9266
rect 12238 9214 12290 9266
rect 14814 9214 14866 9266
rect 16270 9214 16322 9266
rect 25454 9214 25506 9266
rect 28814 9214 28866 9266
rect 29262 9214 29314 9266
rect 30382 9214 30434 9266
rect 49086 9214 49138 9266
rect 49758 9214 49810 9266
rect 49870 9214 49922 9266
rect 51326 9214 51378 9266
rect 52782 9214 52834 9266
rect 57598 9214 57650 9266
rect 57822 9214 57874 9266
rect 58158 9214 58210 9266
rect 5966 9102 6018 9154
rect 7198 9102 7250 9154
rect 8766 9102 8818 9154
rect 8990 9102 9042 9154
rect 9774 9102 9826 9154
rect 16494 9102 16546 9154
rect 18174 9102 18226 9154
rect 29150 9102 29202 9154
rect 40126 9102 40178 9154
rect 41246 9102 41298 9154
rect 43710 9102 43762 9154
rect 48078 9102 48130 9154
rect 49982 9102 50034 9154
rect 52894 9102 52946 9154
rect 56926 9102 56978 9154
rect 6302 8990 6354 9042
rect 8430 8990 8482 9042
rect 9550 8990 9602 9042
rect 10222 8990 10274 9042
rect 12574 8990 12626 9042
rect 14030 8990 14082 9042
rect 15150 8990 15202 9042
rect 16718 8990 16770 9042
rect 17390 8990 17442 9042
rect 20974 8990 21026 9042
rect 29486 8990 29538 9042
rect 36206 8990 36258 9042
rect 36542 8990 36594 9042
rect 42926 8990 42978 9042
rect 46174 8990 46226 9042
rect 48190 8990 48242 9042
rect 48750 8990 48802 9042
rect 48974 8990 49026 9042
rect 49422 8990 49474 9042
rect 50990 8990 51042 9042
rect 51214 8990 51266 9042
rect 51438 8990 51490 9042
rect 51662 8990 51714 9042
rect 53006 8990 53058 9042
rect 53230 8990 53282 9042
rect 53454 8990 53506 9042
rect 53790 8990 53842 9042
rect 54238 8990 54290 9042
rect 54574 8990 54626 9042
rect 55246 8990 55298 9042
rect 55470 8990 55522 9042
rect 56590 8990 56642 9042
rect 12910 8878 12962 8930
rect 13470 8878 13522 8930
rect 14254 8878 14306 8930
rect 15598 8878 15650 8930
rect 20302 8878 20354 8930
rect 20750 8878 20802 8930
rect 33294 8878 33346 8930
rect 35422 8878 35474 8930
rect 37326 8878 37378 8930
rect 39454 8878 39506 8930
rect 45838 8878 45890 8930
rect 52334 8878 52386 8930
rect 7310 8766 7362 8818
rect 12574 8766 12626 8818
rect 20638 8766 20690 8818
rect 40238 8766 40290 8818
rect 41358 8766 41410 8818
rect 46286 8766 46338 8818
rect 54014 8766 54066 8818
rect 54462 8766 54514 8818
rect 54910 8766 54962 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 37998 8430 38050 8482
rect 47182 8430 47234 8482
rect 47630 8430 47682 8482
rect 8654 8318 8706 8370
rect 17278 8318 17330 8370
rect 19406 8318 19458 8370
rect 24222 8318 24274 8370
rect 26462 8318 26514 8370
rect 35086 8318 35138 8370
rect 38110 8318 38162 8370
rect 40462 8318 40514 8370
rect 42142 8318 42194 8370
rect 44270 8318 44322 8370
rect 49758 8318 49810 8370
rect 50318 8318 50370 8370
rect 54014 8318 54066 8370
rect 55246 8318 55298 8370
rect 57374 8318 57426 8370
rect 9214 8206 9266 8258
rect 20190 8206 20242 8258
rect 21310 8206 21362 8258
rect 24782 8206 24834 8258
rect 25566 8206 25618 8258
rect 25790 8206 25842 8258
rect 33966 8206 34018 8258
rect 34750 8206 34802 8258
rect 41470 8206 41522 8258
rect 49982 8206 50034 8258
rect 52894 8206 52946 8258
rect 53902 8206 53954 8258
rect 58046 8206 58098 8258
rect 8766 8094 8818 8146
rect 8990 8094 9042 8146
rect 22094 8094 22146 8146
rect 25902 8094 25954 8146
rect 33854 8094 33906 8146
rect 34190 8094 34242 8146
rect 34414 8094 34466 8146
rect 46846 8094 46898 8146
rect 47518 8094 47570 8146
rect 53118 8094 53170 8146
rect 54462 8094 54514 8146
rect 54910 8094 54962 8146
rect 9662 7982 9714 8034
rect 24558 7982 24610 8034
rect 30270 7982 30322 8034
rect 30606 7982 30658 8034
rect 34974 7982 35026 8034
rect 47070 7982 47122 8034
rect 47630 7982 47682 8034
rect 49646 7982 49698 8034
rect 49870 7982 49922 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 25454 7646 25506 7698
rect 26014 7646 26066 7698
rect 26126 7646 26178 7698
rect 29822 7646 29874 7698
rect 35646 7646 35698 7698
rect 39902 7646 39954 7698
rect 40014 7646 40066 7698
rect 41358 7646 41410 7698
rect 42702 7646 42754 7698
rect 43598 7646 43650 7698
rect 46062 7646 46114 7698
rect 46958 7646 47010 7698
rect 49982 7646 50034 7698
rect 9998 7534 10050 7586
rect 10334 7534 10386 7586
rect 12014 7534 12066 7586
rect 20190 7534 20242 7586
rect 27134 7534 27186 7586
rect 30270 7534 30322 7586
rect 30606 7534 30658 7586
rect 31726 7534 31778 7586
rect 39230 7534 39282 7586
rect 41134 7534 41186 7586
rect 47070 7534 47122 7586
rect 53118 7534 53170 7586
rect 53230 7534 53282 7586
rect 53342 7534 53394 7586
rect 53790 7534 53842 7586
rect 54014 7534 54066 7586
rect 54350 7534 54402 7586
rect 56926 7534 56978 7586
rect 7310 7422 7362 7474
rect 7758 7422 7810 7474
rect 11230 7422 11282 7474
rect 24670 7422 24722 7474
rect 25902 7422 25954 7474
rect 26238 7422 26290 7474
rect 26462 7422 26514 7474
rect 26910 7422 26962 7474
rect 29486 7422 29538 7474
rect 30830 7422 30882 7474
rect 31614 7422 31666 7474
rect 31950 7422 32002 7474
rect 34862 7422 34914 7474
rect 39678 7422 39730 7474
rect 39790 7422 39842 7474
rect 40238 7422 40290 7474
rect 40910 7422 40962 7474
rect 41582 7422 41634 7474
rect 45950 7422 46002 7474
rect 46398 7422 46450 7474
rect 46622 7422 46674 7474
rect 46846 7422 46898 7474
rect 47406 7422 47458 7474
rect 50094 7422 50146 7474
rect 55022 7422 55074 7474
rect 55358 7422 55410 7474
rect 56590 7422 56642 7474
rect 8206 7310 8258 7362
rect 14142 7310 14194 7362
rect 19070 7310 19122 7362
rect 29710 7310 29762 7362
rect 30382 7310 30434 7362
rect 31166 7310 31218 7362
rect 34638 7310 34690 7362
rect 41134 7310 41186 7362
rect 42254 7310 42306 7362
rect 43150 7310 43202 7362
rect 54238 7310 54290 7362
rect 54798 7310 54850 7362
rect 26798 7198 26850 7250
rect 27358 7198 27410 7250
rect 27582 7198 27634 7250
rect 29822 7198 29874 7250
rect 35198 7198 35250 7250
rect 39118 7198 39170 7250
rect 43038 7198 43090 7250
rect 43598 7198 43650 7250
rect 49982 7198 50034 7250
rect 52670 7198 52722 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 43486 6862 43538 6914
rect 48974 6862 49026 6914
rect 50094 6862 50146 6914
rect 53342 6862 53394 6914
rect 53790 6862 53842 6914
rect 5966 6750 6018 6802
rect 16382 6750 16434 6802
rect 16830 6750 16882 6802
rect 19630 6750 19682 6802
rect 21870 6750 21922 6802
rect 21982 6750 22034 6802
rect 22878 6750 22930 6802
rect 27022 6750 27074 6802
rect 29934 6750 29986 6802
rect 32062 6750 32114 6802
rect 33854 6750 33906 6802
rect 43262 6750 43314 6802
rect 45726 6750 45778 6802
rect 46622 6750 46674 6802
rect 52222 6750 52274 6802
rect 53230 6750 53282 6802
rect 54574 6750 54626 6802
rect 55246 6750 55298 6802
rect 8878 6638 8930 6690
rect 13582 6638 13634 6690
rect 17390 6638 17442 6690
rect 19294 6638 19346 6690
rect 19518 6638 19570 6690
rect 19966 6638 20018 6690
rect 21646 6638 21698 6690
rect 22990 6638 23042 6690
rect 23214 6638 23266 6690
rect 24222 6638 24274 6690
rect 24894 6638 24946 6690
rect 29150 6638 29202 6690
rect 33518 6638 33570 6690
rect 35086 6638 35138 6690
rect 35982 6638 36034 6690
rect 42254 6638 42306 6690
rect 42702 6638 42754 6690
rect 43038 6638 43090 6690
rect 43710 6638 43762 6690
rect 44046 6638 44098 6690
rect 45054 6638 45106 6690
rect 45390 6638 45442 6690
rect 45838 6638 45890 6690
rect 47182 6638 47234 6690
rect 49310 6638 49362 6690
rect 49646 6638 49698 6690
rect 53566 6638 53618 6690
rect 57374 6638 57426 6690
rect 58046 6638 58098 6690
rect 8094 6526 8146 6578
rect 14254 6526 14306 6578
rect 22542 6526 22594 6578
rect 22766 6526 22818 6578
rect 34302 6526 34354 6578
rect 35310 6526 35362 6578
rect 36094 6526 36146 6578
rect 37214 6526 37266 6578
rect 46062 6526 46114 6578
rect 46398 6526 46450 6578
rect 49870 6526 49922 6578
rect 50766 6526 50818 6578
rect 51102 6526 51154 6578
rect 52894 6526 52946 6578
rect 16830 6414 16882 6466
rect 16942 6414 16994 6466
rect 17166 6414 17218 6466
rect 19742 6414 19794 6466
rect 36318 6414 36370 6466
rect 42590 6414 42642 6466
rect 43486 6414 43538 6466
rect 45614 6414 45666 6466
rect 46622 6414 46674 6466
rect 49086 6414 49138 6466
rect 50430 6414 50482 6466
rect 53678 6414 53730 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 7982 6078 8034 6130
rect 16270 6078 16322 6130
rect 16830 6078 16882 6130
rect 17950 6078 18002 6130
rect 21310 6078 21362 6130
rect 23550 6078 23602 6130
rect 26014 6078 26066 6130
rect 26686 6078 26738 6130
rect 49646 6078 49698 6130
rect 7870 5966 7922 6018
rect 8094 5966 8146 6018
rect 8542 5966 8594 6018
rect 16382 5966 16434 6018
rect 17390 5966 17442 6018
rect 25230 5966 25282 6018
rect 26462 5966 26514 6018
rect 29150 5966 29202 6018
rect 33854 5966 33906 6018
rect 34974 5966 35026 6018
rect 38222 5966 38274 6018
rect 47854 5966 47906 6018
rect 50094 5966 50146 6018
rect 50206 5966 50258 6018
rect 15710 5854 15762 5906
rect 16046 5854 16098 5906
rect 17614 5854 17666 5906
rect 17838 5854 17890 5906
rect 21646 5854 21698 5906
rect 23774 5854 23826 5906
rect 24446 5854 24498 5906
rect 25454 5854 25506 5906
rect 25790 5854 25842 5906
rect 27134 5854 27186 5906
rect 34414 5854 34466 5906
rect 34638 5854 34690 5906
rect 35310 5854 35362 5906
rect 37550 5854 37602 5906
rect 46174 5854 46226 5906
rect 46958 5854 47010 5906
rect 47406 5854 47458 5906
rect 50318 5854 50370 5906
rect 56030 5854 56082 5906
rect 13358 5742 13410 5794
rect 17726 5742 17778 5794
rect 24334 5742 24386 5794
rect 26574 5742 26626 5794
rect 40350 5742 40402 5794
rect 41134 5742 41186 5794
rect 46510 5742 46562 5794
rect 47966 5742 48018 5794
rect 53118 5742 53170 5794
rect 55246 5742 55298 5794
rect 25790 5630 25842 5682
rect 35310 5630 35362 5682
rect 50766 5630 50818 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 16270 5294 16322 5346
rect 30046 5294 30098 5346
rect 44830 5294 44882 5346
rect 45726 5294 45778 5346
rect 10670 5182 10722 5234
rect 12798 5182 12850 5234
rect 15934 5182 15986 5234
rect 18734 5182 18786 5234
rect 19182 5182 19234 5234
rect 19518 5182 19570 5234
rect 24110 5182 24162 5234
rect 26238 5182 26290 5234
rect 26686 5182 26738 5234
rect 27470 5182 27522 5234
rect 33518 5182 33570 5234
rect 35646 5182 35698 5234
rect 41358 5182 41410 5234
rect 42702 5182 42754 5234
rect 45502 5182 45554 5234
rect 46398 5182 46450 5234
rect 52222 5182 52274 5234
rect 54686 5182 54738 5234
rect 9326 5070 9378 5122
rect 9998 5070 10050 5122
rect 18174 5070 18226 5122
rect 18398 5070 18450 5122
rect 20750 5070 20802 5122
rect 21646 5070 21698 5122
rect 22430 5070 22482 5122
rect 22766 5070 22818 5122
rect 23102 5070 23154 5122
rect 26574 5070 26626 5122
rect 26910 5070 26962 5122
rect 29710 5070 29762 5122
rect 30718 5070 30770 5122
rect 36318 5070 36370 5122
rect 38558 5070 38610 5122
rect 41694 5070 41746 5122
rect 49310 5070 49362 5122
rect 50990 5070 51042 5122
rect 52670 5070 52722 5122
rect 16046 4958 16098 5010
rect 18734 4958 18786 5010
rect 19406 4958 19458 5010
rect 20414 4958 20466 5010
rect 21422 4958 21474 5010
rect 21982 4958 22034 5010
rect 30382 4958 30434 5010
rect 31502 4958 31554 5010
rect 31838 4958 31890 5010
rect 39230 4958 39282 5010
rect 44942 4958 44994 5010
rect 48526 4958 48578 5010
rect 9550 4846 9602 4898
rect 18622 4846 18674 4898
rect 21758 4846 21810 4898
rect 21870 4846 21922 4898
rect 22542 4846 22594 4898
rect 29934 4846 29986 4898
rect 46062 4846 46114 4898
rect 51326 4846 51378 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 33294 4510 33346 4562
rect 34414 4510 34466 4562
rect 34526 4510 34578 4562
rect 47742 4510 47794 4562
rect 54126 4510 54178 4562
rect 10894 4398 10946 4450
rect 14590 4398 14642 4450
rect 19966 4398 20018 4450
rect 22094 4398 22146 4450
rect 26014 4398 26066 4450
rect 30046 4398 30098 4450
rect 33182 4398 33234 4450
rect 34638 4398 34690 4450
rect 36878 4398 36930 4450
rect 41918 4398 41970 4450
rect 47406 4398 47458 4450
rect 48078 4398 48130 4450
rect 52670 4398 52722 4450
rect 53790 4398 53842 4450
rect 57822 4398 57874 4450
rect 10222 4286 10274 4338
rect 13806 4286 13858 4338
rect 20638 4286 20690 4338
rect 21310 4286 21362 4338
rect 25230 4286 25282 4338
rect 29262 4286 29314 4338
rect 36206 4286 36258 4338
rect 41134 4286 41186 4338
rect 44494 4286 44546 4338
rect 53454 4286 53506 4338
rect 58158 4286 58210 4338
rect 13022 4174 13074 4226
rect 16718 4174 16770 4226
rect 17838 4174 17890 4226
rect 24222 4174 24274 4226
rect 28142 4174 28194 4226
rect 32174 4174 32226 4226
rect 39006 4174 39058 4226
rect 44046 4174 44098 4226
rect 48862 4174 48914 4226
rect 50542 4174 50594 4226
rect 57598 4174 57650 4226
rect 45390 4062 45442 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 18846 3614 18898 3666
rect 22094 3614 22146 3666
rect 26126 3614 26178 3666
rect 40798 3614 40850 3666
rect 43150 3614 43202 3666
rect 44382 3614 44434 3666
rect 46510 3614 46562 3666
rect 20078 3502 20130 3554
rect 21086 3502 21138 3554
rect 25230 3502 25282 3554
rect 36654 3502 36706 3554
rect 39790 3502 39842 3554
rect 43710 3502 43762 3554
rect 47406 3502 47458 3554
rect 48974 3390 49026 3442
rect 2942 3278 2994 3330
rect 5518 3278 5570 3330
rect 6974 3278 7026 3330
rect 9326 3278 9378 3330
rect 11006 3278 11058 3330
rect 13134 3278 13186 3330
rect 15038 3278 15090 3330
rect 17054 3278 17106 3330
rect 28366 3278 28418 3330
rect 29150 3278 29202 3330
rect 31166 3278 31218 3330
rect 33182 3278 33234 3330
rect 35198 3278 35250 3330
rect 37662 3278 37714 3330
rect 50318 3278 50370 3330
rect 51326 3278 51378 3330
rect 53342 3278 53394 3330
rect 55358 3278 55410 3330
rect 57374 3278 57426 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
rect 26910 1710 26962 1762
rect 28366 1710 28418 1762
rect 49086 1710 49138 1762
rect 50318 1710 50370 1762
<< metal2 >>
rect 7392 59200 7504 60000
rect 22400 59200 22512 60000
rect 37408 59200 37520 60000
rect 52416 59200 52528 60000
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 7420 55468 7476 59200
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 22428 56308 22484 59200
rect 22652 56308 22708 56318
rect 22428 56306 22708 56308
rect 22428 56254 22430 56306
rect 22482 56254 22654 56306
rect 22706 56254 22708 56306
rect 22428 56252 22708 56254
rect 22428 56242 22484 56252
rect 22652 56242 22708 56252
rect 27020 56306 27076 56318
rect 27020 56254 27022 56306
rect 27074 56254 27076 56306
rect 26684 56082 26740 56094
rect 26684 56030 26686 56082
rect 26738 56030 26740 56082
rect 23100 55972 23156 55982
rect 23100 55878 23156 55916
rect 7420 55412 7588 55468
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 6188 48242 6244 48254
rect 6188 48190 6190 48242
rect 6242 48190 6244 48242
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 6188 47572 6244 48190
rect 6860 48132 6916 48142
rect 6860 48038 6916 48076
rect 6188 47478 6244 47516
rect 6972 47572 7028 47582
rect 6972 46674 7028 47516
rect 6972 46622 6974 46674
rect 7026 46622 7028 46674
rect 6972 46610 7028 46622
rect 4172 46562 4228 46574
rect 4172 46510 4174 46562
rect 4226 46510 4228 46562
rect 4172 45892 4228 46510
rect 6300 46564 6356 46574
rect 6300 46470 6356 46508
rect 7420 46450 7476 46462
rect 7420 46398 7422 46450
rect 7474 46398 7476 46450
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 7196 46004 7252 46014
rect 4172 45826 4228 45836
rect 6748 45892 6804 45902
rect 6748 45798 6804 45836
rect 7196 45890 7252 45948
rect 7308 46004 7364 46014
rect 7420 46004 7476 46398
rect 7308 46002 7476 46004
rect 7308 45950 7310 46002
rect 7362 45950 7476 46002
rect 7308 45948 7476 45950
rect 7308 45938 7364 45948
rect 7196 45838 7198 45890
rect 7250 45838 7252 45890
rect 7196 45826 7252 45838
rect 7420 45556 7476 45566
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 7420 44546 7476 45500
rect 7420 44494 7422 44546
rect 7474 44494 7476 44546
rect 7420 44482 7476 44494
rect 7308 44210 7364 44222
rect 7308 44158 7310 44210
rect 7362 44158 7364 44210
rect 4732 43876 4788 43886
rect 4732 43426 4788 43820
rect 7308 43708 7364 44158
rect 7532 43708 7588 55412
rect 20412 55410 20468 55422
rect 25788 55412 25844 55422
rect 20412 55358 20414 55410
rect 20466 55358 20468 55410
rect 17500 55298 17556 55310
rect 17500 55246 17502 55298
rect 17554 55246 17556 55298
rect 17500 54514 17556 55246
rect 18284 55188 18340 55198
rect 18284 55094 18340 55132
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 17500 54462 17502 54514
rect 17554 54462 17556 54514
rect 17500 52836 17556 54462
rect 18172 54402 18228 54414
rect 18172 54350 18174 54402
rect 18226 54350 18228 54402
rect 18172 53732 18228 54350
rect 20300 54404 20356 54414
rect 20300 54310 20356 54348
rect 20412 54404 20468 55358
rect 20748 55356 21476 55412
rect 20636 54514 20692 54526
rect 20636 54462 20638 54514
rect 20690 54462 20692 54514
rect 20636 54404 20692 54462
rect 20412 54348 20692 54404
rect 18172 53666 18228 53676
rect 20188 53732 20244 53742
rect 20188 53638 20244 53676
rect 20300 53730 20356 53742
rect 20300 53678 20302 53730
rect 20354 53678 20356 53730
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 19068 52948 19124 52958
rect 19124 52892 19236 52948
rect 19068 52854 19124 52892
rect 17500 52770 17556 52780
rect 18060 52276 18116 52286
rect 18060 52182 18116 52220
rect 15260 52162 15316 52174
rect 15260 52110 15262 52162
rect 15314 52110 15316 52162
rect 14364 50482 14420 50494
rect 14364 50430 14366 50482
rect 14418 50430 14420 50482
rect 14252 49812 14308 49822
rect 14364 49812 14420 50430
rect 15260 50428 15316 52110
rect 15932 52052 15988 52062
rect 15932 51958 15988 51996
rect 18844 51268 18900 51278
rect 18396 51266 18900 51268
rect 18396 51214 18846 51266
rect 18898 51214 18900 51266
rect 18396 51212 18900 51214
rect 16156 51156 16212 51166
rect 15260 50372 15428 50428
rect 14028 49810 14364 49812
rect 14028 49758 14254 49810
rect 14306 49758 14364 49810
rect 14028 49756 14364 49758
rect 11340 49698 11396 49710
rect 11340 49646 11342 49698
rect 11394 49646 11396 49698
rect 7980 48914 8036 48926
rect 7980 48862 7982 48914
rect 8034 48862 8036 48914
rect 7756 46674 7812 46686
rect 7756 46622 7758 46674
rect 7810 46622 7812 46674
rect 7644 46564 7700 46574
rect 7644 46470 7700 46508
rect 7756 45556 7812 46622
rect 7980 46004 8036 48862
rect 8092 48804 8148 48814
rect 8092 48710 8148 48748
rect 8316 48802 8372 48814
rect 8316 48750 8318 48802
rect 8370 48750 8372 48802
rect 8316 48356 8372 48750
rect 10444 48804 10500 48814
rect 10500 48748 10612 48804
rect 10444 48738 10500 48748
rect 8316 48290 8372 48300
rect 9548 48356 9604 48366
rect 9548 48262 9604 48300
rect 9772 48354 9828 48366
rect 9772 48302 9774 48354
rect 9826 48302 9828 48354
rect 8988 48130 9044 48142
rect 8988 48078 8990 48130
rect 9042 48078 9044 48130
rect 8988 47684 9044 48078
rect 9660 48132 9716 48142
rect 9660 48038 9716 48076
rect 8764 47628 9044 47684
rect 8764 46786 8820 47628
rect 9772 47348 9828 48302
rect 8764 46734 8766 46786
rect 8818 46734 8820 46786
rect 7980 45892 8036 45948
rect 8540 46450 8596 46462
rect 8540 46398 8542 46450
rect 8594 46398 8596 46450
rect 8204 45892 8260 45902
rect 8540 45892 8596 46398
rect 7980 45890 8260 45892
rect 7980 45838 8206 45890
rect 8258 45838 8260 45890
rect 7980 45836 8260 45838
rect 8204 45826 8260 45836
rect 8316 45890 8596 45892
rect 8316 45838 8542 45890
rect 8594 45838 8596 45890
rect 8316 45836 8596 45838
rect 7756 45490 7812 45500
rect 8204 45108 8260 45118
rect 7644 44436 7700 44446
rect 7644 44342 7700 44380
rect 7868 44324 7924 44334
rect 7868 44230 7924 44268
rect 8204 44210 8260 45052
rect 8316 44324 8372 45836
rect 8540 45826 8596 45836
rect 8428 45668 8484 45678
rect 8764 45668 8820 46734
rect 8876 47292 9828 47348
rect 10444 47458 10500 47470
rect 10444 47406 10446 47458
rect 10498 47406 10500 47458
rect 8876 46562 8932 47292
rect 10444 47236 10500 47406
rect 10220 46676 10276 46686
rect 10220 46674 10388 46676
rect 10220 46622 10222 46674
rect 10274 46622 10388 46674
rect 10220 46620 10388 46622
rect 10220 46610 10276 46620
rect 8876 46510 8878 46562
rect 8930 46510 8932 46562
rect 8876 46498 8932 46510
rect 8428 45666 8820 45668
rect 8428 45614 8430 45666
rect 8482 45614 8820 45666
rect 8428 45612 8820 45614
rect 9548 45892 9604 45902
rect 8428 45220 8484 45612
rect 8540 45220 8596 45230
rect 8428 45164 8540 45220
rect 8540 45154 8596 45164
rect 9548 45106 9604 45836
rect 9660 45220 9716 45230
rect 9660 45126 9716 45164
rect 9548 45054 9550 45106
rect 9602 45054 9604 45106
rect 9548 45042 9604 45054
rect 9884 45108 9940 45118
rect 9884 45014 9940 45052
rect 10220 45106 10276 45118
rect 10220 45054 10222 45106
rect 10274 45054 10276 45106
rect 8316 44258 8372 44268
rect 8540 44436 8596 44446
rect 8204 44158 8206 44210
rect 8258 44158 8260 44210
rect 8204 43876 8260 44158
rect 8428 44210 8484 44222
rect 8428 44158 8430 44210
rect 8482 44158 8484 44210
rect 8428 43988 8484 44158
rect 8540 44098 8596 44380
rect 8876 44322 8932 44334
rect 8876 44270 8878 44322
rect 8930 44270 8932 44322
rect 8876 44212 8932 44270
rect 9660 44324 9716 44334
rect 10108 44324 10164 44334
rect 9660 44322 10164 44324
rect 9660 44270 9662 44322
rect 9714 44270 10110 44322
rect 10162 44270 10164 44322
rect 9660 44268 10164 44270
rect 9660 44258 9716 44268
rect 10108 44258 10164 44268
rect 9100 44212 9156 44222
rect 8876 44210 9156 44212
rect 8876 44158 9102 44210
rect 9154 44158 9156 44210
rect 8876 44156 9156 44158
rect 8540 44046 8542 44098
rect 8594 44046 8596 44098
rect 8540 44034 8596 44046
rect 9100 44100 9156 44156
rect 9436 44210 9492 44222
rect 9436 44158 9438 44210
rect 9490 44158 9492 44210
rect 9100 44034 9156 44044
rect 9212 44098 9268 44110
rect 9212 44046 9214 44098
rect 9266 44046 9268 44098
rect 8428 43922 8484 43932
rect 8204 43810 8260 43820
rect 6860 43652 7364 43708
rect 7420 43652 7588 43708
rect 6860 43650 6916 43652
rect 6860 43598 6862 43650
rect 6914 43598 6916 43650
rect 6860 43586 6916 43598
rect 4732 43374 4734 43426
rect 4786 43374 4788 43426
rect 4732 43362 4788 43374
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 4956 40628 5012 40638
rect 1820 40516 1876 40526
rect 1820 39618 1876 40460
rect 4956 40402 5012 40572
rect 4956 40350 4958 40402
rect 5010 40350 5012 40402
rect 4956 40338 5012 40350
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 1820 39566 1822 39618
rect 1874 39566 1876 39618
rect 1820 38834 1876 39566
rect 4620 39730 4676 39742
rect 4620 39678 4622 39730
rect 4674 39678 4676 39730
rect 2492 39506 2548 39518
rect 2492 39454 2494 39506
rect 2546 39454 2548 39506
rect 2492 38948 2548 39454
rect 4620 38948 4676 39678
rect 5628 39732 5684 39742
rect 5628 39730 5796 39732
rect 5628 39678 5630 39730
rect 5682 39678 5796 39730
rect 5628 39676 5796 39678
rect 5628 39666 5684 39676
rect 5292 39060 5348 39070
rect 5180 38948 5236 38958
rect 4620 38946 5236 38948
rect 4620 38894 5182 38946
rect 5234 38894 5236 38946
rect 4620 38892 5236 38894
rect 2492 38882 2548 38892
rect 1820 38782 1822 38834
rect 1874 38782 1876 38834
rect 1820 38770 1876 38782
rect 2492 38722 2548 38734
rect 2492 38670 2494 38722
rect 2546 38670 2548 38722
rect 2492 38164 2548 38670
rect 4620 38724 4676 38734
rect 4620 38722 5012 38724
rect 4620 38670 4622 38722
rect 4674 38670 5012 38722
rect 4620 38668 5012 38670
rect 4620 38658 4676 38668
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 2492 38098 2548 38108
rect 4956 37604 5012 38668
rect 5068 37828 5124 38892
rect 5180 38882 5236 38892
rect 5292 38946 5348 39004
rect 5292 38894 5294 38946
rect 5346 38894 5348 38946
rect 5292 38882 5348 38894
rect 5740 38946 5796 39676
rect 7308 39396 7364 39406
rect 5964 39060 6020 39070
rect 5964 39058 6468 39060
rect 5964 39006 5966 39058
rect 6018 39006 6468 39058
rect 5964 39004 6468 39006
rect 5964 38994 6020 39004
rect 5740 38894 5742 38946
rect 5794 38894 5796 38946
rect 5628 38834 5684 38846
rect 5628 38782 5630 38834
rect 5682 38782 5684 38834
rect 5180 38610 5236 38622
rect 5180 38558 5182 38610
rect 5234 38558 5236 38610
rect 5180 38500 5236 38558
rect 5180 38434 5236 38444
rect 5628 38052 5684 38782
rect 5740 38836 5796 38894
rect 5740 38770 5796 38780
rect 6188 38834 6244 38846
rect 6188 38782 6190 38834
rect 6242 38782 6244 38834
rect 6188 38500 6244 38782
rect 6300 38836 6356 38846
rect 6300 38742 6356 38780
rect 6412 38834 6468 39004
rect 7308 38946 7364 39340
rect 7308 38894 7310 38946
rect 7362 38894 7364 38946
rect 7308 38882 7364 38894
rect 6748 38836 6804 38846
rect 6412 38782 6414 38834
rect 6466 38782 6468 38834
rect 6412 38770 6468 38782
rect 6636 38780 6748 38836
rect 6188 38434 6244 38444
rect 5852 38164 5908 38174
rect 5852 38070 5908 38108
rect 6076 38108 6580 38164
rect 5628 37986 5684 37996
rect 6076 38050 6132 38108
rect 6076 37998 6078 38050
rect 6130 37998 6132 38050
rect 6076 37986 6132 37998
rect 6524 38050 6580 38108
rect 6524 37998 6526 38050
rect 6578 37998 6580 38050
rect 6524 37986 6580 37998
rect 5740 37938 5796 37950
rect 5740 37886 5742 37938
rect 5794 37886 5796 37938
rect 5180 37828 5236 37838
rect 5068 37772 5180 37828
rect 5180 37762 5236 37772
rect 4956 37548 5572 37604
rect 5516 37492 5572 37548
rect 5516 37490 5684 37492
rect 5516 37438 5518 37490
rect 5570 37438 5684 37490
rect 5516 37436 5684 37438
rect 5516 37426 5572 37436
rect 4956 37380 5012 37390
rect 4844 37378 5012 37380
rect 4844 37326 4958 37378
rect 5010 37326 5012 37378
rect 4844 37324 5012 37326
rect 4732 37268 4788 37278
rect 4284 37266 4788 37268
rect 4284 37214 4734 37266
rect 4786 37214 4788 37266
rect 4284 37212 4788 37214
rect 1820 36482 1876 36494
rect 1820 36430 1822 36482
rect 1874 36430 1876 36482
rect 1820 33348 1876 36430
rect 2492 36372 2548 36382
rect 2492 36278 2548 36316
rect 4172 35812 4228 35822
rect 4172 34804 4228 35756
rect 4284 35698 4340 37212
rect 4732 37202 4788 37212
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4620 36596 4676 36606
rect 4844 36596 4900 37324
rect 4956 37314 5012 37324
rect 4620 36594 4900 36596
rect 4620 36542 4622 36594
rect 4674 36542 4900 36594
rect 4620 36540 4900 36542
rect 4620 36530 4676 36540
rect 4508 36372 4564 36382
rect 4508 35922 4564 36316
rect 4508 35870 4510 35922
rect 4562 35870 4564 35922
rect 4508 35858 4564 35870
rect 4732 36260 4788 36270
rect 4732 35810 4788 36204
rect 4732 35758 4734 35810
rect 4786 35758 4788 35810
rect 4732 35746 4788 35758
rect 4284 35646 4286 35698
rect 4338 35646 4340 35698
rect 4284 35634 4340 35646
rect 4844 35700 4900 36540
rect 5068 37268 5124 37278
rect 5404 37268 5460 37278
rect 5068 37266 5460 37268
rect 5068 37214 5070 37266
rect 5122 37214 5406 37266
rect 5458 37214 5460 37266
rect 5068 37212 5460 37214
rect 5068 35812 5124 37212
rect 5404 37202 5460 37212
rect 5628 36372 5684 37436
rect 5740 37490 5796 37886
rect 6300 37938 6356 37950
rect 6300 37886 6302 37938
rect 6354 37886 6356 37938
rect 6300 37828 6356 37886
rect 6636 37828 6692 38780
rect 6748 38742 6804 38780
rect 7196 38836 7252 38846
rect 7196 38742 7252 38780
rect 6860 38052 6916 38062
rect 6916 37996 7252 38052
rect 6860 37958 6916 37996
rect 6300 37772 6692 37828
rect 6748 37828 6804 37838
rect 6748 37716 6804 37772
rect 5740 37438 5742 37490
rect 5794 37438 5796 37490
rect 5740 37426 5796 37438
rect 6636 37660 6804 37716
rect 5740 36372 5796 36382
rect 5628 36370 5796 36372
rect 5628 36318 5742 36370
rect 5794 36318 5796 36370
rect 5628 36316 5796 36318
rect 5516 36260 5572 36270
rect 5516 36166 5572 36204
rect 5068 35746 5124 35756
rect 4844 35476 4900 35644
rect 4956 35698 5012 35710
rect 4956 35646 4958 35698
rect 5010 35646 5012 35698
rect 4956 35588 5012 35646
rect 5292 35698 5348 35710
rect 5292 35646 5294 35698
rect 5346 35646 5348 35698
rect 4956 35532 5124 35588
rect 4844 35420 5012 35476
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4844 35140 4900 35150
rect 4284 34804 4340 34814
rect 4060 34802 4340 34804
rect 4060 34750 4286 34802
rect 4338 34750 4340 34802
rect 4060 34748 4340 34750
rect 2492 34692 2548 34702
rect 2492 33458 2548 34636
rect 2492 33406 2494 33458
rect 2546 33406 2548 33458
rect 2492 33394 2548 33406
rect 1820 32562 1876 33292
rect 1820 32510 1822 32562
rect 1874 32510 1876 32562
rect 1820 30210 1876 32510
rect 2492 32452 2548 32462
rect 2492 32358 2548 32396
rect 4060 31556 4116 34748
rect 4284 34738 4340 34748
rect 4620 34804 4676 34814
rect 4620 34710 4676 34748
rect 4844 34802 4900 35084
rect 4844 34750 4846 34802
rect 4898 34750 4900 34802
rect 4396 34690 4452 34702
rect 4396 34638 4398 34690
rect 4450 34638 4452 34690
rect 4396 34132 4452 34638
rect 4284 34076 4452 34132
rect 4284 33460 4340 34076
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4620 33460 4676 33470
rect 4284 33458 4676 33460
rect 4284 33406 4622 33458
rect 4674 33406 4676 33458
rect 4284 33404 4676 33406
rect 4620 32788 4676 33404
rect 4844 33124 4900 34750
rect 4956 34802 5012 35420
rect 5068 35364 5124 35532
rect 5068 35298 5124 35308
rect 5292 35140 5348 35646
rect 5516 35700 5572 35710
rect 5516 35606 5572 35644
rect 5740 35698 5796 36316
rect 5740 35646 5742 35698
rect 5794 35646 5796 35698
rect 5740 35634 5796 35646
rect 5852 36370 5908 36382
rect 5852 36318 5854 36370
rect 5906 36318 5908 36370
rect 4956 34750 4958 34802
rect 5010 34750 5012 34802
rect 4956 34738 5012 34750
rect 5068 35084 5348 35140
rect 5852 35140 5908 36318
rect 6076 35812 6132 35822
rect 6076 35718 6132 35756
rect 5964 35588 6020 35598
rect 6636 35588 6692 37660
rect 7196 37490 7252 37996
rect 7196 37438 7198 37490
rect 7250 37438 7252 37490
rect 7196 37426 7252 37438
rect 5964 35586 6692 35588
rect 5964 35534 5966 35586
rect 6018 35534 6692 35586
rect 5964 35532 6692 35534
rect 5964 35522 6020 35532
rect 6076 35252 6132 35262
rect 5964 35140 6020 35150
rect 5852 35084 5964 35140
rect 4956 34018 5012 34030
rect 4956 33966 4958 34018
rect 5010 33966 5012 34018
rect 4956 33348 5012 33966
rect 4956 33282 5012 33292
rect 4844 33068 5012 33124
rect 4620 32722 4676 32732
rect 4172 32564 4228 32574
rect 4172 31778 4228 32508
rect 4844 32562 4900 32574
rect 4844 32510 4846 32562
rect 4898 32510 4900 32562
rect 4620 32450 4676 32462
rect 4620 32398 4622 32450
rect 4674 32398 4676 32450
rect 4620 32340 4676 32398
rect 4172 31726 4174 31778
rect 4226 31726 4228 31778
rect 4172 31714 4228 31726
rect 4284 32284 4676 32340
rect 4284 31892 4340 32284
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4844 32002 4900 32510
rect 4956 32564 5012 33068
rect 5068 32788 5124 35084
rect 5964 35074 6020 35084
rect 5516 34972 5908 35028
rect 5180 34916 5236 34926
rect 5516 34916 5572 34972
rect 5180 34914 5572 34916
rect 5180 34862 5182 34914
rect 5234 34862 5572 34914
rect 5180 34860 5572 34862
rect 5852 34914 5908 34972
rect 6076 34916 6132 35196
rect 5852 34862 5854 34914
rect 5906 34862 5908 34914
rect 5180 34850 5236 34860
rect 5852 34850 5908 34862
rect 5964 34914 6132 34916
rect 5964 34862 6078 34914
rect 6130 34862 6132 34914
rect 5964 34860 6132 34862
rect 5628 34804 5684 34814
rect 5628 34710 5684 34748
rect 5740 34692 5796 34702
rect 5740 34598 5796 34636
rect 5964 33012 6020 34860
rect 6076 34850 6132 34860
rect 6412 33572 6468 33582
rect 6412 33346 6468 33516
rect 6412 33294 6414 33346
rect 6466 33294 6468 33346
rect 6412 33282 6468 33294
rect 6860 33572 6916 33582
rect 5852 32956 6020 33012
rect 6076 33122 6132 33134
rect 6076 33070 6078 33122
rect 6130 33070 6132 33122
rect 5180 32788 5236 32798
rect 5740 32788 5796 32798
rect 5068 32732 5180 32788
rect 5180 32722 5236 32732
rect 5404 32786 5796 32788
rect 5404 32734 5742 32786
rect 5794 32734 5796 32786
rect 5404 32732 5796 32734
rect 5292 32676 5348 32686
rect 5404 32676 5460 32732
rect 5740 32722 5796 32732
rect 5292 32674 5460 32676
rect 5292 32622 5294 32674
rect 5346 32622 5460 32674
rect 5292 32620 5460 32622
rect 5292 32610 5348 32620
rect 4956 32498 5012 32508
rect 5516 32564 5572 32574
rect 5852 32564 5908 32956
rect 5964 32788 6020 32798
rect 5964 32694 6020 32732
rect 5516 32562 5908 32564
rect 5516 32510 5518 32562
rect 5570 32510 5908 32562
rect 5516 32508 5908 32510
rect 5516 32498 5572 32508
rect 5068 32452 5124 32462
rect 5068 32358 5124 32396
rect 4844 31950 4846 32002
rect 4898 31950 4900 32002
rect 4844 31938 4900 31950
rect 5852 31948 5908 32508
rect 6076 32564 6132 33070
rect 6076 32470 6132 32508
rect 5852 31892 6244 31948
rect 4284 31836 4788 31892
rect 4060 31490 4116 31500
rect 4284 31554 4340 31836
rect 4732 31780 4788 31836
rect 4732 31724 4900 31780
rect 4844 31666 4900 31724
rect 4732 31610 4788 31622
rect 4284 31502 4286 31554
rect 4338 31502 4340 31554
rect 1820 30158 1822 30210
rect 1874 30158 1876 30210
rect 1820 30146 1876 30158
rect 2492 30884 2548 30894
rect 2492 30210 2548 30828
rect 4284 30436 4340 31502
rect 4508 31556 4564 31566
rect 4732 31558 4734 31610
rect 4786 31558 4788 31610
rect 4844 31614 4846 31666
rect 4898 31614 4900 31666
rect 4844 31602 4900 31614
rect 4732 31556 4788 31558
rect 4508 31554 4676 31556
rect 4508 31502 4510 31554
rect 4562 31502 4676 31554
rect 4508 31500 4676 31502
rect 4508 31490 4564 31500
rect 4508 31108 4564 31118
rect 4620 31108 4676 31500
rect 4732 31490 4788 31500
rect 5628 31556 5684 31566
rect 5628 31462 5684 31500
rect 5964 31554 6020 31566
rect 5964 31502 5966 31554
rect 6018 31502 6020 31554
rect 5964 31220 6020 31502
rect 5964 31126 6020 31164
rect 4732 31108 4788 31118
rect 4620 31106 4788 31108
rect 4620 31054 4734 31106
rect 4786 31054 4788 31106
rect 4620 31052 4788 31054
rect 4508 31014 4564 31052
rect 4732 31042 4788 31052
rect 5628 31106 5684 31118
rect 5628 31054 5630 31106
rect 5682 31054 5684 31106
rect 5180 30996 5236 31006
rect 5180 30994 5572 30996
rect 5180 30942 5182 30994
rect 5234 30942 5572 30994
rect 5180 30940 5572 30942
rect 5180 30930 5236 30940
rect 4956 30884 5012 30894
rect 4956 30790 5012 30828
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4284 30380 4564 30436
rect 2492 30158 2494 30210
rect 2546 30158 2548 30210
rect 2492 30146 2548 30158
rect 4508 29538 4564 30380
rect 4620 30322 4676 30334
rect 4620 30270 4622 30322
rect 4674 30270 4676 30322
rect 4620 29988 4676 30270
rect 5516 30210 5572 30940
rect 5516 30158 5518 30210
rect 5570 30158 5572 30210
rect 5516 30146 5572 30158
rect 5628 30212 5684 31054
rect 6188 31108 6244 31892
rect 5852 30212 5908 30222
rect 5628 30210 5908 30212
rect 5628 30158 5854 30210
rect 5906 30158 5908 30210
rect 5628 30156 5908 30158
rect 4956 29988 5012 29998
rect 4620 29932 4956 29988
rect 4508 29486 4510 29538
rect 4562 29486 4564 29538
rect 4508 29474 4564 29486
rect 4956 29428 5012 29932
rect 5404 29428 5460 29438
rect 4844 29426 5012 29428
rect 4844 29374 4958 29426
rect 5010 29374 5012 29426
rect 4844 29372 5012 29374
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4844 28868 4900 29372
rect 4956 29362 5012 29372
rect 5068 29426 5460 29428
rect 5068 29374 5406 29426
rect 5458 29374 5460 29426
rect 5068 29372 5460 29374
rect 4396 28812 4900 28868
rect 4396 28530 4452 28812
rect 4396 28478 4398 28530
rect 4450 28478 4452 28530
rect 4396 28466 4452 28478
rect 4508 28530 4564 28542
rect 4508 28478 4510 28530
rect 4562 28478 4564 28530
rect 4172 28418 4228 28430
rect 4172 28366 4174 28418
rect 4226 28366 4228 28418
rect 1820 27858 1876 27870
rect 1820 27806 1822 27858
rect 1874 27806 1876 27858
rect 1820 24724 1876 27806
rect 3836 27860 3892 27870
rect 2492 27748 2548 27758
rect 2492 27654 2548 27692
rect 3836 27074 3892 27804
rect 3948 27748 4004 27758
rect 3948 27186 4004 27692
rect 3948 27134 3950 27186
rect 4002 27134 4004 27186
rect 3948 27122 4004 27134
rect 3836 27022 3838 27074
rect 3890 27022 3892 27074
rect 3836 27010 3892 27022
rect 4172 27074 4228 28366
rect 4508 27636 4564 28478
rect 5068 28084 5124 29372
rect 5404 29362 5460 29372
rect 4620 28082 5124 28084
rect 4620 28030 5070 28082
rect 5122 28030 5124 28082
rect 4620 28028 5124 28030
rect 4620 27746 4676 28028
rect 5068 28018 5124 28028
rect 4844 27860 4900 27870
rect 4844 27766 4900 27804
rect 5180 27860 5236 27870
rect 5628 27860 5684 30156
rect 5852 30146 5908 30156
rect 6188 30098 6244 31052
rect 6188 30046 6190 30098
rect 6242 30046 6244 30098
rect 6188 30034 6244 30046
rect 6524 30098 6580 30110
rect 6524 30046 6526 30098
rect 6578 30046 6580 30098
rect 5740 29988 5796 29998
rect 5740 29894 5796 29932
rect 6524 29876 6580 30046
rect 6524 29810 6580 29820
rect 5852 29652 5908 29662
rect 5852 29558 5908 29596
rect 5180 27858 5684 27860
rect 5180 27806 5182 27858
rect 5234 27806 5684 27858
rect 5180 27804 5684 27806
rect 5964 29538 6020 29550
rect 5964 29486 5966 29538
rect 6018 29486 6020 29538
rect 4620 27694 4622 27746
rect 4674 27694 4676 27746
rect 4620 27636 4676 27694
rect 4956 27636 5012 27646
rect 4620 27580 4900 27636
rect 4508 27570 4564 27580
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4172 27022 4174 27074
rect 4226 27022 4228 27074
rect 4172 27010 4228 27022
rect 4396 26964 4452 26974
rect 4396 26870 4452 26908
rect 4844 26962 4900 27580
rect 4956 27076 5012 27580
rect 4956 26982 5012 27020
rect 4844 26910 4846 26962
rect 4898 26910 4900 26962
rect 4844 26898 4900 26910
rect 4620 26850 4676 26862
rect 4620 26798 4622 26850
rect 4674 26798 4676 26850
rect 3276 26516 3332 26526
rect 3276 26422 3332 26460
rect 3164 26404 3220 26414
rect 3164 26310 3220 26348
rect 3500 26292 3556 26302
rect 3500 26290 3668 26292
rect 3500 26238 3502 26290
rect 3554 26238 3668 26290
rect 3500 26236 3668 26238
rect 3500 26226 3556 26236
rect 3612 25506 3668 26236
rect 4620 26180 4676 26798
rect 4732 26516 4788 26526
rect 4788 26460 4900 26516
rect 4732 26450 4788 26460
rect 4172 26124 4676 26180
rect 3612 25454 3614 25506
rect 3666 25454 3668 25506
rect 3612 25442 3668 25454
rect 4060 25508 4116 25518
rect 4172 25508 4228 26124
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4060 25506 4228 25508
rect 4060 25454 4062 25506
rect 4114 25454 4228 25506
rect 4060 25452 4228 25454
rect 4284 25508 4340 25518
rect 4060 25442 4116 25452
rect 4284 25414 4340 25452
rect 2492 25284 2548 25294
rect 2492 24834 2548 25228
rect 3836 25284 3892 25294
rect 3836 25190 3892 25228
rect 2492 24782 2494 24834
rect 2546 24782 2548 24834
rect 2492 24770 2548 24782
rect 1820 24630 1876 24668
rect 4620 24612 4676 24622
rect 4844 24612 4900 26460
rect 5180 26404 5236 27804
rect 5628 27076 5684 27086
rect 5964 27076 6020 29486
rect 6860 28644 6916 33516
rect 6972 33348 7028 33358
rect 6972 33254 7028 33292
rect 7308 31780 7364 31790
rect 6860 28550 6916 28588
rect 6972 31724 7308 31780
rect 5628 26982 5684 27020
rect 5740 27020 6020 27076
rect 6524 28418 6580 28430
rect 6524 28366 6526 28418
rect 6578 28366 6580 28418
rect 6524 27076 6580 28366
rect 5740 26962 5796 27020
rect 6524 27010 6580 27020
rect 5740 26910 5742 26962
rect 5794 26910 5796 26962
rect 4956 26292 5012 26302
rect 4956 26198 5012 26236
rect 5180 25620 5236 26348
rect 5180 25554 5236 25564
rect 5628 26852 5684 26862
rect 5628 25508 5684 26796
rect 5740 26516 5796 26910
rect 6972 26908 7028 31724
rect 7308 31686 7364 31724
rect 7084 29986 7140 29998
rect 7084 29934 7086 29986
rect 7138 29934 7140 29986
rect 7084 29876 7140 29934
rect 7420 29988 7476 43652
rect 7644 43540 7700 43550
rect 7644 43446 7700 43484
rect 9212 41298 9268 44046
rect 9436 43988 9492 44158
rect 9436 43922 9492 43932
rect 9548 44212 9604 44222
rect 9548 42978 9604 44156
rect 9548 42926 9550 42978
rect 9602 42926 9604 42978
rect 9548 42914 9604 42926
rect 9996 44100 10052 44110
rect 9996 42754 10052 44044
rect 10220 44098 10276 45054
rect 10220 44046 10222 44098
rect 10274 44046 10276 44098
rect 10220 43988 10276 44046
rect 10220 43922 10276 43932
rect 10108 43876 10164 43886
rect 10108 43708 10164 43820
rect 10108 43652 10276 43708
rect 9996 42702 9998 42754
rect 10050 42702 10052 42754
rect 9996 42690 10052 42702
rect 10220 42754 10276 43652
rect 10220 42702 10222 42754
rect 10274 42702 10276 42754
rect 10220 42690 10276 42702
rect 10332 43650 10388 46620
rect 10332 43598 10334 43650
rect 10386 43598 10388 43650
rect 10332 43540 10388 43598
rect 10108 42642 10164 42654
rect 10108 42590 10110 42642
rect 10162 42590 10164 42642
rect 10108 41748 10164 42590
rect 10332 41972 10388 43484
rect 10332 41906 10388 41916
rect 10444 43428 10500 47180
rect 10556 46004 10612 48748
rect 11340 47460 11396 49646
rect 11340 47394 11396 47404
rect 13468 49698 13524 49710
rect 13468 49646 13470 49698
rect 13522 49646 13524 49698
rect 13468 47348 13524 49646
rect 14028 48242 14084 49756
rect 14252 49746 14308 49756
rect 14364 49718 14420 49756
rect 15372 49812 15428 50372
rect 15372 49026 15428 49756
rect 16156 49138 16212 51100
rect 16156 49086 16158 49138
rect 16210 49086 16212 49138
rect 16156 49074 16212 49086
rect 18396 50372 18452 51212
rect 18844 51202 18900 51212
rect 19068 51154 19124 51166
rect 19068 51102 19070 51154
rect 19122 51102 19124 51154
rect 19068 50708 19124 51102
rect 19068 50642 19124 50652
rect 18396 49138 18452 50316
rect 19180 50594 19236 52892
rect 19404 52276 19460 52286
rect 19180 50542 19182 50594
rect 19234 50542 19236 50594
rect 19180 49700 19236 50542
rect 19292 52220 19404 52276
rect 19292 50428 19348 52220
rect 19404 52210 19460 52220
rect 19964 52276 20020 52286
rect 19740 52052 19796 52062
rect 19404 52050 19796 52052
rect 19404 51998 19742 52050
rect 19794 51998 19796 52050
rect 19404 51996 19796 51998
rect 19404 51602 19460 51996
rect 19404 51550 19406 51602
rect 19458 51550 19460 51602
rect 19404 51538 19460 51550
rect 19628 51268 19684 51996
rect 19740 51986 19796 51996
rect 19964 52050 20020 52220
rect 19964 51998 19966 52050
rect 20018 51998 20020 52050
rect 19964 51986 20020 51998
rect 20076 52274 20132 52286
rect 20076 52222 20078 52274
rect 20130 52222 20132 52274
rect 20076 51940 20132 52222
rect 20300 52276 20356 53678
rect 20412 53732 20468 54348
rect 20636 53956 20692 53966
rect 20748 53956 20804 55356
rect 21308 55186 21364 55198
rect 21308 55134 21310 55186
rect 21362 55134 21364 55186
rect 20972 54402 21028 54414
rect 20972 54350 20974 54402
rect 21026 54350 21028 54402
rect 20972 54068 21028 54350
rect 21308 54404 21364 55134
rect 21420 55076 21476 55356
rect 25788 55318 25844 55356
rect 21644 55300 21700 55310
rect 21644 55298 21812 55300
rect 21644 55246 21646 55298
rect 21698 55246 21812 55298
rect 21644 55244 21812 55246
rect 21644 55234 21700 55244
rect 21644 55076 21700 55086
rect 21420 55074 21700 55076
rect 21420 55022 21646 55074
rect 21698 55022 21700 55074
rect 21420 55020 21700 55022
rect 21644 55010 21700 55020
rect 21308 54180 21364 54348
rect 21532 54404 21588 54414
rect 21532 54402 21700 54404
rect 21532 54350 21534 54402
rect 21586 54350 21700 54402
rect 21532 54348 21700 54350
rect 21532 54338 21588 54348
rect 21308 54124 21476 54180
rect 20972 54002 21028 54012
rect 20636 53954 20804 53956
rect 20636 53902 20638 53954
rect 20690 53902 20804 53954
rect 20636 53900 20804 53902
rect 20636 53890 20692 53900
rect 20412 53666 20468 53676
rect 20524 53730 20580 53742
rect 20524 53678 20526 53730
rect 20578 53678 20580 53730
rect 20524 53508 20580 53678
rect 21420 53620 21476 54124
rect 21644 53844 21700 54348
rect 21756 53844 21812 55244
rect 21980 55298 22036 55310
rect 21980 55246 21982 55298
rect 22034 55246 22036 55298
rect 21868 54514 21924 54526
rect 21868 54462 21870 54514
rect 21922 54462 21924 54514
rect 21868 54068 21924 54462
rect 21868 54002 21924 54012
rect 21980 53844 22036 55246
rect 22988 55300 23044 55310
rect 22988 55206 23044 55244
rect 25452 55300 25508 55310
rect 22764 55188 22820 55198
rect 22764 54738 22820 55132
rect 23660 55188 23716 55198
rect 23660 55186 23828 55188
rect 23660 55134 23662 55186
rect 23714 55134 23828 55186
rect 23660 55132 23828 55134
rect 23660 55122 23716 55132
rect 22764 54686 22766 54738
rect 22818 54686 22820 54738
rect 22764 54674 22820 54686
rect 23772 54738 23828 55132
rect 23772 54686 23774 54738
rect 23826 54686 23828 54738
rect 23772 54674 23828 54686
rect 25452 54628 25508 55244
rect 26124 55188 26180 55198
rect 25452 54626 25620 54628
rect 25452 54574 25454 54626
rect 25506 54574 25620 54626
rect 25452 54572 25620 54574
rect 25452 54562 25508 54572
rect 22988 54516 23044 54526
rect 23100 54516 23156 54526
rect 22988 54514 23100 54516
rect 22988 54462 22990 54514
rect 23042 54462 23100 54514
rect 22988 54460 23100 54462
rect 22988 54450 23044 54460
rect 22316 54404 22372 54414
rect 22652 54404 22708 54414
rect 22316 54402 22708 54404
rect 22316 54350 22318 54402
rect 22370 54350 22654 54402
rect 22706 54350 22708 54402
rect 22316 54348 22708 54350
rect 22316 54338 22372 54348
rect 22652 54338 22708 54348
rect 21756 53788 21924 53844
rect 21644 53620 21700 53788
rect 21868 53732 21924 53788
rect 21980 53778 22036 53788
rect 22540 54068 22596 54078
rect 21868 53638 21924 53676
rect 22092 53732 22148 53742
rect 22092 53638 22148 53676
rect 21756 53620 21812 53630
rect 21644 53618 21812 53620
rect 21644 53566 21758 53618
rect 21810 53566 21812 53618
rect 21644 53564 21812 53566
rect 21420 53554 21476 53564
rect 21756 53554 21812 53564
rect 21308 53508 21364 53518
rect 20524 53506 21364 53508
rect 20524 53454 21310 53506
rect 21362 53454 21364 53506
rect 20524 53452 21364 53454
rect 20300 52220 20468 52276
rect 20300 52052 20356 52062
rect 20076 51884 20244 51940
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 20188 51604 20244 51884
rect 19964 51548 20244 51604
rect 19964 51378 20020 51548
rect 20300 51490 20356 51996
rect 20300 51438 20302 51490
rect 20354 51438 20356 51490
rect 20300 51426 20356 51438
rect 19964 51326 19966 51378
rect 20018 51326 20020 51378
rect 19964 51314 20020 51326
rect 20412 51380 20468 52220
rect 19628 50820 19684 51212
rect 20188 51268 20244 51278
rect 20412 51268 20468 51324
rect 20188 51266 20468 51268
rect 20188 51214 20190 51266
rect 20242 51214 20468 51266
rect 20188 51212 20468 51214
rect 20636 51378 20692 51390
rect 20636 51326 20638 51378
rect 20690 51326 20692 51378
rect 20636 51268 20692 51326
rect 21084 51380 21140 51390
rect 21084 51286 21140 51324
rect 20188 51202 20244 51212
rect 20636 51202 20692 51212
rect 19852 51154 19908 51166
rect 19852 51102 19854 51154
rect 19906 51102 19908 51154
rect 19852 51044 19908 51102
rect 20860 51156 20916 51166
rect 21196 51156 21252 51166
rect 20860 51154 21140 51156
rect 20860 51102 20862 51154
rect 20914 51102 21140 51154
rect 20860 51100 21140 51102
rect 20860 51090 20916 51100
rect 19852 50988 20132 51044
rect 19964 50820 20020 50830
rect 19628 50818 20020 50820
rect 19628 50766 19966 50818
rect 20018 50766 20020 50818
rect 19628 50764 20020 50766
rect 19964 50754 20020 50764
rect 19740 50594 19796 50606
rect 19740 50542 19742 50594
rect 19794 50542 19796 50594
rect 19740 50428 19796 50542
rect 20076 50484 20132 50988
rect 20188 50484 20244 50494
rect 20300 50484 20356 50494
rect 20076 50428 20188 50484
rect 20244 50482 20356 50484
rect 20244 50430 20302 50482
rect 20354 50430 20356 50482
rect 20244 50428 20356 50430
rect 21084 50484 21140 51100
rect 21196 51062 21252 51100
rect 21308 50708 21364 53452
rect 21308 50614 21364 50652
rect 21420 50484 21476 50494
rect 21084 50482 21476 50484
rect 21084 50430 21422 50482
rect 21474 50430 21476 50482
rect 21084 50428 21476 50430
rect 19292 50372 19796 50428
rect 19628 49924 19684 50372
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 20188 50036 20244 50428
rect 20300 50418 20356 50428
rect 21420 50418 21476 50428
rect 21980 50484 22036 50494
rect 21532 50372 21588 50382
rect 21532 50278 21588 50316
rect 20076 49980 20244 50036
rect 19628 49868 19796 49924
rect 19628 49700 19684 49710
rect 19180 49698 19684 49700
rect 19180 49646 19630 49698
rect 19682 49646 19684 49698
rect 19180 49644 19684 49646
rect 18956 49140 19012 49150
rect 18396 49086 18398 49138
rect 18450 49086 18452 49138
rect 18396 49074 18452 49086
rect 18620 49084 18956 49140
rect 15372 48974 15374 49026
rect 15426 48974 15428 49026
rect 15372 48962 15428 48974
rect 18620 48354 18676 49084
rect 18956 49074 19012 49084
rect 18620 48302 18622 48354
rect 18674 48302 18676 48354
rect 18620 48290 18676 48302
rect 14028 48190 14030 48242
rect 14082 48190 14084 48242
rect 14028 48178 14084 48190
rect 17836 48242 17892 48254
rect 17836 48190 17838 48242
rect 17890 48190 17892 48242
rect 14700 48132 14756 48142
rect 14700 48038 14756 48076
rect 15932 48132 15988 48142
rect 15932 47570 15988 48076
rect 16828 48130 16884 48142
rect 16828 48078 16830 48130
rect 16882 48078 16884 48130
rect 15932 47518 15934 47570
rect 15986 47518 15988 47570
rect 15932 47506 15988 47518
rect 16044 47684 16100 47694
rect 13468 47282 13524 47292
rect 14588 47460 14644 47470
rect 11004 47236 11060 47246
rect 11340 47236 11396 47246
rect 11060 47234 11396 47236
rect 11060 47182 11342 47234
rect 11394 47182 11396 47234
rect 11060 47180 11396 47182
rect 11004 47170 11060 47180
rect 11340 47170 11396 47180
rect 10892 46564 10948 46574
rect 10892 46562 11396 46564
rect 10892 46510 10894 46562
rect 10946 46510 11396 46562
rect 10892 46508 11396 46510
rect 10892 46498 10948 46508
rect 11340 46114 11396 46508
rect 11340 46062 11342 46114
rect 11394 46062 11396 46114
rect 11340 46050 11396 46062
rect 13020 46562 13076 46574
rect 13020 46510 13022 46562
rect 13074 46510 13076 46562
rect 10556 45948 10724 46004
rect 10556 44996 10612 45006
rect 10556 44902 10612 44940
rect 10668 44436 10724 45948
rect 11340 45890 11396 45902
rect 11340 45838 11342 45890
rect 11394 45838 11396 45890
rect 11340 45556 11396 45838
rect 12012 45890 12068 45902
rect 12012 45838 12014 45890
rect 12066 45838 12068 45890
rect 11676 45780 11732 45790
rect 11676 45686 11732 45724
rect 11340 45490 11396 45500
rect 11228 45108 11284 45118
rect 11228 45014 11284 45052
rect 12012 44996 12068 45838
rect 12236 45890 12292 45902
rect 12236 45838 12238 45890
rect 12290 45838 12292 45890
rect 12236 45108 12292 45838
rect 12572 45780 12628 45790
rect 12572 45686 12628 45724
rect 12460 45666 12516 45678
rect 12460 45614 12462 45666
rect 12514 45614 12516 45666
rect 12460 45332 12516 45614
rect 12684 45668 12740 45678
rect 12684 45574 12740 45612
rect 12460 45266 12516 45276
rect 13020 45332 13076 46510
rect 14588 46114 14644 47404
rect 16044 47458 16100 47628
rect 16044 47406 16046 47458
rect 16098 47406 16100 47458
rect 16044 47394 16100 47406
rect 16492 47460 16548 47470
rect 16716 47460 16772 47470
rect 16492 47458 16772 47460
rect 16492 47406 16494 47458
rect 16546 47406 16718 47458
rect 16770 47406 16772 47458
rect 16492 47404 16772 47406
rect 16492 47394 16548 47404
rect 16716 47394 16772 47404
rect 14924 47346 14980 47358
rect 14924 47294 14926 47346
rect 14978 47294 14980 47346
rect 14924 46562 14980 47294
rect 15260 47348 15316 47358
rect 15260 47254 15316 47292
rect 15820 47348 15876 47358
rect 15820 47254 15876 47292
rect 16268 47236 16324 47246
rect 16828 47236 16884 48078
rect 17612 47684 17668 47694
rect 17612 47590 17668 47628
rect 17052 47460 17108 47470
rect 17052 47366 17108 47404
rect 17500 47460 17556 47470
rect 16940 47236 16996 47246
rect 16828 47180 16940 47236
rect 14924 46510 14926 46562
rect 14978 46510 14980 46562
rect 14924 46498 14980 46510
rect 15036 46786 15092 46798
rect 15036 46734 15038 46786
rect 15090 46734 15092 46786
rect 14588 46062 14590 46114
rect 14642 46062 14644 46114
rect 14252 45780 14308 45790
rect 14252 45686 14308 45724
rect 13020 45266 13076 45276
rect 13244 45668 13300 45678
rect 13244 45330 13300 45612
rect 13244 45278 13246 45330
rect 13298 45278 13300 45330
rect 13244 45266 13300 45278
rect 13916 45666 13972 45678
rect 13916 45614 13918 45666
rect 13970 45614 13972 45666
rect 13916 45556 13972 45614
rect 12236 45042 12292 45052
rect 13020 45108 13076 45118
rect 13020 45014 13076 45052
rect 13356 45108 13412 45118
rect 13356 45014 13412 45052
rect 12012 44930 12068 44940
rect 10668 44322 10724 44380
rect 10668 44270 10670 44322
rect 10722 44270 10724 44322
rect 10668 44258 10724 44270
rect 11116 44882 11172 44894
rect 11116 44830 11118 44882
rect 11170 44830 11172 44882
rect 11116 44100 11172 44830
rect 11116 44034 11172 44044
rect 10108 41682 10164 41692
rect 9212 41246 9214 41298
rect 9266 41246 9268 41298
rect 9212 41234 9268 41246
rect 8428 41186 8484 41198
rect 8428 41134 8430 41186
rect 8482 41134 8484 41186
rect 8316 40516 8372 40526
rect 8316 40422 8372 40460
rect 8428 40516 8484 41134
rect 8428 39618 8484 40460
rect 9660 40628 9716 40638
rect 9660 40404 9716 40572
rect 10444 40628 10500 43372
rect 10668 43988 10724 43998
rect 10668 42642 10724 43932
rect 13580 43538 13636 43550
rect 13580 43486 13582 43538
rect 13634 43486 13636 43538
rect 13580 43428 13636 43486
rect 13580 43362 13636 43372
rect 13804 42756 13860 42766
rect 13916 42756 13972 45500
rect 14588 45444 14644 46062
rect 15036 46452 15092 46734
rect 16268 46786 16324 47180
rect 16940 47142 16996 47180
rect 17388 47236 17444 47246
rect 16268 46734 16270 46786
rect 16322 46734 16324 46786
rect 16268 46722 16324 46734
rect 14924 45892 14980 45902
rect 15036 45892 15092 46396
rect 15260 46450 15316 46462
rect 15260 46398 15262 46450
rect 15314 46398 15316 46450
rect 14924 45890 15204 45892
rect 14924 45838 14926 45890
rect 14978 45838 15204 45890
rect 14924 45836 15204 45838
rect 14924 45826 14980 45836
rect 14700 45668 14756 45678
rect 14700 45574 14756 45612
rect 14588 45388 14756 45444
rect 14364 45332 14420 45342
rect 14364 45238 14420 45276
rect 14700 45332 14756 45388
rect 14700 45266 14756 45276
rect 14588 45220 14644 45230
rect 14588 45126 14644 45164
rect 14700 45108 14756 45118
rect 14700 45014 14756 45052
rect 14812 45106 14868 45118
rect 14812 45054 14814 45106
rect 14866 45054 14868 45106
rect 14252 44436 14308 44446
rect 14812 44436 14868 45054
rect 13804 42754 13972 42756
rect 13804 42702 13806 42754
rect 13858 42702 13972 42754
rect 13804 42700 13972 42702
rect 14140 44324 14196 44334
rect 13804 42690 13860 42700
rect 10668 42590 10670 42642
rect 10722 42590 10724 42642
rect 10668 42578 10724 42590
rect 11004 42642 11060 42654
rect 11004 42590 11006 42642
rect 11058 42590 11060 42642
rect 11004 41748 11060 42590
rect 14140 42642 14196 44268
rect 14252 44322 14308 44380
rect 14252 44270 14254 44322
rect 14306 44270 14308 44322
rect 14252 44258 14308 44270
rect 14476 44380 14868 44436
rect 14364 42756 14420 42766
rect 14364 42662 14420 42700
rect 14140 42590 14142 42642
rect 14194 42590 14196 42642
rect 12684 42532 12740 42542
rect 11340 41972 11396 41982
rect 12012 41972 12068 41982
rect 11396 41916 11508 41972
rect 11340 41906 11396 41916
rect 11340 41748 11396 41758
rect 11004 41692 11340 41748
rect 11340 41298 11396 41692
rect 11340 41246 11342 41298
rect 11394 41246 11396 41298
rect 11340 41234 11396 41246
rect 10444 40562 10500 40572
rect 9660 40402 9828 40404
rect 9660 40350 9662 40402
rect 9714 40350 9828 40402
rect 9660 40348 9828 40350
rect 9660 40338 9716 40348
rect 8428 39566 8430 39618
rect 8482 39566 8484 39618
rect 8428 39554 8484 39566
rect 8988 39564 9492 39620
rect 7756 39508 7812 39518
rect 7532 39506 7812 39508
rect 7532 39454 7758 39506
rect 7810 39454 7812 39506
rect 7532 39452 7812 39454
rect 7532 39058 7588 39452
rect 7756 39442 7812 39452
rect 8876 39506 8932 39518
rect 8876 39454 8878 39506
rect 8930 39454 8932 39506
rect 7532 39006 7534 39058
rect 7586 39006 7588 39058
rect 7532 38994 7588 39006
rect 8540 39172 8596 39182
rect 7644 38834 7700 38846
rect 7644 38782 7646 38834
rect 7698 38782 7700 38834
rect 7532 38724 7588 38734
rect 7532 38050 7588 38668
rect 7644 38274 7700 38782
rect 8540 38834 8596 39116
rect 8876 39060 8932 39454
rect 8988 39506 9044 39564
rect 8988 39454 8990 39506
rect 9042 39454 9044 39506
rect 8988 39442 9044 39454
rect 9212 39396 9268 39406
rect 8876 38994 8932 39004
rect 9100 39394 9268 39396
rect 9100 39342 9214 39394
rect 9266 39342 9268 39394
rect 9100 39340 9268 39342
rect 8540 38782 8542 38834
rect 8594 38782 8596 38834
rect 8540 38770 8596 38782
rect 8764 38834 8820 38846
rect 8764 38782 8766 38834
rect 8818 38782 8820 38834
rect 8204 38724 8260 38734
rect 7644 38222 7646 38274
rect 7698 38222 7700 38274
rect 7644 38210 7700 38222
rect 7756 38612 7812 38622
rect 7532 37998 7534 38050
rect 7586 37998 7588 38050
rect 7532 37986 7588 37998
rect 7644 37828 7700 37838
rect 7756 37828 7812 38556
rect 7644 37826 7812 37828
rect 7644 37774 7646 37826
rect 7698 37774 7812 37826
rect 7644 37772 7812 37774
rect 7532 37266 7588 37278
rect 7532 37214 7534 37266
rect 7586 37214 7588 37266
rect 7532 35700 7588 37214
rect 7644 37044 7700 37772
rect 7644 36978 7700 36988
rect 7980 37042 8036 37054
rect 7980 36990 7982 37042
rect 8034 36990 8036 37042
rect 7756 35812 7812 35822
rect 7756 35718 7812 35756
rect 7868 35812 7924 35822
rect 7980 35812 8036 36990
rect 8092 37042 8148 37054
rect 8092 36990 8094 37042
rect 8146 36990 8148 37042
rect 8092 35924 8148 36990
rect 8092 35858 8148 35868
rect 7868 35810 8036 35812
rect 7868 35758 7870 35810
rect 7922 35758 8036 35810
rect 7868 35756 8036 35758
rect 8204 35810 8260 38668
rect 8764 38274 8820 38782
rect 9100 38834 9156 39340
rect 9212 39330 9268 39340
rect 9324 39396 9380 39406
rect 9436 39396 9492 39564
rect 9660 39506 9716 39518
rect 9660 39454 9662 39506
rect 9714 39454 9716 39506
rect 9548 39396 9604 39406
rect 9436 39394 9604 39396
rect 9436 39342 9550 39394
rect 9602 39342 9604 39394
rect 9436 39340 9604 39342
rect 9324 39302 9380 39340
rect 9100 38782 9102 38834
rect 9154 38782 9156 38834
rect 9100 38770 9156 38782
rect 8876 38724 8932 38734
rect 8876 38630 8932 38668
rect 9548 38722 9604 39340
rect 9548 38670 9550 38722
rect 9602 38670 9604 38722
rect 8764 38222 8766 38274
rect 8818 38222 8820 38274
rect 8764 38210 8820 38222
rect 8876 38052 8932 38062
rect 8876 37958 8932 37996
rect 8764 37828 8820 37838
rect 8204 35758 8206 35810
rect 8258 35758 8260 35810
rect 7868 35746 7924 35756
rect 7532 33572 7588 35644
rect 7756 35476 7812 35486
rect 7756 35474 8148 35476
rect 7756 35422 7758 35474
rect 7810 35422 8148 35474
rect 7756 35420 8148 35422
rect 7756 35410 7812 35420
rect 7532 33506 7588 33516
rect 7756 33234 7812 33246
rect 7756 33182 7758 33234
rect 7810 33182 7812 33234
rect 7756 31890 7812 33182
rect 7756 31838 7758 31890
rect 7810 31838 7812 31890
rect 7756 31826 7812 31838
rect 7868 31668 7924 31678
rect 7868 31574 7924 31612
rect 7644 31556 7700 31566
rect 7644 31554 7812 31556
rect 7644 31502 7646 31554
rect 7698 31502 7812 31554
rect 7644 31500 7812 31502
rect 7644 31490 7700 31500
rect 7532 31220 7588 31230
rect 7532 30994 7588 31164
rect 7756 31218 7812 31500
rect 7756 31166 7758 31218
rect 7810 31166 7812 31218
rect 7756 31154 7812 31166
rect 7532 30942 7534 30994
rect 7586 30942 7588 30994
rect 7532 30930 7588 30942
rect 7420 29922 7476 29932
rect 7868 30770 7924 30782
rect 7868 30718 7870 30770
rect 7922 30718 7924 30770
rect 7084 29810 7140 29820
rect 7756 29876 7812 29886
rect 7532 28644 7588 28654
rect 7588 28588 7700 28644
rect 7532 28578 7588 28588
rect 7644 28530 7700 28588
rect 7644 28478 7646 28530
rect 7698 28478 7700 28530
rect 7644 28466 7700 28478
rect 7756 28084 7812 29820
rect 7868 28756 7924 30718
rect 7868 28690 7924 28700
rect 7980 28532 8036 28542
rect 7980 28438 8036 28476
rect 8092 28196 8148 35420
rect 8204 34804 8260 35758
rect 8316 37826 8820 37828
rect 8316 37774 8766 37826
rect 8818 37774 8820 37826
rect 8316 37772 8820 37774
rect 8316 37266 8372 37772
rect 8764 37762 8820 37772
rect 8316 37214 8318 37266
rect 8370 37214 8372 37266
rect 8316 35922 8372 37214
rect 8540 37268 8596 37278
rect 9548 37268 9604 38670
rect 9660 38052 9716 39454
rect 9660 37986 9716 37996
rect 8540 37266 9604 37268
rect 8540 37214 8542 37266
rect 8594 37214 9604 37266
rect 8540 37212 9604 37214
rect 8540 37202 8596 37212
rect 8652 37044 8708 37054
rect 8652 36950 8708 36988
rect 8764 35980 9492 36036
rect 8316 35870 8318 35922
rect 8370 35870 8372 35922
rect 8316 35308 8372 35870
rect 8540 35924 8596 35934
rect 8764 35924 8820 35980
rect 8540 35922 8820 35924
rect 8540 35870 8542 35922
rect 8594 35870 8820 35922
rect 8540 35868 8820 35870
rect 8540 35858 8596 35868
rect 8876 35812 8932 35822
rect 8764 35700 8820 35710
rect 8764 35606 8820 35644
rect 8316 35252 8484 35308
rect 8428 35026 8484 35252
rect 8428 34974 8430 35026
rect 8482 34974 8484 35026
rect 8428 34962 8484 34974
rect 8204 34748 8596 34804
rect 8540 34354 8596 34748
rect 8540 34302 8542 34354
rect 8594 34302 8596 34354
rect 8540 34290 8596 34302
rect 8204 34132 8260 34142
rect 8764 34132 8820 34142
rect 8204 34038 8260 34076
rect 8428 34130 8820 34132
rect 8428 34078 8766 34130
rect 8818 34078 8820 34130
rect 8428 34076 8820 34078
rect 8204 31780 8260 31790
rect 8204 31686 8260 31724
rect 8204 31220 8260 31230
rect 8204 31126 8260 31164
rect 8428 30996 8484 34076
rect 8764 34066 8820 34076
rect 8876 31948 8932 35756
rect 9100 35700 9156 35710
rect 9324 35700 9380 35710
rect 9100 35698 9324 35700
rect 9100 35646 9102 35698
rect 9154 35646 9324 35698
rect 9100 35644 9324 35646
rect 9100 35634 9156 35644
rect 9324 35634 9380 35644
rect 9436 35698 9492 35980
rect 9436 35646 9438 35698
rect 9490 35646 9492 35698
rect 9436 35634 9492 35646
rect 9660 35586 9716 35598
rect 9660 35534 9662 35586
rect 9714 35534 9716 35586
rect 9660 35028 9716 35534
rect 9660 34962 9716 34972
rect 9660 34132 9716 34142
rect 9772 34132 9828 40348
rect 11452 40402 11508 41916
rect 12012 41878 12068 41916
rect 12684 41970 12740 42476
rect 13916 42532 13972 42542
rect 13916 42438 13972 42476
rect 12684 41918 12686 41970
rect 12738 41918 12740 41970
rect 12684 41906 12740 41918
rect 12796 41074 12852 41086
rect 12796 41022 12798 41074
rect 12850 41022 12852 41074
rect 12684 40964 12740 40974
rect 12124 40962 12740 40964
rect 12124 40910 12686 40962
rect 12738 40910 12740 40962
rect 12124 40908 12740 40910
rect 12124 40514 12180 40908
rect 12684 40898 12740 40908
rect 12124 40462 12126 40514
rect 12178 40462 12180 40514
rect 12124 40450 12180 40462
rect 11452 40350 11454 40402
rect 11506 40350 11508 40402
rect 11452 40338 11508 40350
rect 12796 40292 12852 41022
rect 14140 40404 14196 42590
rect 14476 42084 14532 44380
rect 14588 44268 15092 44324
rect 14588 44098 14644 44268
rect 14588 44046 14590 44098
rect 14642 44046 14644 44098
rect 14588 44034 14644 44046
rect 14700 44098 14756 44110
rect 14700 44046 14702 44098
rect 14754 44046 14756 44098
rect 14700 43652 14756 44046
rect 14812 44100 14868 44110
rect 14812 44006 14868 44044
rect 14700 43586 14756 43596
rect 14476 42018 14532 42028
rect 15036 43428 15092 44268
rect 15148 44322 15204 45836
rect 15260 45780 15316 46398
rect 16156 46452 16212 46462
rect 16156 46358 16212 46396
rect 15260 45714 15316 45724
rect 15484 45332 15540 45342
rect 15372 45108 15428 45118
rect 15372 45014 15428 45052
rect 15148 44270 15150 44322
rect 15202 44270 15204 44322
rect 15148 44258 15204 44270
rect 15484 44322 15540 45276
rect 16044 45218 16100 45230
rect 16044 45166 16046 45218
rect 16098 45166 16100 45218
rect 15820 45108 15876 45118
rect 15820 45106 15988 45108
rect 15820 45054 15822 45106
rect 15874 45054 15988 45106
rect 15820 45052 15988 45054
rect 15820 45042 15876 45052
rect 15484 44270 15486 44322
rect 15538 44270 15540 44322
rect 15484 44258 15540 44270
rect 15932 44210 15988 45052
rect 15932 44158 15934 44210
rect 15986 44158 15988 44210
rect 15932 44146 15988 44158
rect 16044 44100 16100 45166
rect 16604 45108 16660 45118
rect 16492 44994 16548 45006
rect 16492 44942 16494 44994
rect 16546 44942 16548 44994
rect 16268 44324 16324 44334
rect 16268 44230 16324 44268
rect 15372 43652 15428 43662
rect 15372 43558 15428 43596
rect 15596 43540 15652 43550
rect 15484 43538 15652 43540
rect 15484 43486 15598 43538
rect 15650 43486 15652 43538
rect 15484 43484 15652 43486
rect 15484 43428 15540 43484
rect 15596 43474 15652 43484
rect 16044 43538 16100 44044
rect 16380 43652 16436 43662
rect 16380 43558 16436 43596
rect 16044 43486 16046 43538
rect 16098 43486 16100 43538
rect 16044 43474 16100 43486
rect 15036 43372 15540 43428
rect 15820 43426 15876 43438
rect 15820 43374 15822 43426
rect 15874 43374 15876 43426
rect 14812 41860 14868 41870
rect 15036 41860 15092 43372
rect 15820 42756 15876 43374
rect 15820 42690 15876 42700
rect 15820 42084 15876 42094
rect 15372 41972 15428 41982
rect 15372 41878 15428 41916
rect 15260 41860 15316 41870
rect 14812 41858 15316 41860
rect 14812 41806 14814 41858
rect 14866 41806 15262 41858
rect 15314 41806 15316 41858
rect 14812 41804 15316 41806
rect 14812 41794 14868 41804
rect 15260 41794 15316 41804
rect 15820 41186 15876 42028
rect 16492 41298 16548 44942
rect 16604 44210 16660 45052
rect 17388 44322 17444 47180
rect 17500 46898 17556 47404
rect 17836 47236 17892 48190
rect 17948 47460 18004 47498
rect 17948 47394 18004 47404
rect 18172 47458 18228 47470
rect 18172 47406 18174 47458
rect 18226 47406 18228 47458
rect 17948 47236 18004 47246
rect 17836 47180 17948 47236
rect 17948 47170 18004 47180
rect 17500 46846 17502 46898
rect 17554 46846 17556 46898
rect 17500 46834 17556 46846
rect 18172 45668 18228 47406
rect 18620 47460 18676 47470
rect 18620 47234 18676 47404
rect 18620 47182 18622 47234
rect 18674 47182 18676 47234
rect 18620 46788 18676 47182
rect 18620 46722 18676 46732
rect 18732 46676 18788 46686
rect 18620 46116 18676 46126
rect 18620 45890 18676 46060
rect 18620 45838 18622 45890
rect 18674 45838 18676 45890
rect 18620 45826 18676 45838
rect 18284 45668 18340 45678
rect 18172 45666 18340 45668
rect 18172 45614 18286 45666
rect 18338 45614 18340 45666
rect 18172 45612 18340 45614
rect 18284 44436 18340 45612
rect 18284 44370 18340 44380
rect 17388 44270 17390 44322
rect 17442 44270 17444 44322
rect 17388 44258 17444 44270
rect 16604 44158 16606 44210
rect 16658 44158 16660 44210
rect 16604 43764 16660 44158
rect 18172 44210 18228 44222
rect 18172 44158 18174 44210
rect 18226 44158 18228 44210
rect 16604 43698 16660 43708
rect 17948 43764 18004 43774
rect 17948 43670 18004 43708
rect 17388 43652 17444 43662
rect 16492 41246 16494 41298
rect 16546 41246 16548 41298
rect 16492 41234 16548 41246
rect 16604 41746 16660 41758
rect 16604 41694 16606 41746
rect 16658 41694 16660 41746
rect 15820 41134 15822 41186
rect 15874 41134 15876 41186
rect 15260 40628 15316 40638
rect 14252 40404 14308 40414
rect 14140 40348 14252 40404
rect 12796 40226 12852 40236
rect 14252 40290 14308 40348
rect 14252 40238 14254 40290
rect 14306 40238 14308 40290
rect 14252 40226 14308 40238
rect 13468 39618 13524 39630
rect 13468 39566 13470 39618
rect 13522 39566 13524 39618
rect 11004 39172 11060 39182
rect 11004 37938 11060 39116
rect 12460 38836 12516 38846
rect 12572 38836 12628 38846
rect 12460 38834 12572 38836
rect 12460 38782 12462 38834
rect 12514 38782 12572 38834
rect 12460 38780 12572 38782
rect 12460 38770 12516 38780
rect 11676 38724 11732 38734
rect 11676 38630 11732 38668
rect 11004 37886 11006 37938
rect 11058 37886 11060 37938
rect 11004 37874 11060 37886
rect 11340 37938 11396 37950
rect 11340 37886 11342 37938
rect 11394 37886 11396 37938
rect 11340 37492 11396 37886
rect 11900 37826 11956 37838
rect 11900 37774 11902 37826
rect 11954 37774 11956 37826
rect 11676 37492 11732 37502
rect 11900 37492 11956 37774
rect 11116 37436 11676 37492
rect 11732 37436 11956 37492
rect 12348 37492 12404 37502
rect 10556 36932 10612 36942
rect 10556 35924 10612 36876
rect 10108 35922 10612 35924
rect 10108 35870 10558 35922
rect 10610 35870 10612 35922
rect 10108 35868 10612 35870
rect 10108 35810 10164 35868
rect 10556 35858 10612 35868
rect 10108 35758 10110 35810
rect 10162 35758 10164 35810
rect 10108 35746 10164 35758
rect 9884 35700 9940 35710
rect 9884 35606 9940 35644
rect 10556 35028 10612 35038
rect 10556 34934 10612 34972
rect 9716 34076 9828 34132
rect 11116 34468 11172 37436
rect 11676 37266 11732 37436
rect 11676 37214 11678 37266
rect 11730 37214 11732 37266
rect 11676 37202 11732 37214
rect 12124 37154 12180 37166
rect 12124 37102 12126 37154
rect 12178 37102 12180 37154
rect 12124 37044 12180 37102
rect 11340 35252 11396 35262
rect 11340 34914 11396 35196
rect 11340 34862 11342 34914
rect 11394 34862 11396 34914
rect 11340 34850 11396 34862
rect 11788 35252 11844 35262
rect 11116 34412 11732 34468
rect 11116 34130 11172 34412
rect 11116 34078 11118 34130
rect 11170 34078 11172 34130
rect 9660 34038 9716 34076
rect 11116 34066 11172 34078
rect 11340 34242 11396 34254
rect 11340 34190 11342 34242
rect 11394 34190 11396 34242
rect 11340 33572 11396 34190
rect 9884 33458 9940 33470
rect 9884 33406 9886 33458
rect 9938 33406 9940 33458
rect 9884 31948 9940 33406
rect 8540 31892 9940 31948
rect 11340 31948 11396 33516
rect 11676 33458 11732 34412
rect 11788 34130 11844 35196
rect 11788 34078 11790 34130
rect 11842 34078 11844 34130
rect 11788 34066 11844 34078
rect 11676 33406 11678 33458
rect 11730 33406 11732 33458
rect 11676 33394 11732 33406
rect 12124 31948 12180 36988
rect 12348 36594 12404 37436
rect 12348 36542 12350 36594
rect 12402 36542 12404 36594
rect 12348 36530 12404 36542
rect 12572 37268 12628 38780
rect 13468 38836 13524 39566
rect 14252 39508 14308 39518
rect 14252 39506 14756 39508
rect 14252 39454 14254 39506
rect 14306 39454 14756 39506
rect 14252 39452 14756 39454
rect 14252 39442 14308 39452
rect 14700 39058 14756 39452
rect 14700 39006 14702 39058
rect 14754 39006 14756 39058
rect 14700 38994 14756 39006
rect 14812 39396 14868 39406
rect 14812 38946 14868 39340
rect 14812 38894 14814 38946
rect 14866 38894 14868 38946
rect 14812 38882 14868 38894
rect 13468 38770 13524 38780
rect 15260 37492 15316 40572
rect 15820 39956 15876 41134
rect 16380 41188 16436 41198
rect 16380 41094 16436 41132
rect 16604 40628 16660 41694
rect 16604 40562 16660 40572
rect 16156 40404 16212 40414
rect 16156 40310 16212 40348
rect 16380 40402 16436 40414
rect 16380 40350 16382 40402
rect 16434 40350 16436 40402
rect 16380 40068 16436 40350
rect 16604 40404 16660 40414
rect 16604 40310 16660 40348
rect 16828 40402 16884 40414
rect 16828 40350 16830 40402
rect 16882 40350 16884 40402
rect 16492 40292 16548 40302
rect 16828 40292 16884 40350
rect 17276 40292 17332 40302
rect 16828 40236 17276 40292
rect 16492 40198 16548 40236
rect 16380 40012 16548 40068
rect 15820 39900 16436 39956
rect 16380 39732 16436 39900
rect 16492 39844 16548 40012
rect 16492 39788 16884 39844
rect 16380 39730 16772 39732
rect 16380 39678 16382 39730
rect 16434 39678 16772 39730
rect 16380 39676 16772 39678
rect 16380 39666 16436 39676
rect 16716 39618 16772 39676
rect 16716 39566 16718 39618
rect 16770 39566 16772 39618
rect 16716 39554 16772 39566
rect 16828 39508 16884 39788
rect 17164 39620 17220 39630
rect 17164 39526 17220 39564
rect 17276 39618 17332 40236
rect 17276 39566 17278 39618
rect 17330 39566 17332 39618
rect 17276 39554 17332 39566
rect 16940 39508 16996 39518
rect 16828 39452 16940 39508
rect 16940 39414 16996 39452
rect 17052 39396 17108 39406
rect 17052 39302 17108 39340
rect 17052 38612 17108 38622
rect 17052 38162 17108 38556
rect 17052 38110 17054 38162
rect 17106 38110 17108 38162
rect 17052 38098 17108 38110
rect 16380 38052 16436 38062
rect 16380 38050 16548 38052
rect 16380 37998 16382 38050
rect 16434 37998 16548 38050
rect 16380 37996 16548 37998
rect 16380 37986 16436 37996
rect 12572 35252 12628 37212
rect 15036 37436 15316 37492
rect 13244 37154 13300 37166
rect 13244 37102 13246 37154
rect 13298 37102 13300 37154
rect 13244 36260 13300 37102
rect 13244 36194 13300 36204
rect 13468 36652 13748 36708
rect 13356 35924 13412 35934
rect 13356 35830 13412 35868
rect 12572 35186 12628 35196
rect 12684 35700 12740 35710
rect 13468 35700 13524 36652
rect 13580 36482 13636 36494
rect 13580 36430 13582 36482
rect 13634 36430 13636 36482
rect 13580 35924 13636 36430
rect 13692 36482 13748 36652
rect 13692 36430 13694 36482
rect 13746 36430 13748 36482
rect 13692 36418 13748 36430
rect 14140 36482 14196 36494
rect 14140 36430 14142 36482
rect 14194 36430 14196 36482
rect 14140 36372 14196 36430
rect 13916 36316 14140 36372
rect 13804 36260 13860 36270
rect 13804 36166 13860 36204
rect 13692 35924 13748 35934
rect 13580 35922 13748 35924
rect 13580 35870 13694 35922
rect 13746 35870 13748 35922
rect 13580 35868 13748 35870
rect 13692 35858 13748 35868
rect 13804 35924 13860 35934
rect 13916 35924 13972 36316
rect 14140 36306 14196 36316
rect 13804 35922 13972 35924
rect 13804 35870 13806 35922
rect 13858 35870 13972 35922
rect 13804 35868 13972 35870
rect 14252 35924 14308 35934
rect 13804 35858 13860 35868
rect 14252 35830 14308 35868
rect 14924 35924 14980 35934
rect 13580 35700 13636 35710
rect 13468 35644 13580 35700
rect 12460 34018 12516 34030
rect 12460 33966 12462 34018
rect 12514 33966 12516 34018
rect 8540 31778 8596 31892
rect 8540 31726 8542 31778
rect 8594 31726 8596 31778
rect 8540 31714 8596 31726
rect 9996 31890 10052 31902
rect 11340 31892 11508 31948
rect 9996 31838 9998 31890
rect 10050 31838 10052 31890
rect 8652 31668 8708 31678
rect 8652 31574 8708 31612
rect 8764 31556 8820 31566
rect 8764 31554 9044 31556
rect 8764 31502 8766 31554
rect 8818 31502 9044 31554
rect 8764 31500 9044 31502
rect 8764 31490 8820 31500
rect 8540 30996 8596 31006
rect 8428 30994 8596 30996
rect 8428 30942 8542 30994
rect 8594 30942 8596 30994
rect 8428 30940 8596 30942
rect 8428 30324 8484 30334
rect 8092 28130 8148 28140
rect 8316 28530 8372 28542
rect 8316 28478 8318 28530
rect 8370 28478 8372 28530
rect 7532 28082 7812 28084
rect 7532 28030 7758 28082
rect 7810 28030 7812 28082
rect 7532 28028 7812 28030
rect 7308 27076 7364 27086
rect 7196 26964 7252 26974
rect 5740 26450 5796 26460
rect 5964 26850 6020 26862
rect 6972 26852 7140 26908
rect 7196 26870 7252 26908
rect 5964 26798 5966 26850
rect 6018 26798 6020 26850
rect 5628 25414 5684 25452
rect 5964 25506 6020 26798
rect 6636 25732 6692 25742
rect 5964 25454 5966 25506
rect 6018 25454 6020 25506
rect 5964 25442 6020 25454
rect 6300 25730 6692 25732
rect 6300 25678 6638 25730
rect 6690 25678 6692 25730
rect 6300 25676 6692 25678
rect 6300 25506 6356 25676
rect 6636 25666 6692 25676
rect 6300 25454 6302 25506
rect 6354 25454 6356 25506
rect 6300 25442 6356 25454
rect 6524 25508 6580 25518
rect 6524 25414 6580 25452
rect 6636 25396 6692 25406
rect 6636 25302 6692 25340
rect 5964 25284 6020 25294
rect 5740 25282 6020 25284
rect 5740 25230 5966 25282
rect 6018 25230 6020 25282
rect 5740 25228 6020 25230
rect 5068 25172 5124 25182
rect 5068 24724 5124 25116
rect 5740 24834 5796 25228
rect 5964 25218 6020 25228
rect 5740 24782 5742 24834
rect 5794 24782 5796 24834
rect 5740 24770 5796 24782
rect 5068 24630 5124 24668
rect 4620 24610 4900 24612
rect 4620 24558 4622 24610
rect 4674 24558 4900 24610
rect 4620 24556 4900 24558
rect 4620 24546 4676 24556
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 7084 23548 7140 26852
rect 7308 25506 7364 27020
rect 7532 27074 7588 28028
rect 7756 28018 7812 28028
rect 8316 28082 8372 28478
rect 8316 28030 8318 28082
rect 8370 28030 8372 28082
rect 8316 28018 8372 28030
rect 8428 27858 8484 30268
rect 8540 30212 8596 30940
rect 8540 30146 8596 30156
rect 8988 30100 9044 31500
rect 9996 31220 10052 31838
rect 11228 31668 11284 31678
rect 9996 31164 10612 31220
rect 9548 31108 9604 31118
rect 9548 31014 9604 31052
rect 9884 31106 9940 31118
rect 9884 31054 9886 31106
rect 9938 31054 9940 31106
rect 9884 30996 9940 31054
rect 10556 31106 10612 31164
rect 11228 31218 11284 31612
rect 11228 31166 11230 31218
rect 11282 31166 11284 31218
rect 11228 31154 11284 31166
rect 10556 31054 10558 31106
rect 10610 31054 10612 31106
rect 10444 30996 10500 31006
rect 9884 30994 10500 30996
rect 9884 30942 10446 30994
rect 10498 30942 10500 30994
rect 9884 30940 10500 30942
rect 8540 29652 8596 29662
rect 8540 28644 8596 29596
rect 8988 29650 9044 30044
rect 8988 29598 8990 29650
rect 9042 29598 9044 29650
rect 8988 29586 9044 29598
rect 9548 30212 9604 30222
rect 8652 29428 8708 29438
rect 8652 29334 8708 29372
rect 8876 28868 8932 28878
rect 8876 28866 9044 28868
rect 8876 28814 8878 28866
rect 8930 28814 9044 28866
rect 8876 28812 9044 28814
rect 8876 28802 8932 28812
rect 8652 28644 8708 28654
rect 8876 28644 8932 28654
rect 8540 28642 8708 28644
rect 8540 28590 8654 28642
rect 8706 28590 8708 28642
rect 8540 28588 8708 28590
rect 8652 28578 8708 28588
rect 8764 28642 8932 28644
rect 8764 28590 8878 28642
rect 8930 28590 8932 28642
rect 8764 28588 8932 28590
rect 8764 28420 8820 28588
rect 8876 28578 8932 28588
rect 8988 28644 9044 28812
rect 8428 27806 8430 27858
rect 8482 27806 8484 27858
rect 8428 27794 8484 27806
rect 8540 28364 8820 28420
rect 8204 27636 8260 27646
rect 8540 27636 8596 28364
rect 8764 28196 8820 28206
rect 8652 27860 8708 27870
rect 8652 27766 8708 27804
rect 8764 27858 8820 28140
rect 8764 27806 8766 27858
rect 8818 27806 8820 27858
rect 8764 27794 8820 27806
rect 8204 27634 8372 27636
rect 8204 27582 8206 27634
rect 8258 27582 8372 27634
rect 8204 27580 8372 27582
rect 8204 27570 8260 27580
rect 7532 27022 7534 27074
rect 7586 27022 7588 27074
rect 7532 27010 7588 27022
rect 7980 26964 8036 26974
rect 8204 26964 8260 26974
rect 7980 26870 8036 26908
rect 8092 26962 8260 26964
rect 8092 26910 8206 26962
rect 8258 26910 8260 26962
rect 8092 26908 8260 26910
rect 8092 26404 8148 26908
rect 8204 26898 8260 26908
rect 7308 25454 7310 25506
rect 7362 25454 7364 25506
rect 7308 25442 7364 25454
rect 7644 26348 8148 26404
rect 7644 25506 7700 26348
rect 7644 25454 7646 25506
rect 7698 25454 7700 25506
rect 7644 25442 7700 25454
rect 7980 26178 8036 26190
rect 7980 26126 7982 26178
rect 8034 26126 8036 26178
rect 7980 25506 8036 26126
rect 7980 25454 7982 25506
rect 8034 25454 8036 25506
rect 7420 25396 7476 25406
rect 7420 25302 7476 25340
rect 7868 25396 7924 25406
rect 7868 24610 7924 25340
rect 7980 25172 8036 25454
rect 8316 25396 8372 27580
rect 8540 27570 8596 27580
rect 8540 26964 8596 26974
rect 8764 26964 8820 26974
rect 8540 26962 8820 26964
rect 8540 26910 8542 26962
rect 8594 26910 8766 26962
rect 8818 26910 8820 26962
rect 8540 26908 8820 26910
rect 8540 26898 8596 26908
rect 8764 26898 8820 26908
rect 8988 26962 9044 28588
rect 9436 28532 9492 28542
rect 9100 28530 9492 28532
rect 9100 28478 9438 28530
rect 9490 28478 9492 28530
rect 9100 28476 9492 28478
rect 9100 28418 9156 28476
rect 9436 28466 9492 28476
rect 9100 28366 9102 28418
rect 9154 28366 9156 28418
rect 9100 28354 9156 28366
rect 9548 27412 9604 30156
rect 9772 28756 9828 28766
rect 9828 28700 9940 28756
rect 9772 28690 9828 28700
rect 9660 28644 9716 28654
rect 9660 28550 9716 28588
rect 9884 28642 9940 28700
rect 9884 28590 9886 28642
rect 9938 28590 9940 28642
rect 9884 28578 9940 28590
rect 10108 28644 10164 28654
rect 10108 28642 10276 28644
rect 10108 28590 10110 28642
rect 10162 28590 10276 28642
rect 10108 28588 10276 28590
rect 10108 28578 10164 28588
rect 9660 27746 9716 27758
rect 9660 27694 9662 27746
rect 9714 27694 9716 27746
rect 9660 27636 9716 27694
rect 9660 27570 9716 27580
rect 10220 27746 10276 28588
rect 10444 28532 10500 30940
rect 10556 30324 10612 31054
rect 10780 31106 10836 31118
rect 10780 31054 10782 31106
rect 10834 31054 10836 31106
rect 10780 30996 10836 31054
rect 10892 30996 10948 31006
rect 10780 30994 10948 30996
rect 10780 30942 10894 30994
rect 10946 30942 10948 30994
rect 10780 30940 10948 30942
rect 10892 30930 10948 30940
rect 11228 30994 11284 31006
rect 11228 30942 11230 30994
rect 11282 30942 11284 30994
rect 10556 30258 10612 30268
rect 11004 30212 11060 30222
rect 11228 30212 11284 30942
rect 11004 30210 11284 30212
rect 11004 30158 11006 30210
rect 11058 30158 11284 30210
rect 11004 30156 11284 30158
rect 11452 30994 11508 31892
rect 11452 30942 11454 30994
rect 11506 30942 11508 30994
rect 11004 30146 11060 30156
rect 10668 30100 10724 30110
rect 10668 30006 10724 30044
rect 10780 29986 10836 29998
rect 10780 29934 10782 29986
rect 10834 29934 10836 29986
rect 10668 28644 10724 28654
rect 10780 28644 10836 29934
rect 11340 29426 11396 29438
rect 11340 29374 11342 29426
rect 11394 29374 11396 29426
rect 11116 29316 11172 29326
rect 11004 29314 11172 29316
rect 11004 29262 11118 29314
rect 11170 29262 11172 29314
rect 11004 29260 11172 29262
rect 10724 28588 10836 28644
rect 10892 28644 10948 28654
rect 10668 28578 10724 28588
rect 10892 28550 10948 28588
rect 10556 28532 10612 28542
rect 10444 28530 10612 28532
rect 10444 28478 10558 28530
rect 10610 28478 10612 28530
rect 10444 28476 10612 28478
rect 10220 27694 10222 27746
rect 10274 27694 10276 27746
rect 10220 27636 10276 27694
rect 10220 27570 10276 27580
rect 9548 27356 9716 27412
rect 9100 27076 9156 27086
rect 9100 26982 9156 27020
rect 8988 26910 8990 26962
rect 9042 26910 9044 26962
rect 8428 26850 8484 26862
rect 8428 26798 8430 26850
rect 8482 26798 8484 26850
rect 8428 25620 8484 26798
rect 8876 26292 8932 26302
rect 8428 25554 8484 25564
rect 8764 25620 8820 25630
rect 8764 25526 8820 25564
rect 8316 25330 8372 25340
rect 7980 25106 8036 25116
rect 7868 24558 7870 24610
rect 7922 24558 7924 24610
rect 7868 24546 7924 24558
rect 8652 24164 8708 24174
rect 8652 24070 8708 24108
rect 7084 23492 7364 23548
rect 1820 23154 1876 23166
rect 1820 23102 1822 23154
rect 1874 23102 1876 23154
rect 1820 21700 1876 23102
rect 2492 23042 2548 23054
rect 2492 22990 2494 23042
rect 2546 22990 2548 23042
rect 2492 22596 2548 22990
rect 4620 23042 4676 23054
rect 4620 22990 4622 23042
rect 4674 22990 4676 23042
rect 4620 22932 4676 22990
rect 4620 22866 4676 22876
rect 5628 22932 5684 22942
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 2492 22530 2548 22540
rect 4732 22596 4788 22606
rect 4732 22502 4788 22540
rect 3388 22484 3444 22494
rect 3948 22484 4004 22494
rect 3388 22390 3444 22428
rect 3836 22428 3948 22484
rect 3612 22148 3668 22158
rect 1820 20802 1876 21644
rect 1820 20750 1822 20802
rect 1874 20750 1876 20802
rect 1820 17666 1876 20750
rect 3500 22146 3668 22148
rect 3500 22094 3614 22146
rect 3666 22094 3668 22146
rect 3500 22092 3668 22094
rect 2492 20690 2548 20702
rect 2492 20638 2494 20690
rect 2546 20638 2548 20690
rect 2492 20188 2548 20638
rect 2492 20132 3220 20188
rect 3164 19906 3220 20132
rect 3276 20132 3332 20142
rect 3500 20132 3556 22092
rect 3612 22082 3668 22092
rect 3276 20130 3556 20132
rect 3276 20078 3278 20130
rect 3330 20078 3556 20130
rect 3276 20076 3556 20078
rect 3836 20130 3892 22428
rect 3948 22390 4004 22428
rect 4956 22484 5012 22494
rect 4172 22372 4228 22382
rect 4172 22370 4340 22372
rect 4172 22318 4174 22370
rect 4226 22318 4340 22370
rect 4172 22316 4340 22318
rect 4172 22306 4228 22316
rect 4284 21028 4340 22316
rect 4844 22148 4900 22158
rect 4844 22054 4900 22092
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4060 20972 4676 21028
rect 4060 20242 4116 20972
rect 4620 20914 4676 20972
rect 4620 20862 4622 20914
rect 4674 20862 4676 20914
rect 4620 20850 4676 20862
rect 4060 20190 4062 20242
rect 4114 20190 4116 20242
rect 4060 20178 4116 20190
rect 3836 20078 3838 20130
rect 3890 20078 3892 20130
rect 3276 20066 3332 20076
rect 3164 19854 3166 19906
rect 3218 19854 3220 19906
rect 3164 19842 3220 19854
rect 3388 18676 3444 20076
rect 3836 20066 3892 20078
rect 4956 20130 5012 22428
rect 5628 22370 5684 22876
rect 5628 22318 5630 22370
rect 5682 22318 5684 22370
rect 5068 22260 5124 22270
rect 5068 22258 5572 22260
rect 5068 22206 5070 22258
rect 5122 22206 5572 22258
rect 5068 22204 5572 22206
rect 5068 22194 5124 22204
rect 5516 21364 5572 22204
rect 5628 22036 5684 22318
rect 5852 22372 5908 22382
rect 5964 22372 6020 22382
rect 5852 22370 5964 22372
rect 5852 22318 5854 22370
rect 5906 22318 5964 22370
rect 5852 22316 5964 22318
rect 5852 22306 5908 22316
rect 5628 21980 5908 22036
rect 5516 21308 5796 21364
rect 5740 20914 5796 21308
rect 5740 20862 5742 20914
rect 5794 20862 5796 20914
rect 5740 20850 5796 20862
rect 5852 20802 5908 21980
rect 5852 20750 5854 20802
rect 5906 20750 5908 20802
rect 5852 20738 5908 20750
rect 4956 20078 4958 20130
rect 5010 20078 5012 20130
rect 4956 20066 5012 20078
rect 5068 20692 5124 20702
rect 4508 20020 4564 20030
rect 4172 19964 4508 20020
rect 3948 19906 4004 19918
rect 3948 19854 3950 19906
rect 4002 19854 4004 19906
rect 3500 19796 3556 19806
rect 3948 19796 4004 19854
rect 3500 19794 4004 19796
rect 3500 19742 3502 19794
rect 3554 19742 4004 19794
rect 3500 19740 4004 19742
rect 3500 19730 3556 19740
rect 3500 18676 3556 18686
rect 3388 18674 3556 18676
rect 3388 18622 3502 18674
rect 3554 18622 3556 18674
rect 3388 18620 3556 18622
rect 2828 18452 2884 18462
rect 2828 18450 3108 18452
rect 2828 18398 2830 18450
rect 2882 18398 3108 18450
rect 2828 18396 3108 18398
rect 2828 18386 2884 18396
rect 2828 18228 2884 18238
rect 2492 18226 2884 18228
rect 2492 18174 2830 18226
rect 2882 18174 2884 18226
rect 2492 18172 2884 18174
rect 2492 17778 2548 18172
rect 2828 18162 2884 18172
rect 2492 17726 2494 17778
rect 2546 17726 2548 17778
rect 2492 17714 2548 17726
rect 1820 17614 1822 17666
rect 1874 17614 1876 17666
rect 1820 17602 1876 17614
rect 3052 17108 3108 18396
rect 3164 18340 3220 18350
rect 3164 18246 3220 18284
rect 3276 17108 3332 17118
rect 3052 17106 3332 17108
rect 3052 17054 3278 17106
rect 3330 17054 3332 17106
rect 3052 17052 3332 17054
rect 3276 15988 3332 17052
rect 3500 16772 3556 18620
rect 3724 18452 3780 18462
rect 3724 18450 4004 18452
rect 3724 18398 3726 18450
rect 3778 18398 4004 18450
rect 3724 18396 4004 18398
rect 3724 18386 3780 18396
rect 3612 18340 3668 18350
rect 3612 18246 3668 18284
rect 3948 17892 4004 18396
rect 4172 18450 4228 19964
rect 4508 19926 4564 19964
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4172 18398 4174 18450
rect 4226 18398 4228 18450
rect 4172 18386 4228 18398
rect 4508 18340 4564 18350
rect 4508 18246 4564 18284
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 3948 17836 4676 17892
rect 3836 16884 3892 16894
rect 3948 16884 4004 17836
rect 4620 17778 4676 17836
rect 4620 17726 4622 17778
rect 4674 17726 4676 17778
rect 4620 17714 4676 17726
rect 3836 16882 4004 16884
rect 3836 16830 3838 16882
rect 3890 16830 4004 16882
rect 3836 16828 4004 16830
rect 3836 16818 3892 16828
rect 3612 16772 3668 16782
rect 3500 16770 3668 16772
rect 3500 16718 3614 16770
rect 3666 16718 3668 16770
rect 3500 16716 3668 16718
rect 3612 16706 3668 16716
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 3276 15932 3668 15988
rect 3612 15316 3668 15932
rect 3836 15316 3892 15326
rect 3612 15314 3892 15316
rect 3612 15262 3838 15314
rect 3890 15262 3892 15314
rect 3612 15260 3892 15262
rect 3500 15092 3556 15102
rect 3052 15090 3556 15092
rect 3052 15038 3502 15090
rect 3554 15038 3556 15090
rect 3052 15036 3556 15038
rect 1820 14530 1876 14542
rect 1820 14478 1822 14530
rect 1874 14478 1876 14530
rect 1820 12068 1876 14478
rect 2492 14420 2548 14430
rect 2492 14418 2996 14420
rect 2492 14366 2494 14418
rect 2546 14366 2996 14418
rect 2492 14364 2996 14366
rect 2492 14354 2548 14364
rect 2940 13634 2996 14364
rect 2940 13582 2942 13634
rect 2994 13582 2996 13634
rect 2940 13570 2996 13582
rect 3052 13970 3108 15036
rect 3500 15026 3556 15036
rect 3052 13918 3054 13970
rect 3106 13918 3108 13970
rect 3052 13524 3108 13918
rect 3612 13970 3668 15260
rect 3836 15250 3892 15260
rect 4844 15314 4900 15326
rect 4844 15262 4846 15314
rect 4898 15262 4900 15314
rect 4060 15202 4116 15214
rect 4060 15150 4062 15202
rect 4114 15150 4116 15202
rect 4060 15148 4116 15150
rect 3612 13918 3614 13970
rect 3666 13918 3668 13970
rect 3612 13906 3668 13918
rect 3836 15092 4116 15148
rect 3836 13970 3892 15092
rect 4060 14644 4116 15092
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4620 14644 4676 14654
rect 4060 14642 4676 14644
rect 4060 14590 4622 14642
rect 4674 14590 4676 14642
rect 4060 14588 4676 14590
rect 4620 14578 4676 14588
rect 3836 13918 3838 13970
rect 3890 13918 3892 13970
rect 3836 13906 3892 13918
rect 4172 13972 4228 13982
rect 4172 13746 4228 13916
rect 4620 13972 4676 13982
rect 4620 13878 4676 13916
rect 4172 13694 4174 13746
rect 4226 13694 4228 13746
rect 4172 13682 4228 13694
rect 3276 13636 3332 13646
rect 3276 13542 3332 13580
rect 3724 13636 3780 13646
rect 3724 13542 3780 13580
rect 3052 13458 3108 13468
rect 3948 13524 4004 13534
rect 1820 11394 1876 12012
rect 2492 12740 2548 12750
rect 2492 11506 2548 12684
rect 2492 11454 2494 11506
rect 2546 11454 2548 11506
rect 2492 11442 2548 11454
rect 1820 11342 1822 11394
rect 1874 11342 1876 11394
rect 1820 9828 1876 11342
rect 3948 11284 4004 13468
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4508 12850 4564 12862
rect 4508 12798 4510 12850
rect 4562 12798 4564 12850
rect 4284 12740 4340 12750
rect 3948 10612 4004 11228
rect 4060 12738 4340 12740
rect 4060 12686 4286 12738
rect 4338 12686 4340 12738
rect 4060 12684 4340 12686
rect 4060 10836 4116 12684
rect 4284 12674 4340 12684
rect 4396 12740 4452 12750
rect 4396 12646 4452 12684
rect 4508 11956 4564 12798
rect 4844 12292 4900 15262
rect 5068 13972 5124 20636
rect 5628 20580 5684 20590
rect 5964 20580 6020 22316
rect 6748 22370 6804 22382
rect 6748 22318 6750 22370
rect 6802 22318 6804 22370
rect 6188 22148 6244 22158
rect 6188 22054 6244 22092
rect 6412 21700 6468 21710
rect 6748 21700 6804 22318
rect 6468 21644 6804 21700
rect 6860 22148 6916 22158
rect 6412 21606 6468 21644
rect 5628 20578 6020 20580
rect 5628 20526 5630 20578
rect 5682 20526 6020 20578
rect 5628 20524 6020 20526
rect 6300 20802 6356 20814
rect 6300 20750 6302 20802
rect 6354 20750 6356 20802
rect 5628 20514 5684 20524
rect 6300 20130 6356 20750
rect 6300 20078 6302 20130
rect 6354 20078 6356 20130
rect 6300 20020 6356 20078
rect 6636 20468 6692 20478
rect 6636 20130 6692 20412
rect 6636 20078 6638 20130
rect 6690 20078 6692 20130
rect 6636 20066 6692 20078
rect 6300 17666 6356 19964
rect 6636 19122 6692 19134
rect 6636 19070 6638 19122
rect 6690 19070 6692 19122
rect 6300 17614 6302 17666
rect 6354 17614 6356 17666
rect 6300 17602 6356 17614
rect 6412 19010 6468 19022
rect 6412 18958 6414 19010
rect 6466 18958 6468 19010
rect 6412 17556 6468 18958
rect 6524 19010 6580 19022
rect 6524 18958 6526 19010
rect 6578 18958 6580 19010
rect 6524 18564 6580 18958
rect 6636 18788 6692 19070
rect 6636 18732 6804 18788
rect 6636 18564 6692 18574
rect 6524 18562 6692 18564
rect 6524 18510 6638 18562
rect 6690 18510 6692 18562
rect 6524 18508 6692 18510
rect 6636 18498 6692 18508
rect 6636 18340 6692 18350
rect 6636 17666 6692 18284
rect 6748 17778 6804 18732
rect 6748 17726 6750 17778
rect 6802 17726 6804 17778
rect 6748 17714 6804 17726
rect 6860 18228 6916 22092
rect 7308 20692 7364 23492
rect 7420 22260 7476 22270
rect 7420 22258 7700 22260
rect 7420 22206 7422 22258
rect 7474 22206 7700 22258
rect 7420 22204 7700 22206
rect 7420 22194 7476 22204
rect 7308 20598 7364 20636
rect 7644 20690 7700 22204
rect 8876 21812 8932 26236
rect 8988 25956 9044 26910
rect 8988 25890 9044 25900
rect 8988 24164 9044 24174
rect 8988 24162 9604 24164
rect 8988 24110 8990 24162
rect 9042 24110 9604 24162
rect 8988 24108 9604 24110
rect 8988 24098 9044 24108
rect 8428 21810 8932 21812
rect 8428 21758 8878 21810
rect 8930 21758 8932 21810
rect 8428 21756 8932 21758
rect 8428 21586 8484 21756
rect 8428 21534 8430 21586
rect 8482 21534 8484 21586
rect 8428 21522 8484 21534
rect 7644 20638 7646 20690
rect 7698 20638 7700 20690
rect 7644 20626 7700 20638
rect 7980 20692 8036 20702
rect 7980 20690 8372 20692
rect 7980 20638 7982 20690
rect 8034 20638 8372 20690
rect 7980 20636 8372 20638
rect 7980 20626 8036 20636
rect 6972 20578 7028 20590
rect 6972 20526 6974 20578
rect 7026 20526 7028 20578
rect 6972 20468 7028 20526
rect 6972 20402 7028 20412
rect 8316 20132 8372 20636
rect 8652 20356 8708 21756
rect 8876 21746 8932 21756
rect 9212 23938 9268 23950
rect 9212 23886 9214 23938
rect 9266 23886 9268 23938
rect 9212 23716 9268 23886
rect 9548 23940 9604 24108
rect 9660 24162 9716 27356
rect 10556 27076 10612 28476
rect 10668 28420 10724 28430
rect 11004 28420 11060 29260
rect 11116 29250 11172 29260
rect 11340 28642 11396 29374
rect 11340 28590 11342 28642
rect 11394 28590 11396 28642
rect 11340 28578 11396 28590
rect 11452 28644 11508 30942
rect 11900 31892 12180 31948
rect 12348 33572 12404 33582
rect 12348 31948 12404 33516
rect 12460 33458 12516 33966
rect 12460 33406 12462 33458
rect 12514 33406 12516 33458
rect 12460 33394 12516 33406
rect 12684 33346 12740 35644
rect 13580 35606 13636 35644
rect 14588 35700 14644 35710
rect 12684 33294 12686 33346
rect 12738 33294 12740 33346
rect 12684 33282 12740 33294
rect 13916 35252 13972 35262
rect 13916 32564 13972 35196
rect 14588 34018 14644 35644
rect 14924 35364 14980 35868
rect 15036 35588 15092 37436
rect 15708 37380 15764 37390
rect 15148 37378 15764 37380
rect 15148 37326 15710 37378
rect 15762 37326 15764 37378
rect 15148 37324 15764 37326
rect 15148 36372 15204 37324
rect 15708 37314 15764 37324
rect 16044 37266 16100 37278
rect 16044 37214 16046 37266
rect 16098 37214 16100 37266
rect 15372 37156 15428 37166
rect 16044 37156 16100 37214
rect 15372 37154 16100 37156
rect 15372 37102 15374 37154
rect 15426 37102 16100 37154
rect 15372 37100 16100 37102
rect 15372 37090 15428 37100
rect 16044 36484 16100 37100
rect 16492 37268 16548 37996
rect 16044 36418 16100 36428
rect 16380 36594 16436 36606
rect 16380 36542 16382 36594
rect 16434 36542 16436 36594
rect 15148 35812 15204 36316
rect 15372 36260 15428 36270
rect 15148 35718 15204 35756
rect 15260 36258 15428 36260
rect 15260 36206 15374 36258
rect 15426 36206 15428 36258
rect 15260 36204 15428 36206
rect 15260 35700 15316 36204
rect 15372 36194 15428 36204
rect 15708 36258 15764 36270
rect 15708 36206 15710 36258
rect 15762 36206 15764 36258
rect 15708 36036 15764 36206
rect 15708 35980 16212 36036
rect 15372 35924 15428 35934
rect 15372 35922 16100 35924
rect 15372 35870 15374 35922
rect 15426 35870 16100 35922
rect 15372 35868 16100 35870
rect 15372 35858 15428 35868
rect 15372 35700 15428 35710
rect 15260 35698 15428 35700
rect 15260 35646 15374 35698
rect 15426 35646 15428 35698
rect 15260 35644 15428 35646
rect 15372 35588 15428 35644
rect 15036 35532 15204 35588
rect 14924 35298 14980 35308
rect 14588 33966 14590 34018
rect 14642 33966 14644 34018
rect 14588 33954 14644 33966
rect 14700 33124 14756 33134
rect 14700 32674 14756 33068
rect 14700 32622 14702 32674
rect 14754 32622 14756 32674
rect 14700 32610 14756 32622
rect 12908 32562 13972 32564
rect 12908 32510 13918 32562
rect 13970 32510 13972 32562
rect 12908 32508 13972 32510
rect 12348 31892 12516 31948
rect 11564 30324 11620 30334
rect 11564 29650 11620 30268
rect 11564 29598 11566 29650
rect 11618 29598 11620 29650
rect 11564 29586 11620 29598
rect 11676 30100 11732 30110
rect 11676 29540 11732 30044
rect 11676 29538 11844 29540
rect 11676 29486 11678 29538
rect 11730 29486 11844 29538
rect 11676 29484 11844 29486
rect 11676 29474 11732 29484
rect 11564 28644 11620 28654
rect 11452 28642 11620 28644
rect 11452 28590 11566 28642
rect 11618 28590 11620 28642
rect 11452 28588 11620 28590
rect 11564 28578 11620 28588
rect 10668 28418 11060 28420
rect 10668 28366 10670 28418
rect 10722 28366 11060 28418
rect 10668 28364 11060 28366
rect 11116 28530 11172 28542
rect 11116 28478 11118 28530
rect 11170 28478 11172 28530
rect 10668 27636 10724 28364
rect 11116 28196 11172 28478
rect 11340 28420 11396 28430
rect 11340 28326 11396 28364
rect 11116 28140 11508 28196
rect 11452 28082 11508 28140
rect 11452 28030 11454 28082
rect 11506 28030 11508 28082
rect 11452 28018 11508 28030
rect 11228 27970 11284 27982
rect 11228 27918 11230 27970
rect 11282 27918 11284 27970
rect 10668 27570 10724 27580
rect 10892 27860 10948 27870
rect 10556 27010 10612 27020
rect 9772 26292 9828 26302
rect 9772 26198 9828 26236
rect 10892 26178 10948 27804
rect 11116 27858 11172 27870
rect 11116 27806 11118 27858
rect 11170 27806 11172 27858
rect 11116 27076 11172 27806
rect 11228 27860 11284 27918
rect 11788 27970 11844 29484
rect 11900 28308 11956 31892
rect 12124 31668 12180 31678
rect 12124 31574 12180 31612
rect 12124 28756 12180 28766
rect 12124 28662 12180 28700
rect 12012 28644 12068 28654
rect 12012 28550 12068 28588
rect 12236 28642 12292 28654
rect 12236 28590 12238 28642
rect 12290 28590 12292 28642
rect 11900 28252 12068 28308
rect 11788 27918 11790 27970
rect 11842 27918 11844 27970
rect 11788 27906 11844 27918
rect 11900 27970 11956 27982
rect 11900 27918 11902 27970
rect 11954 27918 11956 27970
rect 11228 27794 11284 27804
rect 11900 27860 11956 27918
rect 11900 27794 11956 27804
rect 11116 27010 11172 27020
rect 12012 26908 12068 28252
rect 12124 28084 12180 28094
rect 12236 28084 12292 28590
rect 12460 28642 12516 31892
rect 12908 31778 12964 32508
rect 13916 32498 13972 32508
rect 12908 31726 12910 31778
rect 12962 31726 12964 31778
rect 12908 30996 12964 31726
rect 13020 30996 13076 31006
rect 12908 30994 13076 30996
rect 12908 30942 13022 30994
rect 13074 30942 13076 30994
rect 12908 30940 13076 30942
rect 13020 30930 13076 30940
rect 13804 30882 13860 30894
rect 13804 30830 13806 30882
rect 13858 30830 13860 30882
rect 13804 29652 13860 30830
rect 13804 29586 13860 29596
rect 15148 28980 15204 35532
rect 15372 35522 15428 35532
rect 15708 35698 15764 35710
rect 15708 35646 15710 35698
rect 15762 35646 15764 35698
rect 15148 28914 15204 28924
rect 15484 35364 15540 35374
rect 12460 28590 12462 28642
rect 12514 28590 12516 28642
rect 12460 28578 12516 28590
rect 12124 28082 12292 28084
rect 12124 28030 12126 28082
rect 12178 28030 12292 28082
rect 12124 28028 12292 28030
rect 13020 28420 13076 28430
rect 12124 28018 12180 28028
rect 12012 26852 12180 26908
rect 10892 26126 10894 26178
rect 10946 26126 10948 26178
rect 10892 26114 10948 26126
rect 10892 25956 10948 25966
rect 10892 25618 10948 25900
rect 10892 25566 10894 25618
rect 10946 25566 10948 25618
rect 10892 25554 10948 25566
rect 10108 24724 10164 24734
rect 9772 24612 9828 24622
rect 9772 24610 9940 24612
rect 9772 24558 9774 24610
rect 9826 24558 9940 24610
rect 9772 24556 9940 24558
rect 9772 24546 9828 24556
rect 9660 24110 9662 24162
rect 9714 24110 9716 24162
rect 9660 24098 9716 24110
rect 9772 23940 9828 23950
rect 9548 23938 9828 23940
rect 9548 23886 9774 23938
rect 9826 23886 9828 23938
rect 9548 23884 9828 23886
rect 9660 23716 9716 23726
rect 9212 23660 9660 23716
rect 8428 20132 8484 20142
rect 8316 20130 8484 20132
rect 8316 20078 8430 20130
rect 8482 20078 8484 20130
rect 8316 20076 8484 20078
rect 8428 20066 8484 20076
rect 7420 18452 7476 18462
rect 7420 18358 7476 18396
rect 7756 18340 7812 18350
rect 7756 18246 7812 18284
rect 6636 17614 6638 17666
rect 6690 17614 6692 17666
rect 6636 17602 6692 17614
rect 6860 17666 6916 18172
rect 7980 18228 8036 18238
rect 8316 18228 8372 18238
rect 7980 18134 8036 18172
rect 8092 18226 8372 18228
rect 8092 18174 8318 18226
rect 8370 18174 8372 18226
rect 8092 18172 8372 18174
rect 8092 17780 8148 18172
rect 8316 18162 8372 18172
rect 6860 17614 6862 17666
rect 6914 17614 6916 17666
rect 6860 17602 6916 17614
rect 7756 17724 8148 17780
rect 7756 17666 7812 17724
rect 7756 17614 7758 17666
rect 7810 17614 7812 17666
rect 7756 17602 7812 17614
rect 6412 17490 6468 17500
rect 6748 17556 6804 17566
rect 6748 16098 6804 17500
rect 7420 17556 7476 17566
rect 7420 17462 7476 17500
rect 7308 16156 7812 16212
rect 6748 16046 6750 16098
rect 6802 16046 6804 16098
rect 5516 15876 5572 15886
rect 5516 15426 5572 15820
rect 5516 15374 5518 15426
rect 5570 15374 5572 15426
rect 5516 15362 5572 15374
rect 6748 15428 6804 16046
rect 7196 16100 7252 16110
rect 7308 16100 7364 16156
rect 7196 16098 7364 16100
rect 7196 16046 7198 16098
rect 7250 16046 7364 16098
rect 7196 16044 7364 16046
rect 7196 16034 7252 16044
rect 7420 15988 7476 15998
rect 7420 15986 7588 15988
rect 7420 15934 7422 15986
rect 7474 15934 7588 15986
rect 7420 15932 7588 15934
rect 7420 15922 7476 15932
rect 6972 15876 7028 15886
rect 6972 15782 7028 15820
rect 6748 15362 6804 15372
rect 7420 15428 7476 15438
rect 7420 14532 7476 15372
rect 7532 14756 7588 15932
rect 7644 15202 7700 16156
rect 7756 16098 7812 16156
rect 7756 16046 7758 16098
rect 7810 16046 7812 16098
rect 7756 16034 7812 16046
rect 7980 16100 8036 16110
rect 7980 16006 8036 16044
rect 8092 16098 8148 17724
rect 8540 16100 8596 16110
rect 8092 16046 8094 16098
rect 8146 16046 8148 16098
rect 8092 16034 8148 16046
rect 8428 16044 8540 16100
rect 7980 15428 8036 15438
rect 7980 15314 8036 15372
rect 7980 15262 7982 15314
rect 8034 15262 8036 15314
rect 7980 15250 8036 15262
rect 8316 15314 8372 15326
rect 8316 15262 8318 15314
rect 8370 15262 8372 15314
rect 7644 15150 7646 15202
rect 7698 15150 7700 15202
rect 7644 15148 7700 15150
rect 8204 15204 8260 15242
rect 7644 15092 7812 15148
rect 8204 15138 8260 15148
rect 7756 14980 7812 15092
rect 8316 14980 8372 15262
rect 8428 15316 8484 16044
rect 8540 16034 8596 16044
rect 8540 15874 8596 15886
rect 8540 15822 8542 15874
rect 8594 15822 8596 15874
rect 8540 15764 8596 15822
rect 8540 15698 8596 15708
rect 8652 15540 8708 20300
rect 8988 19908 9044 19918
rect 9212 19908 9268 23660
rect 9660 23622 9716 23660
rect 9660 23380 9716 23390
rect 9772 23380 9828 23884
rect 9884 23716 9940 24556
rect 9884 23650 9940 23660
rect 9660 23378 9828 23380
rect 9660 23326 9662 23378
rect 9714 23326 9828 23378
rect 9660 23324 9828 23326
rect 9660 23314 9716 23324
rect 9548 23042 9604 23054
rect 9548 22990 9550 23042
rect 9602 22990 9604 23042
rect 9548 22482 9604 22990
rect 9548 22430 9550 22482
rect 9602 22430 9604 22482
rect 9548 22418 9604 22430
rect 10108 22370 10164 24668
rect 10780 24724 10836 24734
rect 10780 24630 10836 24668
rect 11452 24612 11508 24622
rect 11452 24518 11508 24556
rect 10220 23716 10276 23726
rect 10220 23622 10276 23660
rect 10108 22318 10110 22370
rect 10162 22318 10164 22370
rect 10108 22306 10164 22318
rect 10780 22258 10836 22270
rect 10780 22206 10782 22258
rect 10834 22206 10836 22258
rect 10780 21812 10836 22206
rect 10780 21746 10836 21756
rect 8988 19906 9268 19908
rect 8988 19854 8990 19906
rect 9042 19854 9268 19906
rect 8988 19852 9268 19854
rect 9660 20018 9716 20030
rect 9660 19966 9662 20018
rect 9714 19966 9716 20018
rect 8764 19796 8820 19806
rect 8764 19702 8820 19740
rect 8988 19012 9044 19852
rect 9212 19012 9268 19022
rect 8988 19010 9268 19012
rect 8988 18958 9214 19010
rect 9266 18958 9268 19010
rect 8988 18956 9268 18958
rect 9212 16548 9268 18956
rect 9660 18452 9716 19966
rect 10332 19908 10388 19918
rect 10332 19814 10388 19852
rect 9996 19796 10052 19806
rect 10052 19740 10164 19796
rect 9996 19730 10052 19740
rect 9660 18386 9716 18396
rect 9212 16482 9268 16492
rect 8876 16210 8932 16222
rect 8876 16158 8878 16210
rect 8930 16158 8932 16210
rect 8876 16100 8932 16158
rect 8876 16034 8932 16044
rect 9548 15764 9604 15774
rect 10108 15764 10164 19740
rect 10220 18452 10276 18462
rect 10220 16996 10276 18396
rect 11004 18340 11060 18350
rect 11004 18246 11060 18284
rect 10220 16994 10388 16996
rect 10220 16942 10222 16994
rect 10274 16942 10388 16994
rect 10220 16940 10388 16942
rect 10220 16930 10276 16940
rect 10332 16100 10388 16940
rect 9604 15708 9716 15764
rect 10108 15708 10276 15764
rect 9548 15698 9604 15708
rect 8652 15484 8820 15540
rect 8540 15316 8596 15326
rect 8428 15314 8596 15316
rect 8428 15262 8542 15314
rect 8594 15262 8596 15314
rect 8428 15260 8596 15262
rect 8540 15250 8596 15260
rect 7756 14924 8372 14980
rect 7532 14700 7700 14756
rect 7644 14642 7700 14700
rect 7644 14590 7646 14642
rect 7698 14590 7700 14642
rect 7644 14578 7700 14590
rect 7532 14532 7588 14542
rect 7420 14530 7588 14532
rect 7420 14478 7534 14530
rect 7586 14478 7588 14530
rect 7420 14476 7588 14478
rect 7532 14466 7588 14476
rect 7756 14530 7812 14924
rect 7756 14478 7758 14530
rect 7810 14478 7812 14530
rect 7756 14466 7812 14478
rect 8204 14530 8260 14542
rect 8204 14478 8206 14530
rect 8258 14478 8260 14530
rect 5068 13906 5124 13916
rect 6636 13972 6692 13982
rect 4844 12226 4900 12236
rect 6300 12962 6356 12974
rect 6300 12910 6302 12962
rect 6354 12910 6356 12962
rect 6300 12292 6356 12910
rect 6300 12198 6356 12236
rect 4508 11900 4900 11956
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4620 11506 4676 11518
rect 4620 11454 4622 11506
rect 4674 11454 4676 11506
rect 4620 11396 4676 11454
rect 4844 11508 4900 11900
rect 4844 11442 4900 11452
rect 5740 11508 5796 11518
rect 6636 11508 6692 13916
rect 5740 11414 5796 11452
rect 6300 11506 6692 11508
rect 6300 11454 6638 11506
rect 6690 11454 6692 11506
rect 6300 11452 6692 11454
rect 5852 11396 5908 11406
rect 4676 11340 4788 11396
rect 4620 11330 4676 11340
rect 4172 10836 4228 10846
rect 4060 10780 4172 10836
rect 4172 10742 4228 10780
rect 4508 10612 4564 10622
rect 3948 10610 4564 10612
rect 3948 10558 4510 10610
rect 4562 10558 4564 10610
rect 3948 10556 4564 10558
rect 4508 10546 4564 10556
rect 4732 10610 4788 11340
rect 5852 11302 5908 11340
rect 6300 11394 6356 11452
rect 6300 11342 6302 11394
rect 6354 11342 6356 11394
rect 5628 11284 5684 11294
rect 5628 11190 5684 11228
rect 5516 10836 5572 10846
rect 5572 10780 5908 10836
rect 5516 10742 5572 10780
rect 4732 10558 4734 10610
rect 4786 10558 4788 10610
rect 4732 10546 4788 10558
rect 5628 10612 5684 10622
rect 5628 10518 5684 10556
rect 5740 10610 5796 10622
rect 5740 10558 5742 10610
rect 5794 10558 5796 10610
rect 5740 10500 5796 10558
rect 5740 10434 5796 10444
rect 5628 10276 5684 10286
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 5068 9940 5124 9950
rect 5628 9940 5684 10220
rect 5068 9938 5684 9940
rect 5068 9886 5070 9938
rect 5122 9886 5630 9938
rect 5682 9886 5684 9938
rect 5068 9884 5684 9886
rect 5068 9874 5124 9884
rect 5628 9874 5684 9884
rect 2156 9828 2212 9838
rect 1820 9826 2212 9828
rect 1820 9774 2158 9826
rect 2210 9774 2212 9826
rect 1820 9772 2212 9774
rect 2156 9762 2212 9772
rect 5852 9826 5908 10780
rect 5852 9774 5854 9826
rect 5906 9774 5908 9826
rect 5852 9762 5908 9774
rect 5964 10612 6020 10622
rect 2940 9714 2996 9726
rect 2940 9662 2942 9714
rect 2994 9662 2996 9714
rect 2940 9268 2996 9662
rect 2940 9202 2996 9212
rect 5964 9154 6020 10556
rect 6188 10612 6244 10622
rect 6300 10612 6356 11342
rect 6636 10834 6692 11452
rect 7084 12850 7140 12862
rect 7084 12798 7086 12850
rect 7138 12798 7140 12850
rect 7084 11508 7140 12798
rect 8204 12628 8260 14478
rect 8204 12562 8260 12572
rect 7084 11442 7140 11452
rect 8316 12404 8372 12414
rect 8316 11394 8372 12348
rect 8652 12180 8708 12190
rect 8428 11508 8484 11518
rect 8428 11414 8484 11452
rect 8316 11342 8318 11394
rect 8370 11342 8372 11394
rect 8316 11330 8372 11342
rect 8652 11394 8708 12124
rect 8652 11342 8654 11394
rect 8706 11342 8708 11394
rect 8652 11330 8708 11342
rect 8764 12178 8820 15484
rect 9660 15314 9716 15708
rect 10108 15540 10164 15550
rect 9660 15262 9662 15314
rect 9714 15262 9716 15314
rect 8764 12126 8766 12178
rect 8818 12126 8820 12178
rect 8764 11172 8820 12126
rect 9212 13074 9268 13086
rect 9660 13076 9716 15262
rect 9996 15428 10052 15438
rect 9996 15314 10052 15372
rect 10108 15426 10164 15484
rect 10108 15374 10110 15426
rect 10162 15374 10164 15426
rect 10108 15362 10164 15374
rect 9996 15262 9998 15314
rect 10050 15262 10052 15314
rect 9996 15250 10052 15262
rect 9772 15204 9828 15242
rect 9772 15138 9828 15148
rect 9212 13022 9214 13074
rect 9266 13022 9268 13074
rect 9212 12180 9268 13022
rect 9436 13020 10052 13076
rect 9436 12404 9492 13020
rect 9996 12962 10052 13020
rect 9996 12910 9998 12962
rect 10050 12910 10052 12962
rect 9996 12898 10052 12910
rect 10220 12964 10276 15708
rect 10332 13746 10388 16044
rect 11676 16100 11732 16110
rect 11676 16006 11732 16044
rect 11004 15986 11060 15998
rect 11004 15934 11006 15986
rect 11058 15934 11060 15986
rect 11004 15540 11060 15934
rect 11004 15474 11060 15484
rect 10556 15428 10612 15438
rect 10556 15334 10612 15372
rect 11116 15204 11172 15214
rect 11116 13858 11172 15148
rect 11116 13806 11118 13858
rect 11170 13806 11172 13858
rect 11116 13794 11172 13806
rect 10332 13694 10334 13746
rect 10386 13694 10388 13746
rect 10332 13682 10388 13694
rect 10332 12964 10388 12974
rect 10220 12962 10388 12964
rect 10220 12910 10334 12962
rect 10386 12910 10388 12962
rect 10220 12908 10388 12910
rect 10108 12850 10164 12862
rect 10108 12798 10110 12850
rect 10162 12798 10164 12850
rect 9548 12740 9604 12750
rect 9548 12738 9940 12740
rect 9548 12686 9550 12738
rect 9602 12686 9940 12738
rect 9548 12684 9940 12686
rect 9548 12674 9604 12684
rect 9548 12404 9604 12414
rect 9492 12402 9604 12404
rect 9492 12350 9550 12402
rect 9602 12350 9604 12402
rect 9492 12348 9604 12350
rect 9436 12310 9492 12348
rect 9548 12338 9604 12348
rect 9212 12114 9268 12124
rect 9772 12180 9828 12190
rect 9772 12086 9828 12124
rect 9660 12066 9716 12078
rect 9660 12014 9662 12066
rect 9714 12014 9716 12066
rect 8988 11618 9044 11630
rect 8988 11566 8990 11618
rect 9042 11566 9044 11618
rect 8876 11396 8932 11406
rect 8988 11396 9044 11566
rect 9660 11618 9716 12014
rect 9660 11566 9662 11618
rect 9714 11566 9716 11618
rect 9660 11554 9716 11566
rect 8876 11394 9044 11396
rect 8876 11342 8878 11394
rect 8930 11342 9044 11394
rect 8876 11340 9044 11342
rect 8876 11330 8932 11340
rect 8764 11106 8820 11116
rect 9324 11172 9380 11182
rect 9324 11078 9380 11116
rect 6636 10782 6638 10834
rect 6690 10782 6692 10834
rect 6636 10770 6692 10782
rect 6188 10610 6356 10612
rect 6188 10558 6190 10610
rect 6242 10558 6356 10610
rect 6188 10556 6356 10558
rect 6188 10546 6244 10556
rect 7308 9938 7364 9950
rect 7308 9886 7310 9938
rect 7362 9886 7364 9938
rect 6860 9826 6916 9838
rect 6860 9774 6862 9826
rect 6914 9774 6916 9826
rect 6188 9716 6244 9726
rect 6188 9622 6244 9660
rect 6860 9716 6916 9774
rect 6916 9660 7252 9716
rect 6860 9650 6916 9660
rect 6636 9602 6692 9614
rect 6636 9550 6638 9602
rect 6690 9550 6692 9602
rect 6076 9268 6132 9278
rect 6076 9174 6132 9212
rect 5964 9102 5966 9154
rect 6018 9102 6020 9154
rect 5964 9090 6020 9102
rect 6300 9044 6356 9054
rect 6300 8950 6356 8988
rect 6636 9044 6692 9550
rect 7196 9154 7252 9660
rect 7196 9102 7198 9154
rect 7250 9102 7252 9154
rect 7196 9090 7252 9102
rect 7308 9266 7364 9886
rect 9436 9716 9492 9726
rect 7308 9214 7310 9266
rect 7362 9214 7364 9266
rect 7308 9156 7364 9214
rect 8652 9714 9492 9716
rect 8652 9662 9438 9714
rect 9490 9662 9492 9714
rect 8652 9660 9492 9662
rect 8652 9266 8708 9660
rect 9436 9650 9492 9660
rect 9660 9268 9716 9278
rect 8652 9214 8654 9266
rect 8706 9214 8708 9266
rect 8652 9202 8708 9214
rect 8988 9266 9716 9268
rect 8988 9214 9662 9266
rect 9714 9214 9716 9266
rect 8988 9212 9716 9214
rect 7308 9090 7364 9100
rect 8764 9156 8820 9166
rect 6636 8978 6692 8988
rect 8428 9044 8484 9054
rect 8428 8950 8484 8988
rect 7308 8818 7364 8830
rect 7308 8766 7310 8818
rect 7362 8766 7364 8818
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 5964 7476 6020 7486
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 5964 6802 6020 7420
rect 7308 7474 7364 8766
rect 8652 8372 8708 8382
rect 8652 8278 8708 8316
rect 7308 7422 7310 7474
rect 7362 7422 7364 7474
rect 7308 7410 7364 7422
rect 7756 8148 7812 8158
rect 7756 7476 7812 8092
rect 8764 8146 8820 9100
rect 8988 9154 9044 9212
rect 9660 9202 9716 9212
rect 8988 9102 8990 9154
rect 9042 9102 9044 9154
rect 8988 9090 9044 9102
rect 9772 9156 9828 9166
rect 9772 9062 9828 9100
rect 9212 9044 9268 9054
rect 9212 8932 9268 8988
rect 9548 9042 9604 9054
rect 9548 8990 9550 9042
rect 9602 8990 9604 9042
rect 9548 8932 9604 8990
rect 9212 8876 9604 8932
rect 9212 8258 9268 8876
rect 9884 8820 9940 12684
rect 10108 12404 10164 12798
rect 9996 12348 10164 12404
rect 10220 12628 10276 12638
rect 9996 12180 10052 12348
rect 9996 12114 10052 12124
rect 10220 12178 10276 12572
rect 10220 12126 10222 12178
rect 10274 12126 10276 12178
rect 10220 12114 10276 12126
rect 10332 11844 10388 12908
rect 10108 11394 10164 11406
rect 10108 11342 10110 11394
rect 10162 11342 10164 11394
rect 10108 9826 10164 11342
rect 10108 9774 10110 9826
rect 10162 9774 10164 9826
rect 10108 9716 10164 9774
rect 10108 9650 10164 9660
rect 10220 9268 10276 9278
rect 10220 9042 10276 9212
rect 10220 8990 10222 9042
rect 10274 8990 10276 9042
rect 10220 8978 10276 8990
rect 9212 8206 9214 8258
rect 9266 8206 9268 8258
rect 9212 8194 9268 8206
rect 9324 8764 9940 8820
rect 8764 8094 8766 8146
rect 8818 8094 8820 8146
rect 8764 8082 8820 8094
rect 8988 8148 9044 8158
rect 8988 8054 9044 8092
rect 7756 7382 7812 7420
rect 5964 6750 5966 6802
rect 6018 6750 6020 6802
rect 5964 6738 6020 6750
rect 8204 7362 8260 7374
rect 8204 7310 8206 7362
rect 8258 7310 8260 7362
rect 8092 6580 8148 6590
rect 7980 6578 8148 6580
rect 7980 6526 8094 6578
rect 8146 6526 8148 6578
rect 7980 6524 8148 6526
rect 7980 6130 8036 6524
rect 8092 6514 8148 6524
rect 7980 6078 7982 6130
rect 8034 6078 8036 6130
rect 7980 6066 8036 6078
rect 7868 6020 7924 6030
rect 7868 5926 7924 5964
rect 8092 6020 8148 6030
rect 8204 6020 8260 7310
rect 8876 6692 8932 6702
rect 8876 6598 8932 6636
rect 8092 6018 8260 6020
rect 8092 5966 8094 6018
rect 8146 5966 8260 6018
rect 8092 5964 8260 5966
rect 8540 6020 8596 6030
rect 8092 5954 8148 5964
rect 8540 5926 8596 5964
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 9324 5122 9380 8764
rect 10332 8372 10388 11788
rect 10780 12068 10836 12078
rect 10780 11506 10836 12012
rect 10780 11454 10782 11506
rect 10834 11454 10836 11506
rect 10780 11442 10836 11454
rect 10668 9268 10724 9278
rect 12124 9268 12180 26852
rect 13020 26402 13076 28364
rect 13020 26350 13022 26402
rect 13074 26350 13076 26402
rect 13020 26338 13076 26350
rect 13916 27858 13972 27870
rect 13916 27806 13918 27858
rect 13970 27806 13972 27858
rect 13804 26292 13860 26302
rect 13916 26292 13972 27806
rect 14700 27748 14756 27758
rect 14700 27654 14756 27692
rect 13804 26290 13972 26292
rect 13804 26238 13806 26290
rect 13858 26238 13972 26290
rect 13804 26236 13972 26238
rect 13804 26226 13860 26236
rect 13916 25394 13972 26236
rect 13916 25342 13918 25394
rect 13970 25342 13972 25394
rect 13916 24724 13972 25342
rect 13916 24630 13972 24668
rect 15036 24724 15092 24734
rect 15092 24668 15316 24724
rect 15036 24658 15092 24668
rect 12348 24612 12404 24622
rect 12348 24162 12404 24556
rect 13580 24612 13636 24622
rect 14700 24612 14756 24622
rect 13580 24610 13860 24612
rect 13580 24558 13582 24610
rect 13634 24558 13860 24610
rect 13580 24556 13860 24558
rect 13580 24546 13636 24556
rect 12348 24110 12350 24162
rect 12402 24110 12404 24162
rect 12348 24098 12404 24110
rect 13804 24052 13860 24556
rect 14700 24518 14756 24556
rect 13804 23996 14308 24052
rect 12348 23938 12404 23950
rect 12348 23886 12350 23938
rect 12402 23886 12404 23938
rect 12348 22932 12404 23886
rect 12684 23828 12740 23838
rect 12684 23734 12740 23772
rect 13916 23156 13972 23996
rect 14252 23938 14308 23996
rect 14252 23886 14254 23938
rect 14306 23886 14308 23938
rect 14252 23874 14308 23886
rect 14588 23940 14644 23950
rect 14588 23846 14644 23884
rect 15036 23940 15092 23950
rect 14140 23828 14196 23838
rect 14140 23734 14196 23772
rect 14028 23714 14084 23726
rect 14028 23662 14030 23714
rect 14082 23662 14084 23714
rect 14028 23380 14084 23662
rect 15036 23714 15092 23884
rect 15036 23662 15038 23714
rect 15090 23662 15092 23714
rect 14028 23324 14196 23380
rect 14028 23156 14084 23166
rect 13916 23154 14084 23156
rect 13916 23102 14030 23154
rect 14082 23102 14084 23154
rect 13916 23100 14084 23102
rect 14028 23090 14084 23100
rect 12348 22372 12404 22876
rect 13468 22932 13524 22942
rect 13468 22838 13524 22876
rect 13804 22932 13860 22942
rect 13804 22838 13860 22876
rect 14140 22932 14196 23324
rect 14140 22866 14196 22876
rect 12908 22484 12964 22494
rect 12908 22482 13412 22484
rect 12908 22430 12910 22482
rect 12962 22430 13412 22482
rect 12908 22428 13412 22430
rect 12908 22418 12964 22428
rect 12348 22306 12404 22316
rect 12796 21812 12852 21822
rect 13356 21812 13412 22428
rect 13468 21812 13524 21822
rect 13356 21756 13468 21812
rect 12796 21718 12852 21756
rect 13468 21718 13524 21756
rect 14700 21812 14756 21822
rect 12684 21698 12740 21710
rect 12684 21646 12686 21698
rect 12738 21646 12740 21698
rect 12684 20804 12740 21646
rect 13244 21588 13300 21598
rect 13244 21494 13300 21532
rect 13916 21586 13972 21598
rect 13916 21534 13918 21586
rect 13970 21534 13972 21586
rect 13356 21474 13412 21486
rect 13356 21422 13358 21474
rect 13410 21422 13412 21474
rect 12908 21364 12964 21374
rect 13356 21364 13412 21422
rect 12908 21362 13412 21364
rect 12908 21310 12910 21362
rect 12962 21310 13412 21362
rect 12908 21308 13412 21310
rect 12908 21298 12964 21308
rect 12684 20738 12740 20748
rect 13132 20804 13188 20814
rect 12908 20580 12964 20590
rect 12908 20020 12964 20524
rect 12460 20018 12964 20020
rect 12460 19966 12910 20018
rect 12962 19966 12964 20018
rect 12460 19964 12964 19966
rect 12460 19906 12516 19964
rect 12908 19954 12964 19964
rect 13132 20018 13188 20748
rect 13468 20804 13524 20814
rect 13468 20710 13524 20748
rect 13580 20804 13636 20814
rect 13580 20802 13860 20804
rect 13580 20750 13582 20802
rect 13634 20750 13860 20802
rect 13580 20748 13860 20750
rect 13580 20738 13636 20748
rect 13692 20580 13748 20590
rect 13692 20486 13748 20524
rect 13580 20356 13636 20366
rect 13636 20300 13748 20356
rect 13580 20290 13636 20300
rect 13580 20132 13636 20142
rect 13132 19966 13134 20018
rect 13186 19966 13188 20018
rect 13132 19954 13188 19966
rect 13468 20020 13524 20030
rect 13580 20020 13636 20076
rect 13468 20018 13636 20020
rect 13468 19966 13470 20018
rect 13522 19966 13636 20018
rect 13468 19964 13636 19966
rect 12460 19854 12462 19906
rect 12514 19854 12516 19906
rect 12460 19842 12516 19854
rect 13468 19234 13524 19964
rect 13692 19572 13748 20300
rect 13804 20130 13860 20748
rect 13916 20692 13972 21534
rect 14476 21588 14532 21598
rect 14476 21494 14532 21532
rect 14700 21586 14756 21756
rect 14700 21534 14702 21586
rect 14754 21534 14756 21586
rect 14700 21522 14756 21534
rect 14140 21362 14196 21374
rect 14140 21310 14142 21362
rect 14194 21310 14196 21362
rect 14140 20804 14196 21310
rect 14140 20738 14196 20748
rect 13916 20690 14084 20692
rect 13916 20638 13918 20690
rect 13970 20638 14084 20690
rect 13916 20636 14084 20638
rect 13916 20626 13972 20636
rect 14028 20356 14084 20636
rect 14028 20300 14196 20356
rect 13804 20078 13806 20130
rect 13858 20078 13860 20130
rect 13804 20066 13860 20078
rect 14028 20132 14084 20142
rect 14028 20038 14084 20076
rect 13916 19908 13972 19918
rect 13916 19814 13972 19852
rect 13692 19516 13860 19572
rect 13468 19182 13470 19234
rect 13522 19182 13524 19234
rect 13468 18676 13524 19182
rect 13580 19012 13636 19022
rect 13580 18918 13636 18956
rect 13692 19010 13748 19022
rect 13692 18958 13694 19010
rect 13746 18958 13748 19010
rect 13468 18620 13636 18676
rect 13468 18452 13524 18462
rect 13132 18396 13468 18452
rect 13132 18338 13188 18396
rect 13468 18358 13524 18396
rect 13132 18286 13134 18338
rect 13186 18286 13188 18338
rect 13132 18274 13188 18286
rect 13580 18228 13636 18620
rect 13692 18452 13748 18958
rect 13692 18386 13748 18396
rect 13692 18228 13748 18238
rect 13580 18226 13748 18228
rect 13580 18174 13694 18226
rect 13746 18174 13748 18226
rect 13580 18172 13748 18174
rect 13692 18162 13748 18172
rect 13804 16884 13860 19516
rect 14140 19234 14196 20300
rect 14924 19348 14980 19358
rect 14924 19254 14980 19292
rect 14140 19182 14142 19234
rect 14194 19182 14196 19234
rect 14028 18452 14084 18462
rect 14028 18358 14084 18396
rect 14140 18228 14196 19182
rect 14252 19012 14308 19022
rect 14308 18956 14420 19012
rect 14252 18946 14308 18956
rect 14364 18562 14420 18956
rect 14364 18510 14366 18562
rect 14418 18510 14420 18562
rect 14364 18498 14420 18510
rect 14700 18452 14756 18490
rect 14700 18386 14756 18396
rect 14476 18340 14532 18350
rect 14476 18246 14532 18284
rect 15036 18228 15092 23662
rect 15260 22370 15316 24668
rect 15260 22318 15262 22370
rect 15314 22318 15316 22370
rect 15260 22306 15316 22318
rect 14140 17554 14196 18172
rect 14700 18172 15092 18228
rect 15148 20468 15204 20478
rect 14364 17668 14420 17678
rect 14140 17502 14142 17554
rect 14194 17502 14196 17554
rect 14140 17490 14196 17502
rect 14252 17666 14420 17668
rect 14252 17614 14366 17666
rect 14418 17614 14420 17666
rect 14252 17612 14420 17614
rect 13804 16790 13860 16828
rect 13804 16100 13860 16110
rect 14252 16100 14308 17612
rect 14364 17602 14420 17612
rect 14700 16212 14756 18172
rect 15036 17556 15092 17566
rect 15148 17556 15204 20412
rect 15036 17554 15204 17556
rect 15036 17502 15038 17554
rect 15090 17502 15204 17554
rect 15036 17500 15204 17502
rect 15036 17490 15092 17500
rect 15148 17108 15204 17500
rect 15148 17042 15204 17052
rect 15372 17554 15428 17566
rect 15372 17502 15374 17554
rect 15426 17502 15428 17554
rect 15260 16884 15316 16894
rect 15260 16790 15316 16828
rect 14700 16118 14756 16156
rect 14812 16660 14868 16670
rect 14476 16100 14532 16110
rect 13804 16098 14476 16100
rect 13804 16046 13806 16098
rect 13858 16046 14254 16098
rect 14306 16046 14476 16098
rect 13804 16044 14476 16046
rect 13804 16034 13860 16044
rect 14252 16034 14308 16044
rect 13468 15874 13524 15886
rect 13468 15822 13470 15874
rect 13522 15822 13524 15874
rect 13244 15314 13300 15326
rect 13244 15262 13246 15314
rect 13298 15262 13300 15314
rect 13244 14532 13300 15262
rect 13356 15204 13412 15242
rect 13356 15138 13412 15148
rect 13244 14466 13300 14476
rect 13468 14530 13524 15822
rect 14476 15538 14532 16044
rect 14476 15486 14478 15538
rect 14530 15486 14532 15538
rect 14476 15474 14532 15486
rect 14812 15426 14868 16604
rect 15372 16660 15428 17502
rect 15372 16594 15428 16604
rect 15484 16212 15540 35308
rect 15708 35252 15764 35646
rect 15708 35186 15764 35196
rect 16044 34692 16100 35868
rect 16156 35700 16212 35980
rect 16268 35812 16324 35822
rect 16268 35718 16324 35756
rect 16156 35606 16212 35644
rect 16380 35698 16436 36542
rect 16380 35646 16382 35698
rect 16434 35646 16436 35698
rect 16380 35252 16436 35646
rect 16380 34804 16436 35196
rect 16492 35026 16548 37212
rect 16604 36484 16660 36494
rect 16604 36390 16660 36428
rect 16716 36482 16772 36494
rect 16716 36430 16718 36482
rect 16770 36430 16772 36482
rect 16716 35700 16772 36430
rect 16716 35634 16772 35644
rect 16492 34974 16494 35026
rect 16546 34974 16548 35026
rect 16492 34962 16548 34974
rect 16828 35474 16884 35486
rect 16828 35422 16830 35474
rect 16882 35422 16884 35474
rect 16380 34748 16548 34804
rect 16044 34636 16324 34692
rect 16268 34130 16324 34636
rect 16268 34078 16270 34130
rect 16322 34078 16324 34130
rect 16268 34066 16324 34078
rect 16380 34354 16436 34366
rect 16380 34302 16382 34354
rect 16434 34302 16436 34354
rect 16380 34132 16436 34302
rect 16380 34066 16436 34076
rect 15708 34018 15764 34030
rect 15708 33966 15710 34018
rect 15762 33966 15764 34018
rect 15708 33908 15764 33966
rect 16492 34020 16548 34748
rect 16828 34244 16884 35422
rect 17388 34916 17444 43596
rect 18060 43538 18116 43550
rect 18060 43486 18062 43538
rect 18114 43486 18116 43538
rect 17500 41298 17556 41310
rect 17500 41246 17502 41298
rect 17554 41246 17556 41298
rect 17500 41188 17556 41246
rect 17500 41122 17556 41132
rect 17612 41300 17668 41310
rect 17500 40628 17556 40638
rect 17612 40628 17668 41244
rect 17500 40626 17668 40628
rect 17500 40574 17502 40626
rect 17554 40574 17668 40626
rect 17500 40572 17668 40574
rect 17500 40404 17556 40572
rect 17500 40338 17556 40348
rect 18060 40068 18116 43486
rect 18172 40292 18228 44158
rect 18732 43652 18788 46620
rect 19628 46676 19684 49644
rect 19740 48804 19796 49868
rect 19964 49140 20020 49150
rect 19964 49046 20020 49084
rect 20076 49028 20132 49980
rect 20076 48972 20244 49028
rect 19740 48738 19796 48748
rect 20076 48804 20132 48842
rect 20076 48738 20132 48748
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 20188 48468 20244 48972
rect 21980 49026 22036 50428
rect 22540 50428 22596 54012
rect 22876 53732 22932 53742
rect 22876 53638 22932 53676
rect 22988 53508 23044 53518
rect 22988 53414 23044 53452
rect 22652 52836 22708 52846
rect 22652 50594 22708 52780
rect 22764 52164 22820 52174
rect 22988 52164 23044 52174
rect 22764 52162 22988 52164
rect 22764 52110 22766 52162
rect 22818 52110 22988 52162
rect 22764 52108 22988 52110
rect 22764 52098 22820 52108
rect 22988 52070 23044 52108
rect 23100 51716 23156 54460
rect 23548 54516 23604 54526
rect 23548 54422 23604 54460
rect 24780 54404 24836 54414
rect 23884 54290 23940 54302
rect 23884 54238 23886 54290
rect 23938 54238 23940 54290
rect 23884 53732 23940 54238
rect 23884 53666 23940 53676
rect 24668 52948 24724 52958
rect 24780 52948 24836 54348
rect 25228 53732 25284 53742
rect 25228 53638 25284 53676
rect 24724 52892 24836 52948
rect 25452 53508 25508 53518
rect 24668 52854 24724 52892
rect 23996 52164 24052 52174
rect 23996 52070 24052 52108
rect 24556 52164 24612 52174
rect 24556 52070 24612 52108
rect 23324 51938 23380 51950
rect 23324 51886 23326 51938
rect 23378 51886 23380 51938
rect 23324 51716 23380 51886
rect 23660 51940 23716 51950
rect 23660 51938 23828 51940
rect 23660 51886 23662 51938
rect 23714 51886 23828 51938
rect 23660 51884 23828 51886
rect 23660 51874 23716 51884
rect 22876 51660 23380 51716
rect 22764 51266 22820 51278
rect 22764 51214 22766 51266
rect 22818 51214 22820 51266
rect 22764 50708 22820 51214
rect 22764 50642 22820 50652
rect 22652 50542 22654 50594
rect 22706 50542 22708 50594
rect 22652 50530 22708 50542
rect 22540 50372 22708 50428
rect 21980 48974 21982 49026
rect 22034 48974 22036 49026
rect 21980 48962 22036 48974
rect 20300 48916 20356 48926
rect 20748 48916 20804 48926
rect 20300 48914 20580 48916
rect 20300 48862 20302 48914
rect 20354 48862 20580 48914
rect 20300 48860 20580 48862
rect 20300 48850 20356 48860
rect 20076 48412 20244 48468
rect 20076 47570 20132 48412
rect 20076 47518 20078 47570
rect 20130 47518 20132 47570
rect 20076 47506 20132 47518
rect 20524 47570 20580 48860
rect 20748 48130 20804 48860
rect 21644 48916 21700 48926
rect 21644 48822 21700 48860
rect 22092 48916 22148 48926
rect 22092 48822 22148 48860
rect 21420 48804 21476 48814
rect 20748 48078 20750 48130
rect 20802 48078 20804 48130
rect 20748 48066 20804 48078
rect 21196 48242 21252 48254
rect 21196 48190 21198 48242
rect 21250 48190 21252 48242
rect 20524 47518 20526 47570
rect 20578 47518 20580 47570
rect 20524 47506 20580 47518
rect 19964 47460 20020 47470
rect 19964 47366 20020 47404
rect 20188 47236 20244 47246
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 20188 46786 20244 47180
rect 21196 47236 21252 48190
rect 21420 47458 21476 48748
rect 21420 47406 21422 47458
rect 21474 47406 21476 47458
rect 21420 47394 21476 47406
rect 21532 48802 21588 48814
rect 22316 48804 22372 48814
rect 21532 48750 21534 48802
rect 21586 48750 21588 48802
rect 21532 47460 21588 48750
rect 22204 48802 22372 48804
rect 22204 48750 22318 48802
rect 22370 48750 22372 48802
rect 22204 48748 22372 48750
rect 21196 47170 21252 47180
rect 21532 47124 21588 47404
rect 21532 47058 21588 47068
rect 21644 48468 21700 48478
rect 20188 46734 20190 46786
rect 20242 46734 20244 46786
rect 20188 46722 20244 46734
rect 19628 46610 19684 46620
rect 21420 46116 21476 46126
rect 21308 46060 21420 46116
rect 19516 45780 19572 45790
rect 19516 45330 19572 45724
rect 20412 45666 20468 45678
rect 20412 45614 20414 45666
rect 20466 45614 20468 45666
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 19516 45278 19518 45330
rect 19570 45278 19572 45330
rect 19516 45266 19572 45278
rect 20412 45220 20468 45614
rect 20636 45220 20692 45230
rect 21196 45220 21252 45230
rect 20300 45218 21252 45220
rect 20300 45166 20638 45218
rect 20690 45166 21198 45218
rect 21250 45166 21252 45218
rect 20300 45164 21252 45166
rect 20076 44996 20132 45006
rect 20300 44996 20356 45164
rect 20636 45154 20692 45164
rect 21196 45154 21252 45164
rect 20076 44994 20356 44996
rect 20076 44942 20078 44994
rect 20130 44942 20356 44994
rect 20076 44940 20356 44942
rect 20748 44996 20804 45006
rect 21308 44996 21364 46060
rect 21420 46050 21476 46060
rect 21644 45890 21700 48412
rect 21980 48132 22036 48142
rect 21868 48130 22036 48132
rect 21868 48078 21982 48130
rect 22034 48078 22036 48130
rect 21868 48076 22036 48078
rect 21868 47570 21924 48076
rect 21980 48066 22036 48076
rect 21868 47518 21870 47570
rect 21922 47518 21924 47570
rect 21868 47506 21924 47518
rect 21756 47458 21812 47470
rect 21756 47406 21758 47458
rect 21810 47406 21812 47458
rect 21756 47236 21812 47406
rect 22092 47460 22148 47470
rect 22204 47460 22260 48748
rect 22316 48738 22372 48748
rect 22540 48468 22596 48478
rect 22092 47458 22260 47460
rect 22092 47406 22094 47458
rect 22146 47406 22260 47458
rect 22092 47404 22260 47406
rect 22316 47458 22372 47470
rect 22316 47406 22318 47458
rect 22370 47406 22372 47458
rect 22092 47394 22148 47404
rect 21756 47170 21812 47180
rect 21644 45838 21646 45890
rect 21698 45838 21700 45890
rect 21644 45826 21700 45838
rect 21756 46002 21812 46014
rect 21756 45950 21758 46002
rect 21810 45950 21812 46002
rect 21756 45892 21812 45950
rect 21756 45826 21812 45836
rect 21980 45780 22036 45790
rect 22316 45780 22372 47406
rect 22540 47346 22596 48412
rect 22540 47294 22542 47346
rect 22594 47294 22596 47346
rect 22540 47282 22596 47294
rect 22652 46900 22708 50372
rect 22876 48804 22932 51660
rect 23660 51492 23716 51502
rect 23436 51490 23716 51492
rect 23436 51438 23662 51490
rect 23714 51438 23716 51490
rect 23436 51436 23716 51438
rect 22988 51380 23044 51390
rect 22988 51286 23044 51324
rect 23324 51268 23380 51278
rect 23324 51174 23380 51212
rect 23436 50706 23492 51436
rect 23660 51426 23716 51436
rect 23772 51380 23828 51884
rect 23772 51314 23828 51324
rect 23996 51378 24052 51390
rect 23996 51326 23998 51378
rect 24050 51326 24052 51378
rect 23996 51268 24052 51326
rect 23996 51202 24052 51212
rect 23436 50654 23438 50706
rect 23490 50654 23492 50706
rect 23436 50642 23492 50654
rect 22876 48738 22932 48748
rect 23324 50372 23380 50382
rect 23324 47458 23380 50316
rect 24556 49812 24612 49822
rect 24556 48466 24612 49756
rect 24556 48414 24558 48466
rect 24610 48414 24612 48466
rect 24556 48402 24612 48414
rect 25340 49700 25396 49710
rect 25340 48466 25396 49644
rect 25452 48692 25508 53452
rect 25564 52164 25620 54572
rect 26124 53842 26180 55132
rect 26684 55188 26740 56030
rect 26684 55122 26740 55132
rect 26908 55074 26964 55086
rect 26908 55022 26910 55074
rect 26962 55022 26964 55074
rect 26908 54292 26964 55022
rect 27020 54740 27076 56254
rect 37436 56308 37492 59200
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 52444 56420 52500 59200
rect 52444 56364 52948 56420
rect 37660 56308 37716 56318
rect 37436 56306 37716 56308
rect 37436 56254 37438 56306
rect 37490 56254 37662 56306
rect 37714 56254 37716 56306
rect 37436 56252 37716 56254
rect 37436 56242 37492 56252
rect 37660 56242 37716 56252
rect 52444 56306 52500 56364
rect 52444 56254 52446 56306
rect 52498 56254 52500 56306
rect 52444 56242 52500 56254
rect 52668 56194 52724 56206
rect 52668 56142 52670 56194
rect 52722 56142 52724 56194
rect 27132 56082 27188 56094
rect 27132 56030 27134 56082
rect 27186 56030 27188 56082
rect 27132 55412 27188 56030
rect 27356 56082 27412 56094
rect 27356 56030 27358 56082
rect 27410 56030 27412 56082
rect 27356 55412 27412 56030
rect 38220 55972 38276 55982
rect 38220 55970 38388 55972
rect 38220 55918 38222 55970
rect 38274 55918 38388 55970
rect 38220 55916 38388 55918
rect 38220 55906 38276 55916
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 27356 55356 27636 55412
rect 27132 55346 27188 55356
rect 27580 55300 27636 55356
rect 29148 55410 29204 55422
rect 29148 55358 29150 55410
rect 29202 55358 29204 55410
rect 27692 55300 27748 55310
rect 27580 55298 27748 55300
rect 27580 55246 27694 55298
rect 27746 55246 27748 55298
rect 27580 55244 27748 55246
rect 27356 55186 27412 55198
rect 27356 55134 27358 55186
rect 27410 55134 27412 55186
rect 27356 55076 27412 55134
rect 27356 55010 27412 55020
rect 27468 55188 27524 55198
rect 27468 54740 27524 55132
rect 27692 55076 27748 55244
rect 27692 55020 28420 55076
rect 27020 54684 27188 54740
rect 26908 54236 27076 54292
rect 26908 54068 26964 54078
rect 26908 53956 26964 54012
rect 26124 53790 26126 53842
rect 26178 53790 26180 53842
rect 26124 53778 26180 53790
rect 26572 53954 26964 53956
rect 26572 53902 26910 53954
rect 26962 53902 26964 53954
rect 26572 53900 26964 53902
rect 25900 53732 25956 53742
rect 25900 53730 26068 53732
rect 25900 53678 25902 53730
rect 25954 53678 26068 53730
rect 25900 53676 26068 53678
rect 25900 53666 25956 53676
rect 26012 53284 26068 53676
rect 26348 53620 26404 53630
rect 26012 53228 26292 53284
rect 26236 53170 26292 53228
rect 26236 53118 26238 53170
rect 26290 53118 26292 53170
rect 25676 52164 25732 52174
rect 25564 52162 25732 52164
rect 25564 52110 25678 52162
rect 25730 52110 25732 52162
rect 25564 52108 25732 52110
rect 25676 52098 25732 52108
rect 25788 52164 25844 52174
rect 25788 51268 25844 52108
rect 26124 51378 26180 51390
rect 26124 51326 26126 51378
rect 26178 51326 26180 51378
rect 26124 51268 26180 51326
rect 25788 51266 26180 51268
rect 25788 51214 25790 51266
rect 25842 51214 26180 51266
rect 25788 51212 26180 51214
rect 25788 51202 25844 51212
rect 25564 50706 25620 50718
rect 25564 50654 25566 50706
rect 25618 50654 25620 50706
rect 25564 50484 25620 50654
rect 25900 50484 25956 50494
rect 25564 50428 25900 50484
rect 25900 50034 25956 50428
rect 25900 49982 25902 50034
rect 25954 49982 25956 50034
rect 25900 49970 25956 49982
rect 25676 49812 25732 49822
rect 25676 49718 25732 49756
rect 25788 49698 25844 49710
rect 25788 49646 25790 49698
rect 25842 49646 25844 49698
rect 25788 49364 25844 49646
rect 25900 49364 25956 49374
rect 25788 49308 25900 49364
rect 25900 49298 25956 49308
rect 25452 48636 25844 48692
rect 25340 48414 25342 48466
rect 25394 48414 25396 48466
rect 25340 48402 25396 48414
rect 23324 47406 23326 47458
rect 23378 47406 23380 47458
rect 23100 47348 23156 47358
rect 22652 46834 22708 46844
rect 22876 47236 22932 47246
rect 20748 44994 21364 44996
rect 20748 44942 20750 44994
rect 20802 44942 21364 44994
rect 20748 44940 21364 44942
rect 21868 45778 22372 45780
rect 21868 45726 21982 45778
rect 22034 45726 22372 45778
rect 21868 45724 22372 45726
rect 22652 45890 22708 45902
rect 22652 45838 22654 45890
rect 22706 45838 22708 45890
rect 20076 44930 20132 44940
rect 19852 44884 19908 44894
rect 19852 44790 19908 44828
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 18732 42866 18788 43596
rect 18732 42814 18734 42866
rect 18786 42814 18788 42866
rect 18732 42802 18788 42814
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 18620 41858 18676 41870
rect 18620 41806 18622 41858
rect 18674 41806 18676 41858
rect 18508 41188 18564 41198
rect 18508 40514 18564 41132
rect 18620 40628 18676 41806
rect 18732 41748 18788 41758
rect 18732 41746 19684 41748
rect 18732 41694 18734 41746
rect 18786 41694 19684 41746
rect 18732 41692 19684 41694
rect 18732 41682 18788 41692
rect 19628 41298 19684 41692
rect 19628 41246 19630 41298
rect 19682 41246 19684 41298
rect 19628 41234 19684 41246
rect 19852 41412 19908 41422
rect 19852 40964 19908 41356
rect 19628 40908 19908 40964
rect 18844 40628 18900 40638
rect 18620 40626 18900 40628
rect 18620 40574 18846 40626
rect 18898 40574 18900 40626
rect 18620 40572 18900 40574
rect 18844 40562 18900 40572
rect 18956 40628 19012 40638
rect 18956 40534 19012 40572
rect 19628 40628 19684 40908
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19628 40534 19684 40572
rect 18508 40462 18510 40514
rect 18562 40462 18564 40514
rect 18508 40450 18564 40462
rect 18732 40404 18788 40414
rect 18732 40402 18900 40404
rect 18732 40350 18734 40402
rect 18786 40350 18900 40402
rect 18732 40348 18900 40350
rect 18732 40338 18788 40348
rect 18172 40226 18228 40236
rect 18620 40292 18676 40302
rect 18060 40012 18564 40068
rect 17836 39620 17892 39630
rect 17836 39526 17892 39564
rect 18508 38946 18564 40012
rect 18620 39508 18676 40236
rect 18732 39508 18788 39518
rect 18620 39506 18788 39508
rect 18620 39454 18734 39506
rect 18786 39454 18788 39506
rect 18620 39452 18788 39454
rect 18732 39442 18788 39452
rect 18844 39508 18900 40348
rect 19068 40402 19124 40414
rect 19068 40350 19070 40402
rect 19122 40350 19124 40402
rect 19068 40292 19124 40350
rect 19068 40226 19124 40236
rect 18844 39284 18900 39452
rect 18508 38894 18510 38946
rect 18562 38894 18564 38946
rect 18508 38836 18564 38894
rect 18508 38770 18564 38780
rect 18732 39228 18900 39284
rect 19068 39394 19124 39406
rect 19068 39342 19070 39394
rect 19122 39342 19124 39394
rect 18732 38834 18788 39228
rect 19068 39060 19124 39342
rect 19628 39394 19684 39406
rect 19628 39342 19630 39394
rect 19682 39342 19684 39394
rect 19628 39060 19684 39342
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19068 39058 19684 39060
rect 19068 39006 19070 39058
rect 19122 39006 19630 39058
rect 19682 39006 19684 39058
rect 19068 39004 19684 39006
rect 19068 38994 19124 39004
rect 18732 38782 18734 38834
rect 18786 38782 18788 38834
rect 18060 38724 18116 38762
rect 18060 38658 18116 38668
rect 17948 38612 18004 38622
rect 17948 38518 18004 38556
rect 18732 37380 18788 38782
rect 18956 38834 19012 38846
rect 18956 38782 18958 38834
rect 19010 38782 19012 38834
rect 18844 38724 18900 38762
rect 18956 38724 19012 38782
rect 19180 38836 19236 38846
rect 19068 38724 19124 38734
rect 18956 38668 19068 38724
rect 18844 38658 18900 38668
rect 19068 38658 19124 38668
rect 19180 38162 19236 38780
rect 19180 38110 19182 38162
rect 19234 38110 19236 38162
rect 19180 38098 19236 38110
rect 18956 37380 19012 37390
rect 18732 37378 19012 37380
rect 18732 37326 18958 37378
rect 19010 37326 19012 37378
rect 18732 37324 19012 37326
rect 18956 37314 19012 37324
rect 19516 37268 19572 37278
rect 19628 37268 19684 39004
rect 20076 38724 20132 38762
rect 20076 38658 20132 38668
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20188 37380 20244 44940
rect 20748 44930 20804 44940
rect 20412 44884 20468 44894
rect 20300 44436 20356 44446
rect 20412 44436 20468 44828
rect 20300 44434 20468 44436
rect 20300 44382 20302 44434
rect 20354 44382 20468 44434
rect 20300 44380 20468 44382
rect 20300 44370 20356 44380
rect 21420 43428 21476 43438
rect 21420 42866 21476 43372
rect 21420 42814 21422 42866
rect 21474 42814 21476 42866
rect 20748 42756 20804 42766
rect 20748 42662 20804 42700
rect 21420 42756 21476 42814
rect 21420 42690 21476 42700
rect 21196 42532 21252 42542
rect 20412 41970 20468 41982
rect 20412 41918 20414 41970
rect 20466 41918 20468 41970
rect 20412 41186 20468 41918
rect 21196 41970 21252 42476
rect 21196 41918 21198 41970
rect 21250 41918 21252 41970
rect 21196 41906 21252 41918
rect 20412 41134 20414 41186
rect 20466 41134 20468 41186
rect 20412 40180 20468 41134
rect 20412 38834 20468 40124
rect 20860 40402 20916 40414
rect 20860 40350 20862 40402
rect 20914 40350 20916 40402
rect 20860 40180 20916 40350
rect 20860 40114 20916 40124
rect 21532 40290 21588 40302
rect 21532 40238 21534 40290
rect 21586 40238 21588 40290
rect 21532 39844 21588 40238
rect 21532 39778 21588 39788
rect 21868 39396 21924 45724
rect 21980 45714 22036 45724
rect 22652 45108 22708 45838
rect 22876 45108 22932 47180
rect 23100 47068 23156 47292
rect 22988 47012 23156 47068
rect 23212 47124 23268 47134
rect 22988 45220 23044 47012
rect 23212 45778 23268 47068
rect 23212 45726 23214 45778
rect 23266 45726 23268 45778
rect 23212 45332 23268 45726
rect 23324 45556 23380 47406
rect 24108 48130 24164 48142
rect 24108 48078 24110 48130
rect 24162 48078 24164 48130
rect 24108 47460 24164 48078
rect 24444 48130 24500 48142
rect 24444 48078 24446 48130
rect 24498 48078 24500 48130
rect 24220 47460 24276 47470
rect 24108 47458 24276 47460
rect 24108 47406 24222 47458
rect 24274 47406 24276 47458
rect 24108 47404 24276 47406
rect 24220 47394 24276 47404
rect 23436 47234 23492 47246
rect 23436 47182 23438 47234
rect 23490 47182 23492 47234
rect 23436 45780 23492 47182
rect 23436 45714 23492 45724
rect 23660 47234 23716 47246
rect 23660 47182 23662 47234
rect 23714 47182 23716 47234
rect 23436 45556 23492 45566
rect 23324 45500 23436 45556
rect 23436 45490 23492 45500
rect 23212 45276 23604 45332
rect 22988 45164 23156 45220
rect 22092 42642 22148 42654
rect 22092 42590 22094 42642
rect 22146 42590 22148 42642
rect 21980 42532 22036 42542
rect 21980 42438 22036 42476
rect 22092 41972 22148 42590
rect 22092 41906 22148 41916
rect 22316 39844 22372 39854
rect 22316 39750 22372 39788
rect 22428 39732 22484 39742
rect 22428 39638 22484 39676
rect 21980 39396 22036 39406
rect 21868 39340 21980 39396
rect 21980 39330 22036 39340
rect 20412 38782 20414 38834
rect 20466 38782 20468 38834
rect 20412 38770 20468 38782
rect 21196 38722 21252 38734
rect 21196 38670 21198 38722
rect 21250 38670 21252 38722
rect 21196 38164 21252 38670
rect 21196 38098 21252 38108
rect 20748 37380 20804 37390
rect 20076 37324 20244 37380
rect 20524 37378 20804 37380
rect 20524 37326 20750 37378
rect 20802 37326 20804 37378
rect 20524 37324 20804 37326
rect 19740 37268 19796 37278
rect 19628 37266 19796 37268
rect 19628 37214 19742 37266
rect 19794 37214 19796 37266
rect 19628 37212 19796 37214
rect 19516 37174 19572 37212
rect 19740 37156 19796 37212
rect 19740 37090 19796 37100
rect 20076 36482 20132 37324
rect 20524 37268 20580 37324
rect 20748 37314 20804 37324
rect 22652 37380 22708 45052
rect 22764 45106 22932 45108
rect 22764 45054 22878 45106
rect 22930 45054 22932 45106
rect 22764 45052 22932 45054
rect 22764 44100 22820 45052
rect 22876 45042 22932 45052
rect 22988 44994 23044 45006
rect 22988 44942 22990 44994
rect 23042 44942 23044 44994
rect 22876 44546 22932 44558
rect 22876 44494 22878 44546
rect 22930 44494 22932 44546
rect 22876 44324 22932 44494
rect 22876 44258 22932 44268
rect 22988 44322 23044 44942
rect 22988 44270 22990 44322
rect 23042 44270 23044 44322
rect 22876 44100 22932 44110
rect 22764 44098 22932 44100
rect 22764 44046 22878 44098
rect 22930 44046 22932 44098
rect 22764 44044 22932 44046
rect 22876 44034 22932 44044
rect 22988 38724 23044 44270
rect 23100 38948 23156 45164
rect 23548 45106 23604 45276
rect 23660 45220 23716 47182
rect 24108 47236 24164 47246
rect 24108 47142 24164 47180
rect 24332 46676 24388 46686
rect 24332 46582 24388 46620
rect 24108 45892 24164 45902
rect 24108 45798 24164 45836
rect 23660 45154 23716 45164
rect 23548 45054 23550 45106
rect 23602 45054 23604 45106
rect 23548 45042 23604 45054
rect 23772 45108 23828 45118
rect 23772 45014 23828 45052
rect 23436 44994 23492 45006
rect 23436 44942 23438 44994
rect 23490 44942 23492 44994
rect 23436 44322 23492 44942
rect 23436 44270 23438 44322
rect 23490 44270 23492 44322
rect 23436 44258 23492 44270
rect 23772 43652 23828 43662
rect 23772 41970 23828 43596
rect 24444 42980 24500 48078
rect 25228 48132 25284 48142
rect 25228 48130 25508 48132
rect 25228 48078 25230 48130
rect 25282 48078 25508 48130
rect 25228 48076 25508 48078
rect 25228 48066 25284 48076
rect 25228 46676 25284 46686
rect 24556 45778 24612 45790
rect 24556 45726 24558 45778
rect 24610 45726 24612 45778
rect 24556 44322 24612 45726
rect 24556 44270 24558 44322
rect 24610 44270 24612 44322
rect 24556 44258 24612 44270
rect 24220 42924 24500 42980
rect 25116 43316 25172 43326
rect 24220 42196 24276 42924
rect 25116 42866 25172 43260
rect 25116 42814 25118 42866
rect 25170 42814 25172 42866
rect 25116 42802 25172 42814
rect 24332 42754 24388 42766
rect 24332 42702 24334 42754
rect 24386 42702 24388 42754
rect 24332 42644 24388 42702
rect 24332 42588 24612 42644
rect 24220 42140 24388 42196
rect 24108 42082 24164 42094
rect 24108 42030 24110 42082
rect 24162 42030 24164 42082
rect 23772 41918 23774 41970
rect 23826 41918 23828 41970
rect 23324 41860 23380 41870
rect 23324 41766 23380 41804
rect 23772 41860 23828 41918
rect 23772 41794 23828 41804
rect 23884 41970 23940 41982
rect 23884 41918 23886 41970
rect 23938 41918 23940 41970
rect 23884 41748 23940 41918
rect 23996 41972 24052 41982
rect 23996 41878 24052 41916
rect 23884 41682 23940 41692
rect 24108 41412 24164 42030
rect 24220 41972 24276 41982
rect 24220 41878 24276 41916
rect 24108 41346 24164 41356
rect 24332 41188 24388 42140
rect 24108 41132 24388 41188
rect 24444 41748 24500 41758
rect 24108 40404 24164 41132
rect 24220 40628 24276 40638
rect 24444 40628 24500 41692
rect 24220 40626 24500 40628
rect 24220 40574 24222 40626
rect 24274 40574 24500 40626
rect 24220 40572 24500 40574
rect 24220 40562 24276 40572
rect 23660 40402 24164 40404
rect 23660 40350 24110 40402
rect 24162 40350 24164 40402
rect 23660 40348 24164 40350
rect 23660 40290 23716 40348
rect 24108 40338 24164 40348
rect 24444 40402 24500 40414
rect 24444 40350 24446 40402
rect 24498 40350 24500 40402
rect 23660 40238 23662 40290
rect 23714 40238 23716 40290
rect 23660 40226 23716 40238
rect 24332 40290 24388 40302
rect 24332 40238 24334 40290
rect 24386 40238 24388 40290
rect 24332 39732 24388 40238
rect 24332 39666 24388 39676
rect 24444 40292 24500 40350
rect 23100 38882 23156 38892
rect 23884 39620 23940 39630
rect 23324 38724 23380 38734
rect 22988 38722 23380 38724
rect 22988 38670 23326 38722
rect 23378 38670 23380 38722
rect 22988 38668 23380 38670
rect 22988 38050 23044 38668
rect 23324 38658 23380 38668
rect 23436 38724 23492 38734
rect 23436 38052 23492 38668
rect 23660 38164 23716 38174
rect 23660 38070 23716 38108
rect 22988 37998 22990 38050
rect 23042 37998 23044 38050
rect 22988 37986 23044 37998
rect 23212 37996 23492 38052
rect 22764 37826 22820 37838
rect 23100 37828 23156 37838
rect 22764 37774 22766 37826
rect 22818 37774 22820 37826
rect 22764 37604 22820 37774
rect 22988 37826 23156 37828
rect 22988 37774 23102 37826
rect 23154 37774 23156 37826
rect 22988 37772 23156 37774
rect 22988 37604 23044 37772
rect 23100 37762 23156 37772
rect 22764 37548 23044 37604
rect 22876 37380 22932 37390
rect 22652 37378 22932 37380
rect 22652 37326 22878 37378
rect 22930 37326 22932 37378
rect 22652 37324 22932 37326
rect 22540 37268 22596 37278
rect 20188 37156 20244 37166
rect 20188 36820 20244 37100
rect 20188 36764 20468 36820
rect 20076 36430 20078 36482
rect 20130 36430 20132 36482
rect 17500 36258 17556 36270
rect 17500 36206 17502 36258
rect 17554 36206 17556 36258
rect 17500 35812 17556 36206
rect 20076 36260 20132 36430
rect 20076 36194 20132 36204
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 17500 35746 17556 35756
rect 19964 35698 20020 35710
rect 19964 35646 19966 35698
rect 20018 35646 20020 35698
rect 17388 34822 17444 34860
rect 19180 34916 19236 34926
rect 19180 34822 19236 34860
rect 19964 34692 20020 35646
rect 19964 34636 20244 34692
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 16492 33954 16548 33964
rect 16604 34188 16884 34244
rect 16044 33908 16100 33918
rect 15708 33852 16044 33908
rect 16044 33814 16100 33852
rect 16380 33906 16436 33918
rect 16380 33854 16382 33906
rect 16434 33854 16436 33906
rect 16380 33796 16436 33854
rect 16604 33796 16660 34188
rect 16380 33740 16660 33796
rect 16604 33234 16660 33246
rect 16604 33182 16606 33234
rect 16658 33182 16660 33234
rect 16380 33122 16436 33134
rect 16380 33070 16382 33122
rect 16434 33070 16436 33122
rect 16380 32788 16436 33070
rect 16492 33124 16548 33134
rect 16492 33030 16548 33068
rect 16604 32788 16660 33182
rect 16156 32732 16380 32788
rect 15932 30882 15988 30894
rect 15932 30830 15934 30882
rect 15986 30830 15988 30882
rect 15932 30212 15988 30830
rect 16156 30434 16212 32732
rect 16380 32722 16436 32732
rect 16492 32732 16660 32788
rect 16828 33012 16884 34188
rect 19516 34132 19572 34142
rect 20188 34132 20244 34636
rect 20412 34244 20468 36764
rect 20524 36482 20580 37212
rect 22428 37212 22540 37268
rect 20524 36430 20526 36482
rect 20578 36430 20580 36482
rect 20524 34468 20580 36430
rect 20636 37156 20692 37166
rect 20636 35810 20692 37100
rect 22428 36484 22484 37212
rect 22540 37174 22596 37212
rect 21980 36428 22484 36484
rect 20636 35758 20638 35810
rect 20690 35758 20692 35810
rect 20636 35746 20692 35758
rect 21196 36260 21252 36270
rect 21420 36260 21476 36270
rect 21252 36258 21476 36260
rect 21252 36206 21422 36258
rect 21474 36206 21476 36258
rect 21252 36204 21476 36206
rect 20860 34916 20916 34926
rect 20524 34412 20692 34468
rect 20524 34244 20580 34254
rect 20412 34188 20524 34244
rect 20524 34178 20580 34188
rect 20300 34132 20356 34142
rect 20188 34076 20300 34132
rect 19516 34038 19572 34076
rect 20300 34038 20356 34076
rect 17388 34020 17444 34030
rect 17388 33926 17444 33964
rect 19516 33908 19572 33918
rect 16828 32956 17780 33012
rect 16492 31892 16548 32732
rect 16828 32676 16884 32956
rect 16492 31826 16548 31836
rect 16604 32620 16884 32676
rect 17388 32788 17444 32798
rect 16604 31668 16660 32620
rect 16828 32452 16884 32462
rect 16828 32450 16996 32452
rect 16828 32398 16830 32450
rect 16882 32398 16996 32450
rect 16828 32396 16996 32398
rect 16828 32386 16884 32396
rect 16828 31892 16884 31902
rect 16828 31798 16884 31836
rect 16716 31668 16772 31678
rect 16604 31666 16772 31668
rect 16604 31614 16718 31666
rect 16770 31614 16772 31666
rect 16604 31612 16772 31614
rect 16716 31602 16772 31612
rect 16940 31554 16996 32396
rect 16940 31502 16942 31554
rect 16994 31502 16996 31554
rect 16156 30382 16158 30434
rect 16210 30382 16212 30434
rect 16156 30370 16212 30382
rect 16492 30884 16548 30894
rect 15932 30146 15988 30156
rect 16380 30212 16436 30222
rect 16380 30118 16436 30156
rect 15820 29988 15876 29998
rect 15820 29986 16100 29988
rect 15820 29934 15822 29986
rect 15874 29934 16100 29986
rect 15820 29932 16100 29934
rect 15820 29922 15876 29932
rect 16044 29426 16100 29932
rect 16268 29652 16324 29662
rect 16268 29558 16324 29596
rect 16380 29540 16436 29550
rect 16492 29540 16548 30828
rect 16716 30212 16772 30222
rect 16716 30118 16772 30156
rect 16380 29538 16548 29540
rect 16380 29486 16382 29538
rect 16434 29486 16548 29538
rect 16380 29484 16548 29486
rect 16828 30098 16884 30110
rect 16828 30046 16830 30098
rect 16882 30046 16884 30098
rect 16380 29474 16436 29484
rect 16044 29374 16046 29426
rect 16098 29374 16100 29426
rect 15932 28868 15988 28878
rect 16044 28868 16100 29374
rect 15932 28866 16548 28868
rect 15932 28814 15934 28866
rect 15986 28814 16548 28866
rect 15932 28812 16548 28814
rect 15932 28802 15988 28812
rect 16156 28642 16212 28654
rect 16156 28590 16158 28642
rect 16210 28590 16212 28642
rect 16156 28532 16212 28590
rect 16492 28642 16548 28812
rect 16492 28590 16494 28642
rect 16546 28590 16548 28642
rect 16492 28578 16548 28590
rect 16380 28532 16436 28542
rect 16156 28476 16380 28532
rect 16380 28466 16436 28476
rect 16716 28532 16772 28542
rect 15596 28420 15652 28430
rect 15596 28418 16212 28420
rect 15596 28366 15598 28418
rect 15650 28366 16212 28418
rect 15596 28364 16212 28366
rect 15596 28354 15652 28364
rect 16156 27076 16212 28364
rect 16604 28418 16660 28430
rect 16604 28366 16606 28418
rect 16658 28366 16660 28418
rect 16268 27748 16324 27758
rect 16268 27298 16324 27692
rect 16268 27246 16270 27298
rect 16322 27246 16324 27298
rect 16268 27234 16324 27246
rect 16604 27298 16660 28366
rect 16716 27748 16772 28476
rect 16828 28196 16884 30046
rect 16940 30100 16996 31502
rect 16940 30034 16996 30044
rect 17164 31554 17220 31566
rect 17164 31502 17166 31554
rect 17218 31502 17220 31554
rect 17164 31220 17220 31502
rect 17164 28642 17220 31164
rect 17388 31218 17444 32732
rect 17724 32562 17780 32956
rect 17724 32510 17726 32562
rect 17778 32510 17780 32562
rect 17724 32498 17780 32510
rect 18956 32562 19012 32574
rect 18956 32510 18958 32562
rect 19010 32510 19012 32562
rect 17948 32450 18004 32462
rect 17948 32398 17950 32450
rect 18002 32398 18004 32450
rect 17388 31166 17390 31218
rect 17442 31166 17444 31218
rect 17388 31154 17444 31166
rect 17836 31220 17892 31230
rect 17836 31126 17892 31164
rect 17612 30994 17668 31006
rect 17612 30942 17614 30994
rect 17666 30942 17668 30994
rect 17500 30884 17556 30894
rect 17500 30790 17556 30828
rect 17612 30212 17668 30942
rect 17612 30146 17668 30156
rect 17948 30100 18004 32398
rect 18956 32228 19012 32510
rect 18956 30994 19012 32172
rect 18956 30942 18958 30994
rect 19010 30942 19012 30994
rect 18956 30930 19012 30942
rect 17948 30034 18004 30044
rect 18732 30210 18788 30222
rect 18732 30158 18734 30210
rect 18786 30158 18788 30210
rect 18508 29876 18564 29886
rect 18396 28756 18452 28766
rect 18396 28662 18452 28700
rect 17164 28590 17166 28642
rect 17218 28590 17220 28642
rect 16828 28140 16996 28196
rect 16828 27748 16884 27758
rect 16716 27746 16884 27748
rect 16716 27694 16830 27746
rect 16882 27694 16884 27746
rect 16716 27692 16884 27694
rect 16828 27682 16884 27692
rect 16604 27246 16606 27298
rect 16658 27246 16660 27298
rect 16604 27234 16660 27246
rect 16268 27076 16324 27086
rect 16156 27074 16324 27076
rect 16156 27022 16270 27074
rect 16322 27022 16324 27074
rect 16156 27020 16324 27022
rect 16156 26178 16212 27020
rect 16268 27010 16324 27020
rect 16604 26292 16660 26302
rect 16940 26292 16996 28140
rect 16604 26290 16996 26292
rect 16604 26238 16606 26290
rect 16658 26238 16996 26290
rect 16604 26236 16996 26238
rect 16604 26226 16660 26236
rect 16156 26126 16158 26178
rect 16210 26126 16212 26178
rect 16156 26114 16212 26126
rect 15820 26066 15876 26078
rect 15820 26014 15822 26066
rect 15874 26014 15876 26066
rect 15820 24162 15876 26014
rect 15820 24110 15822 24162
rect 15874 24110 15876 24162
rect 15820 24098 15876 24110
rect 15932 24612 15988 24622
rect 15932 24050 15988 24556
rect 16828 24610 16884 26236
rect 16828 24558 16830 24610
rect 16882 24558 16884 24610
rect 16828 24546 16884 24558
rect 15932 23998 15934 24050
rect 15986 23998 15988 24050
rect 15932 23986 15988 23998
rect 16044 23716 16100 23726
rect 16716 23716 16772 23726
rect 15932 23714 16772 23716
rect 15932 23662 16046 23714
rect 16098 23662 16718 23714
rect 16770 23662 16772 23714
rect 15932 23660 16772 23662
rect 15820 21586 15876 21598
rect 15820 21534 15822 21586
rect 15874 21534 15876 21586
rect 15820 20468 15876 21534
rect 15820 20402 15876 20412
rect 15932 17444 15988 23660
rect 16044 23650 16100 23660
rect 16716 23650 16772 23660
rect 16716 23156 16772 23166
rect 16044 22260 16100 22270
rect 16044 22258 16548 22260
rect 16044 22206 16046 22258
rect 16098 22206 16548 22258
rect 16044 22204 16548 22206
rect 16044 22194 16100 22204
rect 16156 22036 16212 22046
rect 16156 21810 16212 21980
rect 16156 21758 16158 21810
rect 16210 21758 16212 21810
rect 16156 21746 16212 21758
rect 16492 21474 16548 22204
rect 16716 22036 16772 23100
rect 17164 23156 17220 28590
rect 17724 28642 17780 28654
rect 17724 28590 17726 28642
rect 17778 28590 17780 28642
rect 17724 27748 17780 28590
rect 17724 27682 17780 27692
rect 18060 25506 18116 25518
rect 18060 25454 18062 25506
rect 18114 25454 18116 25506
rect 18060 25284 18116 25454
rect 17836 24612 17892 24622
rect 17836 23938 17892 24556
rect 18060 24610 18116 25228
rect 18060 24558 18062 24610
rect 18114 24558 18116 24610
rect 18060 24164 18116 24558
rect 18060 24108 18340 24164
rect 17836 23886 17838 23938
rect 17890 23886 17892 23938
rect 17388 23380 17444 23390
rect 17388 23378 17780 23380
rect 17388 23326 17390 23378
rect 17442 23326 17780 23378
rect 17388 23324 17780 23326
rect 17388 23314 17444 23324
rect 17164 23090 17220 23100
rect 17612 23154 17668 23166
rect 17612 23102 17614 23154
rect 17666 23102 17668 23154
rect 17500 23042 17556 23054
rect 17500 22990 17502 23042
rect 17554 22990 17556 23042
rect 17500 22148 17556 22990
rect 17612 22596 17668 23102
rect 17612 22530 17668 22540
rect 16716 21970 16772 21980
rect 16828 22092 17556 22148
rect 17724 22372 17780 23324
rect 16604 21698 16660 21710
rect 16604 21646 16606 21698
rect 16658 21646 16660 21698
rect 16604 21588 16660 21646
rect 16828 21698 16884 22092
rect 16828 21646 16830 21698
rect 16882 21646 16884 21698
rect 16828 21634 16884 21646
rect 16604 21522 16660 21532
rect 17388 21588 17444 21598
rect 17388 21494 17444 21532
rect 17724 21586 17780 22316
rect 17724 21534 17726 21586
rect 17778 21534 17780 21586
rect 17724 21522 17780 21534
rect 16492 21422 16494 21474
rect 16546 21422 16548 21474
rect 16492 21410 16548 21422
rect 17836 21140 17892 23886
rect 17948 23156 18004 23166
rect 17948 23062 18004 23100
rect 17948 22596 18004 22606
rect 18004 22540 18228 22596
rect 17948 21586 18004 22540
rect 18172 22482 18228 22540
rect 18172 22430 18174 22482
rect 18226 22430 18228 22482
rect 18172 22418 18228 22430
rect 18284 22260 18340 24108
rect 17948 21534 17950 21586
rect 18002 21534 18004 21586
rect 17948 21522 18004 21534
rect 18172 22204 18340 22260
rect 17724 21084 17892 21140
rect 17724 20188 17780 21084
rect 17948 21028 18004 21038
rect 17836 20916 17892 20926
rect 17948 20916 18004 20972
rect 17836 20914 18004 20916
rect 17836 20862 17838 20914
rect 17890 20862 18004 20914
rect 17836 20860 18004 20862
rect 17836 20850 17892 20860
rect 17612 20132 17668 20142
rect 17724 20132 17892 20188
rect 17500 19906 17556 19918
rect 17500 19854 17502 19906
rect 17554 19854 17556 19906
rect 16604 19796 16660 19806
rect 16492 19348 16548 19358
rect 16492 18676 16548 19292
rect 16492 18582 16548 18620
rect 16044 18450 16100 18462
rect 16044 18398 16046 18450
rect 16098 18398 16100 18450
rect 16044 18228 16100 18398
rect 16604 18450 16660 19740
rect 17388 19796 17444 19806
rect 17388 19702 17444 19740
rect 17500 19460 17556 19854
rect 17052 19404 17556 19460
rect 17052 19346 17108 19404
rect 17052 19294 17054 19346
rect 17106 19294 17108 19346
rect 17052 19282 17108 19294
rect 17612 19012 17668 20076
rect 17724 19236 17780 19246
rect 17836 19236 17892 20132
rect 17724 19234 17892 19236
rect 17724 19182 17726 19234
rect 17778 19182 17892 19234
rect 17724 19180 17892 19182
rect 17724 19170 17780 19180
rect 18172 19012 18228 22204
rect 17612 18956 17780 19012
rect 17388 18676 17444 18686
rect 16604 18398 16606 18450
rect 16658 18398 16660 18450
rect 16604 18386 16660 18398
rect 16716 18562 16772 18574
rect 16716 18510 16718 18562
rect 16770 18510 16772 18562
rect 16716 18452 16772 18510
rect 16716 18386 16772 18396
rect 17388 18450 17444 18620
rect 17388 18398 17390 18450
rect 17442 18398 17444 18450
rect 17388 18386 17444 18398
rect 17612 18452 17668 18462
rect 17612 18358 17668 18396
rect 16044 18162 16100 18172
rect 17724 17668 17780 18956
rect 18172 18946 18228 18956
rect 18284 21028 18340 21038
rect 18284 18676 18340 20972
rect 18508 20188 18564 29820
rect 18732 28532 18788 30158
rect 19292 30100 19348 30110
rect 19292 30006 19348 30044
rect 19068 29876 19124 29886
rect 19068 29650 19124 29820
rect 19068 29598 19070 29650
rect 19122 29598 19124 29650
rect 19068 29586 19124 29598
rect 19404 29652 19460 29662
rect 19404 29558 19460 29596
rect 18732 28466 18788 28476
rect 19292 27748 19348 27758
rect 19292 26290 19348 27692
rect 19292 26238 19294 26290
rect 19346 26238 19348 26290
rect 19180 25284 19236 25294
rect 19180 25190 19236 25228
rect 18620 24612 18676 24622
rect 18620 24518 18676 24556
rect 19292 24612 19348 26238
rect 19292 24546 19348 24556
rect 18620 23828 18676 23838
rect 18620 23826 19348 23828
rect 18620 23774 18622 23826
rect 18674 23774 19348 23826
rect 18620 23772 19348 23774
rect 18620 23762 18676 23772
rect 19292 23266 19348 23772
rect 19292 23214 19294 23266
rect 19346 23214 19348 23266
rect 19292 23202 19348 23214
rect 19404 23156 19460 23166
rect 19516 23156 19572 33852
rect 20300 33236 20356 33246
rect 20300 33142 20356 33180
rect 20188 33124 20244 33134
rect 19628 33122 20244 33124
rect 19628 33070 20190 33122
rect 20242 33070 20244 33122
rect 19628 33068 20244 33070
rect 19628 32674 19684 33068
rect 20188 33058 20244 33068
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19628 32622 19630 32674
rect 19682 32622 19684 32674
rect 19628 32610 19684 32622
rect 20412 31668 20468 31678
rect 20412 31574 20468 31612
rect 20300 31556 20356 31566
rect 20188 31554 20356 31556
rect 20188 31502 20302 31554
rect 20354 31502 20356 31554
rect 20188 31500 20356 31502
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 20188 31220 20244 31500
rect 20300 31490 20356 31500
rect 19740 31164 20244 31220
rect 19740 31106 19796 31164
rect 19740 31054 19742 31106
rect 19794 31054 19796 31106
rect 19740 31042 19796 31054
rect 20412 29986 20468 29998
rect 20412 29934 20414 29986
rect 20466 29934 20468 29986
rect 20412 29876 20468 29934
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20412 29810 20468 29820
rect 19836 29754 20100 29764
rect 19852 29652 19908 29662
rect 19852 29558 19908 29596
rect 20524 29652 20580 29662
rect 20636 29652 20692 34412
rect 20860 33460 20916 34860
rect 20860 33366 20916 33404
rect 20580 29596 20692 29652
rect 20524 29586 20580 29596
rect 20636 28418 20692 28430
rect 20636 28366 20638 28418
rect 20690 28366 20692 28418
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 20636 28084 20692 28366
rect 20972 28084 21028 28094
rect 20636 28028 20972 28084
rect 20972 27858 21028 28028
rect 20972 27806 20974 27858
rect 21026 27806 21028 27858
rect 20972 27794 21028 27806
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 20076 26404 20132 26414
rect 20076 26310 20132 26348
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19404 23154 19516 23156
rect 19404 23102 19406 23154
rect 19458 23102 19516 23154
rect 19404 23100 19516 23102
rect 19628 24164 19684 24174
rect 19628 23156 19684 24108
rect 20748 24052 20804 24062
rect 20748 23958 20804 23996
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19740 23156 19796 23166
rect 19628 23154 19796 23156
rect 19628 23102 19742 23154
rect 19794 23102 19796 23154
rect 19628 23100 19796 23102
rect 19404 23090 19460 23100
rect 19516 23062 19572 23100
rect 19740 23090 19796 23100
rect 19852 23156 19908 23166
rect 19628 22932 19684 22942
rect 19852 22932 19908 23100
rect 19684 22876 19908 22932
rect 20300 23042 20356 23054
rect 20300 22990 20302 23042
rect 20354 22990 20356 23042
rect 20300 22932 20356 22990
rect 19628 22838 19684 22876
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19180 21812 19236 21822
rect 19180 21810 20020 21812
rect 19180 21758 19182 21810
rect 19234 21758 20020 21810
rect 19180 21756 20020 21758
rect 19180 21746 19236 21756
rect 18844 21586 18900 21598
rect 18844 21534 18846 21586
rect 18898 21534 18900 21586
rect 18508 20132 18676 20188
rect 18620 18900 18676 20132
rect 18844 20132 18900 21534
rect 19180 21586 19236 21598
rect 19180 21534 19182 21586
rect 19234 21534 19236 21586
rect 19180 21028 19236 21534
rect 19180 20962 19236 20972
rect 19516 21586 19572 21598
rect 19516 21534 19518 21586
rect 19570 21534 19572 21586
rect 19516 20242 19572 21534
rect 19964 20914 20020 21756
rect 19964 20862 19966 20914
rect 20018 20862 20020 20914
rect 19964 20850 20020 20862
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19516 20190 19518 20242
rect 19570 20190 19572 20242
rect 19516 20178 19572 20190
rect 20300 20188 20356 22876
rect 18844 20066 18900 20076
rect 19404 20132 19460 20142
rect 19404 20038 19460 20076
rect 20188 20132 20356 20188
rect 20748 20802 20804 20814
rect 20748 20750 20750 20802
rect 20802 20750 20804 20802
rect 20524 20132 20580 20142
rect 19628 20018 19684 20030
rect 19628 19966 19630 20018
rect 19682 19966 19684 20018
rect 18620 18844 18900 18900
rect 17948 18564 18004 18574
rect 17948 18450 18004 18508
rect 17948 18398 17950 18450
rect 18002 18398 18004 18450
rect 17948 18386 18004 18398
rect 17836 17668 17892 17678
rect 17724 17612 17836 17668
rect 17836 17574 17892 17612
rect 18060 17556 18116 17566
rect 18060 17462 18116 17500
rect 18284 17554 18340 18620
rect 18396 18564 18452 18574
rect 18396 18450 18452 18508
rect 18396 18398 18398 18450
rect 18450 18398 18452 18450
rect 18396 18386 18452 18398
rect 18620 18562 18676 18574
rect 18620 18510 18622 18562
rect 18674 18510 18676 18562
rect 18284 17502 18286 17554
rect 18338 17502 18340 17554
rect 18284 17490 18340 17502
rect 18396 17666 18452 17678
rect 18396 17614 18398 17666
rect 18450 17614 18452 17666
rect 15932 17378 15988 17388
rect 17388 17444 17444 17454
rect 17388 17442 17892 17444
rect 17388 17390 17390 17442
rect 17442 17390 17892 17442
rect 17388 17388 17892 17390
rect 17388 17378 17444 17388
rect 15708 17108 15764 17118
rect 15708 17014 15764 17052
rect 15148 16210 15540 16212
rect 15148 16158 15486 16210
rect 15538 16158 15540 16210
rect 15148 16156 15540 16158
rect 15036 16100 15092 16110
rect 15036 16006 15092 16044
rect 14812 15374 14814 15426
rect 14866 15374 14868 15426
rect 14812 15362 14868 15374
rect 13580 15314 13636 15326
rect 13580 15262 13582 15314
rect 13634 15262 13636 15314
rect 13580 15148 13636 15262
rect 13804 15314 13860 15326
rect 13804 15262 13806 15314
rect 13858 15262 13860 15314
rect 13580 15092 13748 15148
rect 13468 14478 13470 14530
rect 13522 14478 13524 14530
rect 13244 13636 13300 13646
rect 13244 13542 13300 13580
rect 13468 12628 13524 14478
rect 13692 14308 13748 15092
rect 13804 14644 13860 15262
rect 15148 15148 15204 16156
rect 15484 16146 15540 16156
rect 16044 16994 16100 17006
rect 16044 16942 16046 16994
rect 16098 16942 16100 16994
rect 16044 16772 16100 16942
rect 16044 15876 16100 16716
rect 16828 16884 16884 16894
rect 16044 15820 16436 15876
rect 16380 15148 16436 15820
rect 15148 15092 15428 15148
rect 13916 14644 13972 14654
rect 13804 14642 13972 14644
rect 13804 14590 13918 14642
rect 13970 14590 13972 14642
rect 13804 14588 13972 14590
rect 13916 14578 13972 14588
rect 14028 14532 14084 14542
rect 14028 14438 14084 14476
rect 13804 14308 13860 14318
rect 13692 14306 13860 14308
rect 13692 14254 13806 14306
rect 13858 14254 13860 14306
rect 13692 14252 13860 14254
rect 13580 13746 13636 13758
rect 13580 13694 13582 13746
rect 13634 13694 13636 13746
rect 13580 13636 13636 13694
rect 13692 13748 13748 14252
rect 13804 14242 13860 14252
rect 15260 14308 15316 14318
rect 13692 13654 13748 13692
rect 13580 13570 13636 13580
rect 13468 12562 13524 12572
rect 13916 12628 13972 12638
rect 12572 12348 12964 12404
rect 12572 12290 12628 12348
rect 12572 12238 12574 12290
rect 12626 12238 12628 12290
rect 12572 12226 12628 12238
rect 12236 12180 12292 12190
rect 12236 12086 12292 12124
rect 12796 12178 12852 12190
rect 12796 12126 12798 12178
rect 12850 12126 12852 12178
rect 12348 12068 12404 12078
rect 12348 11974 12404 12012
rect 12796 11508 12852 12126
rect 12796 11442 12852 11452
rect 12908 11506 12964 12348
rect 12908 11454 12910 11506
rect 12962 11454 12964 11506
rect 12908 11396 12964 11454
rect 12908 11330 12964 11340
rect 13468 12180 13524 12190
rect 13468 11394 13524 12124
rect 13580 11508 13636 11518
rect 13580 11414 13636 11452
rect 13468 11342 13470 11394
rect 13522 11342 13524 11394
rect 13468 11330 13524 11342
rect 13692 11396 13748 11406
rect 13692 11302 13748 11340
rect 13916 11282 13972 12572
rect 14252 12290 14308 12302
rect 14252 12238 14254 12290
rect 14306 12238 14308 12290
rect 14252 12180 14308 12238
rect 14924 12292 14980 12302
rect 14252 12114 14308 12124
rect 14588 12180 14644 12190
rect 14924 12180 14980 12236
rect 15260 12290 15316 14252
rect 15260 12238 15262 12290
rect 15314 12238 15316 12290
rect 15260 12226 15316 12238
rect 13916 11230 13918 11282
rect 13970 11230 13972 11282
rect 13916 11218 13972 11230
rect 14028 11844 14084 11854
rect 14028 10610 14084 11788
rect 14476 11396 14532 11406
rect 14476 11284 14532 11340
rect 14588 11394 14644 12124
rect 14812 12178 14980 12180
rect 14812 12126 14926 12178
rect 14978 12126 14980 12178
rect 14812 12124 14980 12126
rect 14588 11342 14590 11394
rect 14642 11342 14644 11394
rect 14588 11330 14644 11342
rect 14700 11844 14756 11854
rect 14364 11282 14532 11284
rect 14364 11230 14478 11282
rect 14530 11230 14532 11282
rect 14364 11228 14532 11230
rect 14252 11172 14308 11182
rect 14028 10558 14030 10610
rect 14082 10558 14084 10610
rect 14028 10546 14084 10558
rect 14140 11170 14308 11172
rect 14140 11118 14254 11170
rect 14306 11118 14308 11170
rect 14140 11116 14308 11118
rect 13580 9716 13636 9726
rect 12236 9268 12292 9278
rect 12124 9266 12628 9268
rect 12124 9214 12238 9266
rect 12290 9214 12628 9266
rect 12124 9212 12628 9214
rect 10668 9174 10724 9212
rect 12236 9202 12292 9212
rect 12572 9044 12628 9212
rect 12572 9042 12740 9044
rect 12572 8990 12574 9042
rect 12626 8990 12740 9042
rect 12572 8988 12740 8990
rect 12572 8978 12628 8988
rect 12572 8820 12628 8830
rect 10332 8306 10388 8316
rect 12348 8818 12628 8820
rect 12348 8766 12574 8818
rect 12626 8766 12628 8818
rect 12348 8764 12628 8766
rect 9660 8036 9716 8046
rect 12348 8036 12404 8764
rect 12572 8754 12628 8764
rect 12684 8148 12740 8988
rect 12908 8932 12964 8942
rect 13468 8932 13524 8942
rect 12908 8930 13524 8932
rect 12908 8878 12910 8930
rect 12962 8878 13470 8930
rect 13522 8878 13524 8930
rect 12908 8876 13524 8878
rect 12908 8866 12964 8876
rect 13468 8866 13524 8876
rect 12684 8082 12740 8092
rect 9660 8034 10052 8036
rect 9660 7982 9662 8034
rect 9714 7982 10052 8034
rect 9660 7980 10052 7982
rect 9660 7970 9716 7980
rect 9996 7586 10052 7980
rect 12012 7980 12404 8036
rect 9996 7534 9998 7586
rect 10050 7534 10052 7586
rect 9996 7522 10052 7534
rect 10332 7588 10388 7598
rect 10332 7586 10724 7588
rect 10332 7534 10334 7586
rect 10386 7534 10724 7586
rect 10332 7532 10724 7534
rect 10332 7522 10388 7532
rect 10668 5234 10724 7532
rect 12012 7586 12068 7980
rect 12012 7534 12014 7586
rect 12066 7534 12068 7586
rect 12012 7522 12068 7534
rect 10668 5182 10670 5234
rect 10722 5182 10724 5234
rect 10668 5170 10724 5182
rect 11228 7474 11284 7486
rect 11228 7422 11230 7474
rect 11282 7422 11284 7474
rect 11228 6692 11284 7422
rect 9324 5070 9326 5122
rect 9378 5070 9380 5122
rect 9324 5058 9380 5070
rect 9996 5124 10052 5134
rect 9996 5122 10164 5124
rect 9996 5070 9998 5122
rect 10050 5070 10164 5122
rect 9996 5068 10164 5070
rect 9996 5058 10052 5068
rect 9548 4900 9604 4910
rect 9548 4806 9604 4844
rect 10108 4340 10164 5068
rect 10892 4900 10948 4910
rect 10892 4450 10948 4844
rect 10892 4398 10894 4450
rect 10946 4398 10948 4450
rect 10892 4386 10948 4398
rect 10220 4340 10276 4350
rect 10108 4284 10220 4340
rect 10220 4246 10276 4284
rect 11228 4340 11284 6636
rect 13580 6690 13636 9660
rect 14028 9042 14084 9054
rect 14028 8990 14030 9042
rect 14082 8990 14084 9042
rect 14028 8708 14084 8990
rect 14140 8932 14196 11116
rect 14252 11106 14308 11116
rect 14364 10836 14420 11228
rect 14476 11218 14532 11228
rect 14252 10780 14420 10836
rect 14252 10722 14308 10780
rect 14252 10670 14254 10722
rect 14306 10670 14308 10722
rect 14252 10658 14308 10670
rect 14364 10610 14420 10622
rect 14364 10558 14366 10610
rect 14418 10558 14420 10610
rect 14252 8932 14308 8942
rect 14140 8930 14308 8932
rect 14140 8878 14254 8930
rect 14306 8878 14308 8930
rect 14140 8876 14308 8878
rect 14252 8866 14308 8876
rect 14364 8708 14420 10558
rect 14700 9268 14756 11788
rect 14812 10610 14868 12124
rect 14924 12114 14980 12124
rect 14924 11954 14980 11966
rect 14924 11902 14926 11954
rect 14978 11902 14980 11954
rect 14924 11508 14980 11902
rect 14924 11442 14980 11452
rect 14812 10558 14814 10610
rect 14866 10558 14868 10610
rect 14812 10546 14868 10558
rect 14924 11172 14980 11182
rect 14924 9826 14980 11116
rect 15036 10612 15092 10622
rect 15260 10612 15316 10622
rect 15036 10610 15316 10612
rect 15036 10558 15038 10610
rect 15090 10558 15262 10610
rect 15314 10558 15316 10610
rect 15036 10556 15316 10558
rect 15036 10546 15092 10556
rect 15260 10546 15316 10556
rect 14924 9774 14926 9826
rect 14978 9774 14980 9826
rect 14812 9268 14868 9278
rect 14700 9266 14868 9268
rect 14700 9214 14814 9266
rect 14866 9214 14868 9266
rect 14700 9212 14868 9214
rect 14812 9202 14868 9212
rect 14028 8652 14420 8708
rect 14140 7362 14196 8652
rect 14140 7310 14142 7362
rect 14194 7310 14196 7362
rect 14140 7298 14196 7310
rect 13580 6638 13582 6690
rect 13634 6638 13636 6690
rect 13580 6626 13636 6638
rect 14252 6580 14308 6590
rect 14252 6486 14308 6524
rect 14924 5908 14980 9774
rect 15372 9268 15428 15092
rect 16268 15092 16436 15148
rect 15484 14532 15540 14542
rect 15484 13972 15540 14476
rect 16156 14420 16212 14430
rect 15484 13878 15540 13916
rect 15596 14418 16212 14420
rect 15596 14366 16158 14418
rect 16210 14366 16212 14418
rect 15596 14364 16212 14366
rect 15596 13970 15652 14364
rect 16156 14354 16212 14364
rect 15596 13918 15598 13970
rect 15650 13918 15652 13970
rect 15596 13906 15652 13918
rect 16268 14306 16324 15092
rect 16716 14644 16772 14654
rect 16268 14254 16270 14306
rect 16322 14254 16324 14306
rect 15932 13858 15988 13870
rect 15932 13806 15934 13858
rect 15986 13806 15988 13858
rect 15708 13748 15764 13758
rect 15596 12180 15652 12190
rect 15596 12086 15652 12124
rect 15708 12178 15764 13692
rect 15708 12126 15710 12178
rect 15762 12126 15764 12178
rect 15708 12114 15764 12126
rect 15932 12404 15988 13806
rect 16268 13860 16324 14254
rect 16492 14308 16548 14318
rect 16492 14214 16548 14252
rect 16380 13972 16436 13982
rect 16716 13972 16772 14588
rect 16380 13878 16436 13916
rect 16492 13970 16772 13972
rect 16492 13918 16718 13970
rect 16770 13918 16772 13970
rect 16492 13916 16772 13918
rect 16268 13794 16324 13804
rect 16492 13412 16548 13916
rect 16716 13906 16772 13916
rect 16828 13748 16884 16828
rect 17052 16212 17108 16222
rect 17052 14644 17108 16156
rect 17836 16098 17892 17388
rect 18284 16772 18340 16782
rect 18396 16772 18452 17614
rect 18620 17668 18676 18510
rect 18620 17602 18676 17612
rect 18340 16716 18452 16772
rect 18284 16706 18340 16716
rect 17836 16046 17838 16098
rect 17890 16046 17892 16098
rect 17836 16034 17892 16046
rect 18172 15874 18228 15886
rect 18172 15822 18174 15874
rect 18226 15822 18228 15874
rect 18172 15426 18228 15822
rect 18172 15374 18174 15426
rect 18226 15374 18228 15426
rect 18172 15362 18228 15374
rect 17500 15314 17556 15326
rect 17500 15262 17502 15314
rect 17554 15262 17556 15314
rect 17500 15148 17556 15262
rect 18844 15148 18900 18844
rect 19068 18676 19124 18686
rect 19628 18676 19684 19966
rect 20076 20020 20132 20030
rect 20076 19926 20132 19964
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19124 18620 19684 18676
rect 19068 18582 19124 18620
rect 18956 18564 19012 18574
rect 18956 18470 19012 18508
rect 19292 18450 19348 18462
rect 19292 18398 19294 18450
rect 19346 18398 19348 18450
rect 19292 17778 19348 18398
rect 19292 17726 19294 17778
rect 19346 17726 19348 17778
rect 19292 17714 19348 17726
rect 20188 18340 20244 20132
rect 20524 20038 20580 20076
rect 20748 19124 20804 20750
rect 21196 20020 21252 36204
rect 21420 36194 21476 36204
rect 21868 34132 21924 34142
rect 21868 33458 21924 34076
rect 21868 33406 21870 33458
rect 21922 33406 21924 33458
rect 21756 32452 21812 32462
rect 21756 32358 21812 32396
rect 21308 32228 21364 32238
rect 21308 29426 21364 32172
rect 21868 32228 21924 33406
rect 21868 32162 21924 32172
rect 21980 32004 22036 36428
rect 22652 35924 22708 37324
rect 22876 37314 22932 37324
rect 22988 37378 23044 37548
rect 23212 37492 23268 37996
rect 23324 37828 23380 37838
rect 23548 37828 23604 37838
rect 23772 37828 23828 37838
rect 23324 37826 23604 37828
rect 23324 37774 23326 37826
rect 23378 37774 23550 37826
rect 23602 37774 23604 37826
rect 23324 37772 23604 37774
rect 23324 37762 23380 37772
rect 23548 37762 23604 37772
rect 23660 37826 23828 37828
rect 23660 37774 23774 37826
rect 23826 37774 23828 37826
rect 23660 37772 23828 37774
rect 22988 37326 22990 37378
rect 23042 37326 23044 37378
rect 22988 37268 23044 37326
rect 22988 37202 23044 37212
rect 23100 37436 23268 37492
rect 22876 35924 22932 35934
rect 22652 35922 22932 35924
rect 22652 35870 22878 35922
rect 22930 35870 22932 35922
rect 22652 35868 22932 35870
rect 22876 35858 22932 35868
rect 22540 34018 22596 34030
rect 22540 33966 22542 34018
rect 22594 33966 22596 34018
rect 22428 33236 22484 33246
rect 22428 32786 22484 33180
rect 22428 32734 22430 32786
rect 22482 32734 22484 32786
rect 22428 32722 22484 32734
rect 22540 32788 22596 33966
rect 22764 32900 22820 32910
rect 22540 32722 22596 32732
rect 22652 32844 22764 32900
rect 22652 32786 22708 32844
rect 22764 32834 22820 32844
rect 23100 32788 23156 37436
rect 23212 37268 23268 37278
rect 23436 37268 23492 37278
rect 23212 37266 23492 37268
rect 23212 37214 23214 37266
rect 23266 37214 23438 37266
rect 23490 37214 23492 37266
rect 23212 37212 23492 37214
rect 23212 37202 23268 37212
rect 23436 37202 23492 37212
rect 23660 37266 23716 37772
rect 23772 37762 23828 37772
rect 23660 37214 23662 37266
rect 23714 37214 23716 37266
rect 23548 37156 23604 37166
rect 23548 37062 23604 37100
rect 23660 35476 23716 37214
rect 23660 35410 23716 35420
rect 23884 34580 23940 39564
rect 24220 39620 24276 39630
rect 23996 37828 24052 37838
rect 23996 37734 24052 37772
rect 24108 37268 24164 37278
rect 24108 37174 24164 37212
rect 24220 36482 24276 39564
rect 24444 39508 24500 40236
rect 24556 40180 24612 42588
rect 24668 41972 24724 41982
rect 24668 40402 24724 41916
rect 25004 40962 25060 40974
rect 25004 40910 25006 40962
rect 25058 40910 25060 40962
rect 24668 40350 24670 40402
rect 24722 40350 24724 40402
rect 24668 40338 24724 40350
rect 24780 40516 24836 40526
rect 24556 39620 24612 40124
rect 24780 39730 24836 40460
rect 25004 40292 25060 40910
rect 25228 40964 25284 46620
rect 25340 45556 25396 45566
rect 25340 45106 25396 45500
rect 25340 45054 25342 45106
rect 25394 45054 25396 45106
rect 25340 45042 25396 45054
rect 25340 44546 25396 44558
rect 25340 44494 25342 44546
rect 25394 44494 25396 44546
rect 25340 42196 25396 44494
rect 25452 43652 25508 48076
rect 25788 46676 25844 48636
rect 25788 46582 25844 46620
rect 25564 45780 25620 45790
rect 25564 45686 25620 45724
rect 26012 44548 26068 51212
rect 26236 50148 26292 53118
rect 26348 53058 26404 53564
rect 26348 53006 26350 53058
rect 26402 53006 26404 53058
rect 26348 52994 26404 53006
rect 26460 53508 26516 53518
rect 26460 52274 26516 53452
rect 26460 52222 26462 52274
rect 26514 52222 26516 52274
rect 26460 52210 26516 52222
rect 26460 51604 26516 51614
rect 26572 51604 26628 53900
rect 26908 53862 26964 53900
rect 27020 53732 27076 54236
rect 27132 53954 27188 54684
rect 27468 54674 27524 54684
rect 28252 54740 28308 54750
rect 27132 53902 27134 53954
rect 27186 53902 27188 53954
rect 27132 53890 27188 53902
rect 28140 53844 28196 53854
rect 27244 53732 27300 53742
rect 27580 53732 27636 53742
rect 27020 53730 27524 53732
rect 27020 53678 27246 53730
rect 27298 53678 27524 53730
rect 27020 53676 27524 53678
rect 27244 53666 27300 53676
rect 27244 53508 27300 53518
rect 27244 53414 27300 53452
rect 27468 53284 27524 53676
rect 27580 53638 27636 53676
rect 27916 53730 27972 53742
rect 27916 53678 27918 53730
rect 27970 53678 27972 53730
rect 27916 53508 27972 53678
rect 27916 53442 27972 53452
rect 27468 53228 28084 53284
rect 28028 53058 28084 53228
rect 28140 53170 28196 53788
rect 28252 53732 28308 54684
rect 28252 53638 28308 53676
rect 28364 53618 28420 55020
rect 29036 54516 29092 54526
rect 29036 54422 29092 54460
rect 28364 53566 28366 53618
rect 28418 53566 28420 53618
rect 28364 53396 28420 53566
rect 28140 53118 28142 53170
rect 28194 53118 28196 53170
rect 28140 53106 28196 53118
rect 28252 53340 28420 53396
rect 28476 53730 28532 53742
rect 28476 53678 28478 53730
rect 28530 53678 28532 53730
rect 28028 53006 28030 53058
rect 28082 53006 28084 53058
rect 28028 52994 28084 53006
rect 26460 51602 26628 51604
rect 26460 51550 26462 51602
rect 26514 51550 26628 51602
rect 26460 51548 26628 51550
rect 26460 51538 26516 51548
rect 28028 51492 28084 51502
rect 28252 51492 28308 53340
rect 28364 52948 28420 52958
rect 28476 52948 28532 53678
rect 28420 52892 28532 52948
rect 29148 52948 29204 55358
rect 36428 55410 36484 55422
rect 36428 55358 36430 55410
rect 36482 55358 36484 55410
rect 32060 55300 32116 55310
rect 32060 55206 32116 55244
rect 33516 55300 33572 55310
rect 33516 55206 33572 55244
rect 34076 55300 34132 55310
rect 29820 55188 29876 55198
rect 29484 53956 29540 53966
rect 29484 53862 29540 53900
rect 29372 53844 29428 53854
rect 29372 53750 29428 53788
rect 29708 53844 29764 53854
rect 29708 53750 29764 53788
rect 29820 53730 29876 55132
rect 31276 55188 31332 55198
rect 31276 55094 31332 55132
rect 31388 55076 31444 55086
rect 31388 54516 31444 55020
rect 29820 53678 29822 53730
rect 29874 53678 29876 53730
rect 29820 53666 29876 53678
rect 30940 54514 31444 54516
rect 30940 54462 31390 54514
rect 31442 54462 31444 54514
rect 30940 54460 31444 54462
rect 30940 53618 30996 54460
rect 31388 54450 31444 54460
rect 31612 54290 31668 54302
rect 31612 54238 31614 54290
rect 31666 54238 31668 54290
rect 30940 53566 30942 53618
rect 30994 53566 30996 53618
rect 30940 53554 30996 53566
rect 31276 53842 31332 53854
rect 31276 53790 31278 53842
rect 31330 53790 31332 53842
rect 30604 53508 30660 53518
rect 29260 52948 29316 52958
rect 29148 52892 29260 52948
rect 28364 52854 28420 52892
rect 28028 51490 28308 51492
rect 28028 51438 28030 51490
rect 28082 51438 28308 51490
rect 28028 51436 28308 51438
rect 28588 52274 28644 52286
rect 28588 52222 28590 52274
rect 28642 52222 28644 52274
rect 27132 50932 27188 50942
rect 26908 50596 26964 50634
rect 26908 50530 26964 50540
rect 27132 50482 27188 50876
rect 27132 50430 27134 50482
rect 27186 50430 27188 50482
rect 27132 50428 27188 50430
rect 26908 50372 27188 50428
rect 26236 50082 26292 50092
rect 26796 50316 26964 50372
rect 26796 50034 26852 50316
rect 26796 49982 26798 50034
rect 26850 49982 26852 50034
rect 26796 49970 26852 49982
rect 26908 50148 26964 50158
rect 26684 49810 26740 49822
rect 26684 49758 26686 49810
rect 26738 49758 26740 49810
rect 26124 49700 26180 49710
rect 26124 49606 26180 49644
rect 26572 49700 26628 49710
rect 26684 49700 26740 49758
rect 26628 49644 26740 49700
rect 26572 49634 26628 49644
rect 26348 49588 26404 49626
rect 26348 49522 26404 49532
rect 26796 49586 26852 49598
rect 26796 49534 26798 49586
rect 26850 49534 26852 49586
rect 26348 49364 26404 49374
rect 26348 49026 26404 49308
rect 26348 48974 26350 49026
rect 26402 48974 26404 49026
rect 26348 48962 26404 48974
rect 26572 48916 26628 48926
rect 26796 48916 26852 49534
rect 26572 48914 26852 48916
rect 26572 48862 26574 48914
rect 26626 48862 26852 48914
rect 26572 48860 26852 48862
rect 26572 48850 26628 48860
rect 26684 48468 26740 48478
rect 26908 48468 26964 50092
rect 27692 49026 27748 49038
rect 27692 48974 27694 49026
rect 27746 48974 27748 49026
rect 26684 48466 26964 48468
rect 26684 48414 26686 48466
rect 26738 48414 26964 48466
rect 26684 48412 26964 48414
rect 26684 48402 26740 48412
rect 26572 48242 26628 48254
rect 26572 48190 26574 48242
rect 26626 48190 26628 48242
rect 26572 47572 26628 48190
rect 26796 48244 26852 48254
rect 26684 48020 26740 48030
rect 26796 48020 26852 48188
rect 26684 48018 26852 48020
rect 26684 47966 26686 48018
rect 26738 47966 26852 48018
rect 26684 47964 26852 47966
rect 26684 47954 26740 47964
rect 26684 47572 26740 47582
rect 26572 47570 26740 47572
rect 26572 47518 26686 47570
rect 26738 47518 26740 47570
rect 26572 47516 26740 47518
rect 26460 46900 26516 46910
rect 26460 46674 26516 46844
rect 26460 46622 26462 46674
rect 26514 46622 26516 46674
rect 26460 46610 26516 46622
rect 26124 46564 26180 46574
rect 26124 46470 26180 46508
rect 26460 46450 26516 46462
rect 26460 46398 26462 46450
rect 26514 46398 26516 46450
rect 26124 45890 26180 45902
rect 26124 45838 26126 45890
rect 26178 45838 26180 45890
rect 26124 44882 26180 45838
rect 26348 45220 26404 45230
rect 26348 45106 26404 45164
rect 26348 45054 26350 45106
rect 26402 45054 26404 45106
rect 26348 45042 26404 45054
rect 26460 45108 26516 46398
rect 26460 45042 26516 45052
rect 26124 44830 26126 44882
rect 26178 44830 26180 44882
rect 26124 44818 26180 44830
rect 26012 44492 26404 44548
rect 25788 44324 25844 44334
rect 25788 44210 25844 44268
rect 25788 44158 25790 44210
rect 25842 44158 25844 44210
rect 25788 44146 25844 44158
rect 25452 43586 25508 43596
rect 25676 43428 25732 43438
rect 25676 43426 25956 43428
rect 25676 43374 25678 43426
rect 25730 43374 25956 43426
rect 25676 43372 25956 43374
rect 25676 43362 25732 43372
rect 25564 43316 25620 43326
rect 25564 43222 25620 43260
rect 25340 42130 25396 42140
rect 25676 42196 25732 42206
rect 25340 41858 25396 41870
rect 25340 41806 25342 41858
rect 25394 41806 25396 41858
rect 25340 41412 25396 41806
rect 25340 41188 25396 41356
rect 25340 41132 25508 41188
rect 25340 40964 25396 40974
rect 25228 40962 25396 40964
rect 25228 40910 25342 40962
rect 25394 40910 25396 40962
rect 25228 40908 25396 40910
rect 25340 40404 25396 40908
rect 25340 40338 25396 40348
rect 25004 40226 25060 40236
rect 24780 39678 24782 39730
rect 24834 39678 24836 39730
rect 24780 39666 24836 39678
rect 24556 39554 24612 39564
rect 25340 39620 25396 39630
rect 25340 39526 25396 39564
rect 24444 39172 24500 39452
rect 24892 39508 24948 39518
rect 24892 39414 24948 39452
rect 24444 39106 24500 39116
rect 24220 36430 24222 36482
rect 24274 36430 24276 36482
rect 24220 36418 24276 36430
rect 25452 36484 25508 41132
rect 25452 36418 25508 36428
rect 25004 36372 25060 36382
rect 25004 36278 25060 36316
rect 25676 34916 25732 42140
rect 25788 41972 25844 41982
rect 25788 41188 25844 41916
rect 25900 41858 25956 43372
rect 25900 41806 25902 41858
rect 25954 41806 25956 41858
rect 25900 41794 25956 41806
rect 26012 42084 26068 42094
rect 26012 41300 26068 42028
rect 26236 41972 26292 41982
rect 26012 41234 26068 41244
rect 26124 41916 26236 41972
rect 26124 41748 26180 41916
rect 26236 41878 26292 41916
rect 26348 41748 26404 44492
rect 26460 44322 26516 44334
rect 26460 44270 26462 44322
rect 26514 44270 26516 44322
rect 26460 44212 26516 44270
rect 26460 44146 26516 44156
rect 26460 42868 26516 42878
rect 26460 42082 26516 42812
rect 26460 42030 26462 42082
rect 26514 42030 26516 42082
rect 26460 42018 26516 42030
rect 25788 41094 25844 41132
rect 26124 41186 26180 41692
rect 26124 41134 26126 41186
rect 26178 41134 26180 41186
rect 26124 41122 26180 41134
rect 26236 41692 26404 41748
rect 25900 40964 25956 40974
rect 25900 40870 25956 40908
rect 26012 40962 26068 40974
rect 26012 40910 26014 40962
rect 26066 40910 26068 40962
rect 26012 40516 26068 40910
rect 26012 40450 26068 40460
rect 26012 39508 26068 39518
rect 26012 39414 26068 39452
rect 26124 36372 26180 36382
rect 26124 35922 26180 36316
rect 26124 35870 26126 35922
rect 26178 35870 26180 35922
rect 26124 35858 26180 35870
rect 26012 35698 26068 35710
rect 26012 35646 26014 35698
rect 26066 35646 26068 35698
rect 26012 35476 26068 35646
rect 26012 35410 26068 35420
rect 25340 34914 25732 34916
rect 25340 34862 25678 34914
rect 25730 34862 25732 34914
rect 25340 34860 25732 34862
rect 23884 34524 24276 34580
rect 24108 32900 24164 32910
rect 23324 32788 23380 32798
rect 22652 32734 22654 32786
rect 22706 32734 22708 32786
rect 22652 32722 22708 32734
rect 22876 32786 23380 32788
rect 22876 32734 23326 32786
rect 23378 32734 23380 32786
rect 22876 32732 23380 32734
rect 22316 32676 22372 32686
rect 22204 32620 22316 32676
rect 21868 31948 22036 32004
rect 22092 32562 22148 32574
rect 22092 32510 22094 32562
rect 22146 32510 22148 32562
rect 22092 32452 22148 32510
rect 21868 31108 21924 31948
rect 21756 31052 21924 31108
rect 21980 31666 22036 31678
rect 21980 31614 21982 31666
rect 22034 31614 22036 31666
rect 21756 30660 21812 31052
rect 21980 30996 22036 31614
rect 22092 31108 22148 32396
rect 22204 31778 22260 32620
rect 22316 32582 22372 32620
rect 22428 32564 22484 32574
rect 22428 32340 22484 32508
rect 22540 32562 22596 32574
rect 22540 32510 22542 32562
rect 22594 32510 22596 32562
rect 22540 32452 22596 32510
rect 22876 32452 22932 32732
rect 23324 32722 23380 32732
rect 23548 32788 23604 32798
rect 23548 32694 23604 32732
rect 24108 32564 24164 32844
rect 24108 32470 24164 32508
rect 24220 32562 24276 34524
rect 24668 34018 24724 34030
rect 24668 33966 24670 34018
rect 24722 33966 24724 34018
rect 24444 32676 24500 32686
rect 24444 32582 24500 32620
rect 24220 32510 24222 32562
rect 24274 32510 24276 32562
rect 22540 32396 22932 32452
rect 23660 32450 23716 32462
rect 23660 32398 23662 32450
rect 23714 32398 23716 32450
rect 22428 32284 22596 32340
rect 22204 31726 22206 31778
rect 22258 31726 22260 31778
rect 22204 31714 22260 31726
rect 22428 31780 22484 31790
rect 22428 31686 22484 31724
rect 22540 31778 22596 32284
rect 23324 32228 23380 32238
rect 23660 32228 23716 32398
rect 24220 32452 24276 32510
rect 24668 32562 24724 33966
rect 25228 33460 25284 33470
rect 25228 33346 25284 33404
rect 25228 33294 25230 33346
rect 25282 33294 25284 33346
rect 25228 33282 25284 33294
rect 24668 32510 24670 32562
rect 24722 32510 24724 32562
rect 24220 32386 24276 32396
rect 24332 32450 24388 32462
rect 24332 32398 24334 32450
rect 24386 32398 24388 32450
rect 24332 32228 24388 32398
rect 23660 32172 24388 32228
rect 22540 31726 22542 31778
rect 22594 31726 22596 31778
rect 22540 31714 22596 31726
rect 22988 31780 23044 31790
rect 22316 31668 22372 31678
rect 22316 31574 22372 31612
rect 22988 31218 23044 31724
rect 23324 31778 23380 32172
rect 24108 32004 24164 32014
rect 24108 31890 24164 31948
rect 24108 31838 24110 31890
rect 24162 31838 24164 31890
rect 24108 31826 24164 31838
rect 23324 31726 23326 31778
rect 23378 31726 23380 31778
rect 23324 31714 23380 31726
rect 22988 31166 22990 31218
rect 23042 31166 23044 31218
rect 22988 31154 23044 31166
rect 22428 31108 22484 31118
rect 22092 31106 22484 31108
rect 22092 31054 22430 31106
rect 22482 31054 22484 31106
rect 22092 31052 22484 31054
rect 22428 31042 22484 31052
rect 21868 30940 22148 30996
rect 21868 30882 21924 30940
rect 21868 30830 21870 30882
rect 21922 30830 21924 30882
rect 21868 30818 21924 30830
rect 22092 30772 22148 30940
rect 22540 30772 22596 30782
rect 22092 30716 22484 30772
rect 21756 30604 21924 30660
rect 21308 29374 21310 29426
rect 21362 29374 21364 29426
rect 21308 29362 21364 29374
rect 21308 27746 21364 27758
rect 21308 27694 21310 27746
rect 21362 27694 21364 27746
rect 21308 27636 21364 27694
rect 21364 27580 21700 27636
rect 21308 27570 21364 27580
rect 21644 27188 21700 27580
rect 21644 27094 21700 27132
rect 21868 26908 21924 30604
rect 22092 29314 22148 29326
rect 22092 29262 22094 29314
rect 22146 29262 22148 29314
rect 22092 28868 22148 29262
rect 22092 28802 22148 28812
rect 22316 28980 22372 28990
rect 22316 28754 22372 28924
rect 22316 28702 22318 28754
rect 22370 28702 22372 28754
rect 22316 28084 22372 28702
rect 22428 28308 22484 30716
rect 22540 30770 22820 30772
rect 22540 30718 22542 30770
rect 22594 30718 22820 30770
rect 22540 30716 22820 30718
rect 22540 30706 22596 30716
rect 22764 28530 22820 30716
rect 24668 30324 24724 32510
rect 25228 32788 25284 32798
rect 25340 32788 25396 34860
rect 25676 34850 25732 34860
rect 26012 34916 26068 34926
rect 26236 34916 26292 41692
rect 26348 41076 26404 41086
rect 26348 40982 26404 41020
rect 26684 41076 26740 47516
rect 26908 47458 26964 48412
rect 27244 48802 27300 48814
rect 27244 48750 27246 48802
rect 27298 48750 27300 48802
rect 27244 48242 27300 48750
rect 27244 48190 27246 48242
rect 27298 48190 27300 48242
rect 27244 48178 27300 48190
rect 27468 48242 27524 48254
rect 27468 48190 27470 48242
rect 27522 48190 27524 48242
rect 27468 47682 27524 48190
rect 27468 47630 27470 47682
rect 27522 47630 27524 47682
rect 27468 47618 27524 47630
rect 27692 47460 27748 48974
rect 28028 49028 28084 51436
rect 28364 51380 28420 51390
rect 28588 51380 28644 52222
rect 28364 51378 28644 51380
rect 28364 51326 28366 51378
rect 28418 51326 28644 51378
rect 28364 51324 28644 51326
rect 28364 51156 28420 51324
rect 28364 51090 28420 51100
rect 28700 50820 28756 50830
rect 28252 50484 28308 50522
rect 28252 50418 28308 50428
rect 28588 50484 28644 50522
rect 28588 50418 28644 50428
rect 28028 48962 28084 48972
rect 27804 48916 27860 48926
rect 27804 47570 27860 48860
rect 27804 47518 27806 47570
rect 27858 47518 27860 47570
rect 27804 47506 27860 47518
rect 28588 47572 28644 47582
rect 28588 47478 28644 47516
rect 26908 47406 26910 47458
rect 26962 47406 26964 47458
rect 26908 47394 26964 47406
rect 27244 47458 27748 47460
rect 27244 47406 27694 47458
rect 27746 47406 27748 47458
rect 27244 47404 27748 47406
rect 26908 46676 26964 46714
rect 26908 46610 26964 46620
rect 26796 46564 26852 46574
rect 26796 45890 26852 46508
rect 26796 45838 26798 45890
rect 26850 45838 26852 45890
rect 26796 45332 26852 45838
rect 26908 46452 26964 46462
rect 26908 45778 26964 46396
rect 26908 45726 26910 45778
rect 26962 45726 26964 45778
rect 26908 45714 26964 45726
rect 27132 45666 27188 45678
rect 27132 45614 27134 45666
rect 27186 45614 27188 45666
rect 26908 45332 26964 45342
rect 26796 45276 26908 45332
rect 26908 45266 26964 45276
rect 27020 45220 27076 45230
rect 27020 44434 27076 45164
rect 27132 45106 27188 45614
rect 27132 45054 27134 45106
rect 27186 45054 27188 45106
rect 27132 45042 27188 45054
rect 27020 44382 27022 44434
rect 27074 44382 27076 44434
rect 27020 44370 27076 44382
rect 27244 42868 27300 47404
rect 27692 47394 27748 47404
rect 28476 47346 28532 47358
rect 28476 47294 28478 47346
rect 28530 47294 28532 47346
rect 28364 46676 28420 46686
rect 28364 45444 28420 46620
rect 28364 45378 28420 45388
rect 27692 45332 27748 45342
rect 27692 44324 27748 45276
rect 27244 42774 27300 42812
rect 27356 44210 27412 44222
rect 27356 44158 27358 44210
rect 27410 44158 27412 44210
rect 26908 42082 26964 42094
rect 26908 42030 26910 42082
rect 26962 42030 26964 42082
rect 26908 41972 26964 42030
rect 26908 41906 26964 41916
rect 27244 41972 27300 41982
rect 27244 41878 27300 41916
rect 26684 41010 26740 41020
rect 26908 40964 26964 40974
rect 26964 40908 27076 40964
rect 26908 40870 26964 40908
rect 26908 39620 26964 39630
rect 26796 38948 26852 38958
rect 26796 38612 26852 38892
rect 26908 38834 26964 39564
rect 26908 38782 26910 38834
rect 26962 38782 26964 38834
rect 26908 38770 26964 38782
rect 27020 38612 27076 40908
rect 26796 38556 26964 38612
rect 26796 36372 26852 36382
rect 26908 36372 26964 38556
rect 27020 37716 27076 38556
rect 27020 37650 27076 37660
rect 27132 36596 27188 36606
rect 27356 36596 27412 44158
rect 27692 43426 27748 44268
rect 27804 44212 27860 44222
rect 27804 44118 27860 44156
rect 27692 43374 27694 43426
rect 27746 43374 27748 43426
rect 27692 43362 27748 43374
rect 27804 42532 27860 42542
rect 27692 42530 27860 42532
rect 27692 42478 27806 42530
rect 27858 42478 27860 42530
rect 27692 42476 27860 42478
rect 27692 42084 27748 42476
rect 27804 42466 27860 42476
rect 27468 41188 27524 41198
rect 27468 41074 27524 41132
rect 27468 41022 27470 41074
rect 27522 41022 27524 41074
rect 27468 41010 27524 41022
rect 27580 38724 27636 38762
rect 27580 38658 27636 38668
rect 27692 38276 27748 42028
rect 27916 41970 27972 41982
rect 27916 41918 27918 41970
rect 27970 41918 27972 41970
rect 27804 40964 27860 40974
rect 27804 40870 27860 40908
rect 27916 40514 27972 41918
rect 28476 41860 28532 47294
rect 28588 46900 28644 46910
rect 28588 46786 28644 46844
rect 28588 46734 28590 46786
rect 28642 46734 28644 46786
rect 28588 46722 28644 46734
rect 28588 45108 28644 45118
rect 28588 45014 28644 45052
rect 28700 44548 28756 50764
rect 29036 48244 29092 48254
rect 29036 48150 29092 48188
rect 29260 47346 29316 52892
rect 30380 51492 30436 51502
rect 30156 50820 30212 50830
rect 29484 50708 29540 50718
rect 29484 50614 29540 50652
rect 30156 50708 30212 50764
rect 30380 50708 30436 51436
rect 30492 51378 30548 51390
rect 30492 51326 30494 51378
rect 30546 51326 30548 51378
rect 30492 50932 30548 51326
rect 30492 50866 30548 50876
rect 30156 50706 30436 50708
rect 30156 50654 30382 50706
rect 30434 50654 30436 50706
rect 30156 50652 30436 50654
rect 29932 50594 29988 50606
rect 29932 50542 29934 50594
rect 29986 50542 29988 50594
rect 29932 50484 29988 50542
rect 29932 50418 29988 50428
rect 30156 50034 30212 50652
rect 30380 50642 30436 50652
rect 30604 50428 30660 53452
rect 31276 52948 31332 53790
rect 31612 53170 31668 54238
rect 31612 53118 31614 53170
rect 31666 53118 31668 53170
rect 31612 53106 31668 53118
rect 31836 54290 31892 54302
rect 31836 54238 31838 54290
rect 31890 54238 31892 54290
rect 31836 53844 31892 54238
rect 31948 54292 32004 54302
rect 31948 54290 33460 54292
rect 31948 54238 31950 54290
rect 32002 54238 33460 54290
rect 31948 54236 33460 54238
rect 31948 54226 32004 54236
rect 31724 53058 31780 53070
rect 31724 53006 31726 53058
rect 31778 53006 31780 53058
rect 31724 52948 31780 53006
rect 31276 52892 31780 52948
rect 31500 52722 31556 52734
rect 31500 52670 31502 52722
rect 31554 52670 31556 52722
rect 31388 52388 31444 52398
rect 31388 52294 31444 52332
rect 31500 52388 31556 52670
rect 31612 52388 31668 52398
rect 31500 52386 31668 52388
rect 31500 52334 31614 52386
rect 31666 52334 31668 52386
rect 31500 52332 31668 52334
rect 31276 51604 31332 51614
rect 31500 51604 31556 52332
rect 31612 52322 31668 52332
rect 31724 52164 31780 52892
rect 31836 52388 31892 53788
rect 33404 53842 33460 54236
rect 33404 53790 33406 53842
rect 33458 53790 33460 53842
rect 33404 53778 33460 53790
rect 31836 52322 31892 52332
rect 34076 53730 34132 55244
rect 34076 53678 34078 53730
rect 34130 53678 34132 53730
rect 34076 53060 34132 53678
rect 34300 55186 34356 55198
rect 34300 55134 34302 55186
rect 34354 55134 34356 55186
rect 34300 53732 34356 55134
rect 36428 54404 36484 55358
rect 37324 55300 37380 55310
rect 37212 55298 37380 55300
rect 37212 55246 37326 55298
rect 37378 55246 37380 55298
rect 37212 55244 37380 55246
rect 36876 54626 36932 54638
rect 36876 54574 36878 54626
rect 36930 54574 36932 54626
rect 36540 54514 36596 54526
rect 36540 54462 36542 54514
rect 36594 54462 36596 54514
rect 36540 54404 36596 54462
rect 35980 54348 36596 54404
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 35868 53844 35924 53854
rect 35980 53844 36036 54348
rect 35868 53842 36036 53844
rect 35868 53790 35870 53842
rect 35922 53790 36036 53842
rect 35868 53788 36036 53790
rect 36428 53844 36484 53854
rect 35868 53778 35924 53788
rect 34300 53666 34356 53676
rect 36092 53732 36148 53742
rect 36092 53730 36260 53732
rect 36092 53678 36094 53730
rect 36146 53678 36260 53730
rect 36092 53676 36260 53678
rect 36092 53666 36148 53676
rect 35868 53508 35924 53518
rect 31612 52108 31780 52164
rect 31836 52162 31892 52174
rect 31836 52110 31838 52162
rect 31890 52110 31892 52162
rect 31612 51716 31668 52108
rect 31724 51940 31780 51950
rect 31724 51846 31780 51884
rect 31612 51660 31780 51716
rect 31276 51602 31556 51604
rect 31276 51550 31278 51602
rect 31330 51550 31556 51602
rect 31276 51548 31556 51550
rect 31276 51538 31332 51548
rect 30828 51492 30884 51502
rect 30828 51398 30884 51436
rect 30156 49982 30158 50034
rect 30210 49982 30212 50034
rect 30156 49970 30212 49982
rect 30380 50372 30660 50428
rect 30716 51380 30772 51390
rect 30716 50484 30772 51324
rect 31612 51378 31668 51390
rect 31612 51326 31614 51378
rect 31666 51326 31668 51378
rect 30716 50418 30772 50428
rect 30828 51156 30884 51166
rect 30380 50034 30436 50372
rect 30380 49982 30382 50034
rect 30434 49982 30436 50034
rect 30380 49970 30436 49982
rect 30716 49812 30772 49822
rect 30716 49718 30772 49756
rect 29932 49700 29988 49710
rect 29932 49026 29988 49644
rect 29932 48974 29934 49026
rect 29986 48974 29988 49026
rect 29932 48962 29988 48974
rect 30268 49028 30324 49038
rect 29820 48916 29876 48926
rect 29820 48822 29876 48860
rect 29708 47460 29764 47470
rect 29708 47458 29876 47460
rect 29708 47406 29710 47458
rect 29762 47406 29876 47458
rect 29708 47404 29876 47406
rect 29708 47394 29764 47404
rect 29260 47294 29262 47346
rect 29314 47294 29316 47346
rect 29260 47236 29316 47294
rect 29036 47180 29316 47236
rect 29708 47234 29764 47246
rect 29708 47182 29710 47234
rect 29762 47182 29764 47234
rect 29036 45892 29092 47180
rect 29484 46676 29540 46686
rect 29372 46674 29540 46676
rect 29372 46622 29486 46674
rect 29538 46622 29540 46674
rect 29372 46620 29540 46622
rect 29260 46562 29316 46574
rect 29260 46510 29262 46562
rect 29314 46510 29316 46562
rect 29148 45892 29204 45902
rect 29036 45890 29204 45892
rect 29036 45838 29150 45890
rect 29202 45838 29204 45890
rect 29036 45836 29204 45838
rect 29148 45826 29204 45836
rect 29260 45780 29316 46510
rect 29372 46002 29428 46620
rect 29484 46610 29540 46620
rect 29708 46676 29764 47182
rect 29708 46610 29764 46620
rect 29484 46116 29540 46126
rect 29820 46116 29876 47404
rect 30268 47458 30324 48972
rect 30268 47406 30270 47458
rect 30322 47406 30324 47458
rect 30268 47394 30324 47406
rect 30380 48242 30436 48254
rect 30380 48190 30382 48242
rect 30434 48190 30436 48242
rect 30380 47572 30436 48190
rect 30828 48130 30884 51100
rect 31276 50932 31332 50942
rect 31612 50932 31668 51326
rect 31332 50876 31668 50932
rect 31164 50706 31220 50718
rect 31164 50654 31166 50706
rect 31218 50654 31220 50706
rect 31164 50596 31220 50654
rect 31164 50530 31220 50540
rect 30940 50484 30996 50494
rect 30940 49922 30996 50428
rect 30940 49870 30942 49922
rect 30994 49870 30996 49922
rect 30940 49858 30996 49870
rect 31276 49922 31332 50876
rect 31724 50428 31780 51660
rect 31836 51604 31892 52110
rect 32396 51938 32452 51950
rect 32396 51886 32398 51938
rect 32450 51886 32452 51938
rect 31948 51604 32004 51614
rect 31836 51602 32004 51604
rect 31836 51550 31950 51602
rect 32002 51550 32004 51602
rect 31836 51548 32004 51550
rect 31948 51538 32004 51548
rect 32396 51492 32452 51886
rect 32396 51426 32452 51436
rect 33292 51940 33348 51950
rect 31836 51380 31892 51390
rect 31836 51286 31892 51324
rect 32284 51378 32340 51390
rect 32284 51326 32286 51378
rect 32338 51326 32340 51378
rect 32284 50596 32340 51326
rect 33180 51266 33236 51278
rect 33180 51214 33182 51266
rect 33234 51214 33236 51266
rect 32284 50530 32340 50540
rect 32956 50596 33012 50606
rect 33180 50596 33236 51214
rect 33292 50706 33348 51884
rect 33292 50654 33294 50706
rect 33346 50654 33348 50706
rect 33292 50642 33348 50654
rect 34076 51380 34132 53004
rect 35196 53060 35252 53070
rect 35196 52966 35252 53004
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 35868 52388 35924 53452
rect 35532 52386 35924 52388
rect 35532 52334 35870 52386
rect 35922 52334 35924 52386
rect 35532 52332 35924 52334
rect 35532 52274 35588 52332
rect 35868 52322 35924 52332
rect 35532 52222 35534 52274
rect 35586 52222 35588 52274
rect 35532 52210 35588 52222
rect 36092 52164 36148 52174
rect 35980 52162 36148 52164
rect 35980 52110 36094 52162
rect 36146 52110 36148 52162
rect 35980 52108 36148 52110
rect 36204 52164 36260 53676
rect 36428 53730 36484 53788
rect 36428 53678 36430 53730
rect 36482 53678 36484 53730
rect 36428 53666 36484 53678
rect 36876 52276 36932 54574
rect 36988 53732 37044 53742
rect 36988 53638 37044 53676
rect 37100 53730 37156 53742
rect 37100 53678 37102 53730
rect 37154 53678 37156 53730
rect 37100 53508 37156 53678
rect 37100 53442 37156 53452
rect 37100 53060 37156 53070
rect 37212 53060 37268 55244
rect 37324 55234 37380 55244
rect 38108 55188 38164 55198
rect 38108 55094 38164 55132
rect 37436 53956 37492 53966
rect 37436 53954 37604 53956
rect 37436 53902 37438 53954
rect 37490 53902 37604 53954
rect 37436 53900 37604 53902
rect 37436 53890 37492 53900
rect 37548 53844 37604 53900
rect 37548 53778 37604 53788
rect 37156 53004 37268 53060
rect 37324 53730 37380 53742
rect 37324 53678 37326 53730
rect 37378 53678 37380 53730
rect 37100 52994 37156 53004
rect 37324 52386 37380 53678
rect 37324 52334 37326 52386
rect 37378 52334 37380 52386
rect 37324 52322 37380 52334
rect 37884 53508 37940 53518
rect 37996 53508 38052 53518
rect 37940 53506 38052 53508
rect 37940 53454 37998 53506
rect 38050 53454 38052 53506
rect 37940 53452 38052 53454
rect 36876 52220 37268 52276
rect 36316 52164 36372 52174
rect 37212 52164 37268 52220
rect 37324 52164 37380 52174
rect 36204 52162 37044 52164
rect 36204 52110 36318 52162
rect 36370 52110 37044 52162
rect 36204 52108 37044 52110
rect 37212 52162 37492 52164
rect 37212 52110 37326 52162
rect 37378 52110 37492 52162
rect 37212 52108 37492 52110
rect 34972 52052 35028 52062
rect 34972 51490 35028 51996
rect 35756 52052 35812 52062
rect 35756 51958 35812 51996
rect 34972 51438 34974 51490
rect 35026 51438 35028 51490
rect 34972 51426 35028 51438
rect 34188 51380 34244 51390
rect 34076 51378 34244 51380
rect 34076 51326 34190 51378
rect 34242 51326 34244 51378
rect 34076 51324 34244 51326
rect 33012 50540 33236 50596
rect 34076 50594 34132 51324
rect 34188 51314 34244 51324
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 35980 50706 36036 52108
rect 36092 52098 36148 52108
rect 36316 52098 36372 52108
rect 36988 52050 37044 52108
rect 37324 52098 37380 52108
rect 36988 51998 36990 52050
rect 37042 51998 37044 52050
rect 36988 51940 37044 51998
rect 36988 51884 37268 51940
rect 37100 51268 37156 51278
rect 35980 50654 35982 50706
rect 36034 50654 36036 50706
rect 35980 50642 36036 50654
rect 36540 51266 37156 51268
rect 36540 51214 37102 51266
rect 37154 51214 37156 51266
rect 36540 51212 37156 51214
rect 34076 50542 34078 50594
rect 34130 50542 34132 50594
rect 31276 49870 31278 49922
rect 31330 49870 31332 49922
rect 31276 49858 31332 49870
rect 31388 50372 31780 50428
rect 31388 49810 31444 50372
rect 31388 49758 31390 49810
rect 31442 49758 31444 49810
rect 31276 49700 31332 49710
rect 31388 49700 31444 49758
rect 31332 49644 31444 49700
rect 31948 49812 32004 49822
rect 31948 49698 32004 49756
rect 31948 49646 31950 49698
rect 32002 49646 32004 49698
rect 31276 49634 31332 49644
rect 31948 48804 32004 49646
rect 31948 48738 32004 48748
rect 32060 48354 32116 48366
rect 32060 48302 32062 48354
rect 32114 48302 32116 48354
rect 30828 48078 30830 48130
rect 30882 48078 30884 48130
rect 30828 48066 30884 48078
rect 31836 48242 31892 48254
rect 31836 48190 31838 48242
rect 31890 48190 31892 48242
rect 30380 47346 30436 47516
rect 30380 47294 30382 47346
rect 30434 47294 30436 47346
rect 30380 47282 30436 47294
rect 30940 48018 30996 48030
rect 30940 47966 30942 48018
rect 30994 47966 30996 48018
rect 30940 46786 30996 47966
rect 31836 47570 31892 48190
rect 32060 47684 32116 48302
rect 32060 47618 32116 47628
rect 32172 48242 32228 48254
rect 32172 48190 32174 48242
rect 32226 48190 32228 48242
rect 31836 47518 31838 47570
rect 31890 47518 31892 47570
rect 31836 47506 31892 47518
rect 30940 46734 30942 46786
rect 30994 46734 30996 46786
rect 30940 46722 30996 46734
rect 31164 47458 31220 47470
rect 31164 47406 31166 47458
rect 31218 47406 31220 47458
rect 29484 46114 29876 46116
rect 29484 46062 29486 46114
rect 29538 46062 29822 46114
rect 29874 46062 29876 46114
rect 29484 46060 29876 46062
rect 29484 46050 29540 46060
rect 29820 46050 29876 46060
rect 29372 45950 29374 46002
rect 29426 45950 29428 46002
rect 29372 45938 29428 45950
rect 31164 46004 31220 47406
rect 31500 46676 31556 46686
rect 31500 46582 31556 46620
rect 31164 46002 31332 46004
rect 31164 45950 31166 46002
rect 31218 45950 31332 46002
rect 31164 45948 31332 45950
rect 31164 45938 31220 45948
rect 29260 45724 29652 45780
rect 29596 45106 29652 45724
rect 29596 45054 29598 45106
rect 29650 45054 29652 45106
rect 29596 45042 29652 45054
rect 29932 45778 29988 45790
rect 29932 45726 29934 45778
rect 29986 45726 29988 45778
rect 29932 45108 29988 45726
rect 29932 45042 29988 45052
rect 30156 44996 30212 45006
rect 30156 44994 30660 44996
rect 30156 44942 30158 44994
rect 30210 44942 30660 44994
rect 30156 44940 30660 44942
rect 30156 44930 30212 44940
rect 28476 41794 28532 41804
rect 28588 44492 28756 44548
rect 30044 44882 30100 44894
rect 30044 44830 30046 44882
rect 30098 44830 30100 44882
rect 27916 40462 27918 40514
rect 27970 40462 27972 40514
rect 27916 39620 27972 40462
rect 28140 41076 28196 41086
rect 28140 39730 28196 41020
rect 28140 39678 28142 39730
rect 28194 39678 28196 39730
rect 28140 39666 28196 39678
rect 27916 39554 27972 39564
rect 28588 38668 28644 44492
rect 29820 43652 29876 43662
rect 30044 43652 30100 44830
rect 30380 44772 30436 44782
rect 30268 44324 30324 44334
rect 30268 44230 30324 44268
rect 29820 43650 30100 43652
rect 29820 43598 29822 43650
rect 29874 43598 30100 43650
rect 29820 43596 30100 43598
rect 29820 43586 29876 43596
rect 29932 42756 29988 42766
rect 30380 42756 30436 44716
rect 30604 44434 30660 44940
rect 30604 44382 30606 44434
rect 30658 44382 30660 44434
rect 30604 44370 30660 44382
rect 30940 44324 30996 44334
rect 30940 44322 31108 44324
rect 30940 44270 30942 44322
rect 30994 44270 31108 44322
rect 30940 44268 31108 44270
rect 30940 44258 30996 44268
rect 30492 44100 30548 44110
rect 30492 44098 30660 44100
rect 30492 44046 30494 44098
rect 30546 44046 30660 44098
rect 30492 44044 30660 44046
rect 30492 44034 30548 44044
rect 30604 43764 30660 44044
rect 30716 44098 30772 44110
rect 30716 44046 30718 44098
rect 30770 44046 30772 44098
rect 30716 43988 30772 44046
rect 30716 43922 30772 43932
rect 30604 43708 30884 43764
rect 30604 43550 30660 43562
rect 30604 43498 30606 43550
rect 30658 43540 30660 43550
rect 30716 43540 30772 43550
rect 30658 43498 30716 43540
rect 30604 43484 30716 43498
rect 30716 43474 30772 43484
rect 30828 43316 30884 43708
rect 30604 42756 30660 42766
rect 30828 42756 30884 43260
rect 30380 42754 30772 42756
rect 30380 42702 30606 42754
rect 30658 42702 30772 42754
rect 30380 42700 30772 42702
rect 29260 42644 29316 42654
rect 29260 42550 29316 42588
rect 29932 42642 29988 42700
rect 30604 42690 30660 42700
rect 29932 42590 29934 42642
rect 29986 42590 29988 42642
rect 29932 42578 29988 42590
rect 29148 42532 29204 42542
rect 29596 42532 29652 42542
rect 28700 42530 29204 42532
rect 28700 42478 29150 42530
rect 29202 42478 29204 42530
rect 28700 42476 29204 42478
rect 28700 42082 28756 42476
rect 29148 42466 29204 42476
rect 29372 42530 29652 42532
rect 29372 42478 29598 42530
rect 29650 42478 29652 42530
rect 29372 42476 29652 42478
rect 28700 42030 28702 42082
rect 28754 42030 28756 42082
rect 28700 42018 28756 42030
rect 29372 41972 29428 42476
rect 29596 42466 29652 42476
rect 30492 42532 30548 42542
rect 29372 41298 29428 41916
rect 29372 41246 29374 41298
rect 29426 41246 29428 41298
rect 29372 41234 29428 41246
rect 30492 41972 30548 42476
rect 29484 41076 29540 41086
rect 29484 40982 29540 41020
rect 30156 41076 30212 41086
rect 30156 40982 30212 41020
rect 30492 41074 30548 41916
rect 30716 41860 30772 42700
rect 31052 42756 31108 44268
rect 31164 43876 31220 43886
rect 31164 43762 31220 43820
rect 31164 43710 31166 43762
rect 31218 43710 31220 43762
rect 31164 43698 31220 43710
rect 31276 43540 31332 45948
rect 32172 45780 32228 48190
rect 31500 45724 32228 45780
rect 32284 48132 32340 48142
rect 31388 45444 31444 45454
rect 31388 44436 31444 45388
rect 31500 45218 31556 45724
rect 31500 45166 31502 45218
rect 31554 45166 31556 45218
rect 31500 45154 31556 45166
rect 32172 45108 32228 45118
rect 32284 45108 32340 48076
rect 32172 45106 32340 45108
rect 32172 45054 32174 45106
rect 32226 45054 32340 45106
rect 32172 45052 32340 45054
rect 32172 45042 32228 45052
rect 32396 44996 32452 45006
rect 32284 44660 32340 44670
rect 32172 44604 32284 44660
rect 31500 44436 31556 44446
rect 31388 44434 31556 44436
rect 31388 44382 31502 44434
rect 31554 44382 31556 44434
rect 31388 44380 31556 44382
rect 31500 43652 31556 44380
rect 32172 43762 32228 44604
rect 32284 44594 32340 44604
rect 32172 43710 32174 43762
rect 32226 43710 32228 43762
rect 32172 43698 32228 43710
rect 32396 43764 32452 44940
rect 32396 43708 32900 43764
rect 31836 43652 31892 43662
rect 31500 43650 31892 43652
rect 31500 43598 31838 43650
rect 31890 43598 31892 43650
rect 31500 43596 31892 43598
rect 31836 43586 31892 43596
rect 31276 43474 31332 43484
rect 32060 43538 32116 43550
rect 32060 43486 32062 43538
rect 32114 43486 32116 43538
rect 32060 43316 32116 43486
rect 31276 42756 31332 42766
rect 31052 42700 31276 42756
rect 30828 42662 30884 42700
rect 31276 42662 31332 42700
rect 30940 42644 30996 42654
rect 30940 42550 30996 42588
rect 31052 42530 31108 42542
rect 31836 42532 31892 42542
rect 31052 42478 31054 42530
rect 31106 42478 31108 42530
rect 31052 42420 31108 42478
rect 31724 42530 31892 42532
rect 31724 42478 31838 42530
rect 31890 42478 31892 42530
rect 31724 42476 31892 42478
rect 31724 42420 31780 42476
rect 31836 42466 31892 42476
rect 31052 42364 31780 42420
rect 30828 41860 30884 41870
rect 30716 41858 30884 41860
rect 30716 41806 30830 41858
rect 30882 41806 30884 41858
rect 30716 41804 30884 41806
rect 30828 41794 30884 41804
rect 31388 41860 31444 41870
rect 31388 41298 31444 41804
rect 31388 41246 31390 41298
rect 31442 41246 31444 41298
rect 31388 41234 31444 41246
rect 30492 41022 30494 41074
rect 30546 41022 30548 41074
rect 30492 41010 30548 41022
rect 28700 40962 28756 40974
rect 28700 40910 28702 40962
rect 28754 40910 28756 40962
rect 28700 40852 28756 40910
rect 28700 40786 28756 40796
rect 29260 40962 29316 40974
rect 29260 40910 29262 40962
rect 29314 40910 29316 40962
rect 29260 40852 29316 40910
rect 29260 40786 29316 40796
rect 29036 40404 29092 40414
rect 29036 40310 29092 40348
rect 29708 39844 29764 39854
rect 29708 39730 29764 39788
rect 29708 39678 29710 39730
rect 29762 39678 29764 39730
rect 29708 39666 29764 39678
rect 30268 39844 30324 39854
rect 29260 39508 29316 39518
rect 29260 39506 29652 39508
rect 29260 39454 29262 39506
rect 29314 39454 29652 39506
rect 29260 39452 29652 39454
rect 29260 39442 29316 39452
rect 29148 39396 29204 39406
rect 29148 39302 29204 39340
rect 29596 38724 29652 39452
rect 30268 38948 30324 39788
rect 30156 38946 30324 38948
rect 30156 38894 30270 38946
rect 30322 38894 30324 38946
rect 30156 38892 30324 38894
rect 29708 38724 29764 38734
rect 29596 38722 29764 38724
rect 29596 38670 29710 38722
rect 29762 38670 29764 38722
rect 29596 38668 29764 38670
rect 28588 38612 28868 38668
rect 29708 38658 29764 38668
rect 27132 36594 27412 36596
rect 27132 36542 27134 36594
rect 27186 36542 27412 36594
rect 27132 36540 27412 36542
rect 27132 36530 27188 36540
rect 27356 36482 27412 36540
rect 27356 36430 27358 36482
rect 27410 36430 27412 36482
rect 27356 36418 27412 36430
rect 27468 38220 27748 38276
rect 26908 36316 27300 36372
rect 26572 36260 26628 36270
rect 26572 35810 26628 36204
rect 26572 35758 26574 35810
rect 26626 35758 26628 35810
rect 26572 35746 26628 35758
rect 26348 35700 26404 35710
rect 26348 35606 26404 35644
rect 26684 35700 26740 35710
rect 26684 35476 26740 35644
rect 26684 35410 26740 35420
rect 26012 34914 26292 34916
rect 26012 34862 26014 34914
rect 26066 34862 26292 34914
rect 26012 34860 26292 34862
rect 26012 34850 26068 34860
rect 25788 34692 25844 34702
rect 25788 34598 25844 34636
rect 26460 34692 26516 34702
rect 26460 34132 26516 34636
rect 26796 34356 26852 36316
rect 27020 35588 27076 35598
rect 27076 35532 27188 35588
rect 27020 35494 27076 35532
rect 26796 34300 26964 34356
rect 26684 34132 26740 34142
rect 26460 34130 26740 34132
rect 26460 34078 26686 34130
rect 26738 34078 26740 34130
rect 26460 34076 26740 34078
rect 26684 34020 26740 34076
rect 26684 33954 26740 33964
rect 26908 33908 26964 34300
rect 25228 32786 25396 32788
rect 25228 32734 25230 32786
rect 25282 32734 25396 32786
rect 25228 32732 25396 32734
rect 26796 33852 26964 33908
rect 25116 30996 25172 31006
rect 25228 30996 25284 32732
rect 25676 32674 25732 32686
rect 25676 32622 25678 32674
rect 25730 32622 25732 32674
rect 25452 32562 25508 32574
rect 25452 32510 25454 32562
rect 25506 32510 25508 32562
rect 25340 32450 25396 32462
rect 25340 32398 25342 32450
rect 25394 32398 25396 32450
rect 25340 32004 25396 32398
rect 25340 31938 25396 31948
rect 25340 30996 25396 31006
rect 25228 30994 25396 30996
rect 25228 30942 25342 30994
rect 25394 30942 25396 30994
rect 25228 30940 25396 30942
rect 25116 30434 25172 30940
rect 25340 30930 25396 30940
rect 25452 30996 25508 32510
rect 25676 31218 25732 32622
rect 26348 32452 26404 32462
rect 26348 32358 26404 32396
rect 26236 31890 26292 31902
rect 26236 31838 26238 31890
rect 26290 31838 26292 31890
rect 26236 31332 26292 31838
rect 26796 31780 26852 33852
rect 26796 31714 26852 31724
rect 25676 31166 25678 31218
rect 25730 31166 25732 31218
rect 25676 31154 25732 31166
rect 25900 31276 26292 31332
rect 25452 30930 25508 30940
rect 25788 30996 25844 31006
rect 25900 30996 25956 31276
rect 25844 30940 25956 30996
rect 26012 30996 26068 31006
rect 26012 30994 26292 30996
rect 26012 30942 26014 30994
rect 26066 30942 26292 30994
rect 26012 30940 26292 30942
rect 25788 30902 25844 30940
rect 26012 30930 26068 30940
rect 25116 30382 25118 30434
rect 25170 30382 25172 30434
rect 25116 30370 25172 30382
rect 24892 30324 24948 30334
rect 24668 30322 24948 30324
rect 24668 30270 24894 30322
rect 24946 30270 24948 30322
rect 24668 30268 24948 30270
rect 24892 30258 24948 30268
rect 26236 30322 26292 30940
rect 26572 30884 26628 30894
rect 26236 30270 26238 30322
rect 26290 30270 26292 30322
rect 24556 30212 24612 30222
rect 23772 30210 24612 30212
rect 23772 30158 24558 30210
rect 24610 30158 24612 30210
rect 23772 30156 24612 30158
rect 23548 28980 23604 28990
rect 22764 28478 22766 28530
rect 22818 28478 22820 28530
rect 22764 28466 22820 28478
rect 23100 28642 23156 28654
rect 23100 28590 23102 28642
rect 23154 28590 23156 28642
rect 22428 28252 22932 28308
rect 22092 28028 22372 28084
rect 22092 27188 22148 28028
rect 22092 27186 22484 27188
rect 22092 27134 22094 27186
rect 22146 27134 22484 27186
rect 22092 27132 22484 27134
rect 22092 27122 22148 27132
rect 22428 26964 22484 27132
rect 22764 27074 22820 27086
rect 22764 27022 22766 27074
rect 22818 27022 22820 27074
rect 22428 26962 22708 26964
rect 22428 26910 22430 26962
rect 22482 26910 22708 26962
rect 22428 26908 22708 26910
rect 21868 26852 22036 26908
rect 22428 26898 22484 26908
rect 21980 23940 22036 26852
rect 22204 26852 22260 26862
rect 22204 26178 22260 26796
rect 22204 26126 22206 26178
rect 22258 26126 22260 26178
rect 22204 26114 22260 26126
rect 22652 25620 22708 26908
rect 22764 26852 22820 27022
rect 22876 26908 22932 28252
rect 23100 28084 23156 28590
rect 23548 28642 23604 28924
rect 23548 28590 23550 28642
rect 23602 28590 23604 28642
rect 23548 28578 23604 28590
rect 23772 28530 23828 30156
rect 24556 30146 24612 30156
rect 26236 30212 26292 30270
rect 26236 30146 26292 30156
rect 26460 30882 26628 30884
rect 26460 30830 26574 30882
rect 26626 30830 26628 30882
rect 26460 30828 26628 30830
rect 24668 30100 24724 30110
rect 24668 30006 24724 30044
rect 26460 30100 26516 30828
rect 26572 30818 26628 30828
rect 27132 30548 27188 35532
rect 27244 34692 27300 36316
rect 27244 34690 27412 34692
rect 27244 34638 27246 34690
rect 27298 34638 27412 34690
rect 27244 34636 27412 34638
rect 27244 34626 27300 34636
rect 27244 34468 27300 34478
rect 27244 34020 27300 34412
rect 27356 34132 27412 34636
rect 27468 34356 27524 38220
rect 28028 38164 28084 38174
rect 28028 38070 28084 38108
rect 27580 38050 27636 38062
rect 27580 37998 27582 38050
rect 27634 37998 27636 38050
rect 27580 37492 27636 37998
rect 28700 37940 28756 37950
rect 28700 37846 28756 37884
rect 28700 37492 28756 37502
rect 27580 37044 27636 37436
rect 28588 37436 28700 37492
rect 28252 37156 28308 37166
rect 27916 37154 28308 37156
rect 27916 37102 28254 37154
rect 28306 37102 28308 37154
rect 27916 37100 28308 37102
rect 27916 37044 27972 37100
rect 28252 37090 28308 37100
rect 27580 36988 27972 37044
rect 27580 36260 27636 36270
rect 27580 36166 27636 36204
rect 27692 36148 27748 36988
rect 28028 36484 28084 36494
rect 28588 36484 28644 37436
rect 28700 37426 28756 37436
rect 28700 37268 28756 37278
rect 28700 37174 28756 37212
rect 28028 36482 28644 36484
rect 28028 36430 28030 36482
rect 28082 36430 28644 36482
rect 28028 36428 28644 36430
rect 28028 36418 28084 36428
rect 27804 36370 27860 36382
rect 27804 36318 27806 36370
rect 27858 36318 27860 36370
rect 27804 36260 27860 36318
rect 28476 36260 28532 36270
rect 27804 36258 28532 36260
rect 27804 36206 28478 36258
rect 28530 36206 28532 36258
rect 27804 36204 28532 36206
rect 27692 36092 27860 36148
rect 27692 35812 27748 35822
rect 27692 35718 27748 35756
rect 27468 34300 27748 34356
rect 27580 34132 27636 34142
rect 27356 34130 27636 34132
rect 27356 34078 27582 34130
rect 27634 34078 27636 34130
rect 27356 34076 27636 34078
rect 27244 34018 27412 34020
rect 27244 33966 27246 34018
rect 27298 33966 27412 34018
rect 27244 33964 27412 33966
rect 27244 33954 27300 33964
rect 27356 30772 27412 33964
rect 27468 33346 27524 33358
rect 27468 33294 27470 33346
rect 27522 33294 27524 33346
rect 27468 31108 27524 33294
rect 27580 33012 27636 34076
rect 27692 33572 27748 34300
rect 27692 33506 27748 33516
rect 27692 33236 27748 33246
rect 27804 33236 27860 36092
rect 28028 35700 28084 35710
rect 28364 35700 28420 35710
rect 28028 35698 28420 35700
rect 28028 35646 28030 35698
rect 28082 35646 28366 35698
rect 28418 35646 28420 35698
rect 28028 35644 28420 35646
rect 28028 35138 28084 35644
rect 28364 35634 28420 35644
rect 28028 35086 28030 35138
rect 28082 35086 28084 35138
rect 28028 35074 28084 35086
rect 28364 35140 28420 35150
rect 28364 35046 28420 35084
rect 27692 33234 27860 33236
rect 27692 33182 27694 33234
rect 27746 33182 27860 33234
rect 27692 33180 27860 33182
rect 27916 34242 27972 34254
rect 27916 34190 27918 34242
rect 27970 34190 27972 34242
rect 27916 34020 27972 34190
rect 28364 34020 28420 34030
rect 27972 34018 28420 34020
rect 27972 33966 28366 34018
rect 28418 33966 28420 34018
rect 27972 33964 28420 33966
rect 27692 33170 27748 33180
rect 27580 32956 27748 33012
rect 27580 32564 27636 32574
rect 27580 32470 27636 32508
rect 27468 31042 27524 31052
rect 27356 30706 27412 30716
rect 27468 30884 27524 30894
rect 27132 30492 27412 30548
rect 24444 29988 24500 29998
rect 24220 29986 24500 29988
rect 24220 29934 24446 29986
rect 24498 29934 24500 29986
rect 24220 29932 24500 29934
rect 24220 29314 24276 29932
rect 24220 29262 24222 29314
rect 24274 29262 24276 29314
rect 24220 29250 24276 29262
rect 24444 29316 24500 29932
rect 26460 29538 26516 30044
rect 26460 29486 26462 29538
rect 26514 29486 26516 29538
rect 26460 29474 26516 29486
rect 27244 29426 27300 29438
rect 27244 29374 27246 29426
rect 27298 29374 27300 29426
rect 24444 28642 24500 29260
rect 25228 29316 25284 29326
rect 25228 29222 25284 29260
rect 25340 29204 25396 29214
rect 26572 29204 26628 29214
rect 26908 29204 26964 29214
rect 25340 29202 26068 29204
rect 25340 29150 25342 29202
rect 25394 29150 26068 29202
rect 25340 29148 26068 29150
rect 25340 29138 25396 29148
rect 26012 28866 26068 29148
rect 26572 29202 26964 29204
rect 26572 29150 26574 29202
rect 26626 29150 26910 29202
rect 26962 29150 26964 29202
rect 26572 29148 26964 29150
rect 26572 29138 26628 29148
rect 26908 29138 26964 29148
rect 26012 28814 26014 28866
rect 26066 28814 26068 28866
rect 26012 28802 26068 28814
rect 26572 28868 26628 28878
rect 24444 28590 24446 28642
rect 24498 28590 24500 28642
rect 24444 28578 24500 28590
rect 26348 28756 26404 28766
rect 26348 28642 26404 28700
rect 26572 28754 26628 28812
rect 27244 28868 27300 29374
rect 27356 29426 27412 30492
rect 27468 29650 27524 30828
rect 27468 29598 27470 29650
rect 27522 29598 27524 29650
rect 27468 29586 27524 29598
rect 27356 29374 27358 29426
rect 27410 29374 27412 29426
rect 27356 29204 27412 29374
rect 27356 29138 27412 29148
rect 27580 29426 27636 29438
rect 27580 29374 27582 29426
rect 27634 29374 27636 29426
rect 27244 28774 27300 28812
rect 26572 28702 26574 28754
rect 26626 28702 26628 28754
rect 26572 28690 26628 28702
rect 27356 28644 27412 28654
rect 27580 28644 27636 29374
rect 26348 28590 26350 28642
rect 26402 28590 26404 28642
rect 26348 28578 26404 28590
rect 26908 28588 27356 28644
rect 27412 28588 27636 28644
rect 23772 28478 23774 28530
rect 23826 28478 23828 28530
rect 23772 28466 23828 28478
rect 23884 28532 23940 28542
rect 23100 28018 23156 28028
rect 23548 28418 23604 28430
rect 23548 28366 23550 28418
rect 23602 28366 23604 28418
rect 22876 26852 23044 26908
rect 23436 26852 23492 26862
rect 22764 26786 22820 26796
rect 22876 26290 22932 26302
rect 22876 26238 22878 26290
rect 22930 26238 22932 26290
rect 22876 25732 22932 26238
rect 22988 26292 23044 26852
rect 23212 26850 23492 26852
rect 23212 26798 23438 26850
rect 23490 26798 23492 26850
rect 23212 26796 23492 26798
rect 23100 26292 23156 26302
rect 22988 26290 23156 26292
rect 22988 26238 23102 26290
rect 23154 26238 23156 26290
rect 22988 26236 23156 26238
rect 23100 26226 23156 26236
rect 22876 25676 23156 25732
rect 22652 25618 23044 25620
rect 22652 25566 22654 25618
rect 22706 25566 23044 25618
rect 22652 25564 23044 25566
rect 22652 25554 22708 25564
rect 22988 25506 23044 25564
rect 22988 25454 22990 25506
rect 23042 25454 23044 25506
rect 22988 25442 23044 25454
rect 22204 25060 22260 25070
rect 22204 24722 22260 25004
rect 22204 24670 22206 24722
rect 22258 24670 22260 24722
rect 22204 24658 22260 24670
rect 22876 24500 22932 24510
rect 21980 23874 22036 23884
rect 22316 24052 22372 24062
rect 22316 23938 22372 23996
rect 22316 23886 22318 23938
rect 22370 23886 22372 23938
rect 22316 23874 22372 23886
rect 22764 23938 22820 23950
rect 22764 23886 22766 23938
rect 22818 23886 22820 23938
rect 22092 23826 22148 23838
rect 22092 23774 22094 23826
rect 22146 23774 22148 23826
rect 21644 23716 21700 23726
rect 21532 23714 21700 23716
rect 21532 23662 21646 23714
rect 21698 23662 21700 23714
rect 21532 23660 21700 23662
rect 21532 23156 21588 23660
rect 21644 23650 21700 23660
rect 22092 23716 22148 23774
rect 22204 23828 22260 23838
rect 22204 23734 22260 23772
rect 22092 23650 22148 23660
rect 21980 23604 22036 23614
rect 21980 23378 22036 23548
rect 21980 23326 21982 23378
rect 22034 23326 22036 23378
rect 21980 23314 22036 23326
rect 21532 23090 21588 23100
rect 21644 23266 21700 23278
rect 21644 23214 21646 23266
rect 21698 23214 21700 23266
rect 21644 22372 21700 23214
rect 22764 23156 22820 23886
rect 22764 22596 22820 23100
rect 22876 23154 22932 24444
rect 23100 24276 23156 25676
rect 23212 25172 23268 26796
rect 23436 26786 23492 26796
rect 23436 25618 23492 25630
rect 23436 25566 23438 25618
rect 23490 25566 23492 25618
rect 23324 25396 23380 25406
rect 23324 25302 23380 25340
rect 23212 25116 23380 25172
rect 23100 24210 23156 24220
rect 23212 24948 23268 24958
rect 22876 23102 22878 23154
rect 22930 23102 22932 23154
rect 22876 23090 22932 23102
rect 23212 23604 23268 24892
rect 23212 23154 23268 23548
rect 23212 23102 23214 23154
rect 23266 23102 23268 23154
rect 23212 23090 23268 23102
rect 23324 23938 23380 25116
rect 23436 24724 23492 25566
rect 23548 24948 23604 28366
rect 23884 27970 23940 28476
rect 26684 28532 26740 28542
rect 26908 28532 26964 28588
rect 27356 28550 27412 28588
rect 26684 28530 26964 28532
rect 26684 28478 26686 28530
rect 26738 28478 26964 28530
rect 26684 28476 26964 28478
rect 26684 28466 26740 28476
rect 25788 28420 25844 28430
rect 25788 28082 25844 28364
rect 26460 28420 26516 28430
rect 26460 28326 26516 28364
rect 27244 28418 27300 28430
rect 27692 28420 27748 32956
rect 27916 31556 27972 33964
rect 28364 33954 28420 33964
rect 28252 33124 28308 33134
rect 28140 33122 28308 33124
rect 28140 33070 28254 33122
rect 28306 33070 28308 33122
rect 28140 33068 28308 33070
rect 28028 31556 28084 31566
rect 27916 31500 28028 31556
rect 28028 31490 28084 31500
rect 27916 31108 27972 31118
rect 28140 31108 28196 33068
rect 28252 33058 28308 33068
rect 28252 32450 28308 32462
rect 28252 32398 28254 32450
rect 28306 32398 28308 32450
rect 28252 32116 28308 32398
rect 28252 32050 28308 32060
rect 28476 31892 28532 36204
rect 28588 35924 28644 36428
rect 28700 35924 28756 35934
rect 28588 35922 28756 35924
rect 28588 35870 28702 35922
rect 28754 35870 28756 35922
rect 28588 35868 28756 35870
rect 28700 35858 28756 35868
rect 27972 31052 28196 31108
rect 28252 31836 28532 31892
rect 28588 34914 28644 34926
rect 28588 34862 28590 34914
rect 28642 34862 28644 34914
rect 27916 30324 27972 31052
rect 27244 28366 27246 28418
rect 27298 28366 27300 28418
rect 27244 28084 27300 28366
rect 27468 28364 27748 28420
rect 27804 28418 27860 28430
rect 27804 28366 27806 28418
rect 27858 28366 27860 28418
rect 25788 28030 25790 28082
rect 25842 28030 25844 28082
rect 25788 28018 25844 28030
rect 27020 28028 27300 28084
rect 27356 28196 27412 28206
rect 27356 28082 27412 28140
rect 27356 28030 27358 28082
rect 27410 28030 27412 28082
rect 23884 27918 23886 27970
rect 23938 27918 23940 27970
rect 23884 27906 23940 27918
rect 26012 27860 26068 27870
rect 26012 27766 26068 27804
rect 26572 27860 26628 27870
rect 24332 27746 24388 27758
rect 24332 27694 24334 27746
rect 24386 27694 24388 27746
rect 23996 27634 24052 27646
rect 23996 27582 23998 27634
rect 24050 27582 24052 27634
rect 23996 27076 24052 27582
rect 23996 27010 24052 27020
rect 24108 27074 24164 27086
rect 24108 27022 24110 27074
rect 24162 27022 24164 27074
rect 24108 26402 24164 27022
rect 24332 26908 24388 27694
rect 25564 27748 25620 27758
rect 25564 27654 25620 27692
rect 25900 27746 25956 27758
rect 25900 27694 25902 27746
rect 25954 27694 25956 27746
rect 24444 27636 24500 27646
rect 24444 27542 24500 27580
rect 25340 27636 25396 27646
rect 25340 27542 25396 27580
rect 25900 27300 25956 27694
rect 25788 27244 25956 27300
rect 26124 27748 26180 27758
rect 25564 27188 25620 27198
rect 25564 26964 25620 27132
rect 25676 26964 25732 26974
rect 25564 26962 25732 26964
rect 25564 26910 25678 26962
rect 25730 26910 25732 26962
rect 25564 26908 25732 26910
rect 24108 26350 24110 26402
rect 24162 26350 24164 26402
rect 24108 26338 24164 26350
rect 24220 26852 24388 26908
rect 25676 26898 25732 26908
rect 24220 26178 24276 26796
rect 25788 26404 25844 27244
rect 25900 27076 25956 27086
rect 25900 26982 25956 27020
rect 26124 27076 26180 27692
rect 25788 26338 25844 26348
rect 26012 26964 26068 26974
rect 24332 26292 24388 26302
rect 25452 26292 25508 26302
rect 24332 26198 24388 26236
rect 25228 26236 25452 26292
rect 24220 26126 24222 26178
rect 24274 26126 24276 26178
rect 24220 26114 24276 26126
rect 25228 25618 25284 26236
rect 25452 26198 25508 26236
rect 25564 26068 25620 26078
rect 25900 26068 25956 26078
rect 25564 26066 25956 26068
rect 25564 26014 25566 26066
rect 25618 26014 25902 26066
rect 25954 26014 25956 26066
rect 25564 26012 25956 26014
rect 25564 26002 25620 26012
rect 25900 26002 25956 26012
rect 26012 25844 26068 26908
rect 26124 26290 26180 27020
rect 26348 26516 26404 26526
rect 26348 26422 26404 26460
rect 26572 26514 26628 27804
rect 26796 27748 26852 27758
rect 27020 27748 27076 28028
rect 27356 28018 27412 28030
rect 26796 27746 27076 27748
rect 26796 27694 26798 27746
rect 26850 27694 27076 27746
rect 26796 27692 27076 27694
rect 26796 27682 26852 27692
rect 26796 27076 26852 27086
rect 26796 26982 26852 27020
rect 27020 26964 27076 27692
rect 27132 27860 27188 27870
rect 27132 27074 27188 27804
rect 27132 27022 27134 27074
rect 27186 27022 27188 27074
rect 27132 27010 27188 27022
rect 27356 27748 27412 27758
rect 27356 26908 27412 27692
rect 27020 26898 27076 26908
rect 26572 26462 26574 26514
rect 26626 26462 26628 26514
rect 26572 26450 26628 26462
rect 27244 26852 27412 26908
rect 27244 26516 27300 26852
rect 27244 26422 27300 26460
rect 26124 26238 26126 26290
rect 26178 26238 26180 26290
rect 26124 26226 26180 26238
rect 26460 26180 26516 26190
rect 26460 26086 26516 26124
rect 27356 26180 27412 26190
rect 25228 25566 25230 25618
rect 25282 25566 25284 25618
rect 25228 25554 25284 25566
rect 25900 25788 26068 25844
rect 23548 24882 23604 24892
rect 24220 25172 24276 25182
rect 24108 24834 24164 24846
rect 24108 24782 24110 24834
rect 24162 24782 24164 24834
rect 24108 24724 24164 24782
rect 23436 24668 24164 24724
rect 24220 24834 24276 25116
rect 24220 24782 24222 24834
rect 24274 24782 24276 24834
rect 23324 23886 23326 23938
rect 23378 23886 23380 23938
rect 23324 22932 23380 23886
rect 23660 24052 23716 24062
rect 23660 23938 23716 23996
rect 23660 23886 23662 23938
rect 23714 23886 23716 23938
rect 23660 23874 23716 23886
rect 22540 22540 22820 22596
rect 23100 22876 23380 22932
rect 23772 23828 23828 23838
rect 23884 23828 23940 24668
rect 24108 24500 24164 24510
rect 24108 24406 24164 24444
rect 23828 23826 23940 23828
rect 23828 23774 23886 23826
rect 23938 23774 23940 23826
rect 23828 23772 23940 23774
rect 21644 22306 21700 22316
rect 22428 22484 22484 22494
rect 22540 22484 22596 22540
rect 22484 22428 22596 22484
rect 22428 21586 22484 22428
rect 22428 21534 22430 21586
rect 22482 21534 22484 21586
rect 22428 21522 22484 21534
rect 22652 22372 22708 22382
rect 22652 22146 22708 22316
rect 23100 22370 23156 22876
rect 23100 22318 23102 22370
rect 23154 22318 23156 22370
rect 23100 22306 23156 22318
rect 23772 22258 23828 23772
rect 23884 23762 23940 23772
rect 23996 24164 24052 24174
rect 23996 23714 24052 24108
rect 24220 23940 24276 24782
rect 23996 23662 23998 23714
rect 24050 23662 24052 23714
rect 23996 23650 24052 23662
rect 24108 23938 24276 23940
rect 24108 23886 24222 23938
rect 24274 23886 24276 23938
rect 24108 23884 24276 23886
rect 24108 23716 24164 23884
rect 24220 23874 24276 23884
rect 23884 23156 23940 23166
rect 23884 23062 23940 23100
rect 23996 22372 24052 22382
rect 24108 22372 24164 23660
rect 23996 22370 24164 22372
rect 23996 22318 23998 22370
rect 24050 22318 24164 22370
rect 23996 22316 24164 22318
rect 24556 23156 24612 23166
rect 23996 22306 24052 22316
rect 23772 22206 23774 22258
rect 23826 22206 23828 22258
rect 23772 22194 23828 22206
rect 22652 22094 22654 22146
rect 22706 22094 22708 22146
rect 22652 21586 22708 22094
rect 23436 22146 23492 22158
rect 23436 22094 23438 22146
rect 23490 22094 23492 22146
rect 23436 21812 23492 22094
rect 23548 21812 23604 21822
rect 23436 21810 23604 21812
rect 23436 21758 23550 21810
rect 23602 21758 23604 21810
rect 23436 21756 23604 21758
rect 22652 21534 22654 21586
rect 22706 21534 22708 21586
rect 22652 21522 22708 21534
rect 22988 21588 23044 21598
rect 22652 21028 22708 21038
rect 22652 20934 22708 20972
rect 22988 20914 23044 21532
rect 22988 20862 22990 20914
rect 23042 20862 23044 20914
rect 22988 20850 23044 20862
rect 23212 21476 23268 21486
rect 23212 21026 23268 21420
rect 23212 20974 23214 21026
rect 23266 20974 23268 21026
rect 22428 20804 22484 20814
rect 22428 20690 22484 20748
rect 23212 20804 23268 20974
rect 23212 20738 23268 20748
rect 23436 21028 23492 21756
rect 23548 21746 23604 21756
rect 24556 21810 24612 23100
rect 25340 23156 25396 23166
rect 25340 23062 25396 23100
rect 24668 23044 24724 23054
rect 24668 23042 24836 23044
rect 24668 22990 24670 23042
rect 24722 22990 24836 23042
rect 24668 22988 24836 22990
rect 24668 22978 24724 22988
rect 24556 21758 24558 21810
rect 24610 21758 24612 21810
rect 24556 21746 24612 21758
rect 24668 22484 24724 22494
rect 22428 20638 22430 20690
rect 22482 20638 22484 20690
rect 22428 20626 22484 20638
rect 21196 19954 21252 19964
rect 22540 20578 22596 20590
rect 22540 20526 22542 20578
rect 22594 20526 22596 20578
rect 22540 19572 22596 20526
rect 23436 20188 23492 20972
rect 23212 20132 23492 20188
rect 23548 21588 23604 21598
rect 23212 19906 23268 20132
rect 23212 19854 23214 19906
rect 23266 19854 23268 19906
rect 23212 19842 23268 19854
rect 23548 20018 23604 21532
rect 23772 21586 23828 21598
rect 23772 21534 23774 21586
rect 23826 21534 23828 21586
rect 23660 21474 23716 21486
rect 23660 21422 23662 21474
rect 23714 21422 23716 21474
rect 23660 20916 23716 21422
rect 23772 21476 23828 21534
rect 24108 21588 24164 21598
rect 24108 21494 24164 21532
rect 23772 21410 23828 21420
rect 23660 20860 24388 20916
rect 23548 19966 23550 20018
rect 23602 19966 23604 20018
rect 22540 19506 22596 19516
rect 22988 19236 23044 19246
rect 20748 19058 20804 19068
rect 22540 19124 22596 19134
rect 21756 19012 21812 19022
rect 21868 19012 21924 19022
rect 21756 19010 21868 19012
rect 21756 18958 21758 19010
rect 21810 18958 21868 19010
rect 21756 18956 21868 18958
rect 21756 18946 21812 18956
rect 19180 17666 19236 17678
rect 19180 17614 19182 17666
rect 19234 17614 19236 17666
rect 19180 17556 19236 17614
rect 19180 16772 19236 17500
rect 19740 17556 19796 17566
rect 20076 17556 20132 17566
rect 19740 17554 20132 17556
rect 19740 17502 19742 17554
rect 19794 17502 20078 17554
rect 20130 17502 20132 17554
rect 19740 17500 20132 17502
rect 19740 17490 19796 17500
rect 20076 17490 20132 17500
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19404 16772 19460 16782
rect 19180 16770 19460 16772
rect 19180 16718 19406 16770
rect 19458 16718 19460 16770
rect 19180 16716 19460 16718
rect 19404 16706 19460 16716
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20188 15428 20244 18284
rect 20412 17780 20468 17790
rect 20412 17778 21588 17780
rect 20412 17726 20414 17778
rect 20466 17726 21588 17778
rect 20412 17724 21588 17726
rect 20412 17714 20468 17724
rect 20300 17554 20356 17566
rect 20300 17502 20302 17554
rect 20354 17502 20356 17554
rect 20300 17444 20356 17502
rect 20412 17444 20468 17454
rect 20300 17388 20412 17444
rect 20412 17378 20468 17388
rect 21420 17444 21476 17454
rect 20188 15362 20244 15372
rect 20300 15204 20356 15214
rect 20300 15202 20468 15204
rect 20300 15150 20302 15202
rect 20354 15150 20468 15202
rect 20300 15148 20468 15150
rect 17500 15092 17668 15148
rect 18844 15092 19124 15148
rect 20300 15138 20356 15148
rect 17052 14642 17556 14644
rect 17052 14590 17054 14642
rect 17106 14590 17556 14642
rect 17052 14588 17556 14590
rect 17052 14578 17108 14588
rect 17388 14418 17444 14430
rect 17388 14366 17390 14418
rect 17442 14366 17444 14418
rect 17388 13972 17444 14366
rect 17500 14418 17556 14588
rect 17500 14366 17502 14418
rect 17554 14366 17556 14418
rect 17500 14354 17556 14366
rect 17388 13906 17444 13916
rect 16828 13682 16884 13692
rect 17612 13636 17668 15092
rect 17724 14420 17780 14430
rect 17724 14326 17780 14364
rect 17612 13570 17668 13580
rect 18172 13748 18228 13758
rect 15932 12178 15988 12348
rect 15932 12126 15934 12178
rect 15986 12126 15988 12178
rect 15932 12114 15988 12126
rect 16156 13356 16548 13412
rect 16156 12178 16212 13356
rect 18172 13074 18228 13692
rect 18172 13022 18174 13074
rect 18226 13022 18228 13074
rect 18172 13010 18228 13022
rect 17500 12404 17556 12414
rect 17500 12310 17556 12348
rect 16156 12126 16158 12178
rect 16210 12126 16212 12178
rect 16156 12114 16212 12126
rect 17612 12068 17668 12078
rect 17612 12066 18340 12068
rect 17612 12014 17614 12066
rect 17666 12014 18340 12066
rect 17612 12012 18340 12014
rect 17612 12002 17668 12012
rect 15484 11732 15540 11742
rect 15484 11394 15540 11676
rect 16156 11508 16212 11518
rect 16156 11414 16212 11452
rect 18284 11506 18340 12012
rect 18284 11454 18286 11506
rect 18338 11454 18340 11506
rect 18284 11442 18340 11454
rect 15484 11342 15486 11394
rect 15538 11342 15540 11394
rect 15484 11330 15540 11342
rect 15372 9202 15428 9212
rect 15596 10722 15652 10734
rect 15596 10670 15598 10722
rect 15650 10670 15652 10722
rect 15596 9156 15652 10670
rect 18956 10610 19012 10622
rect 18956 10558 18958 10610
rect 19010 10558 19012 10610
rect 18508 10498 18564 10510
rect 18508 10446 18510 10498
rect 18562 10446 18564 10498
rect 16716 9940 16772 9950
rect 16716 9380 16772 9884
rect 16268 9324 16772 9380
rect 16268 9266 16324 9324
rect 16268 9214 16270 9266
rect 16322 9214 16324 9266
rect 16268 9202 16324 9214
rect 15596 9090 15652 9100
rect 16492 9154 16548 9166
rect 16492 9102 16494 9154
rect 16546 9102 16548 9154
rect 15148 9044 15204 9054
rect 15148 8950 15204 8988
rect 15708 9044 15764 9054
rect 15596 8932 15652 8942
rect 15708 8932 15764 8988
rect 15596 8930 15764 8932
rect 15596 8878 15598 8930
rect 15650 8878 15764 8930
rect 15596 8876 15764 8878
rect 15596 8866 15652 8876
rect 16492 7028 16548 9102
rect 16716 9042 16772 9324
rect 16716 8990 16718 9042
rect 16770 8990 16772 9042
rect 16716 8978 16772 8990
rect 17388 9716 17444 9726
rect 17388 9042 17444 9660
rect 18172 9156 18228 9166
rect 18172 9062 18228 9100
rect 17388 8990 17390 9042
rect 17442 8990 17444 9042
rect 17388 8978 17444 8990
rect 16156 6972 16548 7028
rect 17276 8370 17332 8382
rect 17276 8318 17278 8370
rect 17330 8318 17332 8370
rect 14924 5842 14980 5852
rect 15708 5908 15764 5918
rect 15708 5814 15764 5852
rect 16044 5908 16100 5918
rect 16156 5908 16212 6972
rect 16380 6802 16436 6814
rect 16828 6804 16884 6814
rect 16380 6750 16382 6802
rect 16434 6750 16436 6802
rect 16268 6580 16324 6590
rect 16268 6130 16324 6524
rect 16380 6468 16436 6750
rect 16380 6402 16436 6412
rect 16492 6802 16884 6804
rect 16492 6750 16830 6802
rect 16882 6750 16884 6802
rect 16492 6748 16884 6750
rect 16268 6078 16270 6130
rect 16322 6078 16324 6130
rect 16268 6066 16324 6078
rect 16380 6020 16436 6030
rect 16492 6020 16548 6748
rect 16828 6738 16884 6748
rect 17276 6692 17332 8318
rect 18508 7364 18564 10446
rect 18956 8484 19012 10558
rect 19068 9940 19124 15092
rect 20188 14420 20244 14430
rect 20188 14326 20244 14364
rect 19740 14308 19796 14318
rect 19628 14252 19740 14308
rect 19180 13636 19236 13646
rect 19180 12178 19236 13580
rect 19628 12404 19684 14252
rect 19740 14242 19796 14252
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20076 12962 20132 12974
rect 20076 12910 20078 12962
rect 20130 12910 20132 12962
rect 20076 12740 20132 12910
rect 20076 12674 20132 12684
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19628 12348 20020 12404
rect 19964 12290 20020 12348
rect 19964 12238 19966 12290
rect 20018 12238 20020 12290
rect 19964 12226 20020 12238
rect 19180 12126 19182 12178
rect 19234 12126 19236 12178
rect 19180 11844 19236 12126
rect 19180 11778 19236 11788
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19628 10500 19684 10510
rect 19628 10498 20020 10500
rect 19628 10446 19630 10498
rect 19682 10446 20020 10498
rect 19628 10444 20020 10446
rect 19628 10434 19684 10444
rect 19964 10050 20020 10444
rect 19964 9998 19966 10050
rect 20018 9998 20020 10050
rect 19964 9986 20020 9998
rect 20300 10164 20356 10174
rect 20300 10050 20356 10108
rect 20300 9998 20302 10050
rect 20354 9998 20356 10050
rect 20300 9986 20356 9998
rect 19068 9826 19124 9884
rect 19068 9774 19070 9826
rect 19122 9774 19124 9826
rect 19068 9762 19124 9774
rect 19404 9604 19460 9614
rect 19404 9510 19460 9548
rect 20076 9604 20132 9642
rect 20076 9538 20132 9548
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 18956 8418 19012 8428
rect 19404 8932 19460 8942
rect 19404 8370 19460 8876
rect 20300 8930 20356 8942
rect 20300 8878 20302 8930
rect 20354 8878 20356 8930
rect 19404 8318 19406 8370
rect 19458 8318 19460 8370
rect 19404 8306 19460 8318
rect 19628 8820 19684 8830
rect 18508 7298 18564 7308
rect 19068 7364 19124 7374
rect 17388 6692 17444 6702
rect 17276 6636 17388 6692
rect 17388 6598 17444 6636
rect 16828 6466 16884 6478
rect 16828 6414 16830 6466
rect 16882 6414 16884 6466
rect 16828 6356 16884 6414
rect 16828 6290 16884 6300
rect 16940 6468 16996 6478
rect 16380 6018 16548 6020
rect 16380 5966 16382 6018
rect 16434 5966 16548 6018
rect 16380 5964 16548 5966
rect 16828 6132 16884 6142
rect 16380 5954 16436 5964
rect 16044 5906 16212 5908
rect 16044 5854 16046 5906
rect 16098 5854 16212 5906
rect 16044 5852 16212 5854
rect 16828 5908 16884 6076
rect 16940 6020 16996 6412
rect 17164 6466 17220 6478
rect 17164 6414 17166 6466
rect 17218 6414 17220 6466
rect 17164 6244 17220 6414
rect 17948 6356 18004 6366
rect 17164 6188 17556 6244
rect 17388 6020 17444 6030
rect 16940 6018 17444 6020
rect 16940 5966 17390 6018
rect 17442 5966 17444 6018
rect 16940 5964 17444 5966
rect 17388 5954 17444 5964
rect 17500 5908 17556 6188
rect 17948 6130 18004 6300
rect 17948 6078 17950 6130
rect 18002 6078 18004 6130
rect 17948 6066 18004 6078
rect 19068 6132 19124 7308
rect 19628 6802 19684 8764
rect 20076 8484 20132 8494
rect 20132 8428 20244 8484
rect 20076 8418 20132 8428
rect 20188 8258 20244 8428
rect 20188 8206 20190 8258
rect 20242 8206 20244 8258
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 20076 7700 20132 7710
rect 20076 7364 20132 7644
rect 20188 7586 20244 8206
rect 20188 7534 20190 7586
rect 20242 7534 20244 7586
rect 20188 7522 20244 7534
rect 20076 7308 20244 7364
rect 19628 6750 19630 6802
rect 19682 6750 19684 6802
rect 19628 6738 19684 6750
rect 19068 6066 19124 6076
rect 19292 6690 19348 6702
rect 19292 6638 19294 6690
rect 19346 6638 19348 6690
rect 19292 6356 19348 6638
rect 19516 6692 19572 6702
rect 19516 6598 19572 6636
rect 19964 6692 20020 6702
rect 19964 6598 20020 6636
rect 19740 6468 19796 6478
rect 19292 6132 19348 6300
rect 17612 5908 17668 5918
rect 17500 5906 17668 5908
rect 17500 5854 17614 5906
rect 17666 5854 17668 5906
rect 17500 5852 17668 5854
rect 13356 5794 13412 5806
rect 13356 5742 13358 5794
rect 13410 5742 13412 5794
rect 11228 4274 11284 4284
rect 12796 5234 12852 5246
rect 12796 5182 12798 5234
rect 12850 5182 12852 5234
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 12796 3556 12852 5182
rect 13356 4340 13412 5742
rect 16044 5348 16100 5852
rect 16828 5842 16884 5852
rect 14588 5236 14644 5246
rect 14588 4450 14644 5180
rect 15932 5236 15988 5246
rect 15932 5142 15988 5180
rect 16044 5010 16100 5292
rect 16268 5796 16324 5806
rect 16268 5346 16324 5740
rect 16268 5294 16270 5346
rect 16322 5294 16324 5346
rect 16268 5282 16324 5294
rect 17612 5236 17668 5852
rect 17836 5906 17892 5918
rect 17836 5854 17838 5906
rect 17890 5854 17892 5906
rect 17724 5796 17780 5806
rect 17724 5702 17780 5740
rect 17612 5170 17668 5180
rect 16044 4958 16046 5010
rect 16098 4958 16100 5010
rect 16044 4946 16100 4958
rect 16716 5124 16772 5134
rect 14588 4398 14590 4450
rect 14642 4398 14644 4450
rect 14588 4386 14644 4398
rect 13804 4340 13860 4350
rect 13412 4338 13860 4340
rect 13412 4286 13806 4338
rect 13858 4286 13860 4338
rect 13412 4284 13860 4286
rect 13356 4246 13412 4284
rect 13804 4274 13860 4284
rect 13020 4228 13076 4238
rect 13020 4134 13076 4172
rect 16716 4226 16772 5068
rect 17836 5124 17892 5854
rect 18732 5236 18788 5246
rect 19180 5236 19236 5246
rect 18732 5234 19236 5236
rect 18732 5182 18734 5234
rect 18786 5182 19182 5234
rect 19234 5182 19236 5234
rect 18732 5180 19236 5182
rect 18732 5170 18788 5180
rect 19180 5170 19236 5180
rect 17836 5058 17892 5068
rect 18172 5124 18228 5134
rect 18172 5030 18228 5068
rect 18396 5124 18452 5134
rect 18396 5030 18452 5068
rect 18732 5012 18788 5022
rect 19292 5012 19348 6076
rect 19628 6466 19796 6468
rect 19628 6414 19742 6466
rect 19794 6414 19796 6466
rect 19628 6412 19796 6414
rect 19628 6020 19684 6412
rect 19740 6402 19796 6412
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19628 5964 19796 6020
rect 18732 5010 19348 5012
rect 18732 4958 18734 5010
rect 18786 4958 19348 5010
rect 18732 4956 19348 4958
rect 19404 5348 19460 5358
rect 19404 5010 19460 5292
rect 19516 5236 19572 5246
rect 19516 5234 19684 5236
rect 19516 5182 19518 5234
rect 19570 5182 19684 5234
rect 19516 5180 19684 5182
rect 19516 5170 19572 5180
rect 19404 4958 19406 5010
rect 19458 4958 19460 5010
rect 18732 4946 18788 4956
rect 19404 4946 19460 4958
rect 16716 4174 16718 4226
rect 16770 4174 16772 4226
rect 16716 4162 16772 4174
rect 17836 4900 17892 4910
rect 17836 4226 17892 4844
rect 18620 4900 18676 4910
rect 18620 4806 18676 4844
rect 19628 4564 19684 5180
rect 19740 5124 19796 5964
rect 19740 5058 19796 5068
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19628 4508 20020 4564
rect 19964 4450 20020 4508
rect 19964 4398 19966 4450
rect 20018 4398 20020 4450
rect 19964 4386 20020 4398
rect 17836 4174 17838 4226
rect 17890 4174 17892 4226
rect 17836 4162 17892 4174
rect 12796 3490 12852 3500
rect 18844 3666 18900 3678
rect 18844 3614 18846 3666
rect 18898 3614 18900 3666
rect 2940 3332 2996 3342
rect 2716 3330 2996 3332
rect 2716 3278 2942 3330
rect 2994 3278 2996 3330
rect 2716 3276 2996 3278
rect 2716 800 2772 3276
rect 2940 3266 2996 3276
rect 4732 3332 4788 3342
rect 4732 800 4788 3276
rect 5516 3332 5572 3342
rect 6972 3332 7028 3342
rect 5516 3238 5572 3276
rect 6748 3330 7028 3332
rect 6748 3278 6974 3330
rect 7026 3278 7028 3330
rect 6748 3276 7028 3278
rect 6748 800 6804 3276
rect 6972 3266 7028 3276
rect 9324 3330 9380 3342
rect 11004 3332 11060 3342
rect 13132 3332 13188 3342
rect 15036 3332 15092 3342
rect 17052 3332 17108 3342
rect 9324 3278 9326 3330
rect 9378 3278 9380 3330
rect 8764 924 9044 980
rect 8764 800 8820 924
rect 2688 0 2800 800
rect 4704 0 4816 800
rect 6720 0 6832 800
rect 8736 0 8848 800
rect 8988 756 9044 924
rect 9324 756 9380 3278
rect 10780 3330 11060 3332
rect 10780 3278 11006 3330
rect 11058 3278 11060 3330
rect 10780 3276 11060 3278
rect 10780 800 10836 3276
rect 11004 3266 11060 3276
rect 12796 3330 13188 3332
rect 12796 3278 13134 3330
rect 13186 3278 13188 3330
rect 12796 3276 13188 3278
rect 12796 800 12852 3276
rect 13132 3266 13188 3276
rect 14812 3330 15092 3332
rect 14812 3278 15038 3330
rect 15090 3278 15092 3330
rect 14812 3276 15092 3278
rect 14812 800 14868 3276
rect 15036 3266 15092 3276
rect 16828 3330 17108 3332
rect 16828 3278 17054 3330
rect 17106 3278 17108 3330
rect 16828 3276 17108 3278
rect 16828 800 16884 3276
rect 17052 3266 17108 3276
rect 18844 800 18900 3614
rect 20076 3556 20132 3566
rect 20188 3556 20244 7308
rect 20300 4116 20356 8878
rect 20412 7924 20468 15148
rect 21420 15148 21476 17388
rect 21532 16994 21588 17724
rect 21532 16942 21534 16994
rect 21586 16942 21588 16994
rect 21532 16930 21588 16942
rect 21420 15092 21588 15148
rect 20524 14532 20580 14542
rect 20748 14532 20804 14542
rect 20524 14530 20692 14532
rect 20524 14478 20526 14530
rect 20578 14478 20692 14530
rect 20524 14476 20692 14478
rect 20524 14466 20580 14476
rect 20524 14308 20580 14318
rect 20524 14214 20580 14252
rect 20636 13636 20692 14476
rect 20748 14438 20804 14476
rect 20636 13580 21364 13636
rect 21308 13186 21364 13580
rect 21308 13134 21310 13186
rect 21362 13134 21364 13186
rect 21308 13122 21364 13134
rect 21420 13076 21476 13086
rect 21420 12982 21476 13020
rect 21308 11732 21364 11742
rect 21308 11394 21364 11676
rect 21532 11508 21588 15092
rect 21868 13748 21924 18956
rect 22316 18340 22372 18350
rect 22316 18246 22372 18284
rect 22540 17668 22596 19068
rect 22988 18450 23044 19180
rect 22988 18398 22990 18450
rect 23042 18398 23044 18450
rect 22988 18386 23044 18398
rect 23212 18452 23268 18462
rect 23548 18452 23604 19966
rect 23772 20692 23828 20702
rect 23772 20018 23828 20636
rect 23772 19966 23774 20018
rect 23826 19966 23828 20018
rect 23772 19954 23828 19966
rect 23884 20692 23940 20702
rect 24108 20692 24164 20702
rect 23884 20690 24164 20692
rect 23884 20638 23886 20690
rect 23938 20638 24110 20690
rect 24162 20638 24164 20690
rect 23884 20636 24164 20638
rect 23212 18450 23492 18452
rect 23212 18398 23214 18450
rect 23266 18398 23492 18450
rect 23212 18396 23492 18398
rect 23212 18386 23268 18396
rect 22764 18340 22820 18350
rect 22764 18246 22820 18284
rect 22652 18226 22708 18238
rect 22652 18174 22654 18226
rect 22706 18174 22708 18226
rect 22652 17892 22708 18174
rect 23436 18228 23492 18396
rect 23548 18386 23604 18396
rect 23884 18450 23940 20636
rect 24108 20626 24164 20636
rect 24220 20188 24276 20860
rect 24332 20802 24388 20860
rect 24332 20750 24334 20802
rect 24386 20750 24388 20802
rect 24332 20738 24388 20750
rect 24108 20132 24276 20188
rect 24444 20578 24500 20590
rect 24444 20526 24446 20578
rect 24498 20526 24500 20578
rect 23884 18398 23886 18450
rect 23938 18398 23940 18450
rect 23884 18386 23940 18398
rect 23996 19794 24052 19806
rect 23996 19742 23998 19794
rect 24050 19742 24052 19794
rect 23436 18226 23604 18228
rect 23436 18174 23438 18226
rect 23490 18174 23604 18226
rect 23436 18172 23604 18174
rect 23436 18162 23492 18172
rect 22652 17836 23492 17892
rect 23436 17778 23492 17836
rect 23436 17726 23438 17778
rect 23490 17726 23492 17778
rect 23436 17714 23492 17726
rect 22652 17668 22708 17678
rect 22316 17666 22708 17668
rect 22316 17614 22654 17666
rect 22706 17614 22708 17666
rect 22316 17612 22708 17614
rect 22316 16882 22372 17612
rect 22652 17602 22708 17612
rect 23548 17556 23604 18172
rect 23436 17500 23604 17556
rect 23324 17108 23380 17118
rect 22316 16830 22318 16882
rect 22370 16830 22372 16882
rect 22316 16818 22372 16830
rect 22988 16994 23044 17006
rect 22988 16942 22990 16994
rect 23042 16942 23044 16994
rect 22988 16660 23044 16942
rect 23324 16994 23380 17052
rect 23324 16942 23326 16994
rect 23378 16942 23380 16994
rect 23324 16930 23380 16942
rect 22988 16594 23044 16604
rect 23436 15876 23492 17500
rect 23884 17108 23940 17118
rect 23884 17014 23940 17052
rect 23436 15810 23492 15820
rect 23884 16098 23940 16110
rect 23884 16046 23886 16098
rect 23938 16046 23940 16098
rect 23660 15428 23716 15438
rect 23548 15426 23716 15428
rect 23548 15374 23662 15426
rect 23714 15374 23716 15426
rect 23548 15372 23716 15374
rect 22764 15092 22820 15102
rect 22764 14532 22820 15036
rect 22988 14644 23044 14682
rect 22988 14578 23044 14588
rect 21868 13682 21924 13692
rect 22540 13860 22596 13870
rect 22092 13076 22148 13086
rect 21980 12740 22036 12750
rect 21980 12646 22036 12684
rect 22092 12066 22148 13020
rect 22540 12740 22596 13804
rect 22652 12964 22708 12974
rect 22764 12964 22820 14476
rect 22876 14530 22932 14542
rect 22876 14478 22878 14530
rect 22930 14478 22932 14530
rect 22876 13076 22932 14478
rect 22876 13010 22932 13020
rect 22988 14420 23044 14430
rect 22652 12962 22820 12964
rect 22652 12910 22654 12962
rect 22706 12910 22820 12962
rect 22652 12908 22820 12910
rect 22988 12962 23044 14364
rect 23324 14418 23380 14430
rect 23324 14366 23326 14418
rect 23378 14366 23380 14418
rect 23324 14196 23380 14366
rect 23548 14196 23604 15372
rect 23660 15362 23716 15372
rect 23772 15314 23828 15326
rect 23772 15262 23774 15314
rect 23826 15262 23828 15314
rect 23660 15092 23716 15102
rect 23660 14998 23716 15036
rect 23324 14140 23604 14196
rect 23548 13860 23604 14140
rect 23772 13972 23828 15262
rect 23884 15204 23940 16046
rect 23884 15138 23940 15148
rect 23996 15148 24052 19742
rect 24108 18450 24164 20132
rect 24444 19236 24500 20526
rect 24444 19170 24500 19180
rect 24556 20580 24612 20590
rect 24668 20580 24724 22428
rect 24556 20578 24724 20580
rect 24556 20526 24558 20578
rect 24610 20526 24724 20578
rect 24556 20524 24724 20526
rect 24780 22370 24836 22988
rect 25676 22484 25732 22494
rect 25676 22390 25732 22428
rect 24780 22318 24782 22370
rect 24834 22318 24836 22370
rect 24780 20802 24836 22318
rect 25340 22258 25396 22270
rect 25340 22206 25342 22258
rect 25394 22206 25396 22258
rect 25340 21476 25396 22206
rect 25340 21410 25396 21420
rect 24780 20750 24782 20802
rect 24834 20750 24836 20802
rect 24108 18398 24110 18450
rect 24162 18398 24164 18450
rect 24108 18386 24164 18398
rect 24220 18450 24276 18462
rect 24220 18398 24222 18450
rect 24274 18398 24276 18450
rect 24108 18228 24164 18238
rect 24220 18228 24276 18398
rect 24444 18452 24500 18462
rect 24556 18452 24612 20524
rect 24780 20188 24836 20750
rect 25900 20188 25956 25788
rect 27356 25618 27412 26124
rect 27356 25566 27358 25618
rect 27410 25566 27412 25618
rect 27356 25554 27412 25566
rect 26572 23154 26628 23166
rect 26572 23102 26574 23154
rect 26626 23102 26628 23154
rect 26348 23044 26404 23054
rect 26572 23044 26628 23102
rect 27020 23154 27076 23166
rect 27020 23102 27022 23154
rect 27074 23102 27076 23154
rect 26348 23042 26628 23044
rect 26348 22990 26350 23042
rect 26402 22990 26628 23042
rect 26348 22988 26628 22990
rect 26796 23044 26852 23054
rect 24444 18450 24612 18452
rect 24444 18398 24446 18450
rect 24498 18398 24612 18450
rect 24444 18396 24612 18398
rect 24668 20132 24836 20188
rect 25676 20132 25956 20188
rect 26012 21476 26068 21486
rect 24444 18386 24500 18396
rect 24668 18228 24724 20132
rect 25228 18452 25284 18462
rect 25228 18358 25284 18396
rect 25340 18340 25396 18350
rect 25340 18338 25620 18340
rect 25340 18286 25342 18338
rect 25394 18286 25620 18338
rect 25340 18284 25620 18286
rect 25340 18274 25396 18284
rect 24220 18172 24724 18228
rect 24108 16882 24164 18172
rect 25340 18116 25396 18126
rect 25340 17106 25396 18060
rect 25564 17778 25620 18284
rect 25564 17726 25566 17778
rect 25618 17726 25620 17778
rect 25564 17714 25620 17726
rect 25340 17054 25342 17106
rect 25394 17054 25396 17106
rect 24668 16996 24724 17006
rect 24668 16902 24724 16940
rect 25340 16996 25396 17054
rect 25340 16930 25396 16940
rect 24108 16830 24110 16882
rect 24162 16830 24164 16882
rect 24108 16818 24164 16830
rect 24332 16660 24388 16670
rect 24332 16100 24388 16604
rect 25564 16212 25620 16222
rect 25676 16212 25732 20132
rect 25900 20020 25956 20030
rect 25900 19926 25956 19964
rect 25788 16770 25844 16782
rect 25788 16718 25790 16770
rect 25842 16718 25844 16770
rect 25788 16548 25844 16718
rect 25788 16482 25844 16492
rect 25564 16210 25732 16212
rect 25564 16158 25566 16210
rect 25618 16158 25732 16210
rect 25564 16156 25732 16158
rect 25564 16146 25620 16156
rect 24332 16006 24388 16044
rect 25004 16100 25060 16110
rect 25004 16006 25060 16044
rect 24332 15876 24388 15886
rect 23996 15092 24164 15148
rect 23772 13906 23828 13916
rect 24108 14530 24164 15092
rect 24108 14478 24110 14530
rect 24162 14478 24164 14530
rect 23660 13860 23716 13870
rect 23548 13804 23660 13860
rect 23436 13748 23492 13758
rect 23436 13654 23492 13692
rect 23660 13074 23716 13804
rect 24108 13858 24164 14478
rect 24108 13806 24110 13858
rect 24162 13806 24164 13858
rect 24108 13794 24164 13806
rect 24332 14418 24388 15820
rect 25676 15316 25732 16156
rect 25676 15250 25732 15260
rect 26012 15148 26068 21420
rect 26348 21476 26404 22988
rect 26796 22950 26852 22988
rect 27020 22484 27076 23102
rect 27020 22418 27076 22428
rect 27244 23154 27300 23166
rect 27244 23102 27246 23154
rect 27298 23102 27300 23154
rect 27244 21810 27300 23102
rect 27244 21758 27246 21810
rect 27298 21758 27300 21810
rect 27244 21746 27300 21758
rect 27356 22484 27412 22494
rect 27356 21810 27412 22428
rect 27356 21758 27358 21810
rect 27410 21758 27412 21810
rect 27356 21746 27412 21758
rect 27132 21588 27188 21598
rect 26908 21586 27188 21588
rect 26908 21534 27134 21586
rect 27186 21534 27188 21586
rect 26908 21532 27188 21534
rect 26348 21410 26404 21420
rect 26796 21476 26852 21486
rect 26908 21476 26964 21532
rect 27132 21522 27188 21532
rect 26852 21420 26964 21476
rect 26796 21382 26852 21420
rect 26796 20916 26852 20926
rect 27244 20916 27300 20926
rect 27468 20916 27524 28364
rect 27804 28196 27860 28366
rect 27804 28130 27860 28140
rect 27580 26964 27636 27002
rect 27916 26908 27972 30268
rect 27580 26898 27636 26908
rect 26124 20914 27524 20916
rect 26124 20862 26798 20914
rect 26850 20862 27246 20914
rect 27298 20862 27524 20914
rect 26124 20860 27524 20862
rect 27692 26852 27972 26908
rect 28028 30772 28084 30782
rect 26124 20188 26180 20860
rect 26796 20850 26852 20860
rect 27244 20850 27300 20860
rect 27692 20804 27748 26852
rect 27916 26178 27972 26190
rect 27916 26126 27918 26178
rect 27970 26126 27972 26178
rect 27916 25396 27972 26126
rect 27916 25330 27972 25340
rect 27804 23044 27860 23054
rect 27804 22482 27860 22988
rect 27804 22430 27806 22482
rect 27858 22430 27860 22482
rect 27804 22418 27860 22430
rect 27916 23044 27972 23054
rect 28028 23044 28084 30716
rect 28140 29314 28196 29326
rect 28140 29262 28142 29314
rect 28194 29262 28196 29314
rect 28140 29204 28196 29262
rect 28140 27748 28196 29148
rect 28140 27682 28196 27692
rect 28252 26404 28308 31836
rect 28476 31556 28532 31566
rect 28364 27860 28420 27870
rect 28364 27766 28420 27804
rect 28476 26908 28532 31500
rect 28588 27970 28644 34862
rect 28700 30884 28756 30894
rect 28700 30790 28756 30828
rect 28588 27918 28590 27970
rect 28642 27918 28644 27970
rect 28588 27524 28644 27918
rect 28700 28420 28756 28430
rect 28700 27970 28756 28364
rect 28700 27918 28702 27970
rect 28754 27918 28756 27970
rect 28700 27906 28756 27918
rect 28700 27524 28756 27534
rect 28588 27468 28700 27524
rect 28700 27458 28756 27468
rect 28140 26292 28196 26302
rect 28140 25506 28196 26236
rect 28140 25454 28142 25506
rect 28194 25454 28196 25506
rect 28140 25284 28196 25454
rect 28140 25218 28196 25228
rect 28252 23380 28308 26348
rect 28364 26852 28532 26908
rect 28364 26068 28420 26852
rect 28364 26002 28420 26012
rect 28812 25732 28868 38612
rect 30044 38610 30100 38622
rect 30044 38558 30046 38610
rect 30098 38558 30100 38610
rect 30044 38050 30100 38558
rect 30156 38164 30212 38892
rect 30268 38882 30324 38892
rect 30604 39396 30660 39406
rect 30604 38834 30660 39340
rect 30604 38782 30606 38834
rect 30658 38782 30660 38834
rect 30604 38770 30660 38782
rect 30380 38724 30436 38762
rect 30380 38658 30436 38668
rect 31612 38724 31668 38734
rect 31724 38724 31780 42364
rect 32060 42194 32116 43260
rect 32284 43538 32340 43550
rect 32284 43486 32286 43538
rect 32338 43486 32340 43538
rect 32284 43316 32340 43486
rect 32284 43250 32340 43260
rect 32396 43538 32452 43550
rect 32396 43486 32398 43538
rect 32450 43486 32452 43538
rect 32060 42142 32062 42194
rect 32114 42142 32116 42194
rect 32060 42130 32116 42142
rect 32284 42084 32340 42094
rect 32284 41990 32340 42028
rect 31836 41970 31892 41982
rect 31836 41918 31838 41970
rect 31890 41918 31892 41970
rect 31836 41860 31892 41918
rect 32396 41972 32452 43486
rect 32396 41878 32452 41916
rect 31836 41794 31892 41804
rect 32284 41860 32340 41870
rect 32284 41766 32340 41804
rect 32508 38948 32564 38958
rect 32508 38854 32564 38892
rect 31668 38668 31780 38724
rect 30156 38098 30212 38108
rect 30828 38610 30884 38622
rect 31612 38612 31780 38668
rect 32508 38612 32564 38622
rect 30828 38558 30830 38610
rect 30882 38558 30884 38610
rect 30604 38052 30660 38062
rect 30044 37998 30046 38050
rect 30098 37998 30100 38050
rect 30044 37986 30100 37998
rect 30380 38050 30660 38052
rect 30380 37998 30606 38050
rect 30658 37998 30660 38050
rect 30380 37996 30660 37998
rect 29260 37940 29316 37950
rect 29036 37828 29092 37838
rect 29036 37734 29092 37772
rect 29260 37604 29316 37884
rect 29260 37538 29316 37548
rect 29372 37940 29428 37950
rect 29708 37940 29764 37950
rect 29372 37938 29764 37940
rect 29372 37886 29374 37938
rect 29426 37886 29710 37938
rect 29762 37886 29764 37938
rect 29372 37884 29764 37886
rect 29148 37492 29204 37502
rect 29036 37434 29092 37446
rect 28924 37378 28980 37390
rect 28924 37326 28926 37378
rect 28978 37326 28980 37378
rect 28924 37268 28980 37326
rect 29036 37382 29038 37434
rect 29090 37382 29092 37434
rect 29036 37380 29092 37382
rect 29148 37380 29204 37436
rect 29372 37380 29428 37884
rect 29708 37874 29764 37884
rect 29036 37324 29428 37380
rect 29820 37826 29876 37838
rect 29820 37774 29822 37826
rect 29874 37774 29876 37826
rect 29484 37268 29540 37278
rect 28924 37212 29484 37268
rect 29484 37174 29540 37212
rect 29820 37156 29876 37774
rect 30156 37156 30212 37166
rect 29820 37100 30156 37156
rect 30156 37062 30212 37100
rect 29036 35924 29092 35934
rect 29036 35830 29092 35868
rect 30044 35812 30100 35822
rect 29484 35810 30100 35812
rect 29484 35758 30046 35810
rect 30098 35758 30100 35810
rect 29484 35756 30100 35758
rect 29372 35476 29428 35486
rect 29484 35476 29540 35756
rect 30044 35746 30100 35756
rect 29372 35474 29540 35476
rect 29372 35422 29374 35474
rect 29426 35422 29540 35474
rect 29372 35420 29540 35422
rect 29596 35586 29652 35598
rect 29596 35534 29598 35586
rect 29650 35534 29652 35586
rect 29372 32788 29428 35420
rect 29596 35140 29652 35534
rect 29596 35074 29652 35084
rect 29708 34916 29764 34926
rect 30380 34916 30436 37996
rect 30604 37986 30660 37996
rect 30828 35812 30884 38558
rect 31388 37938 31444 37950
rect 31388 37886 31390 37938
rect 31442 37886 31444 37938
rect 31388 37492 31444 37886
rect 31388 37426 31444 37436
rect 31612 37266 31668 37278
rect 31612 37214 31614 37266
rect 31666 37214 31668 37266
rect 31276 37156 31332 37166
rect 31612 37156 31668 37214
rect 31276 37154 31668 37156
rect 31276 37102 31278 37154
rect 31330 37102 31668 37154
rect 31276 37100 31668 37102
rect 31276 37044 31332 37100
rect 31276 36978 31332 36988
rect 30828 35746 30884 35756
rect 30492 35588 30548 35598
rect 30492 35026 30548 35532
rect 30492 34974 30494 35026
rect 30546 34974 30548 35026
rect 30492 34962 30548 34974
rect 29372 32722 29428 32732
rect 29596 34914 30436 34916
rect 29596 34862 29710 34914
rect 29762 34862 30436 34914
rect 29596 34860 30436 34862
rect 29596 32564 29652 34860
rect 29708 34850 29764 34860
rect 31164 33572 31220 33582
rect 29708 33348 29764 33358
rect 29932 33348 29988 33358
rect 29764 33346 29988 33348
rect 29764 33294 29934 33346
rect 29986 33294 29988 33346
rect 29764 33292 29988 33294
rect 29708 33254 29764 33292
rect 29932 33282 29988 33292
rect 31164 32900 31220 33516
rect 31612 33236 31668 33246
rect 29260 32452 29316 32462
rect 29148 31892 29204 31902
rect 29148 31798 29204 31836
rect 29260 31890 29316 32396
rect 29260 31838 29262 31890
rect 29314 31838 29316 31890
rect 29260 31826 29316 31838
rect 29484 31780 29540 31790
rect 29596 31780 29652 32508
rect 29540 31724 29652 31780
rect 29820 32788 29876 32798
rect 29484 30994 29540 31724
rect 29484 30942 29486 30994
rect 29538 30942 29540 30994
rect 29484 30930 29540 30942
rect 29820 29652 29876 32732
rect 31164 32786 31220 32844
rect 31164 32734 31166 32786
rect 31218 32734 31220 32786
rect 31164 32722 31220 32734
rect 31500 33180 31612 33236
rect 30940 32676 30996 32686
rect 30716 32562 30772 32574
rect 30716 32510 30718 32562
rect 30770 32510 30772 32562
rect 30380 32452 30436 32462
rect 30716 32452 30772 32510
rect 30380 32450 30772 32452
rect 30380 32398 30382 32450
rect 30434 32398 30772 32450
rect 30380 32396 30772 32398
rect 30380 32386 30436 32396
rect 30156 30884 30212 30894
rect 29932 30212 29988 30222
rect 29932 29988 29988 30156
rect 30156 30210 30212 30828
rect 30156 30158 30158 30210
rect 30210 30158 30212 30210
rect 30156 30146 30212 30158
rect 29932 29922 29988 29932
rect 30268 29986 30324 29998
rect 30268 29934 30270 29986
rect 30322 29934 30324 29986
rect 29260 29596 29876 29652
rect 29036 28644 29092 28654
rect 29036 28550 29092 28588
rect 29260 28530 29316 29596
rect 29596 29426 29652 29438
rect 29596 29374 29598 29426
rect 29650 29374 29652 29426
rect 29260 28478 29262 28530
rect 29314 28478 29316 28530
rect 29260 28466 29316 28478
rect 29372 28530 29428 28542
rect 29372 28478 29374 28530
rect 29426 28478 29428 28530
rect 29372 28420 29428 28478
rect 29372 28354 29428 28364
rect 29596 26292 29652 29374
rect 29820 28754 29876 29596
rect 30268 29540 30324 29934
rect 30380 29540 30436 29550
rect 30268 29538 30436 29540
rect 30268 29486 30382 29538
rect 30434 29486 30436 29538
rect 30268 29484 30436 29486
rect 30380 29474 30436 29484
rect 29820 28702 29822 28754
rect 29874 28702 29876 28754
rect 29820 28690 29876 28702
rect 30492 28532 30548 32396
rect 30828 32340 30884 32350
rect 30828 31666 30884 32284
rect 30828 31614 30830 31666
rect 30882 31614 30884 31666
rect 30828 31602 30884 31614
rect 30940 31332 30996 32620
rect 31276 32562 31332 32574
rect 31276 32510 31278 32562
rect 31330 32510 31332 32562
rect 31052 32452 31108 32462
rect 31052 32358 31108 32396
rect 31276 32340 31332 32510
rect 31276 32274 31332 32284
rect 31500 31780 31556 33180
rect 31612 33170 31668 33180
rect 31500 31686 31556 31724
rect 31164 31556 31220 31566
rect 31164 31554 31556 31556
rect 31164 31502 31166 31554
rect 31218 31502 31556 31554
rect 31164 31500 31556 31502
rect 31164 31490 31220 31500
rect 30716 31276 30996 31332
rect 30716 31218 30772 31276
rect 30716 31166 30718 31218
rect 30770 31166 30772 31218
rect 30716 31154 30772 31166
rect 31500 31108 31556 31500
rect 31724 31220 31780 38612
rect 32284 38556 32508 38612
rect 32060 37492 32116 37502
rect 32060 37398 32116 37436
rect 31948 37266 32004 37278
rect 31948 37214 31950 37266
rect 32002 37214 32004 37266
rect 31948 37044 32004 37214
rect 32284 37266 32340 38556
rect 32508 38546 32564 38556
rect 32284 37214 32286 37266
rect 32338 37214 32340 37266
rect 32284 37202 32340 37214
rect 31948 36978 32004 36988
rect 32396 37156 32452 37166
rect 32396 36708 32452 37100
rect 31948 36484 32004 36494
rect 31836 36482 32004 36484
rect 31836 36430 31950 36482
rect 32002 36430 32004 36482
rect 31836 36428 32004 36430
rect 31836 36258 31892 36428
rect 31948 36418 32004 36428
rect 32396 36482 32452 36652
rect 32396 36430 32398 36482
rect 32450 36430 32452 36482
rect 32396 36418 32452 36430
rect 32620 37044 32676 37054
rect 32620 36482 32676 36988
rect 32620 36430 32622 36482
rect 32674 36430 32676 36482
rect 32620 36418 32676 36430
rect 31836 36206 31838 36258
rect 31890 36206 31892 36258
rect 31836 36148 31892 36206
rect 31836 36082 31892 36092
rect 32508 36258 32564 36270
rect 32508 36206 32510 36258
rect 32562 36206 32564 36258
rect 32508 35810 32564 36206
rect 32508 35758 32510 35810
rect 32562 35758 32564 35810
rect 32508 35746 32564 35758
rect 31948 35700 32004 35710
rect 31948 35606 32004 35644
rect 32172 35698 32228 35710
rect 32172 35646 32174 35698
rect 32226 35646 32228 35698
rect 32060 35588 32116 35598
rect 32060 35494 32116 35532
rect 32172 33572 32228 35646
rect 32620 34692 32676 34702
rect 32172 33506 32228 33516
rect 32284 34636 32620 34692
rect 31948 33236 32004 33246
rect 31948 33142 32004 33180
rect 31836 32900 31892 32910
rect 31836 32786 31892 32844
rect 31836 32734 31838 32786
rect 31890 32734 31892 32786
rect 31836 31668 31892 32734
rect 32284 31890 32340 34636
rect 32620 34626 32676 34636
rect 32732 34690 32788 34702
rect 32732 34638 32734 34690
rect 32786 34638 32788 34690
rect 32732 34356 32788 34638
rect 32732 34290 32788 34300
rect 32284 31838 32286 31890
rect 32338 31838 32340 31890
rect 32284 31826 32340 31838
rect 31836 31602 31892 31612
rect 31724 31126 31780 31164
rect 31052 30996 31108 31006
rect 31052 30902 31108 30940
rect 31500 30994 31556 31052
rect 31500 30942 31502 30994
rect 31554 30942 31556 30994
rect 31500 30930 31556 30942
rect 31948 30996 32004 31006
rect 31948 30902 32004 30940
rect 32172 30994 32228 31006
rect 32172 30942 32174 30994
rect 32226 30942 32228 30994
rect 31836 30884 31892 30894
rect 31836 30790 31892 30828
rect 30604 30212 30660 30222
rect 30604 30118 30660 30156
rect 32172 29316 32228 30942
rect 32508 29316 32564 29326
rect 32172 29314 32564 29316
rect 32172 29262 32510 29314
rect 32562 29262 32564 29314
rect 32172 29260 32564 29262
rect 31052 28756 31108 28766
rect 31052 28662 31108 28700
rect 32508 28756 32564 29260
rect 32508 28690 32564 28700
rect 29932 28476 30548 28532
rect 29932 27298 29988 28476
rect 30940 28418 30996 28430
rect 30940 28366 30942 28418
rect 30994 28366 30996 28418
rect 30268 28084 30324 28094
rect 29932 27246 29934 27298
rect 29986 27246 29988 27298
rect 29932 27234 29988 27246
rect 30044 27748 30100 27758
rect 29820 27076 29876 27086
rect 29820 26982 29876 27020
rect 29596 26226 29652 26236
rect 29708 26850 29764 26862
rect 29708 26798 29710 26850
rect 29762 26798 29764 26850
rect 28812 25666 28868 25676
rect 28588 25508 28644 25518
rect 29372 25508 29428 25518
rect 28588 25506 29428 25508
rect 28588 25454 28590 25506
rect 28642 25454 29374 25506
rect 29426 25454 29428 25506
rect 28588 25452 29428 25454
rect 28588 25442 28644 25452
rect 28588 25284 28644 25294
rect 28252 23324 28420 23380
rect 28252 23154 28308 23166
rect 28252 23102 28254 23154
rect 28306 23102 28308 23154
rect 28252 23044 28308 23102
rect 27916 23042 28308 23044
rect 27916 22990 27918 23042
rect 27970 22990 28308 23042
rect 27916 22988 28308 22990
rect 27804 21586 27860 21598
rect 27804 21534 27806 21586
rect 27858 21534 27860 21586
rect 27804 21474 27860 21534
rect 27804 21422 27806 21474
rect 27858 21422 27860 21474
rect 27804 21410 27860 21422
rect 27356 20748 27748 20804
rect 27132 20578 27188 20590
rect 27132 20526 27134 20578
rect 27186 20526 27188 20578
rect 26124 20132 26292 20188
rect 26236 17108 26292 20132
rect 26460 20020 26516 20030
rect 26460 19926 26516 19964
rect 26908 20020 26964 20030
rect 27132 20020 27188 20526
rect 26964 19964 27188 20020
rect 27356 20018 27412 20748
rect 27916 20132 27972 22988
rect 28252 21812 28308 21822
rect 28364 21812 28420 23324
rect 28588 22372 28644 25228
rect 28812 23156 28868 23166
rect 28812 23062 28868 23100
rect 29148 23044 29204 23054
rect 29148 22950 29204 22988
rect 28588 22370 29204 22372
rect 28588 22318 28590 22370
rect 28642 22318 29204 22370
rect 28588 22316 29204 22318
rect 28588 22306 28644 22316
rect 28252 21810 28420 21812
rect 28252 21758 28254 21810
rect 28306 21758 28420 21810
rect 28252 21756 28420 21758
rect 28252 21362 28308 21756
rect 28252 21310 28254 21362
rect 28306 21310 28308 21362
rect 28252 21298 28308 21310
rect 29148 20802 29204 22316
rect 29148 20750 29150 20802
rect 29202 20750 29204 20802
rect 29148 20738 29204 20750
rect 27916 20066 27972 20076
rect 27356 19966 27358 20018
rect 27410 19966 27412 20018
rect 26908 19926 26964 19964
rect 26348 19908 26404 19918
rect 26348 18676 26404 19852
rect 27356 19460 27412 19966
rect 27692 20020 27748 20030
rect 27692 19926 27748 19964
rect 28252 19908 28308 19918
rect 28252 19814 28308 19852
rect 27356 19394 27412 19404
rect 27692 19572 27748 19582
rect 27356 19236 27412 19246
rect 27356 19142 27412 19180
rect 27692 19234 27748 19516
rect 27692 19182 27694 19234
rect 27746 19182 27748 19234
rect 27692 19170 27748 19182
rect 28252 19234 28308 19246
rect 28252 19182 28254 19234
rect 28306 19182 28308 19234
rect 26572 18676 26628 18686
rect 26348 18674 26628 18676
rect 26348 18622 26350 18674
rect 26402 18622 26574 18674
rect 26626 18622 26628 18674
rect 26348 18620 26628 18622
rect 26348 18610 26404 18620
rect 26572 18610 26628 18620
rect 27020 18338 27076 18350
rect 27020 18286 27022 18338
rect 27074 18286 27076 18338
rect 27020 18228 27076 18286
rect 27020 18162 27076 18172
rect 27580 17556 27636 17566
rect 27804 17556 27860 17566
rect 27580 17462 27636 17500
rect 27692 17554 27860 17556
rect 27692 17502 27806 17554
rect 27858 17502 27860 17554
rect 27692 17500 27860 17502
rect 26236 17042 26292 17052
rect 27692 16772 27748 17500
rect 27804 17490 27860 17500
rect 27916 17556 27972 17566
rect 27916 17462 27972 17500
rect 28140 17444 28196 17454
rect 28028 17442 28196 17444
rect 28028 17390 28142 17442
rect 28194 17390 28196 17442
rect 28028 17388 28196 17390
rect 27916 16996 27972 17006
rect 28028 16996 28084 17388
rect 28140 17378 28196 17388
rect 27916 16994 28084 16996
rect 27916 16942 27918 16994
rect 27970 16942 28084 16994
rect 27916 16940 28084 16942
rect 27916 16930 27972 16940
rect 27356 16716 27748 16772
rect 27020 16548 27076 16558
rect 27020 16210 27076 16492
rect 27020 16158 27022 16210
rect 27074 16158 27076 16210
rect 27020 16146 27076 16158
rect 27356 16210 27412 16716
rect 27356 16158 27358 16210
rect 27410 16158 27412 16210
rect 27356 16146 27412 16158
rect 27804 16548 27860 16558
rect 27804 16098 27860 16492
rect 27804 16046 27806 16098
rect 27858 16046 27860 16098
rect 27804 16034 27860 16046
rect 28140 16210 28196 16222
rect 28140 16158 28142 16210
rect 28194 16158 28196 16210
rect 25564 15092 26068 15148
rect 28140 15428 28196 16158
rect 28140 15092 28196 15372
rect 25004 14532 25060 14542
rect 25004 14530 25396 14532
rect 25004 14478 25006 14530
rect 25058 14478 25396 14530
rect 25004 14476 25396 14478
rect 25004 14466 25060 14476
rect 24332 14366 24334 14418
rect 24386 14366 24388 14418
rect 24332 13746 24388 14366
rect 24668 14420 24724 14430
rect 24668 14326 24724 14364
rect 24780 14306 24836 14318
rect 24780 14254 24782 14306
rect 24834 14254 24836 14306
rect 24668 13972 24724 13982
rect 24668 13878 24724 13916
rect 24332 13694 24334 13746
rect 24386 13694 24388 13746
rect 24332 13682 24388 13694
rect 23660 13022 23662 13074
rect 23714 13022 23716 13074
rect 23660 13010 23716 13022
rect 24780 13076 24836 14254
rect 25228 13972 25284 13982
rect 25228 13858 25284 13916
rect 25340 13970 25396 14476
rect 25340 13918 25342 13970
rect 25394 13918 25396 13970
rect 25340 13906 25396 13918
rect 25228 13806 25230 13858
rect 25282 13806 25284 13858
rect 25228 13794 25284 13806
rect 25452 13860 25508 13870
rect 25452 13766 25508 13804
rect 24780 13010 24836 13020
rect 22988 12910 22990 12962
rect 23042 12910 23044 12962
rect 22652 12898 22708 12908
rect 22988 12898 23044 12910
rect 22876 12852 22932 12862
rect 22764 12796 22876 12852
rect 22764 12740 22820 12796
rect 22876 12786 22932 12796
rect 22540 12738 22820 12740
rect 22540 12686 22766 12738
rect 22818 12686 22820 12738
rect 22540 12684 22820 12686
rect 22764 12674 22820 12684
rect 22092 12014 22094 12066
rect 22146 12014 22148 12066
rect 22092 12002 22148 12014
rect 24220 11508 24276 11518
rect 21532 11442 21588 11452
rect 23660 11506 24276 11508
rect 23660 11454 24222 11506
rect 24274 11454 24276 11506
rect 23660 11452 24276 11454
rect 21308 11342 21310 11394
rect 21362 11342 21364 11394
rect 21308 11330 21364 11342
rect 22092 11282 22148 11294
rect 22092 11230 22094 11282
rect 22146 11230 22148 11282
rect 21756 10498 21812 10510
rect 21756 10446 21758 10498
rect 21810 10446 21812 10498
rect 21756 10388 21812 10446
rect 21756 10322 21812 10332
rect 20748 9940 20804 9950
rect 20748 9846 20804 9884
rect 22092 9938 22148 11230
rect 23660 10836 23716 11452
rect 24220 11442 24276 11452
rect 25116 11508 25172 11518
rect 24780 11394 24836 11406
rect 24780 11342 24782 11394
rect 24834 11342 24836 11394
rect 24780 11172 24836 11342
rect 24780 11106 24836 11116
rect 23100 10834 23716 10836
rect 23100 10782 23662 10834
rect 23714 10782 23716 10834
rect 23100 10780 23716 10782
rect 23100 10722 23156 10780
rect 23660 10770 23716 10780
rect 23100 10670 23102 10722
rect 23154 10670 23156 10722
rect 23100 10658 23156 10670
rect 24108 10724 24164 10734
rect 24108 10630 24164 10668
rect 22540 10610 22596 10622
rect 22540 10558 22542 10610
rect 22594 10558 22596 10610
rect 22204 10500 22260 10510
rect 22204 10050 22260 10444
rect 22204 9998 22206 10050
rect 22258 9998 22260 10050
rect 22204 9986 22260 9998
rect 22540 10052 22596 10558
rect 22540 9986 22596 9996
rect 22652 10610 22708 10622
rect 22652 10558 22654 10610
rect 22706 10558 22708 10610
rect 22652 10388 22708 10558
rect 22876 10612 22932 10622
rect 22876 10518 22932 10556
rect 23436 10610 23492 10622
rect 23436 10558 23438 10610
rect 23490 10558 23492 10610
rect 22092 9886 22094 9938
rect 22146 9886 22148 9938
rect 22092 9874 22148 9886
rect 21868 9826 21924 9838
rect 21868 9774 21870 9826
rect 21922 9774 21924 9826
rect 20972 9604 21028 9614
rect 20972 9042 21028 9548
rect 21868 9604 21924 9774
rect 21868 9538 21924 9548
rect 20972 8990 20974 9042
rect 21026 8990 21028 9042
rect 20748 8932 20804 8942
rect 20748 8838 20804 8876
rect 20636 8820 20692 8830
rect 20636 8726 20692 8764
rect 20412 7858 20468 7868
rect 20636 8484 20692 8494
rect 20412 5124 20468 5134
rect 20412 5010 20468 5068
rect 20412 4958 20414 5010
rect 20466 4958 20468 5010
rect 20412 4946 20468 4958
rect 20636 4340 20692 8428
rect 20972 6692 21028 8990
rect 21308 8484 21364 8494
rect 21308 8258 21364 8428
rect 21308 8206 21310 8258
rect 21362 8206 21364 8258
rect 21308 8194 21364 8206
rect 22092 8148 22148 8158
rect 21868 8146 22148 8148
rect 21868 8094 22094 8146
rect 22146 8094 22148 8146
rect 21868 8092 22148 8094
rect 21868 6802 21924 8092
rect 22092 8082 22148 8092
rect 21868 6750 21870 6802
rect 21922 6750 21924 6802
rect 21868 6738 21924 6750
rect 21980 6804 22036 6814
rect 21980 6710 22036 6748
rect 21644 6692 21700 6702
rect 20972 6690 21700 6692
rect 20972 6638 21646 6690
rect 21698 6638 21700 6690
rect 20972 6636 21700 6638
rect 21644 6626 21700 6636
rect 22540 6580 22596 6590
rect 22652 6580 22708 10332
rect 22764 10498 22820 10510
rect 22764 10446 22766 10498
rect 22818 10446 22820 10498
rect 22764 10164 22820 10446
rect 22764 10098 22820 10108
rect 23436 10052 23492 10558
rect 23884 10612 23940 10622
rect 23772 10500 23828 10510
rect 23772 10406 23828 10444
rect 23212 8036 23268 8046
rect 23436 8036 23492 9996
rect 23268 7980 23492 8036
rect 22876 6804 22932 6814
rect 22876 6710 22932 6748
rect 22988 6692 23044 6702
rect 22988 6598 23044 6636
rect 23212 6690 23268 7980
rect 23212 6638 23214 6690
rect 23266 6638 23268 6690
rect 23212 6626 23268 6638
rect 22540 6578 22708 6580
rect 22540 6526 22542 6578
rect 22594 6526 22708 6578
rect 22540 6524 22708 6526
rect 22764 6580 22820 6590
rect 22540 6514 22596 6524
rect 22764 6486 22820 6524
rect 23548 6580 23604 6590
rect 21756 6468 21812 6478
rect 21308 6132 21364 6142
rect 21308 6038 21364 6076
rect 21644 5908 21700 5918
rect 21756 5908 21812 6412
rect 23548 6130 23604 6524
rect 23884 6580 23940 10556
rect 24220 8372 24276 8382
rect 24108 8370 24276 8372
rect 24108 8318 24222 8370
rect 24274 8318 24276 8370
rect 24108 8316 24276 8318
rect 24108 6692 24164 8316
rect 24220 8306 24276 8316
rect 24780 8258 24836 8270
rect 24780 8206 24782 8258
rect 24834 8206 24836 8258
rect 24556 8036 24612 8046
rect 24556 7942 24612 7980
rect 24668 7474 24724 7486
rect 24668 7422 24670 7474
rect 24722 7422 24724 7474
rect 24668 7364 24724 7422
rect 24668 7298 24724 7308
rect 24780 7476 24836 8206
rect 24108 6626 24164 6636
rect 24220 6690 24276 6702
rect 24220 6638 24222 6690
rect 24274 6638 24276 6690
rect 23884 6514 23940 6524
rect 23548 6078 23550 6130
rect 23602 6078 23604 6130
rect 23548 6066 23604 6078
rect 21644 5906 21812 5908
rect 21644 5854 21646 5906
rect 21698 5854 21812 5906
rect 21644 5852 21812 5854
rect 21644 5842 21700 5852
rect 20748 5124 20804 5134
rect 20748 5030 20804 5068
rect 21644 5124 21700 5134
rect 21756 5124 21812 5852
rect 23772 5906 23828 5918
rect 23772 5854 23774 5906
rect 23826 5854 23828 5906
rect 22764 5348 22820 5358
rect 22428 5124 22484 5134
rect 21756 5068 22036 5124
rect 21644 5030 21700 5068
rect 21420 5010 21476 5022
rect 21420 4958 21422 5010
rect 21474 4958 21476 5010
rect 21420 4900 21476 4958
rect 21980 5010 22036 5068
rect 21980 4958 21982 5010
rect 22034 4958 22036 5010
rect 21980 4946 22036 4958
rect 22092 5122 22484 5124
rect 22092 5070 22430 5122
rect 22482 5070 22484 5122
rect 22092 5068 22484 5070
rect 21420 4834 21476 4844
rect 21756 4898 21812 4910
rect 21756 4846 21758 4898
rect 21810 4846 21812 4898
rect 21756 4676 21812 4846
rect 21868 4900 21924 4910
rect 21868 4806 21924 4844
rect 22092 4676 22148 5068
rect 22428 5058 22484 5068
rect 22764 5122 22820 5292
rect 22764 5070 22766 5122
rect 22818 5070 22820 5122
rect 22764 5058 22820 5070
rect 22876 5236 22932 5246
rect 21756 4620 22148 4676
rect 22540 4898 22596 4910
rect 22540 4846 22542 4898
rect 22594 4846 22596 4898
rect 22540 4564 22596 4846
rect 22092 4508 22596 4564
rect 22092 4450 22148 4508
rect 22092 4398 22094 4450
rect 22146 4398 22148 4450
rect 22092 4386 22148 4398
rect 21308 4340 21364 4350
rect 20636 4338 21364 4340
rect 20636 4286 20638 4338
rect 20690 4286 21310 4338
rect 21362 4286 21364 4338
rect 20636 4284 21364 4286
rect 20636 4274 20692 4284
rect 21308 4274 21364 4284
rect 20300 4050 20356 4060
rect 20076 3554 20244 3556
rect 20076 3502 20078 3554
rect 20130 3502 20244 3554
rect 20076 3500 20244 3502
rect 20860 3668 20916 3678
rect 20076 3490 20132 3500
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20860 800 20916 3612
rect 22092 3668 22148 3678
rect 22092 3574 22148 3612
rect 21084 3556 21140 3566
rect 21084 3462 21140 3500
rect 22876 800 22932 5180
rect 23100 5122 23156 5134
rect 23100 5070 23102 5122
rect 23154 5070 23156 5122
rect 23100 4228 23156 5070
rect 23772 5124 23828 5854
rect 24108 5236 24164 5246
rect 24108 5142 24164 5180
rect 23772 5058 23828 5068
rect 24220 5012 24276 6638
rect 24780 6468 24836 7420
rect 24892 8260 24948 8270
rect 24892 6690 24948 8204
rect 24892 6638 24894 6690
rect 24946 6638 24948 6690
rect 24892 6626 24948 6638
rect 24780 6402 24836 6412
rect 25116 6020 25172 11452
rect 25340 11284 25396 11294
rect 25340 10724 25396 11228
rect 25340 10498 25396 10668
rect 25340 10446 25342 10498
rect 25394 10446 25396 10498
rect 25340 10434 25396 10446
rect 25452 9268 25508 9278
rect 25564 9268 25620 15092
rect 28140 15026 28196 15036
rect 26908 13748 26964 13758
rect 26908 13654 26964 13692
rect 28252 13636 28308 19182
rect 29260 19236 29316 25452
rect 29372 25442 29428 25452
rect 29708 23492 29764 26798
rect 30044 26402 30100 27692
rect 30268 27074 30324 28028
rect 30268 27022 30270 27074
rect 30322 27022 30324 27074
rect 30268 27010 30324 27022
rect 30828 27636 30884 27646
rect 30828 26908 30884 27580
rect 30044 26350 30046 26402
rect 30098 26350 30100 26402
rect 30044 26338 30100 26350
rect 30268 26850 30324 26862
rect 30268 26798 30270 26850
rect 30322 26798 30324 26850
rect 30268 25620 30324 26798
rect 30156 25564 30324 25620
rect 30380 26852 30884 26908
rect 30940 26962 30996 28366
rect 31276 28084 31332 28094
rect 31276 27990 31332 28028
rect 32172 28084 32228 28094
rect 32172 27990 32228 28028
rect 31724 27972 31780 27982
rect 31164 27860 31220 27870
rect 31164 27766 31220 27804
rect 31500 27860 31556 27870
rect 31724 27860 31780 27916
rect 31500 27858 31780 27860
rect 31500 27806 31502 27858
rect 31554 27806 31780 27858
rect 31500 27804 31780 27806
rect 31500 27794 31556 27804
rect 31388 27748 31444 27758
rect 31388 27654 31444 27692
rect 30940 26910 30942 26962
rect 30994 26910 30996 26962
rect 30940 26898 30996 26910
rect 31612 26852 31668 26862
rect 30156 25172 30212 25564
rect 30156 25106 30212 25116
rect 30268 25396 30324 25406
rect 30268 24834 30324 25340
rect 30380 24946 30436 26852
rect 31612 26514 31668 26796
rect 31612 26462 31614 26514
rect 31666 26462 31668 26514
rect 31612 26450 31668 26462
rect 31724 26402 31780 27804
rect 31724 26350 31726 26402
rect 31778 26350 31780 26402
rect 31724 26338 31780 26350
rect 31836 27860 31892 27870
rect 30716 26292 30772 26302
rect 30716 25620 30772 26236
rect 31612 26068 31668 26078
rect 31836 26068 31892 27804
rect 31948 27076 32004 27086
rect 31948 26982 32004 27020
rect 32172 26852 32228 26862
rect 32172 26514 32228 26796
rect 32172 26462 32174 26514
rect 32226 26462 32228 26514
rect 32172 26450 32228 26462
rect 31612 26066 31892 26068
rect 31612 26014 31614 26066
rect 31666 26014 31892 26066
rect 31612 26012 31892 26014
rect 31612 26002 31668 26012
rect 30716 25554 30772 25564
rect 31388 25620 31444 25630
rect 31388 25526 31444 25564
rect 30380 24894 30382 24946
rect 30434 24894 30436 24946
rect 30380 24882 30436 24894
rect 30268 24782 30270 24834
rect 30322 24782 30324 24834
rect 30268 24770 30324 24782
rect 31836 23938 31892 23950
rect 31836 23886 31838 23938
rect 31890 23886 31892 23938
rect 31500 23826 31556 23838
rect 31500 23774 31502 23826
rect 31554 23774 31556 23826
rect 31500 23492 31556 23774
rect 31836 23828 31892 23886
rect 31836 23762 31892 23772
rect 32172 23938 32228 23950
rect 32172 23886 32174 23938
rect 32226 23886 32228 23938
rect 31948 23716 32004 23726
rect 31948 23622 32004 23660
rect 28588 17780 28644 17790
rect 29260 17780 29316 19180
rect 28588 17778 29316 17780
rect 28588 17726 28590 17778
rect 28642 17726 29316 17778
rect 28588 17724 29316 17726
rect 28588 15540 28644 17724
rect 29260 17666 29316 17724
rect 29260 17614 29262 17666
rect 29314 17614 29316 17666
rect 29260 17602 29316 17614
rect 29372 23156 29428 23166
rect 29372 17556 29428 23100
rect 29708 23044 29764 23436
rect 31388 23436 31500 23492
rect 29708 22978 29764 22988
rect 31276 23044 31332 23054
rect 31276 22950 31332 22988
rect 31388 22370 31444 23436
rect 31500 23426 31556 23436
rect 32060 23380 32116 23390
rect 32060 23154 32116 23324
rect 32060 23102 32062 23154
rect 32114 23102 32116 23154
rect 32060 23090 32116 23102
rect 32172 23044 32228 23886
rect 32508 23828 32564 23838
rect 32508 23716 32564 23772
rect 32508 23714 32676 23716
rect 32508 23662 32510 23714
rect 32562 23662 32676 23714
rect 32508 23660 32676 23662
rect 32508 23650 32564 23660
rect 32508 23044 32564 23054
rect 32172 23042 32564 23044
rect 32172 22990 32510 23042
rect 32562 22990 32564 23042
rect 32172 22988 32564 22990
rect 31388 22318 31390 22370
rect 31442 22318 31444 22370
rect 31388 22306 31444 22318
rect 31612 22820 31668 22830
rect 31612 22370 31668 22764
rect 32508 22820 32564 22988
rect 32508 22754 32564 22764
rect 32284 22708 32340 22718
rect 32060 22652 32284 22708
rect 32060 22594 32116 22652
rect 32284 22642 32340 22652
rect 32060 22542 32062 22594
rect 32114 22542 32116 22594
rect 32060 22530 32116 22542
rect 31612 22318 31614 22370
rect 31666 22318 31668 22370
rect 31612 22306 31668 22318
rect 31500 22260 31556 22270
rect 31500 22166 31556 22204
rect 32508 22260 32564 22270
rect 32508 21474 32564 22204
rect 32508 21422 32510 21474
rect 32562 21422 32564 21474
rect 32060 20916 32116 20926
rect 31948 20914 32116 20916
rect 31948 20862 32062 20914
rect 32114 20862 32116 20914
rect 31948 20860 32116 20862
rect 29932 20692 29988 20702
rect 29932 20690 30212 20692
rect 29932 20638 29934 20690
rect 29986 20638 30212 20690
rect 29932 20636 30212 20638
rect 29932 20626 29988 20636
rect 30156 20132 30212 20636
rect 30492 20132 30548 20142
rect 30156 20130 30548 20132
rect 30156 20078 30494 20130
rect 30546 20078 30548 20130
rect 30156 20076 30548 20078
rect 30492 20066 30548 20076
rect 29820 20020 29876 20030
rect 29820 19926 29876 19964
rect 30828 20018 30884 20030
rect 30828 19966 30830 20018
rect 30882 19966 30884 20018
rect 29372 17490 29428 17500
rect 29596 19906 29652 19918
rect 29596 19854 29598 19906
rect 29650 19854 29652 19906
rect 28476 15484 28644 15540
rect 28700 16882 28756 16894
rect 28700 16830 28702 16882
rect 28754 16830 28756 16882
rect 27916 13580 28308 13636
rect 28364 14868 28420 14878
rect 26572 13412 26628 13422
rect 25788 13076 25844 13086
rect 25788 12982 25844 13020
rect 26572 12964 26628 13356
rect 27132 12964 27188 12974
rect 27580 12964 27636 12974
rect 26572 12962 26852 12964
rect 26572 12910 26574 12962
rect 26626 12910 26852 12962
rect 26572 12908 26852 12910
rect 26572 12898 26628 12908
rect 26796 12178 26852 12908
rect 27132 12962 27636 12964
rect 27132 12910 27134 12962
rect 27186 12910 27582 12962
rect 27634 12910 27636 12962
rect 27132 12908 27636 12910
rect 27132 12898 27188 12908
rect 27580 12898 27636 12908
rect 27356 12740 27412 12750
rect 27356 12738 27636 12740
rect 27356 12686 27358 12738
rect 27410 12686 27636 12738
rect 27356 12684 27636 12686
rect 27356 12674 27412 12684
rect 27580 12290 27636 12684
rect 27580 12238 27582 12290
rect 27634 12238 27636 12290
rect 27580 12226 27636 12238
rect 26796 12126 26798 12178
rect 26850 12126 26852 12178
rect 26796 12114 26852 12126
rect 26460 11284 26516 11294
rect 26460 11190 26516 11228
rect 25676 11172 25732 11182
rect 25676 11078 25732 11116
rect 26572 11170 26628 11182
rect 26572 11118 26574 11170
rect 26626 11118 26628 11170
rect 26236 10052 26292 10062
rect 26236 9826 26292 9996
rect 26236 9774 26238 9826
rect 26290 9774 26292 9826
rect 26236 9762 26292 9774
rect 26572 9826 26628 11118
rect 26572 9774 26574 9826
rect 26626 9774 26628 9826
rect 26572 9762 26628 9774
rect 26684 10500 26740 10510
rect 26684 9602 26740 10444
rect 27468 10500 27524 10510
rect 27468 10406 27524 10444
rect 26796 10052 26852 10062
rect 26796 9958 26852 9996
rect 27804 10052 27860 10062
rect 27804 9958 27860 9996
rect 27020 9828 27076 9838
rect 27020 9826 27188 9828
rect 27020 9774 27022 9826
rect 27074 9774 27188 9826
rect 27020 9772 27188 9774
rect 27020 9762 27076 9772
rect 26684 9550 26686 9602
rect 26738 9550 26740 9602
rect 26684 9538 26740 9550
rect 25452 9266 25732 9268
rect 25452 9214 25454 9266
rect 25506 9214 25732 9266
rect 25452 9212 25732 9214
rect 25452 9202 25508 9212
rect 25564 8258 25620 8270
rect 25564 8206 25566 8258
rect 25618 8206 25620 8258
rect 25564 8148 25620 8206
rect 25452 8092 25564 8148
rect 25452 7698 25508 8092
rect 25564 8082 25620 8092
rect 25452 7646 25454 7698
rect 25506 7646 25508 7698
rect 25452 7634 25508 7646
rect 25676 7924 25732 9212
rect 26460 8372 26516 8382
rect 26348 8316 26460 8372
rect 25788 8260 25844 8270
rect 25788 8166 25844 8204
rect 25900 8148 25956 8158
rect 25900 8146 26180 8148
rect 25900 8094 25902 8146
rect 25954 8094 26180 8146
rect 25900 8092 26180 8094
rect 25900 8082 25956 8092
rect 25676 7868 26068 7924
rect 25116 5954 25172 5964
rect 25228 6580 25284 6590
rect 25228 6018 25284 6524
rect 25228 5966 25230 6018
rect 25282 5966 25284 6018
rect 25228 5954 25284 5966
rect 24444 5908 24500 5918
rect 24444 5814 24500 5852
rect 25452 5908 25508 5918
rect 25452 5814 25508 5852
rect 24220 4946 24276 4956
rect 24332 5794 24388 5806
rect 24332 5742 24334 5794
rect 24386 5742 24388 5794
rect 24332 4900 24388 5742
rect 23100 4162 23156 4172
rect 24220 4228 24276 4238
rect 24332 4228 24388 4844
rect 25228 5012 25284 5022
rect 25228 4338 25284 4956
rect 25228 4286 25230 4338
rect 25282 4286 25284 4338
rect 25228 4274 25284 4286
rect 24220 4226 24388 4228
rect 24220 4174 24222 4226
rect 24274 4174 24388 4226
rect 24220 4172 24388 4174
rect 24220 4162 24276 4172
rect 25228 4116 25284 4126
rect 24892 3668 24948 3678
rect 24892 800 24948 3612
rect 25228 3554 25284 4060
rect 25676 3780 25732 7868
rect 26012 7698 26068 7868
rect 26012 7646 26014 7698
rect 26066 7646 26068 7698
rect 26012 7634 26068 7646
rect 26124 7698 26180 8092
rect 26124 7646 26126 7698
rect 26178 7646 26180 7698
rect 26124 7634 26180 7646
rect 25900 7474 25956 7486
rect 25900 7422 25902 7474
rect 25954 7422 25956 7474
rect 25900 6692 25956 7422
rect 26236 7476 26292 7486
rect 26236 7252 26292 7420
rect 26348 7252 26404 8316
rect 26460 8278 26516 8316
rect 26684 7532 26964 7588
rect 26460 7476 26516 7486
rect 26684 7476 26740 7532
rect 26460 7474 26740 7476
rect 26460 7422 26462 7474
rect 26514 7422 26740 7474
rect 26460 7420 26740 7422
rect 26908 7476 26964 7532
rect 27132 7586 27188 9772
rect 27916 9602 27972 13580
rect 28252 13412 28308 13422
rect 28140 13356 28252 13412
rect 28028 13076 28084 13086
rect 28028 12962 28084 13020
rect 28028 12910 28030 12962
rect 28082 12910 28084 12962
rect 28028 12898 28084 12910
rect 28140 10612 28196 13356
rect 28252 13346 28308 13356
rect 28252 13188 28308 13198
rect 28252 12962 28308 13132
rect 28252 12910 28254 12962
rect 28306 12910 28308 12962
rect 28252 12898 28308 12910
rect 28364 12962 28420 14812
rect 28476 13748 28532 15484
rect 28588 15204 28644 15242
rect 28588 14868 28644 15148
rect 28700 15092 28756 16830
rect 29596 16772 29652 19854
rect 30156 19908 30212 19918
rect 30156 19814 30212 19852
rect 30828 19908 30884 19966
rect 31500 20020 31556 20030
rect 31500 19926 31556 19964
rect 31948 20018 32004 20860
rect 32060 20850 32116 20860
rect 32508 20356 32564 21422
rect 32508 20290 32564 20300
rect 31948 19966 31950 20018
rect 32002 19966 32004 20018
rect 30828 19842 30884 19852
rect 31612 19124 31668 19134
rect 31612 19030 31668 19068
rect 31948 19122 32004 19966
rect 32284 19908 32340 19918
rect 32284 19814 32340 19852
rect 31948 19070 31950 19122
rect 32002 19070 32004 19122
rect 31724 19010 31780 19022
rect 31724 18958 31726 19010
rect 31778 18958 31780 19010
rect 31612 18228 31668 18238
rect 31052 18226 31668 18228
rect 31052 18174 31614 18226
rect 31666 18174 31668 18226
rect 31052 18172 31668 18174
rect 30044 17554 30100 17566
rect 30044 17502 30046 17554
rect 30098 17502 30100 17554
rect 30044 17108 30100 17502
rect 30044 17042 30100 17052
rect 30716 17108 30772 17118
rect 30716 16994 30772 17052
rect 30716 16942 30718 16994
rect 30770 16942 30772 16994
rect 30716 16930 30772 16942
rect 31052 16884 31108 18172
rect 31612 18162 31668 18172
rect 31724 17780 31780 18958
rect 31948 18900 32004 19070
rect 32172 19124 32228 19134
rect 32620 19124 32676 23660
rect 32732 22372 32788 22382
rect 32732 22278 32788 22316
rect 32844 19908 32900 43708
rect 32956 32788 33012 50540
rect 34076 50530 34132 50542
rect 35868 50596 35924 50606
rect 35868 50502 35924 50540
rect 36092 50594 36148 50606
rect 36092 50542 36094 50594
rect 36146 50542 36148 50594
rect 35644 50036 35700 50046
rect 35532 49924 35588 49934
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 35420 49028 35476 49038
rect 35532 49028 35588 49868
rect 35420 49026 35588 49028
rect 35420 48974 35422 49026
rect 35474 48974 35588 49026
rect 35420 48972 35588 48974
rect 35420 48962 35476 48972
rect 34860 48914 34916 48926
rect 34860 48862 34862 48914
rect 34914 48862 34916 48914
rect 33628 48804 33684 48814
rect 34860 48804 34916 48862
rect 33628 48802 34916 48804
rect 33628 48750 33630 48802
rect 33682 48750 34916 48802
rect 33628 48748 34916 48750
rect 33628 48738 33684 48748
rect 34636 48580 34692 48590
rect 34636 48466 34692 48524
rect 34636 48414 34638 48466
rect 34690 48414 34692 48466
rect 34412 48244 34468 48254
rect 34412 48150 34468 48188
rect 33292 48132 33348 48142
rect 33292 48038 33348 48076
rect 33628 48130 33684 48142
rect 33628 48078 33630 48130
rect 33682 48078 33684 48130
rect 33628 47572 33684 48078
rect 33964 47572 34020 47582
rect 33628 47516 33964 47572
rect 33964 47478 34020 47516
rect 34524 47458 34580 47470
rect 34524 47406 34526 47458
rect 34578 47406 34580 47458
rect 33068 46788 33124 46798
rect 33068 46694 33124 46732
rect 33180 46788 33236 46798
rect 33740 46788 33796 46798
rect 33180 46786 33348 46788
rect 33180 46734 33182 46786
rect 33234 46734 33348 46786
rect 33180 46732 33348 46734
rect 33180 46722 33236 46732
rect 33292 46116 33348 46732
rect 33740 46694 33796 46732
rect 33404 46676 33460 46686
rect 33404 46582 33460 46620
rect 34188 46564 34244 46574
rect 34524 46564 34580 47406
rect 34188 46562 34580 46564
rect 34188 46510 34190 46562
rect 34242 46510 34580 46562
rect 34188 46508 34580 46510
rect 34188 46452 34244 46508
rect 33292 46050 33348 46060
rect 33852 46396 34244 46452
rect 33068 44994 33124 45006
rect 33068 44942 33070 44994
rect 33122 44942 33124 44994
rect 33068 44660 33124 44942
rect 33740 44996 33796 45006
rect 33740 44902 33796 44940
rect 33180 44884 33236 44894
rect 33180 44882 33684 44884
rect 33180 44830 33182 44882
rect 33234 44830 33684 44882
rect 33180 44828 33684 44830
rect 33180 44818 33236 44828
rect 33068 44594 33124 44604
rect 33628 44434 33684 44828
rect 33628 44382 33630 44434
rect 33682 44382 33684 44434
rect 33628 44370 33684 44382
rect 33628 43764 33684 43774
rect 33180 43426 33236 43438
rect 33180 43374 33182 43426
rect 33234 43374 33236 43426
rect 33180 43316 33236 43374
rect 33180 43250 33236 43260
rect 33628 42754 33684 43708
rect 33628 42702 33630 42754
rect 33682 42702 33684 42754
rect 33628 42690 33684 42702
rect 33068 41860 33124 41870
rect 33068 41766 33124 41804
rect 33628 41860 33684 41870
rect 33628 41766 33684 41804
rect 33180 41748 33236 41758
rect 33180 41746 33572 41748
rect 33180 41694 33182 41746
rect 33234 41694 33572 41746
rect 33180 41692 33572 41694
rect 33180 41682 33236 41692
rect 33516 41298 33572 41692
rect 33516 41246 33518 41298
rect 33570 41246 33572 41298
rect 33516 41234 33572 41246
rect 33516 39508 33572 39518
rect 33740 39508 33796 39518
rect 33516 39506 33796 39508
rect 33516 39454 33518 39506
rect 33570 39454 33742 39506
rect 33794 39454 33796 39506
rect 33516 39452 33796 39454
rect 33516 39442 33572 39452
rect 33740 39442 33796 39452
rect 33180 39394 33236 39406
rect 33180 39342 33182 39394
rect 33234 39342 33236 39394
rect 33180 38612 33236 39342
rect 33404 39394 33460 39406
rect 33404 39342 33406 39394
rect 33458 39342 33460 39394
rect 33404 38948 33460 39342
rect 33404 38668 33460 38892
rect 33404 38612 33572 38668
rect 33180 38546 33236 38556
rect 33516 38162 33572 38612
rect 33516 38110 33518 38162
rect 33570 38110 33572 38162
rect 33516 38098 33572 38110
rect 33180 37154 33236 37166
rect 33180 37102 33182 37154
rect 33234 37102 33236 37154
rect 33180 36708 33236 37102
rect 33180 36642 33236 36652
rect 33516 37044 33572 37054
rect 33516 36482 33572 36988
rect 33516 36430 33518 36482
rect 33570 36430 33572 36482
rect 33516 36418 33572 36430
rect 33068 36258 33124 36270
rect 33068 36206 33070 36258
rect 33122 36206 33124 36258
rect 33068 36148 33124 36206
rect 33292 36260 33348 36270
rect 33292 36166 33348 36204
rect 33404 36258 33460 36270
rect 33404 36206 33406 36258
rect 33458 36206 33460 36258
rect 33124 36092 33236 36148
rect 33068 36082 33124 36092
rect 33180 35922 33236 36092
rect 33180 35870 33182 35922
rect 33234 35870 33236 35922
rect 33180 35858 33236 35870
rect 33068 35700 33124 35710
rect 33068 34914 33124 35644
rect 33404 35252 33460 36206
rect 33852 36148 33908 46396
rect 34412 45220 34468 45230
rect 34412 44324 34468 45164
rect 34636 44548 34692 48414
rect 34748 48356 34804 48366
rect 34748 48242 34804 48300
rect 34748 48190 34750 48242
rect 34802 48190 34804 48242
rect 34748 48178 34804 48190
rect 34636 44482 34692 44492
rect 34412 44322 34692 44324
rect 34412 44270 34414 44322
rect 34466 44270 34692 44322
rect 34412 44268 34692 44270
rect 34412 44258 34468 44268
rect 34636 43764 34692 44268
rect 34636 43538 34692 43708
rect 34636 43486 34638 43538
rect 34690 43486 34692 43538
rect 34636 43474 34692 43486
rect 34300 42642 34356 42654
rect 34300 42590 34302 42642
rect 34354 42590 34356 42642
rect 34300 41972 34356 42590
rect 34300 41906 34356 41916
rect 34300 41186 34356 41198
rect 34300 41134 34302 41186
rect 34354 41134 34356 41186
rect 34300 40404 34356 41134
rect 34300 40338 34356 40348
rect 34524 40290 34580 40302
rect 34524 40238 34526 40290
rect 34578 40238 34580 40290
rect 34524 39842 34580 40238
rect 34860 40068 34916 48748
rect 35084 48244 35140 48254
rect 34972 48188 35084 48244
rect 34972 47570 35028 48188
rect 35084 48150 35140 48188
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 34972 47518 34974 47570
rect 35026 47518 35028 47570
rect 34972 47506 35028 47518
rect 35532 47458 35588 48972
rect 35532 47406 35534 47458
rect 35586 47406 35588 47458
rect 35532 46898 35588 47406
rect 35644 49138 35700 49980
rect 35644 49086 35646 49138
rect 35698 49086 35700 49138
rect 35644 47348 35700 49086
rect 36092 47572 36148 50542
rect 36428 50596 36484 50606
rect 36540 50596 36596 51212
rect 37100 51202 37156 51212
rect 36428 50594 36596 50596
rect 36428 50542 36430 50594
rect 36482 50542 36596 50594
rect 36428 50540 36596 50542
rect 36428 50530 36484 50540
rect 36540 49810 36596 50540
rect 37100 50596 37156 50606
rect 37100 50502 37156 50540
rect 37212 50428 37268 51884
rect 37436 50428 37492 52108
rect 37772 51492 37828 51502
rect 37884 51492 37940 53452
rect 37996 53442 38052 53452
rect 37996 53060 38052 53070
rect 37996 52162 38052 53004
rect 37996 52110 37998 52162
rect 38050 52110 38052 52162
rect 37996 52098 38052 52110
rect 37828 51436 37940 51492
rect 37772 51398 37828 51436
rect 37548 51380 37604 51390
rect 37548 51286 37604 51324
rect 38220 51380 38276 51390
rect 38220 51286 38276 51324
rect 38332 50428 38388 55916
rect 52668 55468 52724 56142
rect 52892 56082 52948 56364
rect 57820 56194 57876 56206
rect 57820 56142 57822 56194
rect 57874 56142 57876 56194
rect 52892 56030 52894 56082
rect 52946 56030 52948 56082
rect 52892 56018 52948 56030
rect 57596 56084 57652 56094
rect 57596 55990 57652 56028
rect 57820 55468 57876 56142
rect 58156 56084 58212 56094
rect 58156 55990 58212 56028
rect 40236 55412 40292 55422
rect 40236 55318 40292 55356
rect 41804 55412 41860 55422
rect 40796 55298 40852 55310
rect 40796 55246 40798 55298
rect 40850 55246 40852 55298
rect 40684 55188 40740 55198
rect 40684 55094 40740 55132
rect 40236 54740 40292 54750
rect 40236 54646 40292 54684
rect 40124 54628 40180 54638
rect 40124 54534 40180 54572
rect 40348 54290 40404 54302
rect 40348 54238 40350 54290
rect 40402 54238 40404 54290
rect 40348 53956 40404 54238
rect 40572 53956 40628 53966
rect 40348 53954 40628 53956
rect 40348 53902 40350 53954
rect 40402 53902 40574 53954
rect 40626 53902 40628 53954
rect 40348 53900 40628 53902
rect 40348 53890 40404 53900
rect 40572 53890 40628 53900
rect 39116 53844 39172 53854
rect 39116 53750 39172 53788
rect 40012 53844 40068 53854
rect 40012 53750 40068 53788
rect 39452 53732 39508 53742
rect 39788 53732 39844 53742
rect 39452 53730 39844 53732
rect 39452 53678 39454 53730
rect 39506 53678 39790 53730
rect 39842 53678 39844 53730
rect 39452 53676 39844 53678
rect 39452 53666 39508 53676
rect 39228 53506 39284 53518
rect 39228 53454 39230 53506
rect 39282 53454 39284 53506
rect 39228 52948 39284 53454
rect 39228 52882 39284 52892
rect 38780 52724 38836 52734
rect 38780 52274 38836 52668
rect 38780 52222 38782 52274
rect 38834 52222 38836 52274
rect 38780 52210 38836 52222
rect 39788 52164 39844 53676
rect 40796 53732 40852 55246
rect 41020 55298 41076 55310
rect 41020 55246 41022 55298
rect 41074 55246 41076 55298
rect 41020 54740 41076 55246
rect 41244 55300 41300 55310
rect 41300 55244 41524 55300
rect 41244 55206 41300 55244
rect 41020 54674 41076 54684
rect 41468 54738 41524 55244
rect 41804 54740 41860 55356
rect 42700 55412 42756 55422
rect 48860 55412 48916 55422
rect 42700 55410 43204 55412
rect 42700 55358 42702 55410
rect 42754 55358 43204 55410
rect 42700 55356 43204 55358
rect 42700 55346 42756 55356
rect 42364 55300 42420 55310
rect 42364 55206 42420 55244
rect 41468 54686 41470 54738
rect 41522 54686 41524 54738
rect 41468 54674 41524 54686
rect 41580 54738 41860 54740
rect 41580 54686 41806 54738
rect 41858 54686 41860 54738
rect 41580 54684 41860 54686
rect 40908 54628 40964 54638
rect 40908 54514 40964 54572
rect 41580 54516 41636 54684
rect 41804 54674 41860 54684
rect 42588 55074 42644 55086
rect 42588 55022 42590 55074
rect 42642 55022 42644 55074
rect 42140 54628 42196 54638
rect 42196 54572 42420 54628
rect 42140 54534 42196 54572
rect 40908 54462 40910 54514
rect 40962 54462 40964 54514
rect 40908 54450 40964 54462
rect 41356 54460 41636 54516
rect 41132 54292 41188 54302
rect 41020 54290 41188 54292
rect 41020 54238 41134 54290
rect 41186 54238 41188 54290
rect 41020 54236 41188 54238
rect 40796 53666 40852 53676
rect 40908 53956 40964 53966
rect 41020 53956 41076 54236
rect 41132 54226 41188 54236
rect 41244 53956 41300 53966
rect 40908 53954 41076 53956
rect 40908 53902 40910 53954
rect 40962 53902 41076 53954
rect 40908 53900 41076 53902
rect 41132 53900 41244 53956
rect 40012 53508 40068 53518
rect 40012 52948 40068 53452
rect 40796 53508 40852 53518
rect 40796 53414 40852 53452
rect 40012 52946 40516 52948
rect 40012 52894 40014 52946
rect 40066 52894 40516 52946
rect 40012 52892 40516 52894
rect 40012 52882 40068 52892
rect 39788 52108 40404 52164
rect 37212 50372 37380 50428
rect 37436 50372 37604 50428
rect 37100 50036 37156 50046
rect 37100 49942 37156 49980
rect 36540 49758 36542 49810
rect 36594 49758 36596 49810
rect 36204 48802 36260 48814
rect 36204 48750 36206 48802
rect 36258 48750 36260 48802
rect 36204 48356 36260 48750
rect 36540 48804 36596 49758
rect 36652 49588 36708 49598
rect 36652 49494 36708 49532
rect 36988 49028 37044 49038
rect 36988 49026 37156 49028
rect 36988 48974 36990 49026
rect 37042 48974 37156 49026
rect 36988 48972 37156 48974
rect 36988 48962 37044 48972
rect 36540 48748 37044 48804
rect 36204 48262 36260 48300
rect 36316 48468 36372 48478
rect 35644 47346 36036 47348
rect 35644 47294 35646 47346
rect 35698 47294 36036 47346
rect 35644 47292 36036 47294
rect 35644 47282 35700 47292
rect 35532 46846 35534 46898
rect 35586 46846 35588 46898
rect 35532 46834 35588 46846
rect 35980 46898 36036 47292
rect 36092 47124 36148 47516
rect 36316 47348 36372 48412
rect 36316 47254 36372 47292
rect 36428 47236 36484 47246
rect 36428 47234 36820 47236
rect 36428 47182 36430 47234
rect 36482 47182 36820 47234
rect 36428 47180 36820 47182
rect 36428 47170 36484 47180
rect 36092 47068 36372 47124
rect 36316 47012 36372 47068
rect 36316 46956 36596 47012
rect 35980 46846 35982 46898
rect 36034 46846 36036 46898
rect 35980 46834 36036 46846
rect 36540 46786 36596 46956
rect 36764 46898 36820 47180
rect 36764 46846 36766 46898
rect 36818 46846 36820 46898
rect 36764 46834 36820 46846
rect 36988 46898 37044 48748
rect 37100 48242 37156 48972
rect 37212 49026 37268 49038
rect 37212 48974 37214 49026
rect 37266 48974 37268 49026
rect 37212 48468 37268 48974
rect 37212 48402 37268 48412
rect 37324 48466 37380 50372
rect 37324 48414 37326 48466
rect 37378 48414 37380 48466
rect 37324 48402 37380 48414
rect 37436 49588 37492 49598
rect 37436 49026 37492 49532
rect 37548 49252 37604 50372
rect 38220 50372 38388 50428
rect 38444 51268 38500 51278
rect 37660 49924 37716 49934
rect 37660 49830 37716 49868
rect 37548 49186 37604 49196
rect 37436 48974 37438 49026
rect 37490 48974 37492 49026
rect 37436 48356 37492 48974
rect 37548 49028 37604 49038
rect 38108 49028 38164 49038
rect 37548 49026 38164 49028
rect 37548 48974 37550 49026
rect 37602 48974 38110 49026
rect 38162 48974 38164 49026
rect 37548 48972 38164 48974
rect 37548 48962 37604 48972
rect 38108 48962 38164 48972
rect 37660 48804 37716 48814
rect 37660 48802 37828 48804
rect 37660 48750 37662 48802
rect 37714 48750 37828 48802
rect 37660 48748 37828 48750
rect 37660 48738 37716 48748
rect 37660 48356 37716 48366
rect 37436 48354 37716 48356
rect 37436 48302 37662 48354
rect 37714 48302 37716 48354
rect 37436 48300 37716 48302
rect 37100 48190 37102 48242
rect 37154 48190 37156 48242
rect 37100 48132 37156 48190
rect 37100 48066 37156 48076
rect 37212 48244 37268 48254
rect 37212 47458 37268 48188
rect 37212 47406 37214 47458
rect 37266 47406 37268 47458
rect 37212 47394 37268 47406
rect 37436 47346 37492 48300
rect 37660 48290 37716 48300
rect 37436 47294 37438 47346
rect 37490 47294 37492 47346
rect 37436 47282 37492 47294
rect 37548 48132 37604 48142
rect 37772 48132 37828 48748
rect 37604 48076 37828 48132
rect 37548 47346 37604 48076
rect 37884 48020 37940 48030
rect 37884 47458 37940 47964
rect 37884 47406 37886 47458
rect 37938 47406 37940 47458
rect 37884 47394 37940 47406
rect 37548 47294 37550 47346
rect 37602 47294 37604 47346
rect 37436 47124 37492 47134
rect 36988 46846 36990 46898
rect 37042 46846 37044 46898
rect 36988 46834 37044 46846
rect 37100 47012 37156 47022
rect 36540 46734 36542 46786
rect 36594 46734 36596 46786
rect 36540 46722 36596 46734
rect 37100 46562 37156 46956
rect 37212 46900 37268 46910
rect 37212 46674 37268 46844
rect 37212 46622 37214 46674
rect 37266 46622 37268 46674
rect 37212 46610 37268 46622
rect 37100 46510 37102 46562
rect 37154 46510 37156 46562
rect 37100 46498 37156 46510
rect 37324 46340 37380 46350
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 36988 46284 37324 46340
rect 36204 46004 36260 46014
rect 36204 45890 36260 45948
rect 36204 45838 36206 45890
rect 36258 45838 36260 45890
rect 36204 45106 36260 45838
rect 36204 45054 36206 45106
rect 36258 45054 36260 45106
rect 36204 45042 36260 45054
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 36316 44210 36372 44222
rect 36316 44158 36318 44210
rect 36370 44158 36372 44210
rect 36204 44100 36260 44110
rect 35420 44098 36260 44100
rect 35420 44046 36206 44098
rect 36258 44046 36260 44098
rect 35420 44044 36260 44046
rect 35420 43650 35476 44044
rect 36204 44034 36260 44044
rect 35420 43598 35422 43650
rect 35474 43598 35476 43650
rect 35420 43586 35476 43598
rect 36316 43652 36372 44158
rect 36316 43586 36372 43596
rect 34524 39790 34526 39842
rect 34578 39790 34580 39842
rect 34524 39778 34580 39790
rect 34636 40012 34916 40068
rect 35084 43428 35140 43438
rect 34076 39506 34132 39518
rect 34076 39454 34078 39506
rect 34130 39454 34132 39506
rect 33964 39394 34020 39406
rect 33964 39342 33966 39394
rect 34018 39342 34020 39394
rect 33964 38836 34020 39342
rect 34076 39284 34132 39454
rect 34076 39218 34132 39228
rect 34524 39394 34580 39406
rect 34524 39342 34526 39394
rect 34578 39342 34580 39394
rect 34524 39284 34580 39342
rect 34524 39218 34580 39228
rect 33964 38668 34020 38780
rect 33964 38612 34132 38668
rect 34076 38162 34132 38612
rect 34188 38276 34244 38286
rect 34412 38276 34468 38286
rect 34188 38274 34468 38276
rect 34188 38222 34190 38274
rect 34242 38222 34414 38274
rect 34466 38222 34468 38274
rect 34188 38220 34468 38222
rect 34188 38210 34244 38220
rect 34412 38210 34468 38220
rect 34076 38110 34078 38162
rect 34130 38110 34132 38162
rect 34076 38098 34132 38110
rect 34636 38164 34692 40012
rect 34636 38098 34692 38108
rect 34748 39842 34804 39854
rect 34748 39790 34750 39842
rect 34802 39790 34804 39842
rect 34748 38836 34804 39790
rect 34860 38948 34916 38958
rect 34860 38854 34916 38892
rect 34748 38162 34804 38780
rect 34972 38834 35028 38846
rect 34972 38782 34974 38834
rect 35026 38782 35028 38834
rect 34972 38274 35028 38782
rect 34972 38222 34974 38274
rect 35026 38222 35028 38274
rect 34972 38210 35028 38222
rect 34748 38110 34750 38162
rect 34802 38110 34804 38162
rect 34748 38098 34804 38110
rect 34188 38052 34244 38062
rect 33964 36260 34020 36270
rect 33964 36166 34020 36204
rect 33852 36082 33908 36092
rect 33404 35196 33684 35252
rect 33068 34862 33070 34914
rect 33122 34862 33124 34914
rect 33068 34850 33124 34862
rect 33180 34916 33236 34926
rect 33180 34356 33236 34860
rect 33628 34914 33684 35196
rect 33628 34862 33630 34914
rect 33682 34862 33684 34914
rect 33628 34850 33684 34862
rect 33516 34802 33572 34814
rect 33516 34750 33518 34802
rect 33570 34750 33572 34802
rect 33292 34692 33348 34702
rect 33292 34598 33348 34636
rect 33516 34356 33572 34750
rect 33628 34356 33684 34366
rect 33516 34354 34132 34356
rect 33516 34302 33630 34354
rect 33682 34302 34132 34354
rect 33516 34300 34132 34302
rect 33180 34242 33236 34300
rect 33628 34290 33684 34300
rect 33180 34190 33182 34242
rect 33234 34190 33236 34242
rect 33180 33124 33236 34190
rect 34076 34242 34132 34300
rect 34076 34190 34078 34242
rect 34130 34190 34132 34242
rect 34076 34178 34132 34190
rect 33740 34020 33796 34030
rect 33740 34018 34132 34020
rect 33740 33966 33742 34018
rect 33794 33966 34132 34018
rect 33740 33964 34132 33966
rect 33740 33954 33796 33964
rect 33292 33906 33348 33918
rect 33292 33854 33294 33906
rect 33346 33854 33348 33906
rect 33292 33572 33348 33854
rect 33292 33506 33348 33516
rect 33180 33058 33236 33068
rect 33852 33124 33908 33134
rect 32956 32732 33460 32788
rect 33180 31220 33236 31230
rect 33180 31126 33236 31164
rect 33180 30324 33236 30334
rect 33180 29650 33236 30268
rect 33180 29598 33182 29650
rect 33234 29598 33236 29650
rect 33180 29586 33236 29598
rect 33292 27860 33348 27870
rect 33292 27766 33348 27804
rect 33068 27634 33124 27646
rect 33068 27582 33070 27634
rect 33122 27582 33124 27634
rect 33068 27188 33124 27582
rect 32956 27076 33012 27086
rect 33068 27076 33124 27132
rect 32956 27074 33124 27076
rect 32956 27022 32958 27074
rect 33010 27022 33124 27074
rect 32956 27020 33124 27022
rect 32956 27010 33012 27020
rect 33068 26290 33124 26302
rect 33068 26238 33070 26290
rect 33122 26238 33124 26290
rect 33068 23380 33124 26238
rect 33180 24276 33236 24286
rect 33180 24050 33236 24220
rect 33180 23998 33182 24050
rect 33234 23998 33236 24050
rect 33180 23986 33236 23998
rect 33180 23716 33236 23726
rect 33236 23660 33348 23716
rect 33180 23650 33236 23660
rect 32956 23324 33068 23380
rect 32956 21588 33012 23324
rect 33068 23314 33124 23324
rect 33292 23378 33348 23660
rect 33292 23326 33294 23378
rect 33346 23326 33348 23378
rect 33292 23314 33348 23326
rect 33068 23154 33124 23166
rect 33068 23102 33070 23154
rect 33122 23102 33124 23154
rect 33068 22708 33124 23102
rect 33180 23044 33236 23054
rect 33180 22950 33236 22988
rect 33068 22642 33124 22652
rect 33180 22820 33236 22830
rect 33180 22148 33236 22764
rect 33404 22260 33460 32732
rect 33852 32562 33908 33068
rect 33852 32510 33854 32562
rect 33906 32510 33908 32562
rect 33852 32498 33908 32510
rect 34076 32564 34132 33964
rect 34188 33012 34244 37996
rect 34636 37828 34692 37838
rect 34300 36596 34356 36606
rect 34300 33908 34356 36540
rect 34636 35308 34692 37772
rect 34412 35252 34468 35262
rect 34412 34468 34468 35196
rect 34412 34402 34468 34412
rect 34524 35252 34692 35308
rect 34972 36372 35028 36382
rect 34972 36258 35028 36316
rect 34972 36206 34974 36258
rect 35026 36206 35028 36258
rect 34972 35252 35028 36206
rect 34300 33814 34356 33852
rect 34188 32946 34244 32956
rect 34524 32900 34580 35252
rect 34972 35186 35028 35196
rect 34636 34914 34692 34926
rect 34636 34862 34638 34914
rect 34690 34862 34692 34914
rect 34636 34356 34692 34862
rect 34748 34916 34804 34954
rect 35084 34916 35140 43372
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 36428 42868 36484 42878
rect 36428 42774 36484 42812
rect 35420 42196 35476 42206
rect 35308 41972 35364 41982
rect 35308 41878 35364 41916
rect 35420 41970 35476 42140
rect 35420 41918 35422 41970
rect 35474 41918 35476 41970
rect 35420 41906 35476 41918
rect 35868 41860 35924 41870
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35756 40404 35812 40414
rect 35756 40310 35812 40348
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35308 39618 35364 39630
rect 35308 39566 35310 39618
rect 35362 39566 35364 39618
rect 35308 39396 35364 39566
rect 35756 39620 35812 39630
rect 35868 39620 35924 41804
rect 36428 41076 36484 41086
rect 36428 40514 36484 41020
rect 36428 40462 36430 40514
rect 36482 40462 36484 40514
rect 36428 40450 36484 40462
rect 36988 40180 37044 46284
rect 37324 46274 37380 46284
rect 37100 46004 37156 46014
rect 37100 45910 37156 45948
rect 37212 41972 37268 41982
rect 37436 41972 37492 47068
rect 37548 43540 37604 47294
rect 38108 47346 38164 47358
rect 38108 47294 38110 47346
rect 38162 47294 38164 47346
rect 38108 47124 38164 47294
rect 38108 47058 38164 47068
rect 38220 46340 38276 50372
rect 38332 48802 38388 48814
rect 38332 48750 38334 48802
rect 38386 48750 38388 48802
rect 38332 48244 38388 48750
rect 38332 48178 38388 48188
rect 38332 47908 38388 47918
rect 38332 47682 38388 47852
rect 38332 47630 38334 47682
rect 38386 47630 38388 47682
rect 38332 47618 38388 47630
rect 38444 46676 38500 51212
rect 40348 50372 40404 52108
rect 38556 49812 38612 49822
rect 38556 49138 38612 49756
rect 39676 49364 39732 49374
rect 39116 49252 39172 49262
rect 39116 49158 39172 49196
rect 38556 49086 38558 49138
rect 38610 49086 38612 49138
rect 38556 49074 38612 49086
rect 39676 49138 39732 49308
rect 39676 49086 39678 49138
rect 39730 49086 39732 49138
rect 39676 49074 39732 49086
rect 39340 49026 39396 49038
rect 39340 48974 39342 49026
rect 39394 48974 39396 49026
rect 38556 48916 38612 48926
rect 39340 48916 39396 48974
rect 39564 49028 39620 49038
rect 39564 48934 39620 48972
rect 40348 49028 40404 50316
rect 40348 48934 40404 48972
rect 38556 48822 38612 48860
rect 38668 48860 39396 48916
rect 38668 48802 38724 48860
rect 38668 48750 38670 48802
rect 38722 48750 38724 48802
rect 38668 48580 38724 48750
rect 39788 48804 39844 48814
rect 38444 46610 38500 46620
rect 38556 48524 38724 48580
rect 38780 48692 38836 48702
rect 38556 47458 38612 48524
rect 38668 47572 38724 47582
rect 38668 47478 38724 47516
rect 38556 47406 38558 47458
rect 38610 47406 38612 47458
rect 38220 46274 38276 46284
rect 37996 46116 38052 46126
rect 38556 46116 38612 47406
rect 38780 47458 38836 48636
rect 39676 48244 39732 48254
rect 39676 48150 39732 48188
rect 39340 48132 39396 48142
rect 39340 48038 39396 48076
rect 38780 47406 38782 47458
rect 38834 47406 38836 47458
rect 38780 47394 38836 47406
rect 39228 48018 39284 48030
rect 39228 47966 39230 48018
rect 39282 47966 39284 48018
rect 39228 46900 39284 47966
rect 39228 46834 39284 46844
rect 37996 46114 38612 46116
rect 37996 46062 37998 46114
rect 38050 46062 38612 46114
rect 37996 46060 38612 46062
rect 39788 46116 39844 48748
rect 40124 48580 40180 48590
rect 40124 48466 40180 48524
rect 40124 48414 40126 48466
rect 40178 48414 40180 48466
rect 40124 48402 40180 48414
rect 39900 48242 39956 48254
rect 39900 48190 39902 48242
rect 39954 48190 39956 48242
rect 39900 47012 39956 48190
rect 40348 48244 40404 48254
rect 40348 48150 40404 48188
rect 40236 48020 40292 48030
rect 40236 47926 40292 47964
rect 39900 46946 39956 46956
rect 40012 46116 40068 46126
rect 39788 46114 40068 46116
rect 39788 46062 40014 46114
rect 40066 46062 40068 46114
rect 39788 46060 40068 46062
rect 37996 46050 38052 46060
rect 40012 46050 40068 46060
rect 40460 46004 40516 52892
rect 40908 52946 40964 53900
rect 41132 53842 41188 53900
rect 41244 53890 41300 53900
rect 41132 53790 41134 53842
rect 41186 53790 41188 53842
rect 41132 53778 41188 53790
rect 41244 53732 41300 53742
rect 40908 52894 40910 52946
rect 40962 52894 40964 52946
rect 40908 52882 40964 52894
rect 41132 52948 41188 52958
rect 41244 52948 41300 53676
rect 41356 53730 41412 54460
rect 41356 53678 41358 53730
rect 41410 53678 41412 53730
rect 41356 53666 41412 53678
rect 41692 53844 41748 53854
rect 41692 53730 41748 53788
rect 41692 53678 41694 53730
rect 41746 53678 41748 53730
rect 41692 53666 41748 53678
rect 41580 53618 41636 53630
rect 41580 53566 41582 53618
rect 41634 53566 41636 53618
rect 41356 52948 41412 52958
rect 41244 52892 41356 52948
rect 41132 52854 41188 52892
rect 41356 52854 41412 52892
rect 41468 52724 41524 52734
rect 41468 52630 41524 52668
rect 40908 52276 40964 52286
rect 41580 52276 41636 53566
rect 42140 53508 42196 53518
rect 42140 53414 42196 53452
rect 40908 52274 41636 52276
rect 40908 52222 40910 52274
rect 40962 52222 41636 52274
rect 40908 52220 41636 52222
rect 40908 52210 40964 52220
rect 41580 52162 41636 52220
rect 41580 52110 41582 52162
rect 41634 52110 41636 52162
rect 41580 52098 41636 52110
rect 42252 52162 42308 52174
rect 42252 52110 42254 52162
rect 42306 52110 42308 52162
rect 41244 51938 41300 51950
rect 41244 51886 41246 51938
rect 41298 51886 41300 51938
rect 41244 50372 41300 51886
rect 42252 51940 42308 52110
rect 42252 51268 42308 51884
rect 42252 51202 42308 51212
rect 41244 50306 41300 50316
rect 41244 50092 41524 50148
rect 40908 49812 40964 49822
rect 40908 49718 40964 49756
rect 41132 49812 41188 49822
rect 41132 49718 41188 49756
rect 41020 49698 41076 49710
rect 41020 49646 41022 49698
rect 41074 49646 41076 49698
rect 41020 49364 41076 49646
rect 40684 49308 41076 49364
rect 40572 48804 40628 48814
rect 40572 48710 40628 48748
rect 40684 48356 40740 49308
rect 40908 49138 40964 49150
rect 41244 49140 41300 50092
rect 41468 50036 41524 50092
rect 41804 50036 41860 50046
rect 41468 50034 41860 50036
rect 41468 49982 41806 50034
rect 41858 49982 41860 50034
rect 41468 49980 41860 49982
rect 41804 49970 41860 49980
rect 40908 49086 40910 49138
rect 40962 49086 40964 49138
rect 40796 49028 40852 49038
rect 40796 48934 40852 48972
rect 40908 48804 40964 49086
rect 41020 49084 41300 49140
rect 41356 49922 41412 49934
rect 41356 49870 41358 49922
rect 41410 49870 41412 49922
rect 41020 49026 41076 49084
rect 41020 48974 41022 49026
rect 41074 48974 41076 49026
rect 41020 48962 41076 48974
rect 41356 49026 41412 49870
rect 41916 49698 41972 49710
rect 41916 49646 41918 49698
rect 41970 49646 41972 49698
rect 41356 48974 41358 49026
rect 41410 48974 41412 49026
rect 41356 48804 41412 48974
rect 41804 49364 41860 49374
rect 40908 48748 41412 48804
rect 41468 48804 41524 48814
rect 41692 48804 41748 48814
rect 41468 48710 41524 48748
rect 41580 48802 41748 48804
rect 41580 48750 41694 48802
rect 41746 48750 41748 48802
rect 41580 48748 41748 48750
rect 40684 48290 40740 48300
rect 41468 48244 41524 48254
rect 41580 48244 41636 48748
rect 41692 48738 41748 48748
rect 41468 48242 41636 48244
rect 41468 48190 41470 48242
rect 41522 48190 41636 48242
rect 41468 48188 41636 48190
rect 41692 48244 41748 48254
rect 41804 48244 41860 49308
rect 41692 48242 41860 48244
rect 41692 48190 41694 48242
rect 41746 48190 41860 48242
rect 41692 48188 41860 48190
rect 41916 48804 41972 49646
rect 42364 49698 42420 54572
rect 42588 54402 42644 55022
rect 42588 54350 42590 54402
rect 42642 54350 42644 54402
rect 42588 53956 42644 54350
rect 42476 52948 42532 52958
rect 42476 52050 42532 52892
rect 42476 51998 42478 52050
rect 42530 51998 42532 52050
rect 42476 51986 42532 51998
rect 42476 51492 42532 51502
rect 42588 51492 42644 53900
rect 43148 53954 43204 55356
rect 48748 55410 48916 55412
rect 48748 55358 48862 55410
rect 48914 55358 48916 55410
rect 48748 55356 48916 55358
rect 45500 55300 45556 55310
rect 45500 54514 45556 55244
rect 46060 55300 46116 55310
rect 46060 55206 46116 55244
rect 46732 55186 46788 55198
rect 46732 55134 46734 55186
rect 46786 55134 46788 55186
rect 46732 54740 46788 55134
rect 46732 54674 46788 54684
rect 47404 54740 47460 54750
rect 47404 54646 47460 54684
rect 45500 54462 45502 54514
rect 45554 54462 45556 54514
rect 45500 54450 45556 54462
rect 46508 54514 46564 54526
rect 46508 54462 46510 54514
rect 46562 54462 46564 54514
rect 43148 53902 43150 53954
rect 43202 53902 43204 53954
rect 43148 53890 43204 53902
rect 43484 54404 43540 54414
rect 43036 53730 43092 53742
rect 43036 53678 43038 53730
rect 43090 53678 43092 53730
rect 43036 53508 43092 53678
rect 43036 52388 43092 53452
rect 43372 53730 43428 53742
rect 43372 53678 43374 53730
rect 43426 53678 43428 53730
rect 43372 52948 43428 53678
rect 43484 53730 43540 54348
rect 44716 54404 44772 54414
rect 44716 54310 44772 54348
rect 43484 53678 43486 53730
rect 43538 53678 43540 53730
rect 43484 53666 43540 53678
rect 46508 53508 46564 54462
rect 46508 53442 46564 53452
rect 46732 54514 46788 54526
rect 46732 54462 46734 54514
rect 46786 54462 46788 54514
rect 43372 52882 43428 52892
rect 45052 53172 45108 53182
rect 43036 52322 43092 52332
rect 43708 52388 43764 52398
rect 43708 52294 43764 52332
rect 45052 52386 45108 53116
rect 46732 53172 46788 54462
rect 47628 54516 47684 54526
rect 46956 54404 47012 54414
rect 47292 54404 47348 54414
rect 46956 54402 47348 54404
rect 46956 54350 46958 54402
rect 47010 54350 47294 54402
rect 47346 54350 47348 54402
rect 46956 54348 47348 54350
rect 46956 54338 47012 54348
rect 47292 54338 47348 54348
rect 46732 53078 46788 53116
rect 45052 52334 45054 52386
rect 45106 52334 45108 52386
rect 45052 52322 45108 52334
rect 45276 52948 45332 52958
rect 45276 52386 45332 52892
rect 46284 52948 46340 52958
rect 45276 52334 45278 52386
rect 45330 52334 45332 52386
rect 45276 52322 45332 52334
rect 45948 52388 46004 52398
rect 45948 52294 46004 52332
rect 46284 52386 46340 52892
rect 46956 52948 47012 52958
rect 46956 52854 47012 52892
rect 46284 52334 46286 52386
rect 46338 52334 46340 52386
rect 46284 52322 46340 52334
rect 44044 52274 44100 52286
rect 44044 52222 44046 52274
rect 44098 52222 44100 52274
rect 42700 52162 42756 52174
rect 42700 52110 42702 52162
rect 42754 52110 42756 52162
rect 42700 51940 42756 52110
rect 44044 52164 44100 52222
rect 44828 52164 44884 52174
rect 45724 52164 45780 52174
rect 44044 52162 44884 52164
rect 44044 52110 44830 52162
rect 44882 52110 44884 52162
rect 44044 52108 44884 52110
rect 44828 52098 44884 52108
rect 45500 52162 45780 52164
rect 45500 52110 45726 52162
rect 45778 52110 45780 52162
rect 45500 52108 45780 52110
rect 45388 52050 45444 52062
rect 45388 51998 45390 52050
rect 45442 51998 45444 52050
rect 42700 51874 42756 51884
rect 43932 51940 43988 51950
rect 43932 51938 45220 51940
rect 43932 51886 43934 51938
rect 43986 51886 45220 51938
rect 43932 51884 45220 51886
rect 43932 51874 43988 51884
rect 42476 51490 42644 51492
rect 42476 51438 42478 51490
rect 42530 51438 42644 51490
rect 42476 51436 42644 51438
rect 42476 51426 42532 51436
rect 43260 51268 43316 51278
rect 43260 51174 43316 51212
rect 42588 51156 42644 51166
rect 42364 49646 42366 49698
rect 42418 49646 42420 49698
rect 42252 49588 42308 49598
rect 42140 49586 42308 49588
rect 42140 49534 42254 49586
rect 42306 49534 42308 49586
rect 42140 49532 42308 49534
rect 42140 49026 42196 49532
rect 42252 49522 42308 49532
rect 42140 48974 42142 49026
rect 42194 48974 42196 49026
rect 42140 48962 42196 48974
rect 42364 49028 42420 49646
rect 42364 48962 42420 48972
rect 42476 51154 42644 51156
rect 42476 51102 42590 51154
rect 42642 51102 42644 51154
rect 42476 51100 42644 51102
rect 42476 49140 42532 51100
rect 42588 51090 42644 51100
rect 42476 49084 43092 49140
rect 42476 49026 42532 49084
rect 42476 48974 42478 49026
rect 42530 48974 42532 49026
rect 42476 48962 42532 48974
rect 43036 49026 43092 49084
rect 43036 48974 43038 49026
rect 43090 48974 43092 49026
rect 43036 48962 43092 48974
rect 43148 49138 43204 49150
rect 44156 49140 44212 51884
rect 45164 50482 45220 51884
rect 45388 51490 45444 51998
rect 45388 51438 45390 51490
rect 45442 51438 45444 51490
rect 45388 51426 45444 51438
rect 45500 51268 45556 52108
rect 45724 52098 45780 52108
rect 46844 51940 46900 51950
rect 46844 51602 46900 51884
rect 47628 51828 47684 54460
rect 48300 54404 48356 54414
rect 48300 54310 48356 54348
rect 48636 53732 48692 53742
rect 48748 53732 48804 55356
rect 48860 55346 48916 55356
rect 52108 55410 52164 55422
rect 52108 55358 52110 55410
rect 52162 55358 52164 55410
rect 49308 55300 49364 55310
rect 49308 55206 49364 55244
rect 51996 55300 52052 55310
rect 49980 55186 50036 55198
rect 49980 55134 49982 55186
rect 50034 55134 50036 55186
rect 49980 53732 50036 55134
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 51996 54626 52052 55244
rect 51996 54574 51998 54626
rect 52050 54574 52052 54626
rect 51996 54562 52052 54574
rect 50764 53956 50820 53966
rect 50764 53954 51492 53956
rect 50764 53902 50766 53954
rect 50818 53902 51492 53954
rect 50764 53900 51492 53902
rect 50764 53890 50820 53900
rect 50540 53842 50596 53854
rect 50540 53790 50542 53842
rect 50594 53790 50596 53842
rect 50428 53732 50484 53742
rect 48636 53730 48916 53732
rect 48636 53678 48638 53730
rect 48690 53678 48916 53730
rect 48636 53676 48916 53678
rect 49980 53730 50484 53732
rect 49980 53678 50430 53730
rect 50482 53678 50484 53730
rect 49980 53676 50484 53678
rect 48636 53666 48692 53676
rect 48748 53508 48804 53518
rect 48748 53414 48804 53452
rect 48076 53172 48132 53182
rect 48076 52500 48132 53116
rect 48076 52444 48580 52500
rect 48076 52162 48132 52444
rect 48076 52110 48078 52162
rect 48130 52110 48132 52162
rect 48076 52098 48132 52110
rect 48188 52276 48244 52286
rect 48188 52050 48244 52220
rect 48412 52164 48468 52174
rect 48412 52070 48468 52108
rect 48524 52162 48580 52444
rect 48524 52110 48526 52162
rect 48578 52110 48580 52162
rect 48524 52098 48580 52110
rect 48860 52276 48916 53676
rect 50428 53666 50484 53676
rect 49644 53508 49700 53518
rect 50540 53508 50596 53790
rect 51436 53842 51492 53900
rect 51436 53790 51438 53842
rect 51490 53790 51492 53842
rect 51436 53778 51492 53790
rect 49700 53452 49812 53508
rect 49644 53442 49700 53452
rect 48860 52162 48916 52220
rect 48860 52110 48862 52162
rect 48914 52110 48916 52162
rect 48860 52098 48916 52110
rect 48972 52332 49700 52388
rect 48188 51998 48190 52050
rect 48242 51998 48244 52050
rect 48188 51986 48244 51998
rect 48860 51938 48916 51950
rect 48860 51886 48862 51938
rect 48914 51886 48916 51938
rect 47628 51772 48356 51828
rect 46844 51550 46846 51602
rect 46898 51550 46900 51602
rect 46844 51538 46900 51550
rect 45500 50594 45556 51212
rect 45500 50542 45502 50594
rect 45554 50542 45556 50594
rect 45500 50530 45556 50542
rect 46060 51378 46116 51390
rect 46060 51326 46062 51378
rect 46114 51326 46116 51378
rect 45164 50430 45166 50482
rect 45218 50430 45220 50482
rect 45164 50418 45220 50430
rect 46060 49476 46116 51326
rect 46508 51378 46564 51390
rect 46508 51326 46510 51378
rect 46562 51326 46564 51378
rect 46172 51156 46228 51166
rect 46172 50706 46228 51100
rect 46508 51156 46564 51326
rect 46508 51090 46564 51100
rect 46172 50654 46174 50706
rect 46226 50654 46228 50706
rect 46172 50642 46228 50654
rect 46060 49410 46116 49420
rect 46956 49476 47012 49486
rect 47012 49420 47124 49476
rect 46956 49410 47012 49420
rect 43148 49086 43150 49138
rect 43202 49086 43204 49138
rect 42588 48916 42644 48926
rect 42588 48914 42756 48916
rect 42588 48862 42590 48914
rect 42642 48862 42756 48914
rect 42588 48860 42756 48862
rect 42588 48850 42644 48860
rect 42252 48804 42308 48814
rect 41916 48802 42308 48804
rect 41916 48750 42254 48802
rect 42306 48750 42308 48802
rect 41916 48748 42308 48750
rect 41468 48178 41524 48188
rect 41692 48178 41748 48188
rect 40796 48020 40852 48030
rect 40684 48018 40852 48020
rect 40684 47966 40798 48018
rect 40850 47966 40852 48018
rect 40684 47964 40852 47966
rect 40684 47570 40740 47964
rect 40796 47954 40852 47964
rect 41244 48020 41300 48030
rect 41244 47926 41300 47964
rect 41916 47908 41972 48748
rect 42252 48738 42308 48748
rect 42364 48804 42420 48814
rect 42364 48580 42420 48748
rect 42700 48804 42756 48860
rect 42700 48738 42756 48748
rect 42364 48524 42868 48580
rect 42476 48356 42532 48366
rect 42476 48242 42532 48300
rect 42812 48354 42868 48524
rect 42812 48302 42814 48354
rect 42866 48302 42868 48354
rect 42812 48290 42868 48302
rect 42476 48190 42478 48242
rect 42530 48190 42532 48242
rect 42476 48178 42532 48190
rect 40684 47518 40686 47570
rect 40738 47518 40740 47570
rect 40684 47506 40740 47518
rect 41692 47852 41972 47908
rect 43036 48020 43092 48030
rect 43148 48020 43204 49086
rect 43932 49138 44212 49140
rect 43932 49086 44158 49138
rect 44210 49086 44212 49138
rect 43932 49084 44212 49086
rect 43596 49028 43652 49038
rect 43372 48916 43428 48926
rect 43372 48822 43428 48860
rect 43596 48466 43652 48972
rect 43932 48468 43988 49084
rect 44156 49074 44212 49084
rect 45388 49028 45444 49038
rect 45388 48934 45444 48972
rect 43596 48414 43598 48466
rect 43650 48414 43652 48466
rect 43596 48402 43652 48414
rect 43708 48466 43988 48468
rect 43708 48414 43934 48466
rect 43986 48414 43988 48466
rect 43708 48412 43988 48414
rect 43260 48244 43316 48254
rect 43484 48244 43540 48254
rect 43708 48244 43764 48412
rect 43932 48402 43988 48412
rect 44044 48916 44100 48926
rect 43316 48188 43428 48244
rect 43260 48150 43316 48188
rect 43036 48018 43204 48020
rect 43036 47966 43038 48018
rect 43090 47966 43204 48018
rect 43036 47964 43204 47966
rect 43036 47908 43092 47964
rect 40796 47234 40852 47246
rect 40796 47182 40798 47234
rect 40850 47182 40852 47234
rect 40796 46676 40852 47182
rect 41132 46788 41188 46798
rect 41132 46694 41188 46732
rect 41020 46676 41076 46686
rect 40796 46674 41076 46676
rect 40796 46622 41022 46674
rect 41074 46622 41076 46674
rect 40796 46620 41076 46622
rect 41020 46610 41076 46620
rect 41580 46676 41636 46686
rect 41580 46582 41636 46620
rect 41692 46452 41748 47852
rect 43036 47842 43092 47852
rect 43372 47684 43428 48188
rect 43484 48242 43764 48244
rect 43484 48190 43486 48242
rect 43538 48190 43764 48242
rect 43484 48188 43764 48190
rect 43820 48244 43876 48254
rect 43484 48178 43540 48188
rect 43820 48150 43876 48188
rect 44044 48132 44100 48860
rect 45164 48914 45220 48926
rect 45164 48862 45166 48914
rect 45218 48862 45220 48914
rect 44268 48802 44324 48814
rect 44268 48750 44270 48802
rect 44322 48750 44324 48802
rect 44268 48692 44324 48750
rect 44268 48626 44324 48636
rect 44156 48468 44212 48478
rect 44156 48466 45108 48468
rect 44156 48414 44158 48466
rect 44210 48414 45108 48466
rect 44156 48412 45108 48414
rect 44156 48402 44212 48412
rect 45052 48354 45108 48412
rect 45052 48302 45054 48354
rect 45106 48302 45108 48354
rect 45052 48290 45108 48302
rect 44492 48242 44548 48254
rect 44492 48190 44494 48242
rect 44546 48190 44548 48242
rect 43932 48076 44100 48132
rect 44268 48132 44324 48142
rect 43484 47684 43540 47694
rect 43372 47682 43540 47684
rect 43372 47630 43486 47682
rect 43538 47630 43540 47682
rect 43372 47628 43540 47630
rect 43484 47618 43540 47628
rect 43596 47348 43652 47358
rect 41580 46396 41748 46452
rect 42028 46674 42084 46686
rect 42028 46622 42030 46674
rect 42082 46622 42084 46674
rect 42028 46564 42084 46622
rect 42700 46564 42756 46574
rect 42028 46562 42756 46564
rect 42028 46510 42702 46562
rect 42754 46510 42756 46562
rect 42028 46508 42756 46510
rect 40572 46004 40628 46014
rect 40516 46002 40628 46004
rect 40516 45950 40574 46002
rect 40626 45950 40628 46002
rect 40516 45948 40628 45950
rect 40460 45910 40516 45948
rect 40572 45938 40628 45948
rect 37884 45780 37940 45790
rect 39900 45780 39956 45790
rect 37548 43426 37604 43484
rect 37548 43374 37550 43426
rect 37602 43374 37604 43426
rect 37548 43362 37604 43374
rect 37660 45778 37940 45780
rect 37660 45726 37886 45778
rect 37938 45726 37940 45778
rect 37660 45724 37940 45726
rect 37660 42868 37716 45724
rect 37884 45714 37940 45724
rect 39564 45778 39956 45780
rect 39564 45726 39902 45778
rect 39954 45726 39956 45778
rect 39564 45724 39956 45726
rect 37772 44436 37828 44446
rect 37772 44342 37828 44380
rect 39564 44436 39620 45724
rect 39900 45714 39956 45724
rect 40572 45332 40628 45342
rect 40124 45220 40180 45230
rect 40124 45126 40180 45164
rect 38220 43652 38276 43662
rect 38444 43652 38500 43662
rect 38220 43558 38276 43596
rect 38332 43596 38444 43652
rect 37548 42756 37604 42766
rect 37660 42756 37716 42812
rect 37548 42754 37716 42756
rect 37548 42702 37550 42754
rect 37602 42702 37716 42754
rect 37548 42700 37716 42702
rect 37996 43538 38052 43550
rect 37996 43486 37998 43538
rect 38050 43486 38052 43538
rect 37996 42756 38052 43486
rect 38108 43538 38164 43550
rect 38108 43486 38110 43538
rect 38162 43486 38164 43538
rect 38108 42980 38164 43486
rect 38108 42914 38164 42924
rect 38332 43538 38388 43596
rect 38444 43586 38500 43596
rect 39340 43652 39396 43662
rect 39340 43558 39396 43596
rect 39564 43650 39620 44380
rect 39900 44210 39956 44222
rect 39900 44158 39902 44210
rect 39954 44158 39956 44210
rect 39900 43762 39956 44158
rect 39900 43710 39902 43762
rect 39954 43710 39956 43762
rect 39900 43698 39956 43710
rect 40572 44212 40628 45276
rect 40908 45220 40964 45230
rect 40908 45106 40964 45164
rect 40908 45054 40910 45106
rect 40962 45054 40964 45106
rect 40908 45042 40964 45054
rect 39564 43598 39566 43650
rect 39618 43598 39620 43650
rect 39564 43586 39620 43598
rect 38332 43486 38334 43538
rect 38386 43486 38388 43538
rect 37996 42754 38164 42756
rect 37996 42702 37998 42754
rect 38050 42702 38164 42754
rect 37996 42700 38164 42702
rect 37548 42690 37604 42700
rect 37996 42690 38052 42700
rect 37660 42530 37716 42542
rect 37660 42478 37662 42530
rect 37714 42478 37716 42530
rect 37660 42420 37716 42478
rect 37548 41972 37604 41982
rect 37436 41970 37604 41972
rect 37436 41918 37550 41970
rect 37602 41918 37604 41970
rect 37436 41916 37604 41918
rect 37660 41972 37716 42364
rect 37772 42530 37828 42542
rect 37772 42478 37774 42530
rect 37826 42478 37828 42530
rect 37772 42196 37828 42478
rect 37884 42532 37940 42542
rect 37884 42438 37940 42476
rect 37772 42130 37828 42140
rect 38108 42196 38164 42700
rect 38332 42420 38388 43486
rect 38556 43540 38612 43550
rect 38892 43540 38948 43550
rect 38556 43446 38612 43484
rect 38780 43538 38948 43540
rect 38780 43486 38894 43538
rect 38946 43486 38948 43538
rect 38780 43484 38948 43486
rect 38668 42532 38724 42542
rect 38668 42438 38724 42476
rect 38332 42354 38388 42364
rect 38108 42194 38612 42196
rect 38108 42142 38110 42194
rect 38162 42142 38612 42194
rect 38108 42140 38612 42142
rect 38108 42130 38164 42140
rect 37772 41972 37828 41982
rect 37660 41970 37828 41972
rect 37660 41918 37774 41970
rect 37826 41918 37828 41970
rect 37660 41916 37828 41918
rect 37212 41878 37268 41916
rect 37548 41748 37604 41916
rect 37772 41906 37828 41916
rect 37996 41972 38052 41982
rect 38556 41972 38612 42140
rect 38780 41972 38836 43484
rect 38892 43474 38948 43484
rect 39116 43538 39172 43550
rect 39116 43486 39118 43538
rect 39170 43486 39172 43538
rect 39004 42980 39060 42990
rect 39004 42530 39060 42924
rect 39004 42478 39006 42530
rect 39058 42478 39060 42530
rect 39004 42196 39060 42478
rect 39116 42532 39172 43486
rect 39228 43426 39284 43438
rect 39228 43374 39230 43426
rect 39282 43374 39284 43426
rect 39228 43316 39284 43374
rect 40012 43426 40068 43438
rect 40012 43374 40014 43426
rect 40066 43374 40068 43426
rect 40012 43316 40068 43374
rect 39228 43260 40068 43316
rect 39788 42532 39844 42542
rect 39116 42530 39844 42532
rect 39116 42478 39790 42530
rect 39842 42478 39844 42530
rect 39116 42476 39844 42478
rect 39004 42130 39060 42140
rect 39564 42308 39620 42318
rect 38556 41916 38836 41972
rect 37884 41858 37940 41870
rect 37884 41806 37886 41858
rect 37938 41806 37940 41858
rect 37772 41748 37828 41758
rect 37548 41692 37772 41748
rect 37772 41682 37828 41692
rect 37884 41524 37940 41806
rect 37212 41468 37940 41524
rect 37212 41298 37268 41468
rect 37212 41246 37214 41298
rect 37266 41246 37268 41298
rect 37212 41234 37268 41246
rect 37324 41300 37380 41310
rect 37100 41076 37156 41086
rect 37100 40982 37156 41020
rect 37324 40404 37380 41244
rect 36988 40124 37268 40180
rect 36988 39956 37044 39966
rect 35756 39618 36484 39620
rect 35756 39566 35758 39618
rect 35810 39566 36484 39618
rect 35756 39564 36484 39566
rect 35756 39554 35812 39564
rect 36428 39508 36484 39564
rect 36428 39452 36820 39508
rect 35308 39330 35364 39340
rect 36316 39396 36372 39406
rect 35756 39060 35812 39070
rect 35756 38946 35812 39004
rect 35756 38894 35758 38946
rect 35810 38894 35812 38946
rect 35756 38882 35812 38894
rect 35756 38722 35812 38734
rect 35756 38670 35758 38722
rect 35810 38670 35812 38722
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35644 38052 35700 38062
rect 35308 37828 35364 37838
rect 35308 37826 35476 37828
rect 35308 37774 35310 37826
rect 35362 37774 35476 37826
rect 35308 37772 35476 37774
rect 35308 37762 35364 37772
rect 35420 37492 35476 37772
rect 35532 37492 35588 37502
rect 35420 37436 35532 37492
rect 35532 37426 35588 37436
rect 35308 37268 35364 37278
rect 35532 37268 35588 37278
rect 35308 37266 35588 37268
rect 35308 37214 35310 37266
rect 35362 37214 35534 37266
rect 35586 37214 35588 37266
rect 35308 37212 35588 37214
rect 35308 37202 35364 37212
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 36484 35252 36494
rect 35532 36484 35588 37212
rect 35644 37268 35700 37996
rect 35644 37202 35700 37212
rect 35756 36596 35812 38670
rect 36316 38668 36372 39340
rect 36652 39284 36708 39294
rect 36652 39060 36708 39228
rect 36652 38834 36708 39004
rect 36652 38782 36654 38834
rect 36706 38782 36708 38834
rect 36652 38770 36708 38782
rect 36316 38612 36708 38668
rect 36316 38052 36372 38062
rect 36316 37958 36372 37996
rect 35980 37828 36036 37838
rect 35756 36530 35812 36540
rect 35868 37826 36036 37828
rect 35868 37774 35982 37826
rect 36034 37774 36036 37826
rect 35868 37772 36036 37774
rect 35868 37044 35924 37772
rect 35980 37762 36036 37772
rect 35980 37604 36036 37614
rect 35980 37490 36036 37548
rect 35980 37438 35982 37490
rect 36034 37438 36036 37490
rect 35980 37426 36036 37438
rect 36092 37492 36148 37502
rect 36092 37490 36596 37492
rect 36092 37438 36094 37490
rect 36146 37438 36596 37490
rect 36092 37436 36596 37438
rect 36092 37426 36148 37436
rect 36540 37378 36596 37436
rect 36540 37326 36542 37378
rect 36594 37326 36596 37378
rect 36540 37314 36596 37326
rect 36204 37268 36260 37278
rect 36204 37174 36260 37212
rect 36428 37268 36484 37278
rect 35196 36482 35588 36484
rect 35196 36430 35198 36482
rect 35250 36430 35588 36482
rect 35196 36428 35588 36430
rect 35868 36482 35924 36988
rect 35868 36430 35870 36482
rect 35922 36430 35924 36482
rect 35196 36372 35252 36428
rect 35868 36418 35924 36430
rect 36316 37156 36372 37166
rect 36316 36596 36372 37100
rect 36316 36482 36372 36540
rect 36316 36430 36318 36482
rect 36370 36430 36372 36482
rect 35196 36306 35252 36316
rect 35644 36372 35700 36382
rect 35644 36278 35700 36316
rect 36316 36372 36372 36430
rect 36316 36306 36372 36316
rect 35756 36258 35812 36270
rect 35756 36206 35758 36258
rect 35810 36206 35812 36258
rect 35756 35812 35812 36206
rect 35868 35812 35924 35822
rect 35756 35810 35924 35812
rect 35756 35758 35870 35810
rect 35922 35758 35924 35810
rect 35756 35756 35924 35758
rect 35868 35746 35924 35756
rect 36204 35698 36260 35710
rect 36204 35646 36206 35698
rect 36258 35646 36260 35698
rect 36204 35476 36260 35646
rect 36428 35700 36484 37212
rect 36428 35606 36484 35644
rect 36204 35410 36260 35420
rect 36316 35586 36372 35598
rect 36316 35534 36318 35586
rect 36370 35534 36372 35586
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 36316 35028 36372 35534
rect 36316 34962 36372 34972
rect 34804 34860 34916 34916
rect 34748 34850 34804 34860
rect 34636 34262 34692 34300
rect 34748 34692 34804 34702
rect 34524 32834 34580 32844
rect 34636 33908 34692 33918
rect 34188 32788 34244 32798
rect 34188 32694 34244 32732
rect 34636 32674 34692 33852
rect 34636 32622 34638 32674
rect 34690 32622 34692 32674
rect 34076 32562 34468 32564
rect 34076 32510 34078 32562
rect 34130 32510 34468 32562
rect 34076 32508 34468 32510
rect 34076 32498 34132 32508
rect 34412 31892 34468 32508
rect 34412 31798 34468 31836
rect 34636 31780 34692 32622
rect 34636 31714 34692 31724
rect 34748 31444 34804 34636
rect 34860 34132 34916 34860
rect 34860 34066 34916 34076
rect 34972 34860 35140 34916
rect 34636 31388 34804 31444
rect 33852 31108 33908 31118
rect 33852 31014 33908 31052
rect 33516 30994 33572 31006
rect 33516 30942 33518 30994
rect 33570 30942 33572 30994
rect 33516 30324 33572 30942
rect 33740 30996 33796 31006
rect 33740 30902 33796 30940
rect 34300 30994 34356 31006
rect 34300 30942 34302 30994
rect 34354 30942 34356 30994
rect 33516 30258 33572 30268
rect 33852 29316 33908 29326
rect 34300 29316 34356 30942
rect 34524 30996 34580 31006
rect 34524 30902 34580 30940
rect 33852 29314 34356 29316
rect 33852 29262 33854 29314
rect 33906 29262 34356 29314
rect 33852 29260 34356 29262
rect 33852 28532 33908 29260
rect 33852 28466 33908 28476
rect 34300 28532 34356 28542
rect 34300 28082 34356 28476
rect 34300 28030 34302 28082
rect 34354 28030 34356 28082
rect 34300 28018 34356 28030
rect 34412 28420 34468 28430
rect 33740 27972 33796 27982
rect 34076 27972 34132 27982
rect 33796 27970 34132 27972
rect 33796 27918 34078 27970
rect 34130 27918 34132 27970
rect 33796 27916 34132 27918
rect 33740 27878 33796 27916
rect 34076 27906 34132 27916
rect 34412 27970 34468 28364
rect 34412 27918 34414 27970
rect 34466 27918 34468 27970
rect 34412 27906 34468 27918
rect 33516 27860 33572 27870
rect 33516 27766 33572 27804
rect 33628 27746 33684 27758
rect 33628 27694 33630 27746
rect 33682 27694 33684 27746
rect 33628 27636 33684 27694
rect 33516 27580 33684 27636
rect 33740 27636 33796 27646
rect 33516 26908 33572 27580
rect 33740 27074 33796 27580
rect 34636 27636 34692 31388
rect 34860 31332 34916 31342
rect 34748 31276 34860 31332
rect 34748 31218 34804 31276
rect 34860 31266 34916 31276
rect 34748 31166 34750 31218
rect 34802 31166 34804 31218
rect 34748 31154 34804 31166
rect 34860 31108 34916 31118
rect 34860 31014 34916 31052
rect 34860 30882 34916 30894
rect 34860 30830 34862 30882
rect 34914 30830 34916 30882
rect 34860 30212 34916 30830
rect 34860 30146 34916 30156
rect 34636 27570 34692 27580
rect 34972 30098 35028 34860
rect 35084 34692 35140 34702
rect 35084 34598 35140 34636
rect 35084 34356 35140 34366
rect 36092 34356 36148 34366
rect 35140 34300 35252 34356
rect 35084 34290 35140 34300
rect 35196 34244 35252 34300
rect 36092 34262 36148 34300
rect 35196 34242 35812 34244
rect 35196 34190 35198 34242
rect 35250 34190 35812 34242
rect 35196 34188 35812 34190
rect 35196 34178 35252 34188
rect 35084 34132 35140 34142
rect 35084 34038 35140 34076
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35532 33572 35588 33582
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 32004 35252 32014
rect 35084 31892 35140 31902
rect 35084 31778 35140 31836
rect 35084 31726 35086 31778
rect 35138 31726 35140 31778
rect 35084 31714 35140 31726
rect 35196 30772 35252 31948
rect 35420 31890 35476 31902
rect 35420 31838 35422 31890
rect 35474 31838 35476 31890
rect 35308 31778 35364 31790
rect 35308 31726 35310 31778
rect 35362 31726 35364 31778
rect 35308 31556 35364 31726
rect 35420 31780 35476 31838
rect 35420 31714 35476 31724
rect 35532 31556 35588 33516
rect 35756 33570 35812 34188
rect 35756 33518 35758 33570
rect 35810 33518 35812 33570
rect 35756 33506 35812 33518
rect 35868 34132 35924 34142
rect 35308 31500 35588 31556
rect 35532 31220 35588 31230
rect 35532 31126 35588 31164
rect 34972 30046 34974 30098
rect 35026 30046 35028 30098
rect 34748 27188 34804 27198
rect 34748 27094 34804 27132
rect 33740 27022 33742 27074
rect 33794 27022 33796 27074
rect 33740 27010 33796 27022
rect 34860 26964 34916 27002
rect 33516 26852 33908 26908
rect 34860 26898 34916 26908
rect 33852 26402 33908 26852
rect 33852 26350 33854 26402
rect 33906 26350 33908 26402
rect 33852 26338 33908 26350
rect 33740 23156 33796 23166
rect 33740 22372 33796 23100
rect 33740 22306 33796 22316
rect 33404 22194 33460 22204
rect 33180 22146 33348 22148
rect 33180 22094 33182 22146
rect 33234 22094 33348 22146
rect 33180 22092 33348 22094
rect 33180 22082 33236 22092
rect 33068 21588 33124 21598
rect 32956 21586 33124 21588
rect 32956 21534 33070 21586
rect 33122 21534 33124 21586
rect 32956 21532 33124 21534
rect 33068 20132 33124 21532
rect 33068 20066 33124 20076
rect 32956 19908 33012 19918
rect 33180 19908 33236 19918
rect 32844 19852 32956 19908
rect 33012 19906 33236 19908
rect 33012 19854 33182 19906
rect 33234 19854 33236 19906
rect 33012 19852 33236 19854
rect 32956 19348 33012 19852
rect 33180 19842 33236 19852
rect 33292 19684 33348 22092
rect 33852 21476 33908 21486
rect 34636 21476 34692 21486
rect 33852 21474 34580 21476
rect 33852 21422 33854 21474
rect 33906 21422 34580 21474
rect 33852 21420 34580 21422
rect 33852 21410 33908 21420
rect 34524 21026 34580 21420
rect 34524 20974 34526 21026
rect 34578 20974 34580 21026
rect 34524 20962 34580 20974
rect 34636 20914 34692 21420
rect 34636 20862 34638 20914
rect 34690 20862 34692 20914
rect 34636 20850 34692 20862
rect 32956 19282 33012 19292
rect 33068 19628 33348 19684
rect 34300 20132 34356 20142
rect 32172 19122 32340 19124
rect 32172 19070 32174 19122
rect 32226 19070 32340 19122
rect 32172 19068 32340 19070
rect 32172 19058 32228 19068
rect 31948 18844 32228 18900
rect 32172 18564 32228 18844
rect 32172 18470 32228 18508
rect 32060 18450 32116 18462
rect 32060 18398 32062 18450
rect 32114 18398 32116 18450
rect 32060 18340 32116 18398
rect 32060 18274 32116 18284
rect 32284 18450 32340 19068
rect 32284 18398 32286 18450
rect 32338 18398 32340 18450
rect 31276 17724 31780 17780
rect 32172 17780 32228 17790
rect 32284 17780 32340 18398
rect 32228 17724 32340 17780
rect 32620 19010 32676 19068
rect 32620 18958 32622 19010
rect 32674 18958 32676 19010
rect 31052 16882 31220 16884
rect 31052 16830 31054 16882
rect 31106 16830 31220 16882
rect 31052 16828 31220 16830
rect 31052 16818 31108 16828
rect 29260 16716 29596 16772
rect 29260 15538 29316 16716
rect 29596 16706 29652 16716
rect 30828 16772 30884 16782
rect 30828 16322 30884 16716
rect 30828 16270 30830 16322
rect 30882 16270 30884 16322
rect 30716 15988 30772 15998
rect 29260 15486 29262 15538
rect 29314 15486 29316 15538
rect 29260 15474 29316 15486
rect 30380 15986 30772 15988
rect 30380 15934 30718 15986
rect 30770 15934 30772 15986
rect 30380 15932 30772 15934
rect 28924 15428 28980 15438
rect 28924 15334 28980 15372
rect 29036 15426 29092 15438
rect 29036 15374 29038 15426
rect 29090 15374 29092 15426
rect 28700 15026 28756 15036
rect 29036 14868 29092 15374
rect 30380 15426 30436 15932
rect 30716 15922 30772 15932
rect 30828 15652 30884 16270
rect 30828 15586 30884 15596
rect 31052 16098 31108 16110
rect 31052 16046 31054 16098
rect 31106 16046 31108 16098
rect 30380 15374 30382 15426
rect 30434 15374 30436 15426
rect 30380 15362 30436 15374
rect 28588 14812 29092 14868
rect 29596 15314 29652 15326
rect 29596 15262 29598 15314
rect 29650 15262 29652 15314
rect 29596 15092 29652 15262
rect 28476 13654 28532 13692
rect 28364 12910 28366 12962
rect 28418 12910 28420 12962
rect 28364 12898 28420 12910
rect 28588 12964 28644 12974
rect 28588 12870 28644 12908
rect 28140 10518 28196 10556
rect 28812 9828 28868 14812
rect 29596 13858 29652 15036
rect 30940 14756 30996 14766
rect 31052 14756 31108 16046
rect 31164 15876 31220 16828
rect 31276 16882 31332 17724
rect 32172 17686 32228 17724
rect 32620 16996 32676 18958
rect 32732 18340 32788 18350
rect 32732 17778 32788 18284
rect 32732 17726 32734 17778
rect 32786 17726 32788 17778
rect 32732 17714 32788 17726
rect 32620 16930 32676 16940
rect 31276 16830 31278 16882
rect 31330 16830 31332 16882
rect 31276 16818 31332 16830
rect 31724 16212 31780 16222
rect 31276 16210 31780 16212
rect 31276 16158 31726 16210
rect 31778 16158 31780 16210
rect 31276 16156 31780 16158
rect 31276 16098 31332 16156
rect 31724 16146 31780 16156
rect 31276 16046 31278 16098
rect 31330 16046 31332 16098
rect 31276 16034 31332 16046
rect 31948 16098 32004 16110
rect 31948 16046 31950 16098
rect 32002 16046 32004 16098
rect 31612 15986 31668 15998
rect 31612 15934 31614 15986
rect 31666 15934 31668 15986
rect 31612 15876 31668 15934
rect 31164 15820 31668 15876
rect 29596 13806 29598 13858
rect 29650 13806 29652 13858
rect 29596 13524 29652 13806
rect 29596 13458 29652 13468
rect 30716 14754 31108 14756
rect 30716 14702 30942 14754
rect 30994 14702 31108 14754
rect 30716 14700 31108 14702
rect 31164 15652 31220 15662
rect 29820 13076 29876 13086
rect 29820 12982 29876 13020
rect 30156 12964 30212 12974
rect 30156 12870 30212 12908
rect 30716 12964 30772 14700
rect 30940 14690 30996 14700
rect 30828 13188 30884 13198
rect 30828 13094 30884 13132
rect 31164 12964 31220 15596
rect 31276 14754 31332 15820
rect 31276 14702 31278 14754
rect 31330 14702 31332 14754
rect 31276 14690 31332 14702
rect 31388 15316 31444 15326
rect 31276 12964 31332 12974
rect 31164 12962 31332 12964
rect 31164 12910 31278 12962
rect 31330 12910 31332 12962
rect 31164 12908 31332 12910
rect 30716 12870 30772 12908
rect 31276 12898 31332 12908
rect 29708 12852 29764 12862
rect 29708 12066 29764 12796
rect 30380 12852 30436 12862
rect 30380 12758 30436 12796
rect 30828 12852 30884 12862
rect 30828 12758 30884 12796
rect 29708 12014 29710 12066
rect 29762 12014 29764 12066
rect 29708 12002 29764 12014
rect 31164 11396 31220 11406
rect 31164 11302 31220 11340
rect 29372 10612 29428 10622
rect 29372 10518 29428 10556
rect 30156 10498 30212 10510
rect 30156 10446 30158 10498
rect 30210 10446 30212 10498
rect 30156 9938 30212 10446
rect 30156 9886 30158 9938
rect 30210 9886 30212 9938
rect 30156 9874 30212 9886
rect 30604 10500 30660 10510
rect 28812 9772 29316 9828
rect 27916 9550 27918 9602
rect 27970 9550 27972 9602
rect 27916 9492 27972 9550
rect 28140 9714 28196 9726
rect 28140 9662 28142 9714
rect 28194 9662 28196 9714
rect 28140 9604 28196 9662
rect 28140 9538 28196 9548
rect 28588 9602 28644 9614
rect 28588 9550 28590 9602
rect 28642 9550 28644 9602
rect 27916 9426 27972 9436
rect 28588 9492 28644 9550
rect 27132 7534 27134 7586
rect 27186 7534 27188 7586
rect 27132 7522 27188 7534
rect 26908 7474 27076 7476
rect 26908 7422 26910 7474
rect 26962 7422 27076 7474
rect 26908 7420 27076 7422
rect 26460 7410 26516 7420
rect 26908 7410 26964 7420
rect 26796 7252 26852 7262
rect 26348 7250 26852 7252
rect 26348 7198 26798 7250
rect 26850 7198 26852 7250
rect 26348 7196 26852 7198
rect 26236 7186 26292 7196
rect 26796 7186 26852 7196
rect 26684 7028 26740 7038
rect 26460 6916 26516 6926
rect 26460 6692 26516 6860
rect 25900 6636 26516 6692
rect 26012 6130 26068 6142
rect 26012 6078 26014 6130
rect 26066 6078 26068 6130
rect 25788 6020 25844 6030
rect 25788 5906 25844 5964
rect 25788 5854 25790 5906
rect 25842 5854 25844 5906
rect 25788 5842 25844 5854
rect 25788 5684 25844 5694
rect 25788 5590 25844 5628
rect 26012 4450 26068 6078
rect 26236 6020 26292 6030
rect 26236 5234 26292 5964
rect 26460 6018 26516 6636
rect 26684 6130 26740 6972
rect 27020 6802 27076 7420
rect 27020 6750 27022 6802
rect 27074 6750 27076 6802
rect 27020 6738 27076 6750
rect 27132 7364 27188 7374
rect 26684 6078 26686 6130
rect 26738 6078 26740 6130
rect 26684 6066 26740 6078
rect 26460 5966 26462 6018
rect 26514 5966 26516 6018
rect 26460 5954 26516 5966
rect 27132 5908 27188 7308
rect 27356 7250 27412 7262
rect 27356 7198 27358 7250
rect 27410 7198 27412 7250
rect 27356 7028 27412 7198
rect 27356 6962 27412 6972
rect 27580 7250 27636 7262
rect 27580 7198 27582 7250
rect 27634 7198 27636 7250
rect 27580 6916 27636 7198
rect 27580 6850 27636 6860
rect 27132 5906 27524 5908
rect 27132 5854 27134 5906
rect 27186 5854 27524 5906
rect 27132 5852 27524 5854
rect 27132 5842 27188 5852
rect 26236 5182 26238 5234
rect 26290 5182 26292 5234
rect 26236 5170 26292 5182
rect 26572 5794 26628 5806
rect 26572 5742 26574 5794
rect 26626 5742 26628 5794
rect 26572 5124 26628 5742
rect 26684 5684 26740 5694
rect 26684 5234 26740 5628
rect 26684 5182 26686 5234
rect 26738 5182 26740 5234
rect 26684 5170 26740 5182
rect 27468 5234 27524 5852
rect 27468 5182 27470 5234
rect 27522 5182 27524 5234
rect 27468 5170 27524 5182
rect 26572 5030 26628 5068
rect 26908 5122 26964 5134
rect 26908 5070 26910 5122
rect 26962 5070 26964 5122
rect 26012 4398 26014 4450
rect 26066 4398 26068 4450
rect 26012 4386 26068 4398
rect 26908 4228 26964 5070
rect 26908 4162 26964 4172
rect 28140 4228 28196 4238
rect 25676 3714 25732 3724
rect 26124 3668 26180 3678
rect 26124 3574 26180 3612
rect 25228 3502 25230 3554
rect 25282 3502 25284 3554
rect 25228 3490 25284 3502
rect 28140 3556 28196 4172
rect 28588 3668 28644 9436
rect 28812 9266 28868 9772
rect 28812 9214 28814 9266
rect 28866 9214 28868 9266
rect 28812 8372 28868 9214
rect 29148 9604 29204 9614
rect 29148 9154 29204 9548
rect 29260 9266 29316 9772
rect 29820 9826 29876 9838
rect 29820 9774 29822 9826
rect 29874 9774 29876 9826
rect 29820 9716 29876 9774
rect 30044 9828 30100 9838
rect 30044 9734 30100 9772
rect 30380 9828 30436 9838
rect 30604 9828 30660 10444
rect 30380 9826 30660 9828
rect 30380 9774 30382 9826
rect 30434 9774 30606 9826
rect 30658 9774 30660 9826
rect 30380 9772 30660 9774
rect 30380 9762 30436 9772
rect 29820 9650 29876 9660
rect 29260 9214 29262 9266
rect 29314 9214 29316 9266
rect 29260 9202 29316 9214
rect 30380 9268 30436 9278
rect 30380 9174 30436 9212
rect 29148 9102 29150 9154
rect 29202 9102 29204 9154
rect 29148 9090 29204 9102
rect 28812 8306 28868 8316
rect 29484 9042 29540 9054
rect 29484 8990 29486 9042
rect 29538 8990 29540 9042
rect 29484 8036 29540 8990
rect 29484 7474 29540 7980
rect 30268 8036 30324 8046
rect 30268 7942 30324 7980
rect 30044 7924 30100 7934
rect 29820 7700 29876 7710
rect 29820 7698 29988 7700
rect 29820 7646 29822 7698
rect 29874 7646 29988 7698
rect 29820 7644 29988 7646
rect 29820 7634 29876 7644
rect 29484 7422 29486 7474
rect 29538 7422 29540 7474
rect 29484 7410 29540 7422
rect 29708 7364 29764 7374
rect 29708 7270 29764 7308
rect 29820 7252 29876 7262
rect 29820 7158 29876 7196
rect 29932 6802 29988 7644
rect 29932 6750 29934 6802
rect 29986 6750 29988 6802
rect 29932 6738 29988 6750
rect 29148 6690 29204 6702
rect 29148 6638 29150 6690
rect 29202 6638 29204 6690
rect 29148 6020 29204 6638
rect 29148 6018 29316 6020
rect 29148 5966 29150 6018
rect 29202 5966 29316 6018
rect 29148 5964 29316 5966
rect 29148 5954 29204 5964
rect 29260 5012 29316 5964
rect 30044 5346 30100 7868
rect 30268 7588 30324 7598
rect 30492 7588 30548 9772
rect 30604 9762 30660 9772
rect 30828 9828 30884 9838
rect 30716 9716 30772 9726
rect 30716 9622 30772 9660
rect 30828 9714 30884 9772
rect 31388 9826 31444 15260
rect 31500 15204 31556 15214
rect 31500 14642 31556 15148
rect 31948 15204 32004 16046
rect 31948 15138 32004 15148
rect 32508 15204 32564 15242
rect 32508 15138 32564 15148
rect 31500 14590 31502 14642
rect 31554 14590 31556 14642
rect 31500 14578 31556 14590
rect 31836 13188 31892 13198
rect 31612 12964 31668 12974
rect 31612 12870 31668 12908
rect 31836 12962 31892 13132
rect 33068 13188 33124 19628
rect 33628 18564 33684 18574
rect 33628 18470 33684 18508
rect 33516 18452 33572 18462
rect 33180 18226 33236 18238
rect 33180 18174 33182 18226
rect 33234 18174 33236 18226
rect 33180 17780 33236 18174
rect 33180 17444 33236 17724
rect 33516 17668 33572 18396
rect 33852 18450 33908 18462
rect 33852 18398 33854 18450
rect 33906 18398 33908 18450
rect 33740 18338 33796 18350
rect 33740 18286 33742 18338
rect 33794 18286 33796 18338
rect 33740 18004 33796 18286
rect 33852 18228 33908 18398
rect 34300 18450 34356 20076
rect 34748 19124 34804 19134
rect 34748 19030 34804 19068
rect 34636 19012 34692 19022
rect 34300 18398 34302 18450
rect 34354 18398 34356 18450
rect 34300 18386 34356 18398
rect 34524 19010 34692 19012
rect 34524 18958 34638 19010
rect 34690 18958 34692 19010
rect 34524 18956 34692 18958
rect 34524 18452 34580 18956
rect 34636 18946 34692 18956
rect 34972 18900 35028 30046
rect 35084 30716 35252 30772
rect 35084 28532 35140 30716
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35084 28466 35140 28476
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35868 26908 35924 34076
rect 35980 33572 36036 33582
rect 35980 33234 36036 33516
rect 36092 33458 36148 33470
rect 36092 33406 36094 33458
rect 36146 33406 36148 33458
rect 36092 33348 36148 33406
rect 36540 33460 36596 33470
rect 36148 33292 36372 33348
rect 36092 33282 36148 33292
rect 35980 33182 35982 33234
rect 36034 33182 36036 33234
rect 35980 33170 36036 33182
rect 35980 31108 36036 31118
rect 35980 31014 36036 31052
rect 36316 30994 36372 33292
rect 36540 30996 36596 33404
rect 36652 31220 36708 38612
rect 36764 34132 36820 39452
rect 36988 39058 37044 39900
rect 36988 39006 36990 39058
rect 37042 39006 37044 39058
rect 36988 38836 37044 39006
rect 37212 39060 37268 40124
rect 37212 38966 37268 39004
rect 36988 38770 37044 38780
rect 37324 38668 37380 40348
rect 37996 39732 38052 41916
rect 38556 41748 38612 41758
rect 38556 40290 38612 41692
rect 38780 40628 38836 41916
rect 38892 40628 38948 40638
rect 38780 40626 38948 40628
rect 38780 40574 38894 40626
rect 38946 40574 38948 40626
rect 38780 40572 38948 40574
rect 38892 40562 38948 40572
rect 39564 40626 39620 42252
rect 39564 40574 39566 40626
rect 39618 40574 39620 40626
rect 39564 40562 39620 40574
rect 38556 40238 38558 40290
rect 38610 40238 38612 40290
rect 38556 40226 38612 40238
rect 39116 40402 39172 40414
rect 39116 40350 39118 40402
rect 39170 40350 39172 40402
rect 39116 40180 39172 40350
rect 38556 39956 38612 39966
rect 38108 39732 38164 39742
rect 37996 39730 38276 39732
rect 37996 39678 38110 39730
rect 38162 39678 38276 39730
rect 37996 39676 38276 39678
rect 38108 39666 38164 39676
rect 37772 39396 37828 39406
rect 36876 38610 36932 38622
rect 36876 38558 36878 38610
rect 36930 38558 36932 38610
rect 36876 38052 36932 38558
rect 36876 37986 36932 37996
rect 37212 38612 37380 38668
rect 37548 39394 37828 39396
rect 37548 39342 37774 39394
rect 37826 39342 37828 39394
rect 37548 39340 37828 39342
rect 37548 38834 37604 39340
rect 37772 39330 37828 39340
rect 37548 38782 37550 38834
rect 37602 38782 37604 38834
rect 37212 38050 37268 38612
rect 37548 38276 37604 38782
rect 37884 39060 37940 39070
rect 37884 38836 37940 39004
rect 37884 38770 37940 38780
rect 38220 39058 38276 39676
rect 38556 39730 38612 39900
rect 38556 39678 38558 39730
rect 38610 39678 38612 39730
rect 38556 39666 38612 39678
rect 38220 39006 38222 39058
rect 38274 39006 38276 39058
rect 38220 38668 38276 39006
rect 37548 38210 37604 38220
rect 37996 38612 38276 38668
rect 38668 39172 38724 39182
rect 38668 38722 38724 39116
rect 38668 38670 38670 38722
rect 38722 38670 38724 38722
rect 38668 38658 38724 38670
rect 37212 37998 37214 38050
rect 37266 37998 37268 38050
rect 37212 37986 37268 37998
rect 37884 37940 37940 37950
rect 37324 37938 37940 37940
rect 37324 37886 37886 37938
rect 37938 37886 37940 37938
rect 37324 37884 37940 37886
rect 37324 37604 37380 37884
rect 37884 37874 37940 37884
rect 36988 37548 37380 37604
rect 37548 37604 37604 37614
rect 36988 37490 37044 37548
rect 36988 37438 36990 37490
rect 37042 37438 37044 37490
rect 36988 37426 37044 37438
rect 37548 37490 37604 37548
rect 37548 37438 37550 37490
rect 37602 37438 37604 37490
rect 37548 37426 37604 37438
rect 36876 37266 36932 37278
rect 36876 37214 36878 37266
rect 36930 37214 36932 37266
rect 36876 37156 36932 37214
rect 37100 37268 37156 37278
rect 37996 37268 38052 38612
rect 38108 37828 38164 37838
rect 38108 37604 38164 37772
rect 38108 37538 38164 37548
rect 37100 37174 37156 37212
rect 37436 37212 38052 37268
rect 36876 37090 36932 37100
rect 37436 36260 37492 37212
rect 38220 37156 38276 37166
rect 38332 37156 38388 37166
rect 38276 37154 38388 37156
rect 38276 37102 38334 37154
rect 38386 37102 38388 37154
rect 38276 37100 38388 37102
rect 37100 34916 37156 34926
rect 37100 34914 37380 34916
rect 37100 34862 37102 34914
rect 37154 34862 37380 34914
rect 37100 34860 37380 34862
rect 37100 34850 37156 34860
rect 36764 34066 36820 34076
rect 36988 33908 37044 33918
rect 36988 31890 37044 33852
rect 36988 31838 36990 31890
rect 37042 31838 37044 31890
rect 36988 31826 37044 31838
rect 37100 33572 37156 33582
rect 36652 31154 36708 31164
rect 36316 30942 36318 30994
rect 36370 30942 36372 30994
rect 36316 30930 36372 30942
rect 36428 30994 36596 30996
rect 36428 30942 36542 30994
rect 36594 30942 36596 30994
rect 36428 30940 36596 30942
rect 36316 30212 36372 30222
rect 36316 30118 36372 30156
rect 36204 29988 36260 29998
rect 35980 29986 36260 29988
rect 35980 29934 36206 29986
rect 36258 29934 36260 29986
rect 35980 29932 36260 29934
rect 35980 29538 36036 29932
rect 36204 29922 36260 29932
rect 35980 29486 35982 29538
rect 36034 29486 36036 29538
rect 35980 29474 36036 29486
rect 36428 27972 36484 30940
rect 36540 30930 36596 30940
rect 36652 30996 36708 31006
rect 36652 29426 36708 30940
rect 36988 30882 37044 30894
rect 36988 30830 36990 30882
rect 37042 30830 37044 30882
rect 36988 29986 37044 30830
rect 36988 29934 36990 29986
rect 37042 29934 37044 29986
rect 36988 29652 37044 29934
rect 36988 29586 37044 29596
rect 36652 29374 36654 29426
rect 36706 29374 36708 29426
rect 36652 29362 36708 29374
rect 36428 27858 36484 27916
rect 36652 28532 36708 28542
rect 36428 27806 36430 27858
rect 36482 27806 36484 27858
rect 36428 27794 36484 27806
rect 36540 27860 36596 27870
rect 36540 27076 36596 27804
rect 36652 27858 36708 28476
rect 37100 28420 37156 33516
rect 37212 33348 37268 33358
rect 37212 32002 37268 33292
rect 37212 31950 37214 32002
rect 37266 31950 37268 32002
rect 37212 31938 37268 31950
rect 37324 31892 37380 34860
rect 37324 30996 37380 31836
rect 37436 31332 37492 36204
rect 37996 36370 38052 36382
rect 37996 36318 37998 36370
rect 38050 36318 38052 36370
rect 37884 35474 37940 35486
rect 37884 35422 37886 35474
rect 37938 35422 37940 35474
rect 37660 35140 37716 35150
rect 37660 33908 37716 35084
rect 37772 35028 37828 35038
rect 37772 34934 37828 34972
rect 37660 33572 37716 33852
rect 37772 33572 37828 33582
rect 37660 33570 37828 33572
rect 37660 33518 37774 33570
rect 37826 33518 37828 33570
rect 37660 33516 37828 33518
rect 37772 33506 37828 33516
rect 37884 33572 37940 35422
rect 37996 35476 38052 36318
rect 37996 35410 38052 35420
rect 38108 36258 38164 36270
rect 38108 36206 38110 36258
rect 38162 36206 38164 36258
rect 37884 33506 37940 33516
rect 38108 33460 38164 36206
rect 38220 35698 38276 37100
rect 38332 37090 38388 37100
rect 38668 37154 38724 37166
rect 38668 37102 38670 37154
rect 38722 37102 38724 37154
rect 38668 36932 38724 37102
rect 38444 36876 38668 36932
rect 38332 36484 38388 36494
rect 38444 36484 38500 36876
rect 38668 36866 38724 36876
rect 38332 36482 38500 36484
rect 38332 36430 38334 36482
rect 38386 36430 38500 36482
rect 38332 36428 38500 36430
rect 38332 36418 38388 36428
rect 38444 35812 38500 36428
rect 38444 35746 38500 35756
rect 38220 35646 38222 35698
rect 38274 35646 38276 35698
rect 38220 34242 38276 35646
rect 38556 35700 38612 35710
rect 39004 35700 39060 35710
rect 38556 35698 39004 35700
rect 38556 35646 38558 35698
rect 38610 35646 39004 35698
rect 38556 35644 39004 35646
rect 38556 35634 38612 35644
rect 39004 35606 39060 35644
rect 38220 34190 38222 34242
rect 38274 34190 38276 34242
rect 38220 34178 38276 34190
rect 38892 35476 38948 35486
rect 38892 34130 38948 35420
rect 38892 34078 38894 34130
rect 38946 34078 38948 34130
rect 38892 34066 38948 34078
rect 38444 33572 38500 33582
rect 38668 33572 38724 33582
rect 38500 33570 38724 33572
rect 38500 33518 38670 33570
rect 38722 33518 38724 33570
rect 38500 33516 38724 33518
rect 38444 33506 38500 33516
rect 38668 33506 38724 33516
rect 39004 33572 39060 33582
rect 39116 33572 39172 40124
rect 39228 38836 39284 38846
rect 39228 38742 39284 38780
rect 39788 37828 39844 42476
rect 40348 40852 40404 40862
rect 40348 40626 40404 40796
rect 40348 40574 40350 40626
rect 40402 40574 40404 40626
rect 40348 40562 40404 40574
rect 39900 40402 39956 40414
rect 39900 40350 39902 40402
rect 39954 40350 39956 40402
rect 39900 40292 39956 40350
rect 39900 40226 39956 40236
rect 40572 39396 40628 44156
rect 40684 44322 40740 44334
rect 40684 44270 40686 44322
rect 40738 44270 40740 44322
rect 40684 43708 40740 44270
rect 40684 43652 40964 43708
rect 40908 41970 40964 43652
rect 40908 41918 40910 41970
rect 40962 41918 40964 41970
rect 40908 41300 40964 41918
rect 40908 41206 40964 41244
rect 40908 40852 40964 40862
rect 40348 39340 40628 39396
rect 40796 40796 40908 40852
rect 40964 40796 41076 40852
rect 40236 38836 40292 38846
rect 39788 37762 39844 37772
rect 40012 38162 40068 38174
rect 40012 38110 40014 38162
rect 40066 38110 40068 38162
rect 40012 36932 40068 38110
rect 40012 36866 40068 36876
rect 39228 36258 39284 36270
rect 39228 36206 39230 36258
rect 39282 36206 39284 36258
rect 39228 36036 39284 36206
rect 39228 35980 39844 36036
rect 39452 35812 39508 35822
rect 39452 35700 39508 35756
rect 39340 35698 39508 35700
rect 39340 35646 39454 35698
rect 39506 35646 39508 35698
rect 39340 35644 39508 35646
rect 39340 34354 39396 35644
rect 39452 35634 39508 35644
rect 39676 35700 39732 35710
rect 39676 35028 39732 35644
rect 39788 35700 39844 35980
rect 40236 35922 40292 38780
rect 40236 35870 40238 35922
rect 40290 35870 40292 35922
rect 40236 35858 40292 35870
rect 39788 35698 40068 35700
rect 39788 35646 39790 35698
rect 39842 35646 40068 35698
rect 39788 35644 40068 35646
rect 39788 35634 39844 35644
rect 39900 35028 39956 35038
rect 39676 35026 39956 35028
rect 39676 34974 39902 35026
rect 39954 34974 39956 35026
rect 39676 34972 39956 34974
rect 39340 34302 39342 34354
rect 39394 34302 39396 34354
rect 39340 34290 39396 34302
rect 39564 34244 39620 34254
rect 39900 34244 39956 34972
rect 39564 34242 39956 34244
rect 39564 34190 39566 34242
rect 39618 34190 39956 34242
rect 39564 34188 39956 34190
rect 39564 34178 39620 34188
rect 39228 33908 39284 33918
rect 39228 33814 39284 33852
rect 39004 33570 39172 33572
rect 39004 33518 39006 33570
rect 39058 33518 39172 33570
rect 39004 33516 39172 33518
rect 39004 33506 39060 33516
rect 38108 33394 38164 33404
rect 37548 33346 37604 33358
rect 37548 33294 37550 33346
rect 37602 33294 37604 33346
rect 37548 32004 37604 33294
rect 38444 33348 38500 33358
rect 38444 33254 38500 33292
rect 38108 33124 38164 33134
rect 38108 33030 38164 33068
rect 37548 31938 37604 31948
rect 38556 32788 38612 32798
rect 37548 31556 37604 31566
rect 37548 31554 37716 31556
rect 37548 31502 37550 31554
rect 37602 31502 37716 31554
rect 37548 31500 37716 31502
rect 37548 31490 37604 31500
rect 37436 31276 37604 31332
rect 37436 30996 37492 31006
rect 37380 30994 37492 30996
rect 37380 30942 37438 30994
rect 37490 30942 37492 30994
rect 37380 30940 37492 30942
rect 37324 30902 37380 30940
rect 37436 30930 37492 30940
rect 37548 30772 37604 31276
rect 37100 28354 37156 28364
rect 37212 30716 37604 30772
rect 36652 27806 36654 27858
rect 36706 27806 36708 27858
rect 36652 27794 36708 27806
rect 35868 26852 36372 26908
rect 35980 26740 36036 26750
rect 35980 26178 36036 26684
rect 35980 26126 35982 26178
rect 36034 26126 36036 26178
rect 35980 26114 36036 26126
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35980 24836 36036 24846
rect 35532 24722 35588 24734
rect 35980 24724 36036 24780
rect 35532 24670 35534 24722
rect 35586 24670 35588 24722
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35532 24164 35588 24670
rect 35308 23828 35364 23838
rect 35308 23734 35364 23772
rect 35308 23380 35364 23390
rect 35308 23266 35364 23324
rect 35308 23214 35310 23266
rect 35362 23214 35364 23266
rect 35308 23202 35364 23214
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35532 22482 35588 24108
rect 35532 22430 35534 22482
rect 35586 22430 35588 22482
rect 35532 22418 35588 22430
rect 35868 24722 36036 24724
rect 35868 24670 35982 24722
rect 36034 24670 36036 24722
rect 35868 24668 36036 24670
rect 35756 22372 35812 22382
rect 35868 22372 35924 24668
rect 35980 24658 36036 24668
rect 36204 24722 36260 24734
rect 36204 24670 36206 24722
rect 36258 24670 36260 24722
rect 36092 24610 36148 24622
rect 36092 24558 36094 24610
rect 36146 24558 36148 24610
rect 35980 23938 36036 23950
rect 35980 23886 35982 23938
rect 36034 23886 36036 23938
rect 35980 23380 36036 23886
rect 36092 23940 36148 24558
rect 36092 23874 36148 23884
rect 36204 24612 36260 24670
rect 35980 23314 36036 23324
rect 35980 22596 36036 22606
rect 36204 22596 36260 24556
rect 35980 22594 36260 22596
rect 35980 22542 35982 22594
rect 36034 22542 36260 22594
rect 35980 22540 36260 22542
rect 35980 22530 36036 22540
rect 35756 22370 35924 22372
rect 35756 22318 35758 22370
rect 35810 22318 35924 22370
rect 35756 22316 35924 22318
rect 36316 22372 36372 26852
rect 36540 26514 36596 27020
rect 36540 26462 36542 26514
rect 36594 26462 36596 26514
rect 36540 26450 36596 26462
rect 36988 27634 37044 27646
rect 36988 27582 36990 27634
rect 37042 27582 37044 27634
rect 36652 26180 36708 26190
rect 36652 26086 36708 26124
rect 36428 26068 36484 26078
rect 36428 25618 36484 26012
rect 36428 25566 36430 25618
rect 36482 25566 36484 25618
rect 36428 25554 36484 25566
rect 36764 24610 36820 24622
rect 36764 24558 36766 24610
rect 36818 24558 36820 24610
rect 36428 23716 36484 23726
rect 36428 22594 36484 23660
rect 36764 23604 36820 24558
rect 36988 23940 37044 27582
rect 37100 27076 37156 27114
rect 37100 27010 37156 27020
rect 37212 26908 37268 30716
rect 37548 30210 37604 30222
rect 37548 30158 37550 30210
rect 37602 30158 37604 30210
rect 37436 30100 37492 30110
rect 37548 30100 37604 30158
rect 37492 30044 37604 30100
rect 37436 30034 37492 30044
rect 37436 29652 37492 29662
rect 37436 29558 37492 29596
rect 37324 27972 37380 27982
rect 37324 27858 37380 27916
rect 37548 27860 37604 30044
rect 37660 29876 37716 31500
rect 38220 30882 38276 30894
rect 38220 30830 38222 30882
rect 38274 30830 38276 30882
rect 38220 30212 38276 30830
rect 38220 30146 38276 30156
rect 37660 29820 38276 29876
rect 37660 29428 37716 29820
rect 37884 29650 37940 29662
rect 37884 29598 37886 29650
rect 37938 29598 37940 29650
rect 37772 29428 37828 29438
rect 37660 29426 37828 29428
rect 37660 29374 37774 29426
rect 37826 29374 37828 29426
rect 37660 29372 37828 29374
rect 37772 29362 37828 29372
rect 37324 27806 37326 27858
rect 37378 27806 37380 27858
rect 37324 27794 37380 27806
rect 37436 27804 37604 27860
rect 37772 29092 37828 29102
rect 37436 26908 37492 27804
rect 37548 27636 37604 27646
rect 37548 27542 37604 27580
rect 37548 27188 37604 27198
rect 37772 27188 37828 29036
rect 37884 28084 37940 29598
rect 37996 29652 38052 29662
rect 37996 29426 38052 29596
rect 37996 29374 37998 29426
rect 38050 29374 38052 29426
rect 37996 29362 38052 29374
rect 38220 28642 38276 29820
rect 38220 28590 38222 28642
rect 38274 28590 38276 28642
rect 38220 28578 38276 28590
rect 38556 28644 38612 32732
rect 40012 32788 40068 35644
rect 40012 32722 40068 32732
rect 40348 31220 40404 39340
rect 40460 39172 40516 39182
rect 40460 35028 40516 39116
rect 40460 34934 40516 34972
rect 40796 34692 40852 40796
rect 40908 40786 40964 40796
rect 41020 40626 41076 40796
rect 41020 40574 41022 40626
rect 41074 40574 41076 40626
rect 41020 40562 41076 40574
rect 41580 40628 41636 46396
rect 41916 45332 41972 45342
rect 42028 45332 42084 46508
rect 42700 46498 42756 46508
rect 41972 45276 42084 45332
rect 43148 46004 43204 46014
rect 41916 45266 41972 45276
rect 41692 44996 41748 45006
rect 43036 44996 43092 45006
rect 41692 44994 41972 44996
rect 41692 44942 41694 44994
rect 41746 44942 41972 44994
rect 41692 44940 41972 44942
rect 41692 44930 41748 44940
rect 41916 44546 41972 44940
rect 41916 44494 41918 44546
rect 41970 44494 41972 44546
rect 41916 44482 41972 44494
rect 42028 44436 42084 44446
rect 42476 44436 42532 44446
rect 42028 44434 42532 44436
rect 42028 44382 42030 44434
rect 42082 44382 42478 44434
rect 42530 44382 42532 44434
rect 42028 44380 42532 44382
rect 42028 44370 42084 44380
rect 42476 44370 42532 44380
rect 42812 44324 42868 44334
rect 42812 44230 42868 44268
rect 43036 44322 43092 44940
rect 43036 44270 43038 44322
rect 43090 44270 43092 44322
rect 43036 44258 43092 44270
rect 43148 44212 43204 45948
rect 43484 45780 43540 45790
rect 43484 44434 43540 45724
rect 43596 45332 43652 47292
rect 43596 45276 43876 45332
rect 43820 44996 43876 45276
rect 43820 44902 43876 44940
rect 43484 44382 43486 44434
rect 43538 44382 43540 44434
rect 43484 44370 43540 44382
rect 43372 44324 43428 44334
rect 42476 44100 42532 44110
rect 42476 44006 42532 44044
rect 42588 44098 42644 44110
rect 42588 44046 42590 44098
rect 42642 44046 42644 44098
rect 42588 43540 42644 44046
rect 42588 43316 42644 43484
rect 42588 43250 42644 43260
rect 41692 41860 41748 41870
rect 41692 41858 42308 41860
rect 41692 41806 41694 41858
rect 41746 41806 42308 41858
rect 41692 41804 42308 41806
rect 41692 41794 41748 41804
rect 41580 40572 41860 40628
rect 41692 40402 41748 40414
rect 41692 40350 41694 40402
rect 41746 40350 41748 40402
rect 40908 40292 40964 40302
rect 40964 40236 41076 40292
rect 40908 40198 40964 40236
rect 41020 39618 41076 40236
rect 41244 40180 41300 40190
rect 41244 40086 41300 40124
rect 41692 40180 41748 40350
rect 41692 40114 41748 40124
rect 41020 39566 41022 39618
rect 41074 39566 41076 39618
rect 41020 39554 41076 39566
rect 41356 39620 41412 39630
rect 41804 39620 41860 40572
rect 42252 40626 42308 41804
rect 43148 41186 43204 44156
rect 43260 44322 43428 44324
rect 43260 44270 43374 44322
rect 43426 44270 43428 44322
rect 43260 44268 43428 44270
rect 43260 44100 43316 44268
rect 43260 44034 43316 44044
rect 43372 43708 43428 44268
rect 43820 44324 43876 44334
rect 43596 44098 43652 44110
rect 43596 44046 43598 44098
rect 43650 44046 43652 44098
rect 43596 43876 43652 44046
rect 43596 43810 43652 43820
rect 43820 44098 43876 44268
rect 43820 44046 43822 44098
rect 43874 44046 43876 44098
rect 43820 43708 43876 44046
rect 43372 43652 43540 43708
rect 43260 43540 43316 43550
rect 43260 43426 43316 43484
rect 43260 43374 43262 43426
rect 43314 43374 43316 43426
rect 43260 42756 43316 43374
rect 43260 42690 43316 42700
rect 43148 41134 43150 41186
rect 43202 41134 43204 41186
rect 42252 40574 42254 40626
rect 42306 40574 42308 40626
rect 42252 40562 42308 40574
rect 42364 40964 42420 40974
rect 41916 40514 41972 40526
rect 41916 40462 41918 40514
rect 41970 40462 41972 40514
rect 41916 40292 41972 40462
rect 42364 40514 42420 40908
rect 43148 40628 43204 41134
rect 43484 41186 43540 43652
rect 43708 43652 43876 43708
rect 43484 41134 43486 41186
rect 43538 41134 43540 41186
rect 43372 40628 43428 40638
rect 43148 40626 43428 40628
rect 43148 40574 43374 40626
rect 43426 40574 43428 40626
rect 43148 40572 43428 40574
rect 43372 40562 43428 40572
rect 42364 40462 42366 40514
rect 42418 40462 42420 40514
rect 42364 40450 42420 40462
rect 41916 40226 41972 40236
rect 42588 40292 42644 40302
rect 41916 39620 41972 39630
rect 41356 39506 41412 39564
rect 41356 39454 41358 39506
rect 41410 39454 41412 39506
rect 41356 39442 41412 39454
rect 41468 39618 41972 39620
rect 41468 39566 41918 39618
rect 41970 39566 41972 39618
rect 41468 39564 41972 39566
rect 41468 39284 41524 39564
rect 41916 39554 41972 39564
rect 42140 39620 42196 39630
rect 42140 39526 42196 39564
rect 42588 39618 42644 40236
rect 43484 40292 43540 41134
rect 43484 40226 43540 40236
rect 43596 42756 43652 42766
rect 42588 39566 42590 39618
rect 42642 39566 42644 39618
rect 42588 39554 42644 39566
rect 43596 39508 43652 42700
rect 43708 41412 43764 43652
rect 43820 41860 43876 41870
rect 43932 41860 43988 48076
rect 44268 48038 44324 48076
rect 44492 47684 44548 48190
rect 44940 48244 44996 48254
rect 44940 48150 44996 48188
rect 44492 47618 44548 47628
rect 45052 47684 45108 47694
rect 45164 47684 45220 48862
rect 45724 48802 45780 48814
rect 45724 48750 45726 48802
rect 45778 48750 45780 48802
rect 45612 48692 45668 48702
rect 45612 48354 45668 48636
rect 45612 48302 45614 48354
rect 45666 48302 45668 48354
rect 45612 48290 45668 48302
rect 45052 47682 45220 47684
rect 45052 47630 45054 47682
rect 45106 47630 45220 47682
rect 45052 47628 45220 47630
rect 45276 48132 45332 48142
rect 45052 47618 45108 47628
rect 44940 47460 44996 47470
rect 45276 47460 45332 48076
rect 44940 47458 45332 47460
rect 44940 47406 44942 47458
rect 44994 47406 45332 47458
rect 44940 47404 45332 47406
rect 44940 47394 44996 47404
rect 45724 46788 45780 48750
rect 46060 48468 46116 48478
rect 46060 48374 46116 48412
rect 46172 48356 46228 48366
rect 46172 48262 46228 48300
rect 45836 48242 45892 48254
rect 45836 48190 45838 48242
rect 45890 48190 45892 48242
rect 45836 47572 45892 48190
rect 46956 48244 47012 48254
rect 46956 48150 47012 48188
rect 45948 48132 46004 48142
rect 45948 48038 46004 48076
rect 46620 48020 46676 48030
rect 45836 47506 45892 47516
rect 46060 48018 46676 48020
rect 46060 47966 46622 48018
rect 46674 47966 46676 48018
rect 46060 47964 46676 47966
rect 45724 46732 46004 46788
rect 45948 46452 46004 46732
rect 46060 46786 46116 47964
rect 46620 47954 46676 47964
rect 46060 46734 46062 46786
rect 46114 46734 46116 46786
rect 46060 46722 46116 46734
rect 47068 47570 47124 49420
rect 48188 49140 48244 49150
rect 47964 49138 48244 49140
rect 47964 49086 48190 49138
rect 48242 49086 48244 49138
rect 47964 49084 48244 49086
rect 47180 48580 47236 48590
rect 47180 48130 47236 48524
rect 47180 48078 47182 48130
rect 47234 48078 47236 48130
rect 47180 47796 47236 48078
rect 47180 47730 47236 47740
rect 47292 48356 47348 48366
rect 47068 47518 47070 47570
rect 47122 47518 47124 47570
rect 46172 46676 46228 46686
rect 46172 46582 46228 46620
rect 46284 46674 46340 46686
rect 46284 46622 46286 46674
rect 46338 46622 46340 46674
rect 46284 46452 46340 46622
rect 46620 46674 46676 46686
rect 46620 46622 46622 46674
rect 46674 46622 46676 46674
rect 46620 46564 46676 46622
rect 46620 46498 46676 46508
rect 45948 46396 46340 46452
rect 47068 45892 47124 47518
rect 47180 45892 47236 45902
rect 47068 45890 47236 45892
rect 47068 45838 47182 45890
rect 47234 45838 47236 45890
rect 47068 45836 47236 45838
rect 44044 45780 44100 45790
rect 44044 45686 44100 45724
rect 44156 45668 44212 45678
rect 44156 45666 44996 45668
rect 44156 45614 44158 45666
rect 44210 45614 44996 45666
rect 44156 45612 44996 45614
rect 44156 45602 44212 45612
rect 44268 45332 44324 45342
rect 44268 45106 44324 45276
rect 44940 45218 44996 45612
rect 44940 45166 44942 45218
rect 44994 45166 44996 45218
rect 44940 45154 44996 45166
rect 45388 45332 45444 45342
rect 44268 45054 44270 45106
rect 44322 45054 44324 45106
rect 44268 45042 44324 45054
rect 44044 44324 44100 44334
rect 44044 44230 44100 44268
rect 44268 43764 44324 43774
rect 44268 43652 44324 43708
rect 44156 43650 44324 43652
rect 44156 43598 44270 43650
rect 44322 43598 44324 43650
rect 44156 43596 44324 43598
rect 43820 41858 44100 41860
rect 43820 41806 43822 41858
rect 43874 41806 44100 41858
rect 43820 41804 44100 41806
rect 43820 41794 43876 41804
rect 43708 41356 43988 41412
rect 43708 41188 43764 41198
rect 43708 41094 43764 41132
rect 43820 40964 43876 40974
rect 43820 40870 43876 40908
rect 43932 40962 43988 41356
rect 44044 41186 44100 41804
rect 44044 41134 44046 41186
rect 44098 41134 44100 41186
rect 44044 41122 44100 41134
rect 43932 40910 43934 40962
rect 43986 40910 43988 40962
rect 43932 40740 43988 40910
rect 43820 40684 43988 40740
rect 43820 39620 43876 40684
rect 43820 39554 43876 39564
rect 43932 40402 43988 40414
rect 43932 40350 43934 40402
rect 43986 40350 43988 40402
rect 43596 39442 43652 39452
rect 40908 39228 41524 39284
rect 42252 39394 42308 39406
rect 42252 39342 42254 39394
rect 42306 39342 42308 39394
rect 40908 38722 40964 39228
rect 42252 38948 42308 39342
rect 42364 39396 42420 39406
rect 42364 39302 42420 39340
rect 43148 39396 43204 39406
rect 40908 38670 40910 38722
rect 40962 38670 40964 38722
rect 40908 38658 40964 38670
rect 41916 38892 42308 38948
rect 41916 38162 41972 38892
rect 43036 38724 43092 38734
rect 42028 38722 43092 38724
rect 42028 38670 43038 38722
rect 43090 38670 43092 38722
rect 42028 38668 43092 38670
rect 42028 38274 42084 38668
rect 43036 38658 43092 38668
rect 43148 38668 43204 39340
rect 43932 39060 43988 40350
rect 44156 40068 44212 43596
rect 44268 43586 44324 43596
rect 45388 43538 45444 45276
rect 47068 45332 47124 45836
rect 47180 45826 47236 45836
rect 47068 45266 47124 45276
rect 47068 44996 47124 45006
rect 47292 44996 47348 48300
rect 47852 48356 47908 48366
rect 47516 48244 47572 48254
rect 47516 48130 47572 48188
rect 47852 48242 47908 48300
rect 47852 48190 47854 48242
rect 47906 48190 47908 48242
rect 47852 48178 47908 48190
rect 47516 48078 47518 48130
rect 47570 48078 47572 48130
rect 47516 48066 47572 48078
rect 47964 46002 48020 49084
rect 48188 49074 48244 49084
rect 48300 48914 48356 51772
rect 48860 51378 48916 51886
rect 48860 51326 48862 51378
rect 48914 51326 48916 51378
rect 48860 51314 48916 51326
rect 48972 51378 49028 52332
rect 49644 52274 49700 52332
rect 49644 52222 49646 52274
rect 49698 52222 49700 52274
rect 49644 52210 49700 52222
rect 49196 52162 49252 52174
rect 49196 52110 49198 52162
rect 49250 52110 49252 52162
rect 49196 52052 49252 52110
rect 49196 51986 49252 51996
rect 49532 52164 49588 52174
rect 49420 51940 49476 51950
rect 49308 51884 49420 51940
rect 48972 51326 48974 51378
rect 49026 51326 49028 51378
rect 48972 49924 49028 51326
rect 49196 51380 49252 51390
rect 49308 51380 49364 51884
rect 49420 51874 49476 51884
rect 49532 51492 49588 52108
rect 49644 51492 49700 51502
rect 49532 51490 49700 51492
rect 49532 51438 49646 51490
rect 49698 51438 49700 51490
rect 49532 51436 49700 51438
rect 49644 51426 49700 51436
rect 49196 51378 49364 51380
rect 49196 51326 49198 51378
rect 49250 51326 49364 51378
rect 49196 51324 49364 51326
rect 49196 51314 49252 51324
rect 49308 51154 49364 51166
rect 49308 51102 49310 51154
rect 49362 51102 49364 51154
rect 48972 49810 49028 49868
rect 48972 49758 48974 49810
rect 49026 49758 49028 49810
rect 48972 49746 49028 49758
rect 49196 50708 49252 50718
rect 49196 49810 49252 50652
rect 49196 49758 49198 49810
rect 49250 49758 49252 49810
rect 49196 49746 49252 49758
rect 48748 49700 48804 49710
rect 48524 49698 48804 49700
rect 48524 49646 48750 49698
rect 48802 49646 48804 49698
rect 48524 49644 48804 49646
rect 48524 49250 48580 49644
rect 48748 49634 48804 49644
rect 49308 49588 49364 51102
rect 49756 51044 49812 53452
rect 50428 53452 50596 53508
rect 50876 53732 50932 53742
rect 50428 53172 50484 53452
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 50652 53172 50708 53182
rect 50876 53172 50932 53676
rect 51660 53732 51716 53742
rect 52108 53732 52164 55358
rect 51660 53730 52164 53732
rect 51660 53678 51662 53730
rect 51714 53678 52164 53730
rect 51660 53676 52164 53678
rect 52220 55412 52724 55468
rect 55580 55412 55636 55422
rect 51324 53620 51380 53630
rect 50428 53116 50596 53172
rect 49980 53060 50036 53070
rect 49980 52966 50036 53004
rect 50092 52948 50148 52958
rect 50092 52854 50148 52892
rect 50204 52948 50260 52958
rect 50204 52946 50372 52948
rect 50204 52894 50206 52946
rect 50258 52894 50372 52946
rect 50204 52892 50372 52894
rect 50204 52882 50260 52892
rect 50316 52276 50372 52892
rect 50316 52220 50484 52276
rect 49308 49522 49364 49532
rect 49532 50988 49812 51044
rect 49868 52164 49924 52174
rect 50204 52164 50260 52174
rect 49868 52162 50260 52164
rect 49868 52110 49870 52162
rect 49922 52110 50206 52162
rect 50258 52110 50260 52162
rect 49868 52108 50260 52110
rect 49532 50818 49588 50988
rect 49532 50766 49534 50818
rect 49586 50766 49588 50818
rect 48524 49198 48526 49250
rect 48578 49198 48580 49250
rect 48524 49186 48580 49198
rect 48300 48862 48302 48914
rect 48354 48862 48356 48914
rect 48300 48850 48356 48862
rect 48076 48356 48132 48366
rect 48076 48262 48132 48300
rect 49532 48356 49588 50766
rect 49644 50820 49700 50830
rect 49868 50820 49924 52108
rect 50204 51378 50260 52108
rect 50316 52052 50372 52062
rect 50316 51958 50372 51996
rect 50428 51828 50484 52220
rect 50540 51940 50596 53116
rect 50652 53170 50932 53172
rect 50652 53118 50654 53170
rect 50706 53118 50932 53170
rect 50652 53116 50932 53118
rect 50988 53618 51380 53620
rect 50988 53566 51326 53618
rect 51378 53566 51380 53618
rect 50988 53564 51380 53566
rect 50652 53106 50708 53116
rect 50540 51874 50596 51884
rect 50204 51326 50206 51378
rect 50258 51326 50260 51378
rect 50204 51314 50260 51326
rect 50316 51772 50484 51828
rect 50556 51772 50820 51782
rect 49644 50818 49924 50820
rect 49644 50766 49646 50818
rect 49698 50766 49924 50818
rect 49644 50764 49924 50766
rect 50092 50820 50148 50830
rect 49644 50754 49700 50764
rect 50092 50726 50148 50764
rect 50204 50820 50260 50830
rect 50316 50820 50372 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 50204 50818 50372 50820
rect 50204 50766 50206 50818
rect 50258 50766 50372 50818
rect 50204 50764 50372 50766
rect 50652 51378 50708 51390
rect 50652 51326 50654 51378
rect 50706 51326 50708 51378
rect 50652 50818 50708 51326
rect 50652 50766 50654 50818
rect 50706 50766 50708 50818
rect 50204 50754 50260 50764
rect 49980 50708 50036 50718
rect 49868 50596 49924 50606
rect 49980 50596 50036 50652
rect 50652 50708 50708 50766
rect 50652 50642 50708 50652
rect 50764 51380 50820 51390
rect 49868 50594 50036 50596
rect 49868 50542 49870 50594
rect 49922 50542 50036 50594
rect 49868 50540 50036 50542
rect 49868 50530 49924 50540
rect 50540 50484 50596 50494
rect 50316 50482 50596 50484
rect 50316 50430 50542 50482
rect 50594 50430 50596 50482
rect 50316 50428 50596 50430
rect 50204 49924 50260 49934
rect 50204 49830 50260 49868
rect 50316 49922 50372 50428
rect 50540 50418 50596 50428
rect 50764 50484 50820 51324
rect 50988 51268 51044 53564
rect 51324 53554 51380 53564
rect 51660 53060 51716 53676
rect 51212 52052 51268 52062
rect 51212 52050 51380 52052
rect 51212 51998 51214 52050
rect 51266 51998 51380 52050
rect 51212 51996 51380 51998
rect 51212 51986 51268 51996
rect 51100 51938 51156 51950
rect 51100 51886 51102 51938
rect 51154 51886 51156 51938
rect 51100 51492 51156 51886
rect 51212 51492 51268 51502
rect 51100 51490 51268 51492
rect 51100 51438 51214 51490
rect 51266 51438 51268 51490
rect 51100 51436 51268 51438
rect 50988 51266 51156 51268
rect 50988 51214 50990 51266
rect 51042 51214 51156 51266
rect 50988 51212 51156 51214
rect 50988 51202 51044 51212
rect 50988 50484 51044 50494
rect 50764 50418 50820 50428
rect 50876 50482 51044 50484
rect 50876 50430 50990 50482
rect 51042 50430 51044 50482
rect 50876 50428 51044 50430
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 50540 50036 50596 50046
rect 50876 50036 50932 50428
rect 50988 50418 51044 50428
rect 51100 50372 51156 51212
rect 51212 50820 51268 51436
rect 51324 51268 51380 51996
rect 51660 51492 51716 53004
rect 51660 51436 51940 51492
rect 51660 51268 51716 51278
rect 51324 51266 51716 51268
rect 51324 51214 51662 51266
rect 51714 51214 51716 51266
rect 51324 51212 51716 51214
rect 51212 50594 51268 50764
rect 51436 50596 51492 50606
rect 51212 50542 51214 50594
rect 51266 50542 51268 50594
rect 51212 50530 51268 50542
rect 51324 50594 51492 50596
rect 51324 50542 51438 50594
rect 51490 50542 51492 50594
rect 51324 50540 51492 50542
rect 51324 50372 51380 50540
rect 51436 50530 51492 50540
rect 51548 50594 51604 50606
rect 51548 50542 51550 50594
rect 51602 50542 51604 50594
rect 51548 50484 51604 50542
rect 51548 50418 51604 50428
rect 51100 50316 51380 50372
rect 50540 50034 50932 50036
rect 50540 49982 50542 50034
rect 50594 49982 50932 50034
rect 50540 49980 50932 49982
rect 50988 50260 51044 50270
rect 50988 50034 51044 50204
rect 50988 49982 50990 50034
rect 51042 49982 51044 50034
rect 50540 49970 50596 49980
rect 50988 49970 51044 49982
rect 50316 49870 50318 49922
rect 50370 49870 50372 49922
rect 50316 48468 50372 49870
rect 51548 49588 51604 49598
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 49532 48290 49588 48300
rect 50204 48412 50372 48468
rect 49980 48132 50036 48142
rect 50204 48132 50260 48412
rect 51548 48354 51604 49532
rect 51548 48302 51550 48354
rect 51602 48302 51604 48354
rect 51548 48290 51604 48302
rect 49980 48130 50260 48132
rect 49980 48078 49982 48130
rect 50034 48078 50260 48130
rect 49980 48076 50260 48078
rect 50316 48242 50372 48254
rect 50316 48190 50318 48242
rect 50370 48190 50372 48242
rect 49868 47348 49924 47358
rect 49868 46676 49924 47292
rect 49756 46674 49924 46676
rect 49756 46622 49870 46674
rect 49922 46622 49924 46674
rect 49756 46620 49924 46622
rect 49644 46452 49700 46462
rect 49644 46358 49700 46396
rect 47964 45950 47966 46002
rect 48018 45950 48020 46002
rect 47964 45938 48020 45950
rect 49420 45668 49476 45678
rect 47068 44994 47348 44996
rect 47068 44942 47070 44994
rect 47122 44942 47348 44994
rect 47068 44940 47348 44942
rect 48188 44996 48244 45006
rect 45388 43486 45390 43538
rect 45442 43486 45444 43538
rect 45388 43474 45444 43486
rect 45500 44322 45556 44334
rect 45500 44270 45502 44322
rect 45554 44270 45556 44322
rect 44716 43428 44772 43438
rect 44716 43334 44772 43372
rect 45500 43428 45556 44270
rect 47068 44324 47124 44940
rect 47068 44258 47124 44268
rect 45500 43362 45556 43372
rect 46060 43428 46116 43438
rect 46060 43426 46340 43428
rect 46060 43374 46062 43426
rect 46114 43374 46340 43426
rect 46060 43372 46340 43374
rect 46060 43362 46116 43372
rect 46284 42978 46340 43372
rect 48188 43426 48244 44940
rect 49084 44996 49140 45006
rect 49084 44902 49140 44940
rect 49420 44994 49476 45612
rect 49756 45220 49812 46620
rect 49868 46610 49924 46620
rect 49980 46452 50036 48076
rect 50316 46900 50372 48190
rect 50876 48244 50932 48254
rect 50876 48242 51044 48244
rect 50876 48190 50878 48242
rect 50930 48190 51044 48242
rect 50876 48188 51044 48190
rect 50876 48178 50932 48188
rect 50652 47572 50708 47582
rect 50652 47458 50708 47516
rect 50652 47406 50654 47458
rect 50706 47406 50708 47458
rect 50652 47394 50708 47406
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 50316 46844 50484 46900
rect 50092 46674 50148 46686
rect 50092 46622 50094 46674
rect 50146 46622 50148 46674
rect 50092 46452 50148 46622
rect 50316 46676 50372 46686
rect 50316 46582 50372 46620
rect 49868 46396 50148 46452
rect 50204 46562 50260 46574
rect 50204 46510 50206 46562
rect 50258 46510 50260 46562
rect 49868 45444 49924 46396
rect 50204 46228 50260 46510
rect 49868 45378 49924 45388
rect 49980 46172 50260 46228
rect 49980 45332 50036 46172
rect 50092 46004 50148 46014
rect 50428 46004 50484 46844
rect 50092 46002 50484 46004
rect 50092 45950 50094 46002
rect 50146 45950 50484 46002
rect 50092 45948 50484 45950
rect 50092 45938 50148 45948
rect 50428 45890 50484 45948
rect 50428 45838 50430 45890
rect 50482 45838 50484 45890
rect 50428 45826 50484 45838
rect 50540 46676 50596 46686
rect 50540 45668 50596 46620
rect 50540 45602 50596 45612
rect 50876 46674 50932 46686
rect 50876 46622 50878 46674
rect 50930 46622 50932 46674
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50316 45332 50372 45342
rect 49980 45276 50260 45332
rect 49756 45164 50148 45220
rect 50092 45106 50148 45164
rect 50092 45054 50094 45106
rect 50146 45054 50148 45106
rect 49420 44942 49422 44994
rect 49474 44942 49476 44994
rect 48188 43374 48190 43426
rect 48242 43374 48244 43426
rect 48188 43362 48244 43374
rect 49420 43540 49476 44942
rect 49756 44996 49812 45006
rect 49756 44994 50036 44996
rect 49756 44942 49758 44994
rect 49810 44942 50036 44994
rect 49756 44940 50036 44942
rect 49756 44930 49812 44940
rect 49756 44436 49812 44446
rect 49756 44342 49812 44380
rect 46284 42926 46286 42978
rect 46338 42926 46340 42978
rect 46284 42914 46340 42926
rect 46732 42980 46788 42990
rect 46732 42886 46788 42924
rect 49420 42980 49476 43484
rect 49420 42914 49476 42924
rect 46284 42754 46340 42766
rect 46284 42702 46286 42754
rect 46338 42702 46340 42754
rect 45500 42644 45556 42654
rect 44940 42532 44996 42542
rect 44828 42196 44884 42206
rect 44828 42102 44884 42140
rect 44380 42084 44436 42094
rect 44268 42028 44380 42084
rect 44268 40628 44324 42028
rect 44380 42018 44436 42028
rect 44492 41858 44548 41870
rect 44492 41806 44494 41858
rect 44546 41806 44548 41858
rect 44492 41188 44548 41806
rect 44492 41122 44548 41132
rect 44268 40626 44548 40628
rect 44268 40574 44270 40626
rect 44322 40574 44548 40626
rect 44268 40572 44548 40574
rect 44268 40562 44324 40572
rect 44492 40516 44548 40572
rect 44828 40516 44884 40526
rect 44492 40514 44884 40516
rect 44492 40462 44830 40514
rect 44882 40462 44884 40514
rect 44492 40460 44884 40462
rect 44828 40450 44884 40460
rect 44940 40514 44996 42476
rect 45276 42196 45332 42206
rect 45276 42102 45332 42140
rect 45500 42194 45556 42588
rect 46172 42644 46228 42654
rect 46172 42550 46228 42588
rect 45948 42532 46004 42542
rect 45500 42142 45502 42194
rect 45554 42142 45556 42194
rect 45500 42130 45556 42142
rect 45724 42530 46116 42532
rect 45724 42478 45950 42530
rect 46002 42478 46116 42530
rect 45724 42476 46116 42478
rect 45164 42084 45220 42094
rect 45164 41990 45220 42028
rect 45164 41188 45220 41198
rect 44940 40462 44942 40514
rect 44994 40462 44996 40514
rect 44156 40002 44212 40012
rect 44940 39394 44996 40462
rect 44940 39342 44942 39394
rect 44994 39342 44996 39394
rect 44940 39284 44996 39342
rect 43820 38834 43876 38846
rect 43820 38782 43822 38834
rect 43874 38782 43876 38834
rect 43148 38612 43652 38668
rect 42028 38222 42030 38274
rect 42082 38222 42084 38274
rect 42028 38210 42084 38222
rect 41916 38110 41918 38162
rect 41970 38110 41972 38162
rect 41916 38098 41972 38110
rect 43596 38164 43652 38612
rect 43596 38050 43652 38108
rect 43596 37998 43598 38050
rect 43650 37998 43652 38050
rect 43596 37986 43652 37998
rect 43708 38500 43764 38510
rect 43708 38162 43764 38444
rect 43708 38110 43710 38162
rect 43762 38110 43764 38162
rect 42028 37604 42084 37614
rect 42028 37266 42084 37548
rect 43484 37380 43540 37390
rect 42028 37214 42030 37266
rect 42082 37214 42084 37266
rect 41580 36482 41636 36494
rect 41580 36430 41582 36482
rect 41634 36430 41636 36482
rect 41580 36372 41636 36430
rect 41468 36316 41580 36372
rect 41244 35140 41300 35150
rect 41244 35046 41300 35084
rect 41468 34916 41524 36316
rect 41580 36306 41636 36316
rect 41804 35810 41860 35822
rect 41804 35758 41806 35810
rect 41858 35758 41860 35810
rect 41580 35700 41636 35710
rect 41580 35138 41636 35644
rect 41580 35086 41582 35138
rect 41634 35086 41636 35138
rect 41580 35074 41636 35086
rect 41692 35140 41748 35150
rect 41468 34860 41636 34916
rect 40908 34692 40964 34702
rect 41468 34692 41524 34702
rect 40796 34690 41524 34692
rect 40796 34638 40910 34690
rect 40962 34638 41470 34690
rect 41522 34638 41524 34690
rect 40796 34636 41524 34638
rect 40348 31154 40404 31164
rect 40460 32116 40516 32126
rect 40348 30996 40404 31006
rect 40348 30882 40404 30940
rect 40348 30830 40350 30882
rect 40402 30830 40404 30882
rect 40348 30818 40404 30830
rect 39452 30324 39508 30334
rect 39340 30212 39396 30222
rect 39340 30118 39396 30156
rect 39452 30210 39508 30268
rect 39452 30158 39454 30210
rect 39506 30158 39508 30210
rect 39452 30146 39508 30158
rect 39900 29988 39956 29998
rect 39900 28754 39956 29932
rect 39900 28702 39902 28754
rect 39954 28702 39956 28754
rect 39900 28690 39956 28702
rect 38556 28588 38724 28644
rect 38556 28420 38612 28430
rect 38332 28418 38612 28420
rect 38332 28366 38558 28418
rect 38610 28366 38612 28418
rect 38332 28364 38612 28366
rect 37884 28028 38052 28084
rect 37548 27186 37828 27188
rect 37548 27134 37550 27186
rect 37602 27134 37828 27186
rect 37548 27132 37828 27134
rect 37884 27634 37940 27646
rect 37884 27582 37886 27634
rect 37938 27582 37940 27634
rect 37548 27122 37604 27132
rect 37884 26908 37940 27582
rect 37100 26852 37268 26908
rect 37324 26852 37492 26908
rect 37660 26852 37940 26908
rect 37100 26516 37156 26852
rect 37100 26422 37156 26460
rect 37324 26292 37380 26852
rect 37212 26236 37380 26292
rect 37436 26290 37492 26302
rect 37436 26238 37438 26290
rect 37490 26238 37492 26290
rect 37212 23940 37268 26236
rect 37436 26180 37492 26238
rect 37436 26114 37492 26124
rect 37324 26068 37380 26078
rect 37324 25508 37380 26012
rect 37324 25506 37492 25508
rect 37324 25454 37326 25506
rect 37378 25454 37492 25506
rect 37324 25452 37492 25454
rect 37324 25442 37380 25452
rect 37436 24946 37492 25452
rect 37436 24894 37438 24946
rect 37490 24894 37492 24946
rect 37436 24724 37492 24894
rect 37548 24724 37604 24734
rect 37436 24722 37604 24724
rect 37436 24670 37550 24722
rect 37602 24670 37604 24722
rect 37436 24668 37604 24670
rect 37548 24658 37604 24668
rect 37436 23940 37492 23950
rect 36988 23884 37156 23940
rect 37212 23884 37380 23940
rect 36876 23828 36932 23838
rect 36876 23734 36932 23772
rect 36988 23714 37044 23726
rect 36988 23662 36990 23714
rect 37042 23662 37044 23714
rect 36988 23604 37044 23662
rect 36764 23548 37044 23604
rect 36428 22542 36430 22594
rect 36482 22542 36484 22594
rect 36428 22530 36484 22542
rect 36876 23156 36932 23548
rect 36316 22316 36820 22372
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 34524 18386 34580 18396
rect 34748 18844 35028 18900
rect 35084 20804 35140 20814
rect 33852 18162 33908 18172
rect 33740 17948 34244 18004
rect 33628 17668 33684 17678
rect 33516 17666 33684 17668
rect 33516 17614 33630 17666
rect 33682 17614 33684 17666
rect 33516 17612 33684 17614
rect 33628 17602 33684 17612
rect 34188 17666 34244 17948
rect 34188 17614 34190 17666
rect 34242 17614 34244 17666
rect 34188 17602 34244 17614
rect 33740 17444 33796 17454
rect 33180 17442 33796 17444
rect 33180 17390 33742 17442
rect 33794 17390 33796 17442
rect 33180 17388 33796 17390
rect 33740 17378 33796 17388
rect 33964 17442 34020 17454
rect 33964 17390 33966 17442
rect 34018 17390 34020 17442
rect 33964 17332 34020 17390
rect 34300 17442 34356 17454
rect 34300 17390 34302 17442
rect 34354 17390 34356 17442
rect 34300 17332 34356 17390
rect 33964 17276 34356 17332
rect 34524 17442 34580 17454
rect 34524 17390 34526 17442
rect 34578 17390 34580 17442
rect 33740 15596 34356 15652
rect 33628 15428 33684 15438
rect 33516 15426 33684 15428
rect 33516 15374 33630 15426
rect 33682 15374 33684 15426
rect 33516 15372 33684 15374
rect 33404 15204 33460 15214
rect 33516 15204 33572 15372
rect 33628 15362 33684 15372
rect 33740 15426 33796 15596
rect 33740 15374 33742 15426
rect 33794 15374 33796 15426
rect 33740 15362 33796 15374
rect 34300 15428 34356 15596
rect 34412 15428 34468 15438
rect 34524 15428 34580 17390
rect 34300 15426 34580 15428
rect 34300 15374 34414 15426
rect 34466 15374 34580 15426
rect 34300 15372 34580 15374
rect 34412 15362 34468 15372
rect 33460 15148 33572 15204
rect 34076 15314 34132 15326
rect 34076 15262 34078 15314
rect 34130 15262 34132 15314
rect 34076 15204 34132 15262
rect 33404 15138 33460 15148
rect 34076 15138 34132 15148
rect 34300 15202 34356 15214
rect 34300 15150 34302 15202
rect 34354 15150 34356 15202
rect 34300 15148 34356 15150
rect 33628 15092 33684 15102
rect 34300 15092 34468 15148
rect 33516 15090 33684 15092
rect 33516 15038 33630 15090
rect 33682 15038 33684 15090
rect 33516 15036 33684 15038
rect 33516 14420 33572 15036
rect 33628 15026 33684 15036
rect 33516 14354 33572 14364
rect 34076 13916 34356 13972
rect 33852 13860 33908 13870
rect 34076 13860 34132 13916
rect 33852 13858 34132 13860
rect 33852 13806 33854 13858
rect 33906 13806 34132 13858
rect 33852 13804 34132 13806
rect 34300 13858 34356 13916
rect 34300 13806 34302 13858
rect 34354 13806 34356 13858
rect 33852 13794 33908 13804
rect 33068 13122 33124 13132
rect 33516 13634 33572 13646
rect 33516 13582 33518 13634
rect 33570 13582 33572 13634
rect 31836 12910 31838 12962
rect 31890 12910 31892 12962
rect 31836 12898 31892 12910
rect 33516 12852 33572 13582
rect 34300 13524 34356 13806
rect 34412 13748 34468 15092
rect 34412 13682 34468 13692
rect 34300 13458 34356 13468
rect 33852 12964 33908 12974
rect 33852 12870 33908 12908
rect 34636 12964 34692 12974
rect 34636 12870 34692 12908
rect 33516 12786 33572 12796
rect 33964 12850 34020 12862
rect 33964 12798 33966 12850
rect 34018 12798 34020 12850
rect 31724 12738 31780 12750
rect 31724 12686 31726 12738
rect 31778 12686 31780 12738
rect 31724 11508 31780 12686
rect 31836 11508 31892 11518
rect 31724 11506 31892 11508
rect 31724 11454 31838 11506
rect 31890 11454 31892 11506
rect 31724 11452 31892 11454
rect 31836 11442 31892 11452
rect 33964 11506 34020 12798
rect 34748 12740 34804 18844
rect 35084 18676 35140 20748
rect 35756 20692 35812 22316
rect 36316 21586 36372 21598
rect 36316 21534 36318 21586
rect 36370 21534 36372 21586
rect 35980 21476 36036 21486
rect 36316 21476 36372 21534
rect 35980 21474 36372 21476
rect 35980 21422 35982 21474
rect 36034 21422 36372 21474
rect 35980 21420 36372 21422
rect 35980 20804 36036 21420
rect 35980 20738 36036 20748
rect 35756 20626 35812 20636
rect 35980 20580 36036 20590
rect 36428 20580 36484 22316
rect 36764 21810 36820 22316
rect 36764 21758 36766 21810
rect 36818 21758 36820 21810
rect 36764 21746 36820 21758
rect 36540 21588 36596 21598
rect 36540 21494 36596 21532
rect 36652 21476 36708 21486
rect 36652 21382 36708 21420
rect 35980 20578 36484 20580
rect 35980 20526 35982 20578
rect 36034 20526 36484 20578
rect 35980 20524 36484 20526
rect 35980 20514 36036 20524
rect 35980 20356 36036 20366
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 34860 18620 35140 18676
rect 34860 15148 34916 18620
rect 35084 18340 35140 18350
rect 35084 18246 35140 18284
rect 34972 18228 35028 18238
rect 34972 17892 35028 18172
rect 35532 18228 35588 18238
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35420 17892 35476 17902
rect 34972 17890 35476 17892
rect 34972 17838 35422 17890
rect 35474 17838 35476 17890
rect 34972 17836 35476 17838
rect 35420 17826 35476 17836
rect 35532 17778 35588 18172
rect 35532 17726 35534 17778
rect 35586 17726 35588 17778
rect 35532 17714 35588 17726
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35980 16210 36036 20300
rect 36092 18340 36148 18350
rect 36092 17890 36148 18284
rect 36092 17838 36094 17890
rect 36146 17838 36148 17890
rect 36092 17826 36148 17838
rect 36204 17780 36260 17790
rect 36204 17686 36260 17724
rect 35980 16158 35982 16210
rect 36034 16158 36036 16210
rect 35980 16100 36036 16158
rect 35980 16034 36036 16044
rect 36428 15988 36484 15998
rect 36428 15894 36484 15932
rect 36092 15876 36148 15886
rect 35308 15428 35364 15438
rect 34860 15092 35140 15148
rect 35084 14420 35140 15092
rect 35308 15090 35364 15372
rect 35308 15038 35310 15090
rect 35362 15038 35364 15090
rect 35308 15026 35364 15038
rect 35532 15316 35588 15326
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35532 14530 35588 15260
rect 35980 15314 36036 15326
rect 35980 15262 35982 15314
rect 36034 15262 36036 15314
rect 35980 15148 36036 15262
rect 35532 14478 35534 14530
rect 35586 14478 35588 14530
rect 35532 14466 35588 14478
rect 35868 15092 36036 15148
rect 35196 14420 35252 14430
rect 35756 14420 35812 14430
rect 35084 14418 35252 14420
rect 35084 14366 35198 14418
rect 35250 14366 35252 14418
rect 35084 14364 35252 14366
rect 34972 14308 35028 14318
rect 34972 14214 35028 14252
rect 34860 13860 34916 13870
rect 34860 13746 34916 13804
rect 34860 13694 34862 13746
rect 34914 13694 34916 13746
rect 34860 13682 34916 13694
rect 35084 12962 35140 14364
rect 35196 14354 35252 14364
rect 35644 14418 35812 14420
rect 35644 14366 35758 14418
rect 35810 14366 35812 14418
rect 35644 14364 35812 14366
rect 35308 14308 35364 14318
rect 35308 14306 35588 14308
rect 35308 14254 35310 14306
rect 35362 14254 35588 14306
rect 35308 14252 35588 14254
rect 35308 14242 35364 14252
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35084 12910 35086 12962
rect 35138 12910 35140 12962
rect 35084 12898 35140 12910
rect 35532 12964 35588 14252
rect 35644 13860 35700 14364
rect 35756 14354 35812 14364
rect 35756 13972 35812 13982
rect 35868 13972 35924 15092
rect 35980 14532 36036 14542
rect 36092 14532 36148 15820
rect 35980 14530 36148 14532
rect 35980 14478 35982 14530
rect 36034 14478 36148 14530
rect 35980 14476 36148 14478
rect 36316 15764 36372 15774
rect 36316 14530 36372 15708
rect 36316 14478 36318 14530
rect 36370 14478 36372 14530
rect 35980 14466 36036 14476
rect 36316 14466 36372 14478
rect 36428 15314 36484 15326
rect 36428 15262 36430 15314
rect 36482 15262 36484 15314
rect 35756 13970 35924 13972
rect 35756 13918 35758 13970
rect 35810 13918 35924 13970
rect 35756 13916 35924 13918
rect 36092 14306 36148 14318
rect 36092 14254 36094 14306
rect 36146 14254 36148 14306
rect 35756 13906 35812 13916
rect 35644 13748 35700 13804
rect 35980 13748 36036 13758
rect 35644 13692 35924 13748
rect 35532 12898 35588 12908
rect 35756 13524 35812 13534
rect 35756 12962 35812 13468
rect 35756 12910 35758 12962
rect 35810 12910 35812 12962
rect 35756 12898 35812 12910
rect 35868 13074 35924 13692
rect 35980 13654 36036 13692
rect 35868 13022 35870 13074
rect 35922 13022 35924 13074
rect 34748 12674 34804 12684
rect 33964 11454 33966 11506
rect 34018 11454 34020 11506
rect 33964 11442 34020 11454
rect 34636 12066 34692 12078
rect 34636 12014 34638 12066
rect 34690 12014 34692 12066
rect 34636 11396 34692 12014
rect 35196 11956 35252 11966
rect 34524 10612 34580 10622
rect 34636 10612 34692 11340
rect 35084 11900 35196 11956
rect 35084 10724 35140 11900
rect 35196 11890 35252 11900
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35868 10836 35924 13022
rect 36092 13076 36148 14254
rect 36204 14308 36260 14318
rect 36204 13524 36260 14252
rect 36204 13458 36260 13468
rect 36092 13010 36148 13020
rect 36092 12852 36148 12862
rect 36428 12852 36484 15262
rect 36652 15316 36708 15326
rect 36652 15222 36708 15260
rect 36876 15148 36932 23100
rect 36988 21588 37044 21598
rect 37100 21588 37156 23884
rect 37212 23716 37268 23726
rect 37212 23622 37268 23660
rect 37212 23380 37268 23390
rect 37212 22370 37268 23324
rect 37212 22318 37214 22370
rect 37266 22318 37268 22370
rect 37212 22306 37268 22318
rect 37324 21812 37380 23884
rect 37436 23846 37492 23884
rect 36988 21586 37156 21588
rect 36988 21534 36990 21586
rect 37042 21534 37156 21586
rect 36988 21532 37156 21534
rect 36988 21522 37044 21532
rect 37100 21364 37156 21532
rect 37100 21298 37156 21308
rect 37212 21756 37380 21812
rect 36988 20690 37044 20702
rect 36988 20638 36990 20690
rect 37042 20638 37044 20690
rect 36988 20580 37044 20638
rect 37100 20580 37156 20590
rect 36988 20524 37100 20580
rect 37100 20514 37156 20524
rect 37212 20356 37268 21756
rect 37436 21700 37492 21710
rect 37324 21588 37380 21598
rect 37324 21474 37380 21532
rect 37324 21422 37326 21474
rect 37378 21422 37380 21474
rect 37324 20802 37380 21422
rect 37324 20750 37326 20802
rect 37378 20750 37380 20802
rect 37324 20738 37380 20750
rect 36092 12850 36484 12852
rect 36092 12798 36094 12850
rect 36146 12798 36484 12850
rect 36092 12796 36484 12798
rect 36540 15092 36932 15148
rect 36988 20300 37268 20356
rect 36988 15148 37044 20300
rect 37436 19796 37492 21644
rect 37660 21588 37716 26852
rect 37772 26402 37828 26414
rect 37772 26350 37774 26402
rect 37826 26350 37828 26402
rect 37772 24724 37828 26350
rect 37884 26404 37940 26414
rect 37884 25620 37940 26348
rect 37884 25526 37940 25564
rect 37996 25060 38052 28028
rect 38332 27636 38388 28364
rect 38556 28354 38612 28364
rect 38556 27972 38612 27982
rect 38556 27858 38612 27916
rect 38556 27806 38558 27858
rect 38610 27806 38612 27858
rect 38556 27794 38612 27806
rect 38668 27860 38724 28588
rect 39228 28642 39284 28654
rect 39228 28590 39230 28642
rect 39282 28590 39284 28642
rect 38780 27860 38836 27870
rect 38668 27858 38836 27860
rect 38668 27806 38782 27858
rect 38834 27806 38836 27858
rect 38668 27804 38836 27806
rect 38220 27580 38388 27636
rect 38108 26516 38164 26526
rect 38108 26422 38164 26460
rect 38108 25060 38164 25070
rect 37996 25004 38108 25060
rect 38108 24994 38164 25004
rect 38220 24948 38276 27580
rect 38332 27188 38388 27198
rect 38668 27188 38724 27804
rect 38780 27794 38836 27804
rect 39116 27636 39172 27646
rect 39116 27542 39172 27580
rect 38332 27186 38724 27188
rect 38332 27134 38334 27186
rect 38386 27134 38724 27186
rect 38332 27132 38724 27134
rect 38332 27122 38388 27132
rect 38780 26962 38836 26974
rect 38780 26910 38782 26962
rect 38834 26910 38836 26962
rect 38780 26908 38836 26910
rect 38668 26852 38836 26908
rect 39228 26852 39284 28590
rect 38556 26180 38612 26190
rect 38668 26180 38724 26852
rect 38612 26124 38724 26180
rect 38892 26796 39228 26852
rect 38556 25284 38612 26124
rect 38668 25508 38724 25518
rect 38892 25508 38948 26796
rect 39228 26786 39284 26796
rect 39004 26516 39060 26526
rect 39004 26422 39060 26460
rect 39676 26180 39732 26190
rect 39676 26178 40068 26180
rect 39676 26126 39678 26178
rect 39730 26126 40068 26178
rect 39676 26124 40068 26126
rect 39676 26114 39732 26124
rect 39564 26068 39620 26078
rect 39340 26066 39620 26068
rect 39340 26014 39566 26066
rect 39618 26014 39620 26066
rect 39340 26012 39620 26014
rect 39340 25618 39396 26012
rect 39564 26002 39620 26012
rect 39340 25566 39342 25618
rect 39394 25566 39396 25618
rect 39340 25554 39396 25566
rect 38668 25506 38948 25508
rect 38668 25454 38670 25506
rect 38722 25454 38948 25506
rect 38668 25452 38948 25454
rect 38668 25442 38724 25452
rect 38556 25218 38612 25228
rect 39564 25284 39620 25294
rect 38220 24882 38276 24892
rect 39116 25060 39172 25070
rect 37996 24836 38052 24846
rect 37996 24742 38052 24780
rect 38332 24836 38388 24846
rect 37772 24658 37828 24668
rect 38220 24724 38276 24734
rect 38332 24724 38388 24780
rect 38220 24722 38388 24724
rect 38220 24670 38222 24722
rect 38274 24670 38388 24722
rect 38220 24668 38388 24670
rect 38668 24724 38724 24734
rect 38108 24610 38164 24622
rect 38108 24558 38110 24610
rect 38162 24558 38164 24610
rect 38108 23940 38164 24558
rect 38220 24612 38276 24668
rect 38220 24546 38276 24556
rect 38108 23874 38164 23884
rect 38556 23826 38612 23838
rect 38556 23774 38558 23826
rect 38610 23774 38612 23826
rect 38444 23716 38500 23726
rect 37996 23714 38500 23716
rect 37996 23662 38446 23714
rect 38498 23662 38500 23714
rect 37996 23660 38500 23662
rect 37996 22482 38052 23660
rect 38444 23650 38500 23660
rect 37996 22430 37998 22482
rect 38050 22430 38052 22482
rect 37996 22418 38052 22430
rect 38444 23492 38500 23502
rect 38108 21810 38164 21822
rect 38108 21758 38110 21810
rect 38162 21758 38164 21810
rect 37996 21700 38052 21710
rect 38108 21700 38164 21758
rect 38052 21644 38164 21700
rect 37996 21634 38052 21644
rect 37324 19460 37380 19470
rect 37436 19460 37492 19740
rect 37380 19404 37492 19460
rect 37548 21532 37716 21588
rect 37324 19394 37380 19404
rect 37548 19348 37604 21532
rect 37660 21364 37716 21374
rect 37660 20802 37716 21308
rect 37660 20750 37662 20802
rect 37714 20750 37716 20802
rect 37660 20738 37716 20750
rect 37436 19292 37604 19348
rect 37884 20580 37940 20590
rect 37100 19124 37156 19134
rect 37100 17780 37156 19068
rect 37212 18338 37268 18350
rect 37212 18286 37214 18338
rect 37266 18286 37268 18338
rect 37212 18228 37268 18286
rect 37212 18162 37268 18172
rect 37324 17780 37380 17790
rect 37100 17778 37380 17780
rect 37100 17726 37326 17778
rect 37378 17726 37380 17778
rect 37100 17724 37380 17726
rect 37324 17714 37380 17724
rect 37436 15148 37492 19292
rect 37884 18676 37940 20524
rect 37996 20578 38052 20590
rect 37996 20526 37998 20578
rect 38050 20526 38052 20578
rect 37996 19460 38052 20526
rect 37996 19394 38052 19404
rect 38444 19236 38500 23436
rect 38556 22596 38612 23774
rect 38668 23716 38724 24668
rect 38668 23650 38724 23660
rect 38556 22540 39060 22596
rect 38780 21812 38836 21822
rect 38780 21718 38836 21756
rect 39004 21810 39060 22540
rect 39004 21758 39006 21810
rect 39058 21758 39060 21810
rect 39004 21746 39060 21758
rect 39116 21810 39172 25004
rect 39340 24724 39396 24734
rect 39340 24630 39396 24668
rect 39116 21758 39118 21810
rect 39170 21758 39172 21810
rect 38892 21586 38948 21598
rect 38892 21534 38894 21586
rect 38946 21534 38948 21586
rect 38892 21476 38948 21534
rect 39116 21588 39172 21758
rect 39340 22484 39396 22494
rect 39340 21698 39396 22428
rect 39340 21646 39342 21698
rect 39394 21646 39396 21698
rect 39340 21634 39396 21646
rect 39116 21522 39172 21532
rect 38892 21410 38948 21420
rect 39228 20916 39284 20926
rect 39228 20802 39284 20860
rect 39228 20750 39230 20802
rect 39282 20750 39284 20802
rect 39228 20738 39284 20750
rect 39340 20580 39396 20590
rect 39340 20486 39396 20524
rect 38444 19170 38500 19180
rect 38556 19460 38612 19470
rect 37996 19124 38052 19134
rect 37996 19030 38052 19068
rect 38220 19012 38276 19022
rect 38108 19010 38276 19012
rect 38108 18958 38222 19010
rect 38274 18958 38276 19010
rect 38108 18956 38276 18958
rect 38108 18676 38164 18956
rect 38220 18946 38276 18956
rect 38332 19010 38388 19022
rect 38332 18958 38334 19010
rect 38386 18958 38388 19010
rect 38332 18900 38388 18958
rect 38444 19012 38500 19022
rect 38444 18918 38500 18956
rect 38556 19010 38612 19404
rect 38556 18958 38558 19010
rect 38610 18958 38612 19010
rect 38332 18834 38388 18844
rect 38556 18788 38612 18958
rect 37772 18620 38164 18676
rect 38444 18732 38612 18788
rect 37548 18450 37604 18462
rect 37548 18398 37550 18450
rect 37602 18398 37604 18450
rect 37548 18228 37604 18398
rect 37548 18162 37604 18172
rect 37772 18450 37828 18620
rect 37772 18398 37774 18450
rect 37826 18398 37828 18450
rect 37660 16884 37716 16894
rect 36988 15092 37156 15148
rect 36092 12786 36148 12796
rect 35868 10770 35924 10780
rect 35196 10724 35252 10734
rect 35084 10722 35252 10724
rect 35084 10670 35198 10722
rect 35250 10670 35252 10722
rect 35084 10668 35252 10670
rect 35196 10658 35252 10668
rect 34524 10610 34692 10612
rect 34524 10558 34526 10610
rect 34578 10558 34692 10610
rect 34524 10556 34692 10558
rect 34524 10546 34580 10556
rect 31388 9774 31390 9826
rect 31442 9774 31444 9826
rect 30828 9662 30830 9714
rect 30882 9662 30884 9714
rect 30604 8034 30660 8046
rect 30604 7982 30606 8034
rect 30658 7982 30660 8034
rect 30604 7924 30660 7982
rect 30604 7858 30660 7868
rect 30828 7700 30884 9662
rect 30940 9716 30996 9726
rect 30940 9622 30996 9660
rect 31388 9268 31444 9774
rect 31388 9202 31444 9212
rect 31724 10500 31780 10510
rect 30268 7586 30548 7588
rect 30268 7534 30270 7586
rect 30322 7534 30548 7586
rect 30268 7532 30548 7534
rect 30604 7644 30884 7700
rect 30604 7586 30660 7644
rect 30604 7534 30606 7586
rect 30658 7534 30660 7586
rect 30268 7522 30324 7532
rect 30380 7364 30436 7374
rect 30380 7270 30436 7308
rect 30604 7028 30660 7534
rect 31724 7586 31780 10444
rect 32284 10500 32340 10510
rect 32284 10406 32340 10444
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 33964 9716 34020 9726
rect 33964 9622 34020 9660
rect 34300 9714 34356 9726
rect 36540 9716 36596 15092
rect 36988 14644 37044 14654
rect 36988 14550 37044 14588
rect 37100 13748 37156 15092
rect 37324 15092 37492 15148
rect 37548 16100 37604 16110
rect 37100 13692 37268 13748
rect 37100 13076 37156 13086
rect 37100 12982 37156 13020
rect 36988 12738 37044 12750
rect 36988 12686 36990 12738
rect 37042 12686 37044 12738
rect 36988 11956 37044 12686
rect 36988 11890 37044 11900
rect 34300 9662 34302 9714
rect 34354 9662 34356 9714
rect 34188 9604 34244 9614
rect 34076 9602 34244 9604
rect 34076 9550 34190 9602
rect 34242 9550 34244 9602
rect 34076 9548 34244 9550
rect 33292 8932 33348 8942
rect 33292 8838 33348 8876
rect 33964 8260 34020 8270
rect 33964 8166 34020 8204
rect 31724 7534 31726 7586
rect 31778 7534 31780 7586
rect 31724 7522 31780 7534
rect 33852 8146 33908 8158
rect 33852 8094 33854 8146
rect 33906 8094 33908 8146
rect 30828 7476 30884 7486
rect 30828 7382 30884 7420
rect 31612 7476 31668 7486
rect 31948 7476 32004 7486
rect 31164 7364 31220 7374
rect 31164 7270 31220 7308
rect 30044 5294 30046 5346
rect 30098 5294 30100 5346
rect 30044 5282 30100 5294
rect 30380 6972 30660 7028
rect 30716 7028 30772 7038
rect 29708 5124 29764 5134
rect 29708 5030 29764 5068
rect 30380 5124 30436 6972
rect 29260 4338 29316 4956
rect 30380 5010 30436 5068
rect 30716 5124 30772 6972
rect 31612 6804 31668 7420
rect 31836 7474 32004 7476
rect 31836 7422 31950 7474
rect 32002 7422 32004 7474
rect 31836 7420 32004 7422
rect 31836 7028 31892 7420
rect 31948 7410 32004 7420
rect 33852 7364 33908 8094
rect 34076 8148 34132 9548
rect 34188 9538 34244 9548
rect 34300 8932 34356 9662
rect 35644 9660 36596 9716
rect 35420 8932 35476 8942
rect 34188 8148 34244 8158
rect 34076 8146 34244 8148
rect 34076 8094 34190 8146
rect 34242 8094 34244 8146
rect 34076 8092 34244 8094
rect 34300 8148 34356 8876
rect 35084 8930 35476 8932
rect 35084 8878 35422 8930
rect 35474 8878 35476 8930
rect 35084 8876 35476 8878
rect 35084 8370 35140 8876
rect 35420 8866 35476 8876
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35084 8318 35086 8370
rect 35138 8318 35140 8370
rect 35084 8306 35140 8318
rect 34748 8260 34804 8270
rect 34748 8166 34804 8204
rect 34412 8148 34468 8158
rect 34300 8146 34468 8148
rect 34300 8094 34414 8146
rect 34466 8094 34468 8146
rect 34300 8092 34468 8094
rect 34188 7364 34244 8092
rect 34412 8036 34468 8092
rect 34412 7980 34804 8036
rect 34748 7476 34804 7980
rect 34972 8034 35028 8046
rect 34972 7982 34974 8034
rect 35026 7982 35028 8034
rect 34972 7924 35028 7982
rect 34860 7476 34916 7486
rect 34748 7474 34916 7476
rect 34748 7422 34862 7474
rect 34914 7422 34916 7474
rect 34748 7420 34916 7422
rect 34860 7410 34916 7420
rect 34636 7364 34692 7374
rect 34188 7362 34692 7364
rect 34188 7310 34638 7362
rect 34690 7310 34692 7362
rect 34188 7308 34692 7310
rect 31836 6962 31892 6972
rect 33740 7028 33796 7038
rect 32060 6804 32116 6814
rect 31612 6802 32116 6804
rect 31612 6750 32062 6802
rect 32114 6750 32116 6802
rect 31612 6748 32116 6750
rect 32060 6738 32116 6748
rect 33516 6692 33572 6702
rect 33516 5234 33572 6636
rect 33740 6020 33796 6972
rect 33852 6802 33908 7308
rect 33852 6750 33854 6802
rect 33906 6750 33908 6802
rect 33852 6738 33908 6750
rect 34636 6804 34692 7308
rect 34636 6738 34692 6748
rect 34300 6580 34356 6590
rect 34300 6578 34916 6580
rect 34300 6526 34302 6578
rect 34354 6526 34916 6578
rect 34300 6524 34916 6526
rect 34300 6514 34356 6524
rect 34636 6356 34692 6366
rect 34524 6300 34636 6356
rect 33852 6020 33908 6030
rect 33740 6018 33908 6020
rect 33740 5966 33854 6018
rect 33906 5966 33908 6018
rect 33740 5964 33908 5966
rect 33852 5954 33908 5964
rect 33516 5182 33518 5234
rect 33570 5182 33572 5234
rect 33516 5170 33572 5182
rect 34412 5906 34468 5918
rect 34412 5854 34414 5906
rect 34466 5854 34468 5906
rect 30716 5122 31556 5124
rect 30716 5070 30718 5122
rect 30770 5070 31556 5122
rect 30716 5068 31556 5070
rect 30716 5058 30772 5068
rect 30380 4958 30382 5010
rect 30434 4958 30436 5010
rect 30380 4946 30436 4958
rect 31500 5010 31556 5068
rect 31500 4958 31502 5010
rect 31554 4958 31556 5010
rect 31500 4946 31556 4958
rect 31836 5012 31892 5022
rect 31836 5010 32228 5012
rect 31836 4958 31838 5010
rect 31890 4958 32228 5010
rect 31836 4956 32228 4958
rect 31836 4946 31892 4956
rect 29932 4898 29988 4910
rect 29932 4846 29934 4898
rect 29986 4846 29988 4898
rect 29932 4452 29988 4846
rect 30044 4452 30100 4462
rect 29932 4450 30100 4452
rect 29932 4398 30046 4450
rect 30098 4398 30100 4450
rect 29932 4396 30100 4398
rect 30044 4386 30100 4396
rect 32172 4452 32228 4956
rect 33292 4564 33348 4574
rect 33292 4470 33348 4508
rect 34412 4564 34468 5854
rect 34524 5684 34580 6300
rect 34636 6290 34692 6300
rect 34860 6020 34916 6524
rect 34972 6356 35028 7868
rect 35644 7700 35700 9660
rect 36204 9044 36260 9054
rect 36540 9044 36596 9054
rect 36204 9042 36596 9044
rect 36204 8990 36206 9042
rect 36258 8990 36542 9042
rect 36594 8990 36596 9042
rect 36204 8988 36596 8990
rect 35644 7698 36148 7700
rect 35644 7646 35646 7698
rect 35698 7646 36148 7698
rect 35644 7644 36148 7646
rect 35644 7634 35700 7644
rect 35196 7252 35252 7262
rect 34972 6290 35028 6300
rect 35084 7250 35252 7252
rect 35084 7198 35198 7250
rect 35250 7198 35252 7250
rect 35084 7196 35252 7198
rect 35084 6690 35140 7196
rect 35196 7186 35252 7196
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35084 6638 35086 6690
rect 35138 6638 35140 6690
rect 34972 6020 35028 6030
rect 34860 6018 35028 6020
rect 34860 5966 34974 6018
rect 35026 5966 35028 6018
rect 34860 5964 35028 5966
rect 34972 5954 35028 5964
rect 34636 5906 34692 5918
rect 34636 5854 34638 5906
rect 34690 5854 34692 5906
rect 34636 5796 34692 5854
rect 35084 5796 35140 6638
rect 35308 6916 35364 6926
rect 35308 6578 35364 6860
rect 35980 6916 36036 6926
rect 35980 6690 36036 6860
rect 35980 6638 35982 6690
rect 36034 6638 36036 6690
rect 35980 6626 36036 6638
rect 35308 6526 35310 6578
rect 35362 6526 35364 6578
rect 35308 6514 35364 6526
rect 36092 6578 36148 7644
rect 36092 6526 36094 6578
rect 36146 6526 36148 6578
rect 36092 6514 36148 6526
rect 35196 6356 35252 6366
rect 35252 6300 35364 6356
rect 35196 6290 35252 6300
rect 35308 5906 35364 6300
rect 36204 6244 36260 8988
rect 36540 8978 36596 8988
rect 37212 7812 37268 13692
rect 37324 10612 37380 15092
rect 37548 13076 37604 16044
rect 37660 15988 37716 16828
rect 37660 15314 37716 15932
rect 37772 15876 37828 18398
rect 37996 18450 38052 18462
rect 37996 18398 37998 18450
rect 38050 18398 38052 18450
rect 37884 18338 37940 18350
rect 37884 18286 37886 18338
rect 37938 18286 37940 18338
rect 37884 17780 37940 18286
rect 37996 18340 38052 18398
rect 37996 18274 38052 18284
rect 38108 18450 38164 18462
rect 38108 18398 38110 18450
rect 38162 18398 38164 18450
rect 38108 17780 38164 18398
rect 38444 17780 38500 18732
rect 38556 18564 38612 18574
rect 38556 18470 38612 18508
rect 39116 18340 39172 18350
rect 39116 18246 39172 18284
rect 38668 18228 38724 18238
rect 38668 18226 39060 18228
rect 38668 18174 38670 18226
rect 38722 18174 39060 18226
rect 38668 18172 39060 18174
rect 38668 18162 38724 18172
rect 39004 18004 39060 18172
rect 39004 17948 39508 18004
rect 38108 17724 38500 17780
rect 37884 17714 37940 17724
rect 38332 16100 38388 16110
rect 38332 16006 38388 16044
rect 37772 15810 37828 15820
rect 37884 15986 37940 15998
rect 37884 15934 37886 15986
rect 37938 15934 37940 15986
rect 37660 15262 37662 15314
rect 37714 15262 37716 15314
rect 37660 15250 37716 15262
rect 37884 14644 37940 15934
rect 38108 15876 38164 15886
rect 38108 15782 38164 15820
rect 38220 15876 38276 15886
rect 38220 15874 38388 15876
rect 38220 15822 38222 15874
rect 38274 15822 38388 15874
rect 38220 15820 38388 15822
rect 38220 15810 38276 15820
rect 38332 15428 38388 15820
rect 38444 15874 38500 17724
rect 39452 17778 39508 17948
rect 39452 17726 39454 17778
rect 39506 17726 39508 17778
rect 39452 17714 39508 17726
rect 38444 15822 38446 15874
rect 38498 15822 38500 15874
rect 38444 15764 38500 15822
rect 38444 15698 38500 15708
rect 38444 15428 38500 15438
rect 38332 15426 38500 15428
rect 38332 15374 38446 15426
rect 38498 15374 38500 15426
rect 38332 15372 38500 15374
rect 38444 15362 38500 15372
rect 38556 15092 38612 15102
rect 38556 15090 39172 15092
rect 38556 15038 38558 15090
rect 38610 15038 39172 15090
rect 38556 15036 39172 15038
rect 38556 15026 38612 15036
rect 37772 13860 37828 13870
rect 37884 13860 37940 14588
rect 39116 14642 39172 15036
rect 39116 14590 39118 14642
rect 39170 14590 39172 14642
rect 39116 14578 39172 14590
rect 37772 13858 37940 13860
rect 37772 13806 37774 13858
rect 37826 13806 37940 13858
rect 37772 13804 37940 13806
rect 37996 14420 38052 14430
rect 37772 13794 37828 13804
rect 37996 13746 38052 14364
rect 37996 13694 37998 13746
rect 38050 13694 38052 13746
rect 37996 13682 38052 13694
rect 37884 13188 37940 13198
rect 37884 13094 37940 13132
rect 39116 13188 39172 13198
rect 37660 13076 37716 13086
rect 37548 13020 37660 13076
rect 37660 12982 37716 13020
rect 38668 13076 38724 13086
rect 38668 12982 38724 13020
rect 39116 13074 39172 13132
rect 39116 13022 39118 13074
rect 39170 13022 39172 13074
rect 38220 12738 38276 12750
rect 38220 12686 38222 12738
rect 38274 12686 38276 12738
rect 37996 12180 38052 12190
rect 37996 11506 38052 12124
rect 38220 11844 38276 12686
rect 38220 11778 38276 11788
rect 37996 11454 37998 11506
rect 38050 11454 38052 11506
rect 37996 11442 38052 11454
rect 38220 11172 38276 11182
rect 37436 10836 37492 10846
rect 37436 10742 37492 10780
rect 38220 10834 38276 11116
rect 38220 10782 38222 10834
rect 38274 10782 38276 10834
rect 38220 10770 38276 10782
rect 39004 11172 39060 11182
rect 37324 10546 37380 10556
rect 37996 10612 38052 10622
rect 37996 9940 38052 10556
rect 39004 10610 39060 11116
rect 39004 10558 39006 10610
rect 39058 10558 39060 10610
rect 39004 10546 39060 10558
rect 39116 9940 39172 13022
rect 37996 9938 38388 9940
rect 37996 9886 37998 9938
rect 38050 9886 38388 9938
rect 37996 9884 38388 9886
rect 37996 9874 38052 9884
rect 37660 9828 37716 9838
rect 37660 9734 37716 9772
rect 38332 9826 38388 9884
rect 39116 9874 39172 9884
rect 39228 11956 39284 11966
rect 38332 9774 38334 9826
rect 38386 9774 38388 9826
rect 38332 9762 38388 9774
rect 39228 9828 39284 11900
rect 39340 10612 39396 10622
rect 39340 10518 39396 10556
rect 39228 9734 39284 9772
rect 39452 10386 39508 10398
rect 39452 10334 39454 10386
rect 39506 10334 39508 10386
rect 39452 9826 39508 10334
rect 39564 10052 39620 25228
rect 39676 24948 39732 24958
rect 39676 24722 39732 24892
rect 40012 24946 40068 26124
rect 40348 25284 40404 25294
rect 40012 24894 40014 24946
rect 40066 24894 40068 24946
rect 40012 24882 40068 24894
rect 40124 25060 40180 25070
rect 40124 24946 40180 25004
rect 40124 24894 40126 24946
rect 40178 24894 40180 24946
rect 40124 24882 40180 24894
rect 40348 24834 40404 25228
rect 40348 24782 40350 24834
rect 40402 24782 40404 24834
rect 40348 24770 40404 24782
rect 39676 24670 39678 24722
rect 39730 24670 39732 24722
rect 39676 21812 39732 24670
rect 39900 24724 39956 24734
rect 39900 24630 39956 24668
rect 39788 23154 39844 23166
rect 39788 23102 39790 23154
rect 39842 23102 39844 23154
rect 39788 23044 39844 23102
rect 40236 23044 40292 23054
rect 39788 23042 40292 23044
rect 39788 22990 40238 23042
rect 40290 22990 40292 23042
rect 39788 22988 40292 22990
rect 39676 21746 39732 21756
rect 39788 21476 39844 21486
rect 39788 21382 39844 21420
rect 39788 20916 39844 20926
rect 39788 20822 39844 20860
rect 39900 14532 39956 14542
rect 39900 14438 39956 14476
rect 40012 13412 40068 22988
rect 40236 22978 40292 22988
rect 40124 22820 40180 22830
rect 40124 22484 40180 22764
rect 40124 22390 40180 22428
rect 40460 19908 40516 32060
rect 40908 32116 40964 34636
rect 41468 34626 41524 34636
rect 41580 34356 41636 34860
rect 40908 32050 40964 32060
rect 41132 34300 41636 34356
rect 41132 31780 41188 34300
rect 41580 34132 41636 34142
rect 41692 34132 41748 35084
rect 41804 34804 41860 35758
rect 41804 34738 41860 34748
rect 41916 34914 41972 34926
rect 41916 34862 41918 34914
rect 41970 34862 41972 34914
rect 41244 34130 41748 34132
rect 41244 34078 41582 34130
rect 41634 34078 41748 34130
rect 41244 34076 41748 34078
rect 41804 34356 41860 34366
rect 41916 34356 41972 34862
rect 41804 34354 41972 34356
rect 41804 34302 41806 34354
rect 41858 34302 41972 34354
rect 41804 34300 41972 34302
rect 41244 33124 41300 34076
rect 41580 34066 41636 34076
rect 41804 33572 41860 34300
rect 41692 33516 41860 33572
rect 41244 33058 41300 33068
rect 41356 33460 41412 33470
rect 41356 32674 41412 33404
rect 41356 32622 41358 32674
rect 41410 32622 41412 32674
rect 41356 32610 41412 32622
rect 41692 33348 41748 33516
rect 41916 33460 41972 33498
rect 41916 33394 41972 33404
rect 41804 33348 41860 33358
rect 41692 33346 41860 33348
rect 41692 33294 41806 33346
rect 41858 33294 41860 33346
rect 41692 33292 41860 33294
rect 41468 32452 41524 32462
rect 41468 32358 41524 32396
rect 41132 31714 41188 31724
rect 41580 31668 41636 31678
rect 40348 19012 40404 19022
rect 39900 13356 40012 13412
rect 39900 13076 39956 13356
rect 40012 13346 40068 13356
rect 40124 18340 40180 18350
rect 39676 13074 39956 13076
rect 39676 13022 39902 13074
rect 39954 13022 39956 13074
rect 39676 13020 39956 13022
rect 39676 12178 39732 13020
rect 39900 13010 39956 13020
rect 40124 12740 40180 18284
rect 40236 17666 40292 17678
rect 40236 17614 40238 17666
rect 40290 17614 40292 17666
rect 40236 14532 40292 17614
rect 40236 14466 40292 14476
rect 40348 13748 40404 18956
rect 40460 18676 40516 19852
rect 40460 18450 40516 18620
rect 40460 18398 40462 18450
rect 40514 18398 40516 18450
rect 40460 18386 40516 18398
rect 40684 31220 40740 31230
rect 40684 20916 40740 31164
rect 41356 31220 41412 31230
rect 41356 31126 41412 31164
rect 41580 31218 41636 31612
rect 41580 31166 41582 31218
rect 41634 31166 41636 31218
rect 41580 31154 41636 31166
rect 41692 31220 41748 33292
rect 41804 33282 41860 33292
rect 42028 33348 42084 37214
rect 42588 37268 42644 37278
rect 42588 37266 42756 37268
rect 42588 37214 42590 37266
rect 42642 37214 42756 37266
rect 42588 37212 42756 37214
rect 42588 37202 42644 37212
rect 42700 37156 42756 37212
rect 43036 37156 43092 37166
rect 42700 37154 43092 37156
rect 42700 37102 43038 37154
rect 43090 37102 43092 37154
rect 42700 37100 43092 37102
rect 42476 36482 42532 36494
rect 42476 36430 42478 36482
rect 42530 36430 42532 36482
rect 42140 36260 42196 36270
rect 42140 36258 42308 36260
rect 42140 36206 42142 36258
rect 42194 36206 42308 36258
rect 42140 36204 42308 36206
rect 42140 36194 42196 36204
rect 42140 35700 42196 35710
rect 42140 35606 42196 35644
rect 42252 35588 42308 36204
rect 42364 35588 42420 35598
rect 42252 35532 42364 35588
rect 42364 35522 42420 35532
rect 42140 35028 42196 35038
rect 42140 34914 42196 34972
rect 42140 34862 42142 34914
rect 42194 34862 42196 34914
rect 42140 34850 42196 34862
rect 42364 34804 42420 34814
rect 42252 34692 42308 34702
rect 42252 34598 42308 34636
rect 42028 33254 42084 33292
rect 42140 34580 42196 34590
rect 42140 33124 42196 34524
rect 42252 33348 42308 33358
rect 42364 33348 42420 34748
rect 42476 33460 42532 36430
rect 42700 36372 42756 37100
rect 43036 37090 43092 37100
rect 43372 36596 43428 36606
rect 43372 36502 43428 36540
rect 42588 35588 42644 35598
rect 42588 35494 42644 35532
rect 42588 34804 42644 34814
rect 42588 34710 42644 34748
rect 42588 34580 42644 34590
rect 42700 34580 42756 36316
rect 43036 36260 43092 36270
rect 43036 35476 43092 36204
rect 43260 35586 43316 35598
rect 43260 35534 43262 35586
rect 43314 35534 43316 35586
rect 43260 35476 43316 35534
rect 42924 35420 43316 35476
rect 43372 35588 43428 35598
rect 42924 35308 42980 35420
rect 42924 35252 43092 35308
rect 42644 34524 42756 34580
rect 42588 34514 42644 34524
rect 42476 33404 42644 33460
rect 42252 33346 42420 33348
rect 42252 33294 42254 33346
rect 42306 33294 42420 33346
rect 42252 33292 42420 33294
rect 42252 33282 42308 33292
rect 42140 33068 42308 33124
rect 41804 32562 41860 32574
rect 41804 32510 41806 32562
rect 41858 32510 41860 32562
rect 41804 31892 41860 32510
rect 41804 31798 41860 31836
rect 41692 31218 42196 31220
rect 41692 31166 41694 31218
rect 41746 31166 42196 31218
rect 41692 31164 42196 31166
rect 41692 31154 41748 31164
rect 41132 30996 41188 31006
rect 41132 30902 41188 30940
rect 42140 30994 42196 31164
rect 42140 30942 42142 30994
rect 42194 30942 42196 30994
rect 42140 30930 42196 30942
rect 40908 30884 40964 30894
rect 40908 30210 40964 30828
rect 41468 30882 41524 30894
rect 41468 30830 41470 30882
rect 41522 30830 41524 30882
rect 41468 30324 41524 30830
rect 41468 30258 41524 30268
rect 41916 30434 41972 30446
rect 41916 30382 41918 30434
rect 41970 30382 41972 30434
rect 40908 30158 40910 30210
rect 40962 30158 40964 30210
rect 40908 30146 40964 30158
rect 41916 30210 41972 30382
rect 41916 30158 41918 30210
rect 41970 30158 41972 30210
rect 41916 30146 41972 30158
rect 40796 29988 40852 29998
rect 40796 29894 40852 29932
rect 42028 28756 42084 28766
rect 42028 28662 42084 28700
rect 41020 27860 41076 27870
rect 41020 27858 41188 27860
rect 41020 27806 41022 27858
rect 41074 27806 41188 27858
rect 41020 27804 41188 27806
rect 41020 27794 41076 27804
rect 41132 26908 41188 27804
rect 41692 27748 41748 27758
rect 41692 27654 41748 27692
rect 41020 26852 41188 26908
rect 41020 26786 41076 26796
rect 41132 26402 41188 26852
rect 41132 26350 41134 26402
rect 41186 26350 41188 26402
rect 40908 25060 40964 25070
rect 40964 25004 41076 25060
rect 40908 24994 40964 25004
rect 40796 24948 40852 24958
rect 40796 23938 40852 24892
rect 41020 24052 41076 25004
rect 41132 24724 41188 26350
rect 41468 25618 41524 25630
rect 41468 25566 41470 25618
rect 41522 25566 41524 25618
rect 41468 25284 41524 25566
rect 41468 25218 41524 25228
rect 41132 24722 41412 24724
rect 41132 24670 41134 24722
rect 41186 24670 41412 24722
rect 41132 24668 41412 24670
rect 41132 24658 41188 24668
rect 41020 23996 41300 24052
rect 40796 23886 40798 23938
rect 40850 23886 40852 23938
rect 40796 23874 40852 23886
rect 41244 23938 41300 23996
rect 41244 23886 41246 23938
rect 41298 23886 41300 23938
rect 41244 23874 41300 23886
rect 41132 23828 41188 23838
rect 41132 23734 41188 23772
rect 41020 23714 41076 23726
rect 41020 23662 41022 23714
rect 41074 23662 41076 23714
rect 40908 21812 40964 21822
rect 40908 21586 40964 21756
rect 40908 21534 40910 21586
rect 40962 21534 40964 21586
rect 40908 21522 40964 21534
rect 40684 19346 40740 20860
rect 40684 19294 40686 19346
rect 40738 19294 40740 19346
rect 40684 18452 40740 19294
rect 41020 20356 41076 23662
rect 41356 22370 41412 24668
rect 41804 24610 41860 24622
rect 41804 24558 41806 24610
rect 41858 24558 41860 24610
rect 41468 24500 41524 24510
rect 41468 23938 41524 24444
rect 41804 24162 41860 24558
rect 41804 24110 41806 24162
rect 41858 24110 41860 24162
rect 41804 24098 41860 24110
rect 41468 23886 41470 23938
rect 41522 23886 41524 23938
rect 41468 23874 41524 23886
rect 41692 23828 41748 23838
rect 41916 23828 41972 23838
rect 41748 23826 41972 23828
rect 41748 23774 41918 23826
rect 41970 23774 41972 23826
rect 41748 23772 41972 23774
rect 41692 23762 41748 23772
rect 41916 23762 41972 23772
rect 41916 23044 41972 23054
rect 41356 22318 41358 22370
rect 41410 22318 41412 22370
rect 41356 22306 41412 22318
rect 41468 23042 41972 23044
rect 41468 22990 41918 23042
rect 41970 22990 41972 23042
rect 41468 22988 41972 22990
rect 41244 21812 41300 21822
rect 41468 21812 41524 22988
rect 41916 22978 41972 22988
rect 42028 22932 42084 22942
rect 42028 22930 42196 22932
rect 42028 22878 42030 22930
rect 42082 22878 42196 22930
rect 42028 22876 42196 22878
rect 42028 22866 42084 22876
rect 41244 21810 41524 21812
rect 41244 21758 41246 21810
rect 41298 21758 41524 21810
rect 41244 21756 41524 21758
rect 41580 22484 41636 22494
rect 41244 21746 41300 21756
rect 41580 21698 41636 22428
rect 42140 22482 42196 22876
rect 42140 22430 42142 22482
rect 42194 22430 42196 22482
rect 42140 22418 42196 22430
rect 41580 21646 41582 21698
rect 41634 21646 41636 21698
rect 41580 21634 41636 21646
rect 42252 21700 42308 33068
rect 42364 32228 42420 33292
rect 42476 33236 42532 33246
rect 42476 33142 42532 33180
rect 42588 32676 42644 33404
rect 42700 33348 42756 33358
rect 42924 33348 42980 33358
rect 42756 33346 42980 33348
rect 42756 33294 42926 33346
rect 42978 33294 42980 33346
rect 42756 33292 42980 33294
rect 42700 33282 42756 33292
rect 42924 33282 42980 33292
rect 42588 32620 42756 32676
rect 42588 32452 42644 32462
rect 42588 32358 42644 32396
rect 42364 32172 42644 32228
rect 42364 31780 42420 31790
rect 42364 31218 42420 31724
rect 42364 31166 42366 31218
rect 42418 31166 42420 31218
rect 42364 30434 42420 31166
rect 42588 31220 42644 32172
rect 42588 31126 42644 31164
rect 42700 31668 42756 32620
rect 42476 30884 42532 30894
rect 42476 30790 42532 30828
rect 42364 30382 42366 30434
rect 42418 30382 42420 30434
rect 42364 30370 42420 30382
rect 42700 30324 42756 31612
rect 42476 30268 42756 30324
rect 42812 30994 42868 31006
rect 42812 30942 42814 30994
rect 42866 30942 42868 30994
rect 42364 30100 42420 30110
rect 42476 30100 42532 30268
rect 42364 30098 42532 30100
rect 42364 30046 42366 30098
rect 42418 30046 42532 30098
rect 42364 30044 42532 30046
rect 42364 30034 42420 30044
rect 42812 28756 42868 30942
rect 42812 28690 42868 28700
rect 43036 28532 43092 35252
rect 43260 34916 43316 34954
rect 43260 34850 43316 34860
rect 43148 34802 43204 34814
rect 43148 34750 43150 34802
rect 43202 34750 43204 34802
rect 43148 34692 43204 34750
rect 43148 34626 43204 34636
rect 43372 34468 43428 35532
rect 42700 28476 43092 28532
rect 43148 34412 43428 34468
rect 42588 27636 42644 27646
rect 42476 21700 42532 21710
rect 42252 21644 42476 21700
rect 41132 21586 41188 21598
rect 41132 21534 41134 21586
rect 41186 21534 41188 21586
rect 41132 20580 41188 21534
rect 41356 21588 41412 21598
rect 41356 21494 41412 21532
rect 42476 21586 42532 21644
rect 42476 21534 42478 21586
rect 42530 21534 42532 21586
rect 42476 21522 42532 21534
rect 42588 20804 42644 27580
rect 42140 20748 42644 20804
rect 41916 20580 41972 20590
rect 41132 20578 41972 20580
rect 41132 20526 41918 20578
rect 41970 20526 41972 20578
rect 41132 20524 41972 20526
rect 41020 20300 41636 20356
rect 41020 19012 41076 20300
rect 41580 20130 41636 20300
rect 41580 20078 41582 20130
rect 41634 20078 41636 20130
rect 41580 20066 41636 20078
rect 41020 18946 41076 18956
rect 41244 19012 41300 19022
rect 41580 19012 41636 19022
rect 41244 19010 41636 19012
rect 41244 18958 41246 19010
rect 41298 18958 41582 19010
rect 41634 18958 41636 19010
rect 41244 18956 41636 18958
rect 40684 18386 40740 18396
rect 41244 18450 41300 18956
rect 41244 18398 41246 18450
rect 41298 18398 41300 18450
rect 41244 18386 41300 18398
rect 41020 17780 41076 17790
rect 40908 17668 40964 17678
rect 41020 17668 41076 17724
rect 41468 17668 41524 18956
rect 41580 18946 41636 18956
rect 41692 18452 41748 18462
rect 41692 18358 41748 18396
rect 41804 18116 41860 20524
rect 41916 20514 41972 20524
rect 41916 20132 41972 20142
rect 41916 20038 41972 20076
rect 42140 19572 42196 20748
rect 42252 20578 42308 20590
rect 42252 20526 42254 20578
rect 42306 20526 42308 20578
rect 42252 20356 42308 20526
rect 42700 20578 42756 28476
rect 42924 25396 42980 25406
rect 42700 20526 42702 20578
rect 42754 20526 42756 20578
rect 42700 20356 42756 20526
rect 42252 20300 42756 20356
rect 42364 20132 42420 20142
rect 42364 20038 42420 20076
rect 42588 19796 42644 19806
rect 42140 19516 42420 19572
rect 42140 19348 42196 19358
rect 42140 19254 42196 19292
rect 41916 18676 41972 18686
rect 41916 18452 41972 18620
rect 42252 18676 42308 18686
rect 42028 18452 42084 18462
rect 41916 18450 42084 18452
rect 41916 18398 42030 18450
rect 42082 18398 42084 18450
rect 41916 18396 42084 18398
rect 42028 18386 42084 18396
rect 42252 18450 42308 18620
rect 42252 18398 42254 18450
rect 42306 18398 42308 18450
rect 42252 18386 42308 18398
rect 42364 18452 42420 19516
rect 42588 19346 42644 19740
rect 42700 19684 42756 20300
rect 42812 25340 42924 25396
rect 42812 20130 42868 25340
rect 42924 25302 42980 25340
rect 42812 20078 42814 20130
rect 42866 20078 42868 20130
rect 42812 19908 42868 20078
rect 42924 21476 42980 21486
rect 42924 20020 42980 21420
rect 43148 20132 43204 34412
rect 43260 34132 43316 34142
rect 43484 34132 43540 37324
rect 43260 34130 43540 34132
rect 43260 34078 43262 34130
rect 43314 34078 43540 34130
rect 43260 34076 43540 34078
rect 43260 34066 43316 34076
rect 43484 28756 43540 28766
rect 43484 28662 43540 28700
rect 43708 28084 43764 38110
rect 43820 38388 43876 38782
rect 43932 38836 43988 39004
rect 43932 38770 43988 38780
rect 44716 39228 44996 39284
rect 45052 41186 45220 41188
rect 45052 41134 45166 41186
rect 45218 41134 45220 41186
rect 45052 41132 45220 41134
rect 43820 37380 43876 38332
rect 44268 38164 44324 38174
rect 44268 38070 44324 38108
rect 43820 37314 43876 37324
rect 44716 36596 44772 39228
rect 45052 38388 45108 41132
rect 45164 41122 45220 41132
rect 45724 40964 45780 42476
rect 45948 42466 46004 42476
rect 46060 42420 46116 42476
rect 46284 42420 46340 42702
rect 46060 42364 46340 42420
rect 46956 42754 47012 42766
rect 46956 42702 46958 42754
rect 47010 42702 47012 42754
rect 45948 41076 46004 41086
rect 45164 40404 45220 40414
rect 45500 40404 45556 40414
rect 45164 40402 45556 40404
rect 45164 40350 45166 40402
rect 45218 40350 45502 40402
rect 45554 40350 45556 40402
rect 45164 40348 45556 40350
rect 45164 40338 45220 40348
rect 45500 40338 45556 40348
rect 45612 40404 45668 40414
rect 45724 40404 45780 40908
rect 45836 41074 46004 41076
rect 45836 41022 45950 41074
rect 46002 41022 46004 41074
rect 45836 41020 46004 41022
rect 45836 40514 45892 41020
rect 45948 41010 46004 41020
rect 45836 40462 45838 40514
rect 45890 40462 45892 40514
rect 45836 40450 45892 40462
rect 45612 40402 45780 40404
rect 45612 40350 45614 40402
rect 45666 40350 45780 40402
rect 45612 40348 45780 40350
rect 46060 40404 46116 40414
rect 45388 39844 45444 39854
rect 45612 39844 45668 40348
rect 46060 40310 46116 40348
rect 46284 40292 46340 40302
rect 46284 40198 46340 40236
rect 46620 40292 46676 40302
rect 45444 39788 45668 39844
rect 45388 39730 45444 39788
rect 45388 39678 45390 39730
rect 45442 39678 45444 39730
rect 45388 39666 45444 39678
rect 45388 39060 45444 39070
rect 45388 39058 46004 39060
rect 45388 39006 45390 39058
rect 45442 39006 46004 39058
rect 45388 39004 46004 39006
rect 45388 38994 45444 39004
rect 45724 38836 45780 38846
rect 45724 38742 45780 38780
rect 45948 38834 46004 39004
rect 46620 39058 46676 40236
rect 46956 40292 47012 42702
rect 49756 42756 49812 42766
rect 47852 42252 48132 42308
rect 47852 42196 47908 42252
rect 47516 42140 47908 42196
rect 48076 42194 48132 42252
rect 48076 42142 48078 42194
rect 48130 42142 48132 42194
rect 47516 42084 47572 42140
rect 48076 42130 48132 42142
rect 47404 42028 47572 42084
rect 47964 42084 48020 42094
rect 46956 40226 47012 40236
rect 47180 41860 47236 41870
rect 47404 41860 47460 42028
rect 47964 41990 48020 42028
rect 47628 41972 47684 41982
rect 48972 41972 49028 41982
rect 47628 41970 47908 41972
rect 47628 41918 47630 41970
rect 47682 41918 47908 41970
rect 47628 41916 47908 41918
rect 47628 41906 47684 41916
rect 47180 41858 47460 41860
rect 47180 41806 47182 41858
rect 47234 41806 47460 41858
rect 47180 41804 47460 41806
rect 47516 41860 47572 41870
rect 46620 39006 46622 39058
rect 46674 39006 46676 39058
rect 46620 38948 46676 39006
rect 46620 38882 46676 38892
rect 46844 39060 46900 39070
rect 45948 38782 45950 38834
rect 46002 38782 46004 38834
rect 45836 38722 45892 38734
rect 45836 38670 45838 38722
rect 45890 38670 45892 38722
rect 45836 38668 45892 38670
rect 45052 38162 45108 38332
rect 45052 38110 45054 38162
rect 45106 38110 45108 38162
rect 45052 38098 45108 38110
rect 45612 38612 45892 38668
rect 45948 38668 46004 38782
rect 46284 38836 46340 38846
rect 46284 38742 46340 38780
rect 46844 38834 46900 39004
rect 46844 38782 46846 38834
rect 46898 38782 46900 38834
rect 46844 38770 46900 38782
rect 45948 38612 46116 38668
rect 45612 37378 45668 38612
rect 45612 37326 45614 37378
rect 45666 37326 45668 37378
rect 45612 37314 45668 37326
rect 45948 37828 46004 37838
rect 44940 37266 44996 37278
rect 44940 37214 44942 37266
rect 44994 37214 44996 37266
rect 44716 36530 44772 36540
rect 44828 36708 44884 36718
rect 44828 36594 44884 36652
rect 44828 36542 44830 36594
rect 44882 36542 44884 36594
rect 44828 36530 44884 36542
rect 43820 36482 43876 36494
rect 43820 36430 43822 36482
rect 43874 36430 43876 36482
rect 43820 36260 43876 36430
rect 44940 36484 44996 37214
rect 45948 36594 46004 37772
rect 45948 36542 45950 36594
rect 46002 36542 46004 36594
rect 45948 36530 46004 36542
rect 43876 36204 44212 36260
rect 43820 36194 43876 36204
rect 44156 35922 44212 36204
rect 44156 35870 44158 35922
rect 44210 35870 44212 35922
rect 44156 35858 44212 35870
rect 43932 34916 43988 34926
rect 43932 34242 43988 34860
rect 43932 34190 43934 34242
rect 43986 34190 43988 34242
rect 43932 34178 43988 34190
rect 44716 33236 44772 33246
rect 44716 32452 44772 33180
rect 44716 32358 44772 32396
rect 44940 33236 44996 36428
rect 45276 36482 45332 36494
rect 45276 36430 45278 36482
rect 45330 36430 45332 36482
rect 45276 35588 45332 36430
rect 45612 35588 45668 35598
rect 45332 35586 45668 35588
rect 45332 35534 45614 35586
rect 45666 35534 45668 35586
rect 45332 35532 45668 35534
rect 45276 35522 45332 35532
rect 45612 35522 45668 35532
rect 46060 35028 46116 38612
rect 47180 37828 47236 41804
rect 47516 41746 47572 41804
rect 47516 41694 47518 41746
rect 47570 41694 47572 41746
rect 47516 40404 47572 41694
rect 47852 41412 47908 41916
rect 48972 41878 49028 41916
rect 49644 41860 49700 41870
rect 49420 41858 49700 41860
rect 49420 41806 49646 41858
rect 49698 41806 49700 41858
rect 49420 41804 49700 41806
rect 48076 41748 48132 41758
rect 48076 41654 48132 41692
rect 49084 41748 49140 41758
rect 47852 41356 48132 41412
rect 48076 41298 48132 41356
rect 49084 41410 49140 41692
rect 49084 41358 49086 41410
rect 49138 41358 49140 41410
rect 49084 41346 49140 41358
rect 48076 41246 48078 41298
rect 48130 41246 48132 41298
rect 48076 41234 48132 41246
rect 49420 41298 49476 41804
rect 49644 41794 49700 41804
rect 49644 41412 49700 41422
rect 49756 41412 49812 42700
rect 49644 41410 49812 41412
rect 49644 41358 49646 41410
rect 49698 41358 49812 41410
rect 49644 41356 49812 41358
rect 49644 41346 49700 41356
rect 49420 41246 49422 41298
rect 49474 41246 49476 41298
rect 49420 41234 49476 41246
rect 49868 41188 49924 41198
rect 49756 41186 49924 41188
rect 49756 41134 49870 41186
rect 49922 41134 49924 41186
rect 49756 41132 49924 41134
rect 49308 41074 49364 41086
rect 49308 41022 49310 41074
rect 49362 41022 49364 41074
rect 48748 40964 48804 40974
rect 48748 40870 48804 40908
rect 49308 40964 49364 41022
rect 49308 40898 49364 40908
rect 49756 40626 49812 41132
rect 49868 41122 49924 41132
rect 49756 40574 49758 40626
rect 49810 40574 49812 40626
rect 49420 40404 49476 40414
rect 47516 40338 47572 40348
rect 49308 40402 49476 40404
rect 49308 40350 49422 40402
rect 49474 40350 49476 40402
rect 49308 40348 49476 40350
rect 48748 39844 48804 39854
rect 48524 39506 48580 39518
rect 48524 39454 48526 39506
rect 48578 39454 48580 39506
rect 47404 39394 47460 39406
rect 47404 39342 47406 39394
rect 47458 39342 47460 39394
rect 47404 38500 47460 39342
rect 48524 39396 48580 39454
rect 48636 39396 48692 39406
rect 48524 39394 48692 39396
rect 48524 39342 48638 39394
rect 48690 39342 48692 39394
rect 48524 39340 48692 39342
rect 48636 39330 48692 39340
rect 47852 39284 47908 39294
rect 47516 38948 47572 38958
rect 47516 38834 47572 38892
rect 47516 38782 47518 38834
rect 47570 38782 47572 38834
rect 47516 38770 47572 38782
rect 47740 38724 47796 38734
rect 47740 38630 47796 38668
rect 47404 38434 47460 38444
rect 47180 37762 47236 37772
rect 47740 37156 47796 37166
rect 47852 37156 47908 39228
rect 48748 39284 48804 39788
rect 48860 39394 48916 39406
rect 48860 39342 48862 39394
rect 48914 39342 48916 39394
rect 48860 39284 48916 39342
rect 49084 39396 49140 39406
rect 49308 39396 49364 40348
rect 49420 40338 49476 40348
rect 49756 40292 49812 40574
rect 49756 40226 49812 40236
rect 49980 39844 50036 44940
rect 50092 43652 50148 45054
rect 50204 44324 50260 45276
rect 50204 44258 50260 44268
rect 50092 43586 50148 43596
rect 50316 43426 50372 45276
rect 50876 45332 50932 46622
rect 50876 45266 50932 45276
rect 50988 45220 51044 48188
rect 50988 45154 51044 45164
rect 51100 47572 51156 47582
rect 51100 45106 51156 47516
rect 51324 45892 51380 45902
rect 51100 45054 51102 45106
rect 51154 45054 51156 45106
rect 51100 44996 51156 45054
rect 50540 44940 51156 44996
rect 51212 45890 51380 45892
rect 51212 45838 51326 45890
rect 51378 45838 51380 45890
rect 51212 45836 51380 45838
rect 50316 43374 50318 43426
rect 50370 43374 50372 43426
rect 50316 43362 50372 43374
rect 50428 44436 50484 44446
rect 50540 44436 50596 44940
rect 50484 44434 50596 44436
rect 50484 44382 50542 44434
rect 50594 44382 50596 44434
rect 50484 44380 50596 44382
rect 49980 39778 50036 39788
rect 50092 40516 50148 40526
rect 49084 39394 49364 39396
rect 49084 39342 49086 39394
rect 49138 39342 49364 39394
rect 49084 39340 49364 39342
rect 49420 39396 49476 39406
rect 48860 39228 49028 39284
rect 47964 38834 48020 38846
rect 47964 38782 47966 38834
rect 48018 38782 48020 38834
rect 47964 38500 48020 38782
rect 47964 38434 48020 38444
rect 48188 38834 48244 38846
rect 48188 38782 48190 38834
rect 48242 38782 48244 38834
rect 48188 37492 48244 38782
rect 48748 38834 48804 39228
rect 48748 38782 48750 38834
rect 48802 38782 48804 38834
rect 48748 38770 48804 38782
rect 48860 38836 48916 38846
rect 48860 38742 48916 38780
rect 48972 38834 49028 39228
rect 49084 39060 49140 39340
rect 49084 38994 49140 39004
rect 48972 38782 48974 38834
rect 49026 38782 49028 38834
rect 48748 38052 48804 38062
rect 48188 37426 48244 37436
rect 48636 37996 48748 38052
rect 47740 37154 47908 37156
rect 47740 37102 47742 37154
rect 47794 37102 47908 37154
rect 47740 37100 47908 37102
rect 48188 37156 48244 37166
rect 48300 37156 48356 37166
rect 48188 37154 48300 37156
rect 48188 37102 48190 37154
rect 48242 37102 48300 37154
rect 48188 37100 48300 37102
rect 47740 37090 47796 37100
rect 48188 37090 48244 37100
rect 46284 36482 46340 36494
rect 46284 36430 46286 36482
rect 46338 36430 46340 36482
rect 46284 36372 46340 36430
rect 46284 36306 46340 36316
rect 46844 36372 46900 36382
rect 46844 36278 46900 36316
rect 47180 36260 47236 36270
rect 47180 35922 47236 36204
rect 47180 35870 47182 35922
rect 47234 35870 47236 35922
rect 47180 35858 47236 35870
rect 47852 35810 47908 35822
rect 47852 35758 47854 35810
rect 47906 35758 47908 35810
rect 46844 35698 46900 35710
rect 46844 35646 46846 35698
rect 46898 35646 46900 35698
rect 46844 35140 46900 35646
rect 47516 35700 47572 35710
rect 47516 35606 47572 35644
rect 47852 35364 47908 35758
rect 47852 35298 47908 35308
rect 46844 35074 46900 35084
rect 43820 31780 43876 31790
rect 44380 31780 44436 31790
rect 43820 31778 44380 31780
rect 43820 31726 43822 31778
rect 43874 31726 44380 31778
rect 43820 31724 44380 31726
rect 43820 31714 43876 31724
rect 44380 31686 44436 31724
rect 44940 31778 44996 33180
rect 45948 34972 46116 35028
rect 44940 31726 44942 31778
rect 44994 31726 44996 31778
rect 44940 31714 44996 31726
rect 45836 31892 45892 31902
rect 45612 31668 45668 31678
rect 45500 31666 45668 31668
rect 45500 31614 45614 31666
rect 45666 31614 45668 31666
rect 45500 31612 45668 31614
rect 45500 31106 45556 31612
rect 45612 31602 45668 31612
rect 45500 31054 45502 31106
rect 45554 31054 45556 31106
rect 45500 31042 45556 31054
rect 45836 30994 45892 31836
rect 45948 31108 46004 34972
rect 46060 34804 46116 34814
rect 46060 34244 46116 34748
rect 46396 34244 46452 34254
rect 46060 34242 46452 34244
rect 46060 34190 46398 34242
rect 46450 34190 46452 34242
rect 46060 34188 46452 34190
rect 46060 34018 46116 34188
rect 46396 34178 46452 34188
rect 47628 34132 47684 34142
rect 47516 34130 47684 34132
rect 47516 34078 47630 34130
rect 47682 34078 47684 34130
rect 47516 34076 47684 34078
rect 47292 34020 47348 34030
rect 47516 34020 47572 34076
rect 47628 34066 47684 34076
rect 46060 33966 46062 34018
rect 46114 33966 46116 34018
rect 46060 33954 46116 33966
rect 47068 34018 47572 34020
rect 47068 33966 47294 34018
rect 47346 33966 47572 34018
rect 47068 33964 47572 33966
rect 46508 33906 46564 33918
rect 46508 33854 46510 33906
rect 46562 33854 46564 33906
rect 46508 32116 46564 33854
rect 47068 33796 47124 33964
rect 47292 33954 47348 33964
rect 47628 33908 47684 33918
rect 46620 33346 46676 33358
rect 46620 33294 46622 33346
rect 46674 33294 46676 33346
rect 46620 33236 46676 33294
rect 46620 33170 46676 33180
rect 46508 32050 46564 32060
rect 46956 31108 47012 31118
rect 45948 31052 46228 31108
rect 45836 30942 45838 30994
rect 45890 30942 45892 30994
rect 45836 30930 45892 30942
rect 45612 30884 45668 30894
rect 45612 30790 45668 30828
rect 46060 30884 46116 30894
rect 45948 30770 46004 30782
rect 45948 30718 45950 30770
rect 46002 30718 46004 30770
rect 45724 30436 45780 30446
rect 45948 30436 46004 30718
rect 45724 30434 46004 30436
rect 45724 30382 45726 30434
rect 45778 30382 46004 30434
rect 45724 30380 46004 30382
rect 45724 30370 45780 30380
rect 45612 30324 45668 30334
rect 45388 30100 45444 30110
rect 45388 30098 45556 30100
rect 45388 30046 45390 30098
rect 45442 30046 45556 30098
rect 45388 30044 45556 30046
rect 45388 30034 45444 30044
rect 44044 29538 44100 29550
rect 44044 29486 44046 29538
rect 44098 29486 44100 29538
rect 43708 28018 43764 28028
rect 43820 29426 43876 29438
rect 43820 29374 43822 29426
rect 43874 29374 43876 29426
rect 43820 28642 43876 29374
rect 44044 28868 44100 29486
rect 44044 28802 44100 28812
rect 44492 29314 44548 29326
rect 44492 29262 44494 29314
rect 44546 29262 44548 29314
rect 44492 28756 44548 29262
rect 45052 29316 45108 29326
rect 45052 29314 45220 29316
rect 45052 29262 45054 29314
rect 45106 29262 45220 29314
rect 45052 29260 45220 29262
rect 45052 29250 45108 29260
rect 44604 29204 44660 29214
rect 44604 29110 44660 29148
rect 44492 28690 44548 28700
rect 44940 28756 44996 28766
rect 43820 28590 43822 28642
rect 43874 28590 43876 28642
rect 43708 27860 43764 27870
rect 43372 25506 43428 25518
rect 43372 25454 43374 25506
rect 43426 25454 43428 25506
rect 43372 25396 43428 25454
rect 43708 25506 43764 27804
rect 43820 27746 43876 28590
rect 44268 28644 44324 28654
rect 44268 28550 44324 28588
rect 44940 28642 44996 28700
rect 44940 28590 44942 28642
rect 44994 28590 44996 28642
rect 43820 27694 43822 27746
rect 43874 27694 43876 27746
rect 43820 27682 43876 27694
rect 44044 27858 44100 27870
rect 44044 27806 44046 27858
rect 44098 27806 44100 27858
rect 43708 25454 43710 25506
rect 43762 25454 43764 25506
rect 43708 25442 43764 25454
rect 43820 26962 43876 26974
rect 43820 26910 43822 26962
rect 43874 26910 43876 26962
rect 43820 26908 43876 26910
rect 44044 26908 44100 27806
rect 44380 27860 44436 27870
rect 44380 27766 44436 27804
rect 44716 27860 44772 27870
rect 44940 27860 44996 28590
rect 45164 28642 45220 29260
rect 45500 28868 45556 30044
rect 45612 30098 45668 30268
rect 45612 30046 45614 30098
rect 45666 30046 45668 30098
rect 45612 30034 45668 30046
rect 46060 29428 46116 30828
rect 45724 29372 46116 29428
rect 45612 28868 45668 28878
rect 45164 28590 45166 28642
rect 45218 28590 45220 28642
rect 45052 28530 45108 28542
rect 45052 28478 45054 28530
rect 45106 28478 45108 28530
rect 45052 28308 45108 28478
rect 45052 28242 45108 28252
rect 44716 27858 44996 27860
rect 44716 27806 44718 27858
rect 44770 27806 44996 27858
rect 44716 27804 44996 27806
rect 45052 27858 45108 27870
rect 45052 27806 45054 27858
rect 45106 27806 45108 27858
rect 44716 27794 44772 27804
rect 44268 27746 44324 27758
rect 44268 27694 44270 27746
rect 44322 27694 44324 27746
rect 44268 27636 44324 27694
rect 45052 27636 45108 27806
rect 44268 27580 45108 27636
rect 45164 26908 45220 28590
rect 45276 28866 45668 28868
rect 45276 28814 45614 28866
rect 45666 28814 45668 28866
rect 45276 28812 45668 28814
rect 45276 27858 45332 28812
rect 45612 28802 45668 28812
rect 45724 28644 45780 29372
rect 46060 29204 46116 29214
rect 46060 28866 46116 29148
rect 46172 29092 46228 31052
rect 46956 30324 47012 31052
rect 46172 29026 46228 29036
rect 46396 29428 46452 29438
rect 46060 28814 46062 28866
rect 46114 28814 46116 28866
rect 46060 28802 46116 28814
rect 45276 27806 45278 27858
rect 45330 27806 45332 27858
rect 45276 27794 45332 27806
rect 45500 28588 45780 28644
rect 46396 28756 46452 29372
rect 46956 29426 47012 30268
rect 46956 29374 46958 29426
rect 47010 29374 47012 29426
rect 46956 29362 47012 29374
rect 46396 28642 46452 28700
rect 46396 28590 46398 28642
rect 46450 28590 46452 28642
rect 45500 27858 45556 28588
rect 46396 28578 46452 28590
rect 46620 29316 46676 29326
rect 46172 28420 46228 28430
rect 46172 28326 46228 28364
rect 45500 27806 45502 27858
rect 45554 27806 45556 27858
rect 45388 27074 45444 27086
rect 45388 27022 45390 27074
rect 45442 27022 45444 27074
rect 45388 26908 45444 27022
rect 43820 26852 44100 26908
rect 44828 26852 45220 26908
rect 45276 26852 45444 26908
rect 43372 25330 43428 25340
rect 43372 21700 43428 21710
rect 43372 21606 43428 21644
rect 43204 20076 43428 20132
rect 43148 20066 43204 20076
rect 42924 19964 43092 20020
rect 42812 19842 42868 19852
rect 43036 19684 43092 19964
rect 43148 19908 43204 19918
rect 43204 19852 43316 19908
rect 43148 19842 43204 19852
rect 42700 19628 42868 19684
rect 42588 19294 42590 19346
rect 42642 19294 42644 19346
rect 42588 19236 42644 19294
rect 42588 19170 42644 19180
rect 42700 18562 42756 18574
rect 42700 18510 42702 18562
rect 42754 18510 42756 18562
rect 42364 18450 42532 18452
rect 42364 18398 42366 18450
rect 42418 18398 42532 18450
rect 42364 18396 42532 18398
rect 42364 18386 42420 18396
rect 40908 17666 41076 17668
rect 40908 17614 40910 17666
rect 40962 17614 41076 17666
rect 40908 17612 41076 17614
rect 40908 17602 40964 17612
rect 41020 17106 41076 17612
rect 41132 17666 41524 17668
rect 41132 17614 41470 17666
rect 41522 17614 41524 17666
rect 41132 17612 41524 17614
rect 41132 17554 41188 17612
rect 41468 17602 41524 17612
rect 41692 18060 41860 18116
rect 42476 18228 42532 18396
rect 41132 17502 41134 17554
rect 41186 17502 41188 17554
rect 41132 17490 41188 17502
rect 41020 17054 41022 17106
rect 41074 17054 41076 17106
rect 41020 17042 41076 17054
rect 41468 16884 41524 16894
rect 41468 16790 41524 16828
rect 41692 16100 41748 18060
rect 41916 17780 41972 17790
rect 41804 17778 41972 17780
rect 41804 17726 41918 17778
rect 41970 17726 41972 17778
rect 41804 17724 41972 17726
rect 41804 16884 41860 17724
rect 41916 17714 41972 17724
rect 42476 17778 42532 18172
rect 42476 17726 42478 17778
rect 42530 17726 42532 17778
rect 42476 17220 42532 17726
rect 42028 17164 42532 17220
rect 41804 16818 41860 16828
rect 41916 16996 41972 17006
rect 41916 16882 41972 16940
rect 41916 16830 41918 16882
rect 41970 16830 41972 16882
rect 41916 16818 41972 16830
rect 42028 16210 42084 17164
rect 42028 16158 42030 16210
rect 42082 16158 42084 16210
rect 42028 16146 42084 16158
rect 42252 16994 42308 17006
rect 42252 16942 42254 16994
rect 42306 16942 42308 16994
rect 41804 16100 41860 16110
rect 41692 16044 41804 16100
rect 41132 15202 41188 15214
rect 41132 15150 41134 15202
rect 41186 15150 41188 15202
rect 41132 15148 41188 15150
rect 40908 15092 41188 15148
rect 40908 14532 40964 15092
rect 40908 14438 40964 14476
rect 40460 14418 40516 14430
rect 40460 14366 40462 14418
rect 40514 14366 40516 14418
rect 40460 14084 40516 14366
rect 41692 14418 41748 14430
rect 41692 14366 41694 14418
rect 41746 14366 41748 14418
rect 40572 14308 40628 14318
rect 41692 14308 41748 14366
rect 40572 14306 41748 14308
rect 40572 14254 40574 14306
rect 40626 14254 41748 14306
rect 40572 14252 41748 14254
rect 40572 14242 40628 14252
rect 40684 14140 41636 14196
rect 40684 14084 40740 14140
rect 40460 14028 40740 14084
rect 41580 13970 41636 14140
rect 41580 13918 41582 13970
rect 41634 13918 41636 13970
rect 41580 13906 41636 13918
rect 41692 13972 41748 13982
rect 41692 13878 41748 13916
rect 40348 13682 40404 13692
rect 41356 13746 41412 13758
rect 41356 13694 41358 13746
rect 41410 13694 41412 13746
rect 40908 13524 40964 13534
rect 40572 12740 40628 12750
rect 40124 12738 40628 12740
rect 40124 12686 40574 12738
rect 40626 12686 40628 12738
rect 40124 12684 40628 12686
rect 39676 12126 39678 12178
rect 39730 12126 39732 12178
rect 39676 12114 39732 12126
rect 40460 12516 40516 12526
rect 40012 12068 40068 12078
rect 40012 11974 40068 12012
rect 40124 11954 40180 11966
rect 40124 11902 40126 11954
rect 40178 11902 40180 11954
rect 40124 11506 40180 11902
rect 40124 11454 40126 11506
rect 40178 11454 40180 11506
rect 40124 11442 40180 11454
rect 40012 10612 40068 10622
rect 40012 10518 40068 10556
rect 39564 9996 39732 10052
rect 39452 9774 39454 9826
rect 39506 9774 39508 9826
rect 39452 9716 39508 9774
rect 39452 9650 39508 9660
rect 39564 9826 39620 9838
rect 39564 9774 39566 9826
rect 39618 9774 39620 9826
rect 38108 9604 38164 9614
rect 37324 8932 37380 8942
rect 37324 8930 38052 8932
rect 37324 8878 37326 8930
rect 37378 8878 38052 8930
rect 37324 8876 38052 8878
rect 37324 8866 37380 8876
rect 37996 8482 38052 8876
rect 37996 8430 37998 8482
rect 38050 8430 38052 8482
rect 37996 8418 38052 8430
rect 38108 8370 38164 9548
rect 38668 9604 38724 9614
rect 39116 9604 39172 9614
rect 38668 9602 39172 9604
rect 38668 9550 38670 9602
rect 38722 9550 39118 9602
rect 39170 9550 39172 9602
rect 38668 9548 39172 9550
rect 38668 9538 38724 9548
rect 39116 9492 39172 9548
rect 39340 9604 39396 9614
rect 39340 9510 39396 9548
rect 39116 9426 39172 9436
rect 39564 9156 39620 9774
rect 39452 8932 39508 8942
rect 39564 8932 39620 9100
rect 39452 8930 39620 8932
rect 39452 8878 39454 8930
rect 39506 8878 39620 8930
rect 39452 8876 39620 8878
rect 39452 8866 39508 8876
rect 39676 8820 39732 9996
rect 40236 9716 40292 9726
rect 40292 9660 40404 9716
rect 40236 9650 40292 9660
rect 40124 9156 40180 9166
rect 40124 9062 40180 9100
rect 38108 8318 38110 8370
rect 38162 8318 38164 8370
rect 38108 8306 38164 8318
rect 39564 8764 39732 8820
rect 40236 8820 40292 8830
rect 37324 7812 37380 7822
rect 37212 7756 37324 7812
rect 37324 7746 37380 7756
rect 39228 7700 39284 7710
rect 39228 7586 39284 7644
rect 39228 7534 39230 7586
rect 39282 7534 39284 7586
rect 39228 7522 39284 7534
rect 38220 7252 38276 7262
rect 37212 6578 37268 6590
rect 37212 6526 37214 6578
rect 37266 6526 37268 6578
rect 36316 6468 36372 6478
rect 36316 6466 36932 6468
rect 36316 6414 36318 6466
rect 36370 6414 36932 6466
rect 36316 6412 36932 6414
rect 36316 6402 36372 6412
rect 36316 6244 36372 6254
rect 36204 6188 36316 6244
rect 35308 5854 35310 5906
rect 35362 5854 35364 5906
rect 35308 5842 35364 5854
rect 34636 5740 35140 5796
rect 35308 5684 35364 5694
rect 34524 5628 34692 5684
rect 34412 4470 34468 4508
rect 34524 5012 34580 5022
rect 34524 4562 34580 4956
rect 34524 4510 34526 4562
rect 34578 4510 34580 4562
rect 34524 4498 34580 4510
rect 29260 4286 29262 4338
rect 29314 4286 29316 4338
rect 29260 4274 29316 4286
rect 32172 4226 32228 4396
rect 33180 4452 33236 4462
rect 33180 4358 33236 4396
rect 34636 4450 34692 5628
rect 35308 5682 35700 5684
rect 35308 5630 35310 5682
rect 35362 5630 35700 5682
rect 35308 5628 35700 5630
rect 35308 5618 35364 5628
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35644 5234 35700 5628
rect 35644 5182 35646 5234
rect 35698 5182 35700 5234
rect 35644 5170 35700 5182
rect 34636 4398 34638 4450
rect 34690 4398 34692 4450
rect 34636 4386 34692 4398
rect 36316 5122 36372 6188
rect 36316 5070 36318 5122
rect 36370 5070 36372 5122
rect 36204 4340 36260 4350
rect 36316 4340 36372 5070
rect 36876 4450 36932 6412
rect 37212 6244 37268 6526
rect 37212 6178 37268 6188
rect 38220 6018 38276 7196
rect 39116 7252 39172 7262
rect 39116 7158 39172 7196
rect 38220 5966 38222 6018
rect 38274 5966 38276 6018
rect 38220 5954 38276 5966
rect 37548 5908 37604 5918
rect 37548 5814 37604 5852
rect 38556 5908 38612 5918
rect 38556 5122 38612 5852
rect 38556 5070 38558 5122
rect 38610 5070 38612 5122
rect 38556 5058 38612 5070
rect 39228 5012 39284 5022
rect 39228 4918 39284 4956
rect 36876 4398 36878 4450
rect 36930 4398 36932 4450
rect 36876 4386 36932 4398
rect 39564 4452 39620 8764
rect 40236 8726 40292 8764
rect 40348 8596 40404 9660
rect 40012 8540 40348 8596
rect 39900 7700 39956 7710
rect 39900 7606 39956 7644
rect 40012 7698 40068 8540
rect 40348 8502 40404 8540
rect 40460 8372 40516 12460
rect 40572 11956 40628 12684
rect 40908 12516 40964 13468
rect 41356 13300 41412 13694
rect 40908 12450 40964 12460
rect 41020 13244 41356 13300
rect 41020 12402 41076 13244
rect 41356 13234 41412 13244
rect 41468 13748 41524 13758
rect 41356 13074 41412 13086
rect 41356 13022 41358 13074
rect 41410 13022 41412 13074
rect 41356 12628 41412 13022
rect 41356 12562 41412 12572
rect 41020 12350 41022 12402
rect 41074 12350 41076 12402
rect 41020 12338 41076 12350
rect 41356 12404 41412 12414
rect 41356 12310 41412 12348
rect 40572 11890 40628 11900
rect 41132 12178 41188 12190
rect 41468 12180 41524 13692
rect 41132 12126 41134 12178
rect 41186 12126 41188 12178
rect 41132 11956 41188 12126
rect 41356 12124 41524 12180
rect 41580 12180 41636 12190
rect 41244 12068 41300 12078
rect 41244 11974 41300 12012
rect 41132 11890 41188 11900
rect 40908 11394 40964 11406
rect 40908 11342 40910 11394
rect 40962 11342 40964 11394
rect 40908 10724 40964 11342
rect 40908 10658 40964 10668
rect 41020 9828 41076 9838
rect 41356 9828 41412 12124
rect 41580 12086 41636 12124
rect 41804 11172 41860 16044
rect 42252 15148 42308 16942
rect 42476 16882 42532 17164
rect 42476 16830 42478 16882
rect 42530 16830 42532 16882
rect 42476 16818 42532 16830
rect 42028 15092 42308 15148
rect 41916 13860 41972 13870
rect 41916 13766 41972 13804
rect 42028 13300 42084 15092
rect 42028 13234 42084 13244
rect 42140 13972 42196 13982
rect 41916 12628 41972 12638
rect 41916 12290 41972 12572
rect 42140 12404 42196 13916
rect 42700 13972 42756 18510
rect 42812 15428 42868 19628
rect 42812 15362 42868 15372
rect 42924 19628 43092 19684
rect 42700 13906 42756 13916
rect 42588 13636 42644 13646
rect 41916 12238 41918 12290
rect 41970 12238 41972 12290
rect 41916 12226 41972 12238
rect 42028 12348 42140 12404
rect 41916 11956 41972 11966
rect 41916 11394 41972 11900
rect 41916 11342 41918 11394
rect 41970 11342 41972 11394
rect 41916 11330 41972 11342
rect 42028 11396 42084 12348
rect 42140 12310 42196 12348
rect 42252 13634 42644 13636
rect 42252 13582 42590 13634
rect 42642 13582 42644 13634
rect 42252 13580 42644 13582
rect 42252 12402 42308 13580
rect 42588 13570 42644 13580
rect 42700 13524 42756 13534
rect 42700 13430 42756 13468
rect 42476 13300 42532 13310
rect 42252 12350 42254 12402
rect 42306 12350 42308 12402
rect 42252 12338 42308 12350
rect 42364 12404 42420 12414
rect 42364 12310 42420 12348
rect 42476 12402 42532 13244
rect 42476 12350 42478 12402
rect 42530 12350 42532 12402
rect 42476 11956 42532 12350
rect 42924 12404 42980 19628
rect 43036 19236 43092 19246
rect 43036 19142 43092 19180
rect 43260 19234 43316 19852
rect 43260 19182 43262 19234
rect 43314 19182 43316 19234
rect 43036 18676 43092 18686
rect 43036 18450 43092 18620
rect 43036 18398 43038 18450
rect 43090 18398 43092 18450
rect 43036 18386 43092 18398
rect 43260 18452 43316 19182
rect 43260 18386 43316 18396
rect 43260 18116 43316 18126
rect 43260 16996 43316 18060
rect 43036 12404 43092 12414
rect 42980 12402 43092 12404
rect 42980 12350 43038 12402
rect 43090 12350 43092 12402
rect 42980 12348 43092 12350
rect 42924 12310 42980 12348
rect 43036 12338 43092 12348
rect 42476 11890 42532 11900
rect 42812 11508 42868 11518
rect 42364 11506 42868 11508
rect 42364 11454 42814 11506
rect 42866 11454 42868 11506
rect 42364 11452 42868 11454
rect 42028 11340 42308 11396
rect 42252 11282 42308 11340
rect 42252 11230 42254 11282
rect 42306 11230 42308 11282
rect 42252 11218 42308 11230
rect 42028 11172 42084 11182
rect 41804 11170 42084 11172
rect 41804 11118 42030 11170
rect 42082 11118 42084 11170
rect 41804 11116 42084 11118
rect 41020 9826 41412 9828
rect 41020 9774 41022 9826
rect 41074 9774 41412 9826
rect 41020 9772 41412 9774
rect 41580 10724 41636 10734
rect 41020 9762 41076 9772
rect 41468 9716 41524 9726
rect 41468 9622 41524 9660
rect 40012 7646 40014 7698
rect 40066 7646 40068 7698
rect 40012 7634 40068 7646
rect 40124 8370 40516 8372
rect 40124 8318 40462 8370
rect 40514 8318 40516 8370
rect 40124 8316 40516 8318
rect 39676 7476 39732 7486
rect 39676 7382 39732 7420
rect 39788 7476 39844 7486
rect 40124 7476 40180 8316
rect 40460 8306 40516 8316
rect 40908 9602 40964 9614
rect 40908 9550 40910 9602
rect 40962 9550 40964 9602
rect 40908 9492 40964 9550
rect 39788 7474 40180 7476
rect 39788 7422 39790 7474
rect 39842 7422 40180 7474
rect 39788 7420 40180 7422
rect 40236 7474 40292 7486
rect 40236 7422 40238 7474
rect 40290 7422 40292 7474
rect 39788 7410 39844 7420
rect 40236 6580 40292 7422
rect 40908 7476 40964 9436
rect 41132 9602 41188 9614
rect 41132 9550 41134 9602
rect 41186 9550 41188 9602
rect 41132 9156 41188 9550
rect 41244 9604 41300 9614
rect 41244 9510 41300 9548
rect 41244 9156 41300 9166
rect 41132 9154 41300 9156
rect 41132 9102 41246 9154
rect 41298 9102 41300 9154
rect 41132 9100 41300 9102
rect 41244 9090 41300 9100
rect 41356 8818 41412 8830
rect 41356 8766 41358 8818
rect 41410 8766 41412 8818
rect 41244 8596 41300 8606
rect 41244 7700 41300 8540
rect 41356 8372 41412 8766
rect 41356 8306 41412 8316
rect 41468 8260 41524 8270
rect 41580 8260 41636 10668
rect 41468 8258 41636 8260
rect 41468 8206 41470 8258
rect 41522 8206 41636 8258
rect 41468 8204 41636 8206
rect 41468 8194 41524 8204
rect 41916 8036 41972 11116
rect 42028 11106 42084 11116
rect 42140 11170 42196 11182
rect 42140 11118 42142 11170
rect 42194 11118 42196 11170
rect 42140 11060 42196 11118
rect 42364 11060 42420 11452
rect 42812 11442 42868 11452
rect 42140 11004 42420 11060
rect 42476 11282 42532 11294
rect 42476 11230 42478 11282
rect 42530 11230 42532 11282
rect 42476 10836 42532 11230
rect 42924 11172 42980 11182
rect 42924 11170 43092 11172
rect 42924 11118 42926 11170
rect 42978 11118 43092 11170
rect 42924 11116 43092 11118
rect 42924 11106 42980 11116
rect 42476 10770 42532 10780
rect 42924 10724 42980 10734
rect 42588 10052 42644 10062
rect 42252 9940 42308 9950
rect 42252 9716 42308 9884
rect 42588 9826 42644 9996
rect 42588 9774 42590 9826
rect 42642 9774 42644 9826
rect 42588 9762 42644 9774
rect 42252 9714 42532 9716
rect 42252 9662 42254 9714
rect 42306 9662 42532 9714
rect 42252 9660 42532 9662
rect 42252 9650 42308 9660
rect 42476 8708 42532 9660
rect 42924 9042 42980 10668
rect 43036 9156 43092 11116
rect 43036 9090 43092 9100
rect 42924 8990 42926 9042
rect 42978 8990 42980 9042
rect 42924 8978 42980 8990
rect 43260 9044 43316 16940
rect 43372 9268 43428 20076
rect 43596 19122 43652 19134
rect 43596 19070 43598 19122
rect 43650 19070 43652 19122
rect 43484 19012 43540 19022
rect 43484 18918 43540 18956
rect 43484 15876 43540 15886
rect 43484 15782 43540 15820
rect 43484 13524 43540 13534
rect 43484 12962 43540 13468
rect 43484 12910 43486 12962
rect 43538 12910 43540 12962
rect 43484 12898 43540 12910
rect 43596 10052 43652 19070
rect 43820 18116 43876 26852
rect 44268 25396 44324 25406
rect 44268 25394 44772 25396
rect 44268 25342 44270 25394
rect 44322 25342 44772 25394
rect 44268 25340 44772 25342
rect 44268 25330 44324 25340
rect 44716 24834 44772 25340
rect 44716 24782 44718 24834
rect 44770 24782 44772 24834
rect 44716 24770 44772 24782
rect 43932 24610 43988 24622
rect 43932 24558 43934 24610
rect 43986 24558 43988 24610
rect 43932 24500 43988 24558
rect 43932 24434 43988 24444
rect 44268 22484 44324 22494
rect 44268 22390 44324 22428
rect 44604 21588 44660 21598
rect 44156 20580 44212 20590
rect 43932 19012 43988 19022
rect 43932 18450 43988 18956
rect 44156 18788 44212 20524
rect 44604 20018 44660 21532
rect 44828 20580 44884 26852
rect 45052 25508 45108 25518
rect 45052 25506 45220 25508
rect 45052 25454 45054 25506
rect 45106 25454 45220 25506
rect 45052 25452 45220 25454
rect 45052 25442 45108 25452
rect 44940 24612 44996 24622
rect 44996 24556 45108 24612
rect 44940 24518 44996 24556
rect 45052 23826 45108 24556
rect 45052 23774 45054 23826
rect 45106 23774 45108 23826
rect 45052 23762 45108 23774
rect 45164 23716 45220 25452
rect 45276 24946 45332 26852
rect 45276 24894 45278 24946
rect 45330 24894 45332 24946
rect 45276 24882 45332 24894
rect 45276 23940 45332 23950
rect 45276 23846 45332 23884
rect 45500 23828 45556 27806
rect 45612 27748 45668 27758
rect 45612 27654 45668 27692
rect 46620 26908 46676 29260
rect 45612 26852 45668 26862
rect 46620 26852 46788 26908
rect 45612 26850 45780 26852
rect 45612 26798 45614 26850
rect 45666 26798 45780 26850
rect 45612 26796 45780 26798
rect 45612 26786 45668 26796
rect 45724 25618 45780 26796
rect 46172 26292 46228 26302
rect 46620 26292 46676 26302
rect 46172 26290 46620 26292
rect 46172 26238 46174 26290
rect 46226 26238 46620 26290
rect 46172 26236 46620 26238
rect 46172 26226 46228 26236
rect 46620 26198 46676 26236
rect 45724 25566 45726 25618
rect 45778 25566 45780 25618
rect 45724 25554 45780 25566
rect 46732 24388 46788 26852
rect 46620 24332 46788 24388
rect 45948 23940 46004 23950
rect 45948 23846 46004 23884
rect 46396 23940 46452 23950
rect 46396 23846 46452 23884
rect 45724 23828 45780 23838
rect 45500 23772 45724 23828
rect 45724 23734 45780 23772
rect 45164 23660 45332 23716
rect 45276 23492 45332 23660
rect 45276 23436 45444 23492
rect 45388 22482 45444 23436
rect 45388 22430 45390 22482
rect 45442 22430 45444 22482
rect 45388 21588 45444 22430
rect 46060 23044 46116 23054
rect 46060 21698 46116 22988
rect 46060 21646 46062 21698
rect 46114 21646 46116 21698
rect 46060 21634 46116 21646
rect 45388 21494 45444 21532
rect 44828 20524 44996 20580
rect 44604 19966 44606 20018
rect 44658 19966 44660 20018
rect 44604 19954 44660 19966
rect 44716 19348 44772 19358
rect 44940 19348 44996 20524
rect 44772 19292 44996 19348
rect 44492 19236 44548 19246
rect 44268 19012 44324 19022
rect 44268 18918 44324 18956
rect 44156 18732 44324 18788
rect 43932 18398 43934 18450
rect 43986 18398 43988 18450
rect 43932 18386 43988 18398
rect 44156 18562 44212 18574
rect 44156 18510 44158 18562
rect 44210 18510 44212 18562
rect 43820 18050 43876 18060
rect 44156 17556 44212 18510
rect 44156 17490 44212 17500
rect 44268 17106 44324 18732
rect 44268 17054 44270 17106
rect 44322 17054 44324 17106
rect 44268 17042 44324 17054
rect 44492 17106 44548 19180
rect 44716 18450 44772 19292
rect 44940 19234 44996 19292
rect 44940 19182 44942 19234
rect 44994 19182 44996 19234
rect 44940 19170 44996 19182
rect 45388 19906 45444 19918
rect 45388 19854 45390 19906
rect 45442 19854 45444 19906
rect 44828 19122 44884 19134
rect 44828 19070 44830 19122
rect 44882 19070 44884 19122
rect 44828 18676 44884 19070
rect 45276 19012 45332 19022
rect 45164 18676 45220 18686
rect 44828 18674 45220 18676
rect 44828 18622 45166 18674
rect 45218 18622 45220 18674
rect 44828 18620 45220 18622
rect 45164 18610 45220 18620
rect 44716 18398 44718 18450
rect 44770 18398 44772 18450
rect 44716 18386 44772 18398
rect 45052 18452 45108 18462
rect 45276 18452 45332 18956
rect 45388 18674 45444 19854
rect 46620 19460 46676 24332
rect 47068 24276 47124 33740
rect 47404 33906 47684 33908
rect 47404 33854 47630 33906
rect 47682 33854 47684 33906
rect 47404 33852 47684 33854
rect 47404 33458 47460 33852
rect 47628 33842 47684 33852
rect 47964 33908 48020 33918
rect 47964 33906 48244 33908
rect 47964 33854 47966 33906
rect 48018 33854 48244 33906
rect 47964 33852 48244 33854
rect 47964 33842 48020 33852
rect 47404 33406 47406 33458
rect 47458 33406 47460 33458
rect 47404 33394 47460 33406
rect 48188 32674 48244 33852
rect 48188 32622 48190 32674
rect 48242 32622 48244 32674
rect 48188 32610 48244 32622
rect 47740 32564 47796 32574
rect 47740 32470 47796 32508
rect 47292 32450 47348 32462
rect 47292 32398 47294 32450
rect 47346 32398 47348 32450
rect 47292 32004 47348 32398
rect 47740 32116 47796 32126
rect 47796 32060 47908 32116
rect 47740 32050 47796 32060
rect 47292 31938 47348 31948
rect 47740 31892 47796 31902
rect 47404 31890 47796 31892
rect 47404 31838 47742 31890
rect 47794 31838 47796 31890
rect 47404 31836 47796 31838
rect 47404 31108 47460 31836
rect 47740 31826 47796 31836
rect 47516 31220 47572 31230
rect 47516 31126 47572 31164
rect 47404 31014 47460 31052
rect 47404 29538 47460 29550
rect 47404 29486 47406 29538
rect 47458 29486 47460 29538
rect 47180 29428 47236 29438
rect 47180 29334 47236 29372
rect 47180 28644 47236 28654
rect 47180 28550 47236 28588
rect 47404 28530 47460 29486
rect 47516 29426 47572 29438
rect 47516 29374 47518 29426
rect 47570 29374 47572 29426
rect 47516 29316 47572 29374
rect 47516 29250 47572 29260
rect 47852 28644 47908 32060
rect 48188 31666 48244 31678
rect 48188 31614 48190 31666
rect 48242 31614 48244 31666
rect 47964 31556 48020 31566
rect 47964 29650 48020 31500
rect 48188 31220 48244 31614
rect 48188 31154 48244 31164
rect 47964 29598 47966 29650
rect 48018 29598 48020 29650
rect 47964 29586 48020 29598
rect 48188 30772 48244 30782
rect 47404 28478 47406 28530
rect 47458 28478 47460 28530
rect 47180 27860 47236 27870
rect 47180 26962 47236 27804
rect 47180 26910 47182 26962
rect 47234 26910 47236 26962
rect 47180 26898 47236 26910
rect 47404 26908 47460 28478
rect 47516 28642 47908 28644
rect 47516 28590 47854 28642
rect 47906 28590 47908 28642
rect 47516 28588 47908 28590
rect 47516 28082 47572 28588
rect 47852 28578 47908 28588
rect 48188 28530 48244 30716
rect 48188 28478 48190 28530
rect 48242 28478 48244 28530
rect 47628 28418 47684 28430
rect 47628 28366 47630 28418
rect 47682 28366 47684 28418
rect 47628 28308 47684 28366
rect 47628 28242 47684 28252
rect 47516 28030 47518 28082
rect 47570 28030 47572 28082
rect 47516 28018 47572 28030
rect 47740 27860 47796 27870
rect 47740 27766 47796 27804
rect 48188 27858 48244 28478
rect 48188 27806 48190 27858
rect 48242 27806 48244 27858
rect 48188 27794 48244 27806
rect 47628 27748 47684 27758
rect 47628 27654 47684 27692
rect 47404 26852 47572 26908
rect 47516 26850 47572 26852
rect 47516 26798 47518 26850
rect 47570 26798 47572 26850
rect 47516 25620 47572 26798
rect 47852 25620 47908 25630
rect 47516 25618 47908 25620
rect 47516 25566 47854 25618
rect 47906 25566 47908 25618
rect 47516 25564 47908 25566
rect 47852 25554 47908 25564
rect 48300 25620 48356 37100
rect 48412 34692 48468 34702
rect 48636 34692 48692 37996
rect 48748 37958 48804 37996
rect 48748 37604 48804 37614
rect 48748 37378 48804 37548
rect 48860 37492 48916 37502
rect 48860 37398 48916 37436
rect 48748 37326 48750 37378
rect 48802 37326 48804 37378
rect 48748 37314 48804 37326
rect 48972 37266 49028 38782
rect 49308 38948 49364 38958
rect 49420 38948 49476 39340
rect 49308 38946 49476 38948
rect 49308 38894 49310 38946
rect 49362 38894 49476 38946
rect 49308 38892 49476 38894
rect 49308 37378 49364 38892
rect 49980 38724 50036 38734
rect 50092 38724 50148 40460
rect 50428 40404 50484 44380
rect 50540 44370 50596 44380
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 51212 43876 51268 45836
rect 51324 45826 51380 45836
rect 51436 45780 51492 45790
rect 51660 45780 51716 51212
rect 51772 51268 51828 51278
rect 51772 50370 51828 51212
rect 51772 50318 51774 50370
rect 51826 50318 51828 50370
rect 51772 50306 51828 50318
rect 51436 45778 51716 45780
rect 51436 45726 51438 45778
rect 51490 45726 51716 45778
rect 51436 45724 51716 45726
rect 51324 45666 51380 45678
rect 51324 45614 51326 45666
rect 51378 45614 51380 45666
rect 51324 44548 51380 45614
rect 51324 44482 51380 44492
rect 50556 43866 50820 43876
rect 50988 43820 51268 43876
rect 50988 43708 51044 43820
rect 51436 43708 51492 45724
rect 51884 45668 51940 51436
rect 51660 45612 51940 45668
rect 51996 47236 52052 47246
rect 50876 43652 51044 43708
rect 51212 43652 51492 43708
rect 51548 45332 51604 45342
rect 51548 44322 51604 45276
rect 51548 44270 51550 44322
rect 51602 44270 51604 44322
rect 50764 43540 50820 43550
rect 50764 43446 50820 43484
rect 50764 42756 50820 42766
rect 50876 42756 50932 43652
rect 50764 42754 50932 42756
rect 50764 42702 50766 42754
rect 50818 42702 50932 42754
rect 50764 42700 50932 42702
rect 50764 42690 50820 42700
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 50764 41860 50820 41870
rect 50876 41860 50932 42700
rect 50988 42756 51044 42766
rect 51212 42756 51268 43652
rect 51548 42978 51604 44270
rect 51660 43708 51716 45612
rect 51884 45220 51940 45230
rect 51772 44324 51828 44334
rect 51772 44230 51828 44268
rect 51660 43652 51828 43708
rect 51548 42926 51550 42978
rect 51602 42926 51604 42978
rect 51548 42914 51604 42926
rect 50988 42754 51268 42756
rect 50988 42702 50990 42754
rect 51042 42702 51268 42754
rect 50988 42700 51268 42702
rect 51324 42866 51380 42878
rect 51324 42814 51326 42866
rect 51378 42814 51380 42866
rect 51324 42756 51380 42814
rect 50988 42690 51044 42700
rect 51324 42690 51380 42700
rect 51772 42754 51828 43652
rect 51772 42702 51774 42754
rect 51826 42702 51828 42754
rect 51772 42644 51828 42702
rect 51772 42578 51828 42588
rect 50820 41804 50932 41860
rect 51548 42084 51604 42094
rect 50764 41794 50820 41804
rect 51212 41188 51268 41198
rect 51212 41094 51268 41132
rect 51548 41186 51604 42028
rect 51884 41972 51940 45164
rect 51996 44434 52052 47180
rect 52108 46788 52164 46798
rect 52108 46694 52164 46732
rect 51996 44382 51998 44434
rect 52050 44382 52052 44434
rect 51996 44370 52052 44382
rect 52108 44548 52164 44558
rect 52108 44322 52164 44492
rect 52108 44270 52110 44322
rect 52162 44270 52164 44322
rect 52108 43708 52164 44270
rect 51996 43652 52164 43708
rect 51996 43538 52052 43652
rect 51996 43486 51998 43538
rect 52050 43486 52052 43538
rect 51996 43474 52052 43486
rect 52220 42196 52276 55412
rect 55356 55410 55636 55412
rect 55356 55358 55582 55410
rect 55634 55358 55636 55410
rect 55356 55356 55636 55358
rect 52668 55300 52724 55310
rect 52668 55206 52724 55244
rect 53452 55188 53508 55198
rect 53452 55094 53508 55132
rect 54460 55188 54516 55198
rect 54460 54738 54516 55132
rect 54460 54686 54462 54738
rect 54514 54686 54516 54738
rect 54460 54674 54516 54686
rect 54572 54626 54628 54638
rect 54572 54574 54574 54626
rect 54626 54574 54628 54626
rect 52892 54514 52948 54526
rect 52892 54462 52894 54514
rect 52946 54462 52948 54514
rect 52892 54404 52948 54462
rect 54572 54516 54628 54574
rect 54572 54450 54628 54460
rect 52780 53844 52836 53854
rect 52780 53750 52836 53788
rect 52892 50596 52948 54348
rect 54348 54290 54404 54302
rect 54348 54238 54350 54290
rect 54402 54238 54404 54290
rect 54236 53956 54292 53966
rect 53676 53844 53732 53854
rect 53228 53730 53284 53742
rect 53228 53678 53230 53730
rect 53282 53678 53284 53730
rect 53228 53620 53284 53678
rect 53676 53730 53732 53788
rect 53676 53678 53678 53730
rect 53730 53678 53732 53730
rect 53676 53666 53732 53678
rect 54236 53730 54292 53900
rect 54348 53844 54404 54238
rect 54348 53778 54404 53788
rect 54908 53956 54964 53966
rect 54236 53678 54238 53730
rect 54290 53678 54292 53730
rect 54236 53666 54292 53678
rect 53228 53554 53284 53564
rect 54012 53620 54068 53630
rect 52556 50594 52948 50596
rect 52556 50542 52894 50594
rect 52946 50542 52948 50594
rect 52556 50540 52948 50542
rect 52556 50034 52612 50540
rect 52892 50530 52948 50540
rect 53004 52164 53060 52174
rect 52556 49982 52558 50034
rect 52610 49982 52612 50034
rect 52444 47796 52500 47806
rect 52444 46898 52500 47740
rect 52556 47572 52612 49982
rect 53004 49140 53060 52108
rect 53788 51268 53844 51278
rect 53788 51174 53844 51212
rect 54012 49364 54068 53564
rect 54908 53058 54964 53900
rect 55356 53956 55412 55356
rect 55580 55346 55636 55356
rect 57596 55412 57652 55422
rect 57708 55412 57876 55468
rect 57596 55410 57764 55412
rect 57596 55358 57598 55410
rect 57650 55358 57764 55410
rect 57596 55356 57764 55358
rect 57596 55346 57652 55356
rect 57484 55074 57540 55086
rect 57484 55022 57486 55074
rect 57538 55022 57540 55074
rect 54908 53006 54910 53058
rect 54962 53006 54964 53058
rect 54908 52994 54964 53006
rect 55020 53732 55076 53742
rect 55020 53058 55076 53676
rect 55356 53730 55412 53900
rect 55356 53678 55358 53730
rect 55410 53678 55412 53730
rect 55356 53666 55412 53678
rect 56252 54628 56308 54638
rect 55580 53618 55636 53630
rect 55580 53566 55582 53618
rect 55634 53566 55636 53618
rect 55244 53508 55300 53518
rect 55244 53414 55300 53452
rect 55580 53172 55636 53566
rect 55020 53006 55022 53058
rect 55074 53006 55076 53058
rect 55020 52994 55076 53006
rect 55244 53116 55636 53172
rect 55916 53506 55972 53518
rect 55916 53454 55918 53506
rect 55970 53454 55972 53506
rect 54796 52948 54852 52958
rect 54796 52854 54852 52892
rect 55244 52948 55300 53116
rect 55244 52276 55300 52892
rect 55468 52948 55524 52958
rect 55468 52854 55524 52892
rect 55244 52182 55300 52220
rect 55916 51940 55972 53454
rect 56252 53506 56308 54572
rect 56252 53454 56254 53506
rect 56306 53454 56308 53506
rect 55916 51874 55972 51884
rect 56140 52276 56196 52286
rect 54572 51378 54628 51390
rect 54572 51326 54574 51378
rect 54626 51326 54628 51378
rect 54572 50484 54628 51326
rect 55356 51380 55412 51390
rect 55692 51380 55748 51390
rect 55412 51378 55748 51380
rect 55412 51326 55694 51378
rect 55746 51326 55748 51378
rect 55412 51324 55748 51326
rect 55356 51286 55412 51324
rect 55692 51314 55748 51324
rect 55916 51266 55972 51278
rect 55916 51214 55918 51266
rect 55970 51214 55972 51266
rect 54572 50418 54628 50428
rect 55244 50484 55300 50494
rect 53788 49308 54068 49364
rect 53004 49138 53172 49140
rect 53004 49086 53006 49138
rect 53058 49086 53172 49138
rect 53004 49084 53172 49086
rect 53004 49074 53060 49084
rect 52556 47506 52612 47516
rect 52780 47236 52836 47246
rect 52780 47142 52836 47180
rect 52892 47234 52948 47246
rect 52892 47182 52894 47234
rect 52946 47182 52948 47234
rect 52444 46846 52446 46898
rect 52498 46846 52500 46898
rect 52444 46834 52500 46846
rect 52780 46676 52836 46686
rect 52780 45890 52836 46620
rect 52780 45838 52782 45890
rect 52834 45838 52836 45890
rect 52780 45826 52836 45838
rect 52892 45556 52948 47182
rect 52892 45490 52948 45500
rect 53004 47234 53060 47246
rect 53004 47182 53006 47234
rect 53058 47182 53060 47234
rect 53004 46788 53060 47182
rect 52780 45220 52836 45230
rect 52780 45126 52836 45164
rect 53004 44434 53060 46732
rect 53004 44382 53006 44434
rect 53058 44382 53060 44434
rect 53004 44370 53060 44382
rect 53116 46452 53172 49084
rect 53452 48804 53508 48814
rect 53452 48802 53732 48804
rect 53452 48750 53454 48802
rect 53506 48750 53732 48802
rect 53452 48748 53732 48750
rect 53452 48738 53508 48748
rect 53676 48130 53732 48748
rect 53676 48078 53678 48130
rect 53730 48078 53732 48130
rect 52780 44322 52836 44334
rect 52780 44270 52782 44322
rect 52834 44270 52836 44322
rect 52444 43652 52500 43662
rect 52444 43538 52500 43596
rect 52444 43486 52446 43538
rect 52498 43486 52500 43538
rect 52444 43474 52500 43486
rect 52780 42978 52836 44270
rect 53116 43538 53172 46396
rect 53340 47458 53396 47470
rect 53340 47406 53342 47458
rect 53394 47406 53396 47458
rect 53340 45780 53396 47406
rect 53676 47458 53732 48078
rect 53676 47406 53678 47458
rect 53730 47406 53732 47458
rect 53676 47394 53732 47406
rect 53788 47012 53844 49308
rect 55244 49026 55300 50428
rect 55804 49924 55860 49934
rect 55244 48974 55246 49026
rect 55298 48974 55300 49026
rect 55244 48962 55300 48974
rect 55580 49810 55636 49822
rect 55580 49758 55582 49810
rect 55634 49758 55636 49810
rect 55244 47570 55300 47582
rect 55244 47518 55246 47570
rect 55298 47518 55300 47570
rect 54124 47460 54180 47470
rect 55244 47460 55300 47518
rect 54124 47458 55300 47460
rect 54124 47406 54126 47458
rect 54178 47406 55300 47458
rect 54124 47404 55300 47406
rect 54124 47394 54180 47404
rect 53900 47348 53956 47358
rect 53900 47254 53956 47292
rect 53564 46956 53844 47012
rect 54012 47234 54068 47246
rect 54012 47182 54014 47234
rect 54066 47182 54068 47234
rect 53452 45892 53508 45902
rect 53452 45798 53508 45836
rect 53340 45714 53396 45724
rect 53564 45444 53620 46956
rect 54012 45890 54068 47182
rect 54236 47234 54292 47246
rect 54236 47182 54238 47234
rect 54290 47182 54292 47234
rect 54236 47012 54292 47182
rect 55244 47068 55300 47404
rect 55580 47348 55636 49758
rect 55804 49810 55860 49868
rect 55804 49758 55806 49810
rect 55858 49758 55860 49810
rect 55804 49746 55860 49758
rect 55916 49140 55972 51214
rect 56028 51154 56084 51166
rect 56028 51102 56030 51154
rect 56082 51102 56084 51154
rect 56028 49922 56084 51102
rect 56028 49870 56030 49922
rect 56082 49870 56084 49922
rect 56028 49858 56084 49870
rect 56028 49140 56084 49150
rect 55916 49138 56084 49140
rect 55916 49086 56030 49138
rect 56082 49086 56084 49138
rect 55916 49084 56084 49086
rect 56028 49074 56084 49084
rect 55580 47282 55636 47292
rect 55244 47012 55524 47068
rect 54236 46946 54292 46956
rect 54012 45838 54014 45890
rect 54066 45838 54068 45890
rect 54012 45826 54068 45838
rect 54124 46786 54180 46798
rect 54124 46734 54126 46786
rect 54178 46734 54180 46786
rect 53900 45780 53956 45790
rect 53900 45686 53956 45724
rect 54124 45778 54180 46734
rect 55468 46788 55524 47012
rect 55468 46694 55524 46732
rect 55692 47012 55748 47022
rect 54684 46676 54740 46686
rect 55020 46676 55076 46686
rect 54124 45726 54126 45778
rect 54178 45726 54180 45778
rect 54124 45714 54180 45726
rect 54236 46674 54740 46676
rect 54236 46622 54686 46674
rect 54738 46622 54740 46674
rect 54236 46620 54740 46622
rect 53564 44322 53620 45388
rect 53564 44270 53566 44322
rect 53618 44270 53620 44322
rect 53564 44258 53620 44270
rect 53676 45668 53732 45678
rect 53676 44434 53732 45612
rect 54012 45556 54068 45566
rect 54068 45500 54180 45556
rect 54012 45490 54068 45500
rect 53676 44382 53678 44434
rect 53730 44382 53732 44434
rect 53116 43486 53118 43538
rect 53170 43486 53172 43538
rect 53116 43474 53172 43486
rect 52780 42926 52782 42978
rect 52834 42926 52836 42978
rect 52780 42914 52836 42926
rect 52892 42756 52948 42766
rect 53228 42756 53284 42766
rect 52948 42754 53284 42756
rect 52948 42702 53230 42754
rect 53282 42702 53284 42754
rect 52948 42700 53284 42702
rect 52892 42662 52948 42700
rect 53228 42690 53284 42700
rect 52780 42644 52836 42654
rect 52780 42550 52836 42588
rect 53340 42642 53396 42654
rect 53340 42590 53342 42642
rect 53394 42590 53396 42642
rect 51884 41906 51940 41916
rect 52108 42140 52276 42196
rect 51772 41860 51828 41870
rect 51772 41766 51828 41804
rect 51548 41134 51550 41186
rect 51602 41134 51604 41186
rect 51548 41122 51604 41134
rect 51660 41188 51716 41198
rect 51660 41074 51716 41132
rect 51660 41022 51662 41074
rect 51714 41022 51716 41074
rect 51660 41010 51716 41022
rect 51884 40964 51940 40974
rect 51884 40870 51940 40908
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 50428 40338 50484 40348
rect 51884 40404 51940 40414
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 49980 38722 50148 38724
rect 49980 38670 49982 38722
rect 50034 38670 50148 38722
rect 49980 38668 50148 38670
rect 49756 37604 49812 37614
rect 49980 37604 50036 38668
rect 50540 38052 50596 38062
rect 50540 37958 50596 37996
rect 51884 38052 51940 40348
rect 52108 39956 52164 42140
rect 52220 41970 52276 41982
rect 52220 41918 52222 41970
rect 52274 41918 52276 41970
rect 52220 40180 52276 41918
rect 52892 41860 52948 41870
rect 53340 41860 53396 42590
rect 52892 41858 53060 41860
rect 52892 41806 52894 41858
rect 52946 41806 53060 41858
rect 52892 41804 53060 41806
rect 52892 41794 52948 41804
rect 52332 41188 52388 41198
rect 52388 41132 52500 41188
rect 52332 41122 52388 41132
rect 52332 40628 52388 40638
rect 52332 40534 52388 40572
rect 52220 40114 52276 40124
rect 52108 39890 52164 39900
rect 52444 39620 52500 41132
rect 52668 41186 52724 41198
rect 52668 41134 52670 41186
rect 52722 41134 52724 41186
rect 52556 40964 52612 40974
rect 52556 40180 52612 40908
rect 52668 40404 52724 41134
rect 52668 40338 52724 40348
rect 52780 40628 52836 40638
rect 52780 40402 52836 40572
rect 53004 40514 53060 41804
rect 53340 41794 53396 41804
rect 53004 40462 53006 40514
rect 53058 40462 53060 40514
rect 53004 40450 53060 40462
rect 53676 40516 53732 44382
rect 53900 45108 53956 45118
rect 53900 43426 53956 45052
rect 54124 44884 54180 45500
rect 54236 45108 54292 46620
rect 54684 46610 54740 46620
rect 54908 46674 55076 46676
rect 54908 46622 55022 46674
rect 55074 46622 55076 46674
rect 54908 46620 55076 46622
rect 54348 45892 54404 45902
rect 54348 45332 54404 45836
rect 54460 45890 54516 45902
rect 54460 45838 54462 45890
rect 54514 45838 54516 45890
rect 54460 45444 54516 45838
rect 54796 45780 54852 45790
rect 54572 45668 54628 45678
rect 54572 45574 54628 45612
rect 54796 45666 54852 45724
rect 54796 45614 54798 45666
rect 54850 45614 54852 45666
rect 54796 45602 54852 45614
rect 54572 45444 54628 45454
rect 54460 45388 54572 45444
rect 54572 45378 54628 45388
rect 54908 45332 54964 46620
rect 55020 46610 55076 46620
rect 55244 46676 55300 46686
rect 55244 46582 55300 46620
rect 55692 46676 55748 46956
rect 55692 46674 55860 46676
rect 55692 46622 55694 46674
rect 55746 46622 55860 46674
rect 55692 46620 55860 46622
rect 55692 46610 55748 46620
rect 55356 46564 55412 46574
rect 55356 46470 55412 46508
rect 55692 45890 55748 45902
rect 55692 45838 55694 45890
rect 55746 45838 55748 45890
rect 54348 45276 54516 45332
rect 54236 45042 54292 45052
rect 54124 44828 54404 44884
rect 54348 44322 54404 44828
rect 54348 44270 54350 44322
rect 54402 44270 54404 44322
rect 54348 44258 54404 44270
rect 54460 44210 54516 45276
rect 54684 45276 54964 45332
rect 55580 45778 55636 45790
rect 55580 45726 55582 45778
rect 55634 45726 55636 45778
rect 54684 44322 54740 45276
rect 55244 45220 55300 45230
rect 54684 44270 54686 44322
rect 54738 44270 54740 44322
rect 54684 44258 54740 44270
rect 54908 45108 54964 45118
rect 54460 44158 54462 44210
rect 54514 44158 54516 44210
rect 54460 44146 54516 44158
rect 53900 43374 53902 43426
rect 53954 43374 53956 43426
rect 53900 43362 53956 43374
rect 54460 43876 54516 43886
rect 54460 43314 54516 43820
rect 54572 43764 54628 43774
rect 54572 43538 54628 43708
rect 54908 43650 54964 45052
rect 55244 44322 55300 45164
rect 55244 44270 55246 44322
rect 55298 44270 55300 44322
rect 55244 44258 55300 44270
rect 55580 44100 55636 45726
rect 54908 43598 54910 43650
rect 54962 43598 54964 43650
rect 54908 43586 54964 43598
rect 55020 44044 55636 44100
rect 55020 43650 55076 44044
rect 55468 43876 55524 43886
rect 55020 43598 55022 43650
rect 55074 43598 55076 43650
rect 55020 43586 55076 43598
rect 55132 43764 55188 43774
rect 54572 43486 54574 43538
rect 54626 43486 54628 43538
rect 54572 43474 54628 43486
rect 54460 43262 54462 43314
rect 54514 43262 54516 43314
rect 54236 40628 54292 40638
rect 54236 40534 54292 40572
rect 53676 40450 53732 40460
rect 52780 40350 52782 40402
rect 52834 40350 52836 40402
rect 52668 40180 52724 40190
rect 52556 40178 52724 40180
rect 52556 40126 52670 40178
rect 52722 40126 52724 40178
rect 52556 40124 52724 40126
rect 52668 40114 52724 40124
rect 52668 39732 52724 39742
rect 52668 39620 52724 39676
rect 52444 39618 52724 39620
rect 52444 39566 52670 39618
rect 52722 39566 52724 39618
rect 52444 39564 52724 39566
rect 52668 39554 52724 39564
rect 52668 39060 52724 39070
rect 52108 38724 52164 38734
rect 52108 38630 52164 38668
rect 49812 37548 50036 37604
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 49756 37538 49812 37548
rect 49308 37326 49310 37378
rect 49362 37326 49364 37378
rect 49308 37314 49364 37326
rect 48972 37214 48974 37266
rect 49026 37214 49028 37266
rect 48972 37156 49028 37214
rect 48972 37090 49028 37100
rect 49756 37154 49812 37166
rect 49756 37102 49758 37154
rect 49810 37102 49812 37154
rect 49644 37044 49700 37054
rect 49420 37042 49700 37044
rect 49420 36990 49646 37042
rect 49698 36990 49700 37042
rect 49420 36988 49700 36990
rect 49420 36594 49476 36988
rect 49644 36978 49700 36988
rect 49420 36542 49422 36594
rect 49474 36542 49476 36594
rect 49420 36530 49476 36542
rect 48748 36484 48804 36494
rect 48804 36428 49028 36484
rect 48748 36390 48804 36428
rect 48972 35812 49028 36428
rect 48972 35718 49028 35756
rect 49644 36260 49700 36270
rect 49644 34914 49700 36204
rect 49756 35026 49812 37102
rect 51884 37044 51940 37996
rect 51884 36988 52276 37044
rect 51548 36594 51604 36606
rect 51548 36542 51550 36594
rect 51602 36542 51604 36594
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 51212 35812 51268 35822
rect 49756 34974 49758 35026
rect 49810 34974 49812 35026
rect 49756 34962 49812 34974
rect 49980 35364 50036 35374
rect 49644 34862 49646 34914
rect 49698 34862 49700 34914
rect 49644 34850 49700 34862
rect 49980 34914 50036 35308
rect 49980 34862 49982 34914
rect 50034 34862 50036 34914
rect 49980 34850 50036 34862
rect 50204 34916 50260 34926
rect 50204 34822 50260 34860
rect 50764 34916 50820 34926
rect 50820 34860 50932 34916
rect 50764 34850 50820 34860
rect 48412 34690 48692 34692
rect 48412 34638 48414 34690
rect 48466 34638 48692 34690
rect 48412 34636 48692 34638
rect 49196 34692 49252 34702
rect 49756 34692 49812 34702
rect 49196 34690 49812 34692
rect 49196 34638 49198 34690
rect 49250 34638 49758 34690
rect 49810 34638 49812 34690
rect 49196 34636 49812 34638
rect 48412 31780 48468 34636
rect 49196 34132 49252 34636
rect 49756 34626 49812 34636
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 48972 34076 49196 34132
rect 48412 31714 48468 31724
rect 48636 32564 48692 32574
rect 48636 31778 48692 32508
rect 48636 31726 48638 31778
rect 48690 31726 48692 31778
rect 48636 31714 48692 31726
rect 48748 32452 48804 32462
rect 48748 31778 48804 32396
rect 48748 31726 48750 31778
rect 48802 31726 48804 31778
rect 48748 31714 48804 31726
rect 48412 31554 48468 31566
rect 48412 31502 48414 31554
rect 48466 31502 48468 31554
rect 48412 30996 48468 31502
rect 48412 30930 48468 30940
rect 48524 31554 48580 31566
rect 48524 31502 48526 31554
rect 48578 31502 48580 31554
rect 48524 30212 48580 31502
rect 48972 31332 49028 34076
rect 49196 34066 49252 34076
rect 49532 33458 49588 33470
rect 49532 33406 49534 33458
rect 49586 33406 49588 33458
rect 49532 33236 49588 33406
rect 50764 33460 50820 33470
rect 50876 33460 50932 34860
rect 51212 34130 51268 35756
rect 51548 34916 51604 36542
rect 52108 36596 52164 36606
rect 52108 36502 52164 36540
rect 51996 36258 52052 36270
rect 51996 36206 51998 36258
rect 52050 36206 52052 36258
rect 51604 34860 51716 34916
rect 51548 34850 51604 34860
rect 51212 34078 51214 34130
rect 51266 34078 51268 34130
rect 51212 34066 51268 34078
rect 50764 33458 50932 33460
rect 50764 33406 50766 33458
rect 50818 33406 50932 33458
rect 50764 33404 50932 33406
rect 50764 33394 50820 33404
rect 49980 33236 50036 33246
rect 49532 33234 50036 33236
rect 49532 33182 49982 33234
rect 50034 33182 50036 33234
rect 49532 33180 50036 33182
rect 49196 32676 49252 32686
rect 49532 32676 49588 33180
rect 49980 33170 50036 33180
rect 50316 33236 50372 33246
rect 49196 32674 49588 32676
rect 49196 32622 49198 32674
rect 49250 32622 49588 32674
rect 49196 32620 49588 32622
rect 50316 32674 50372 33180
rect 50876 33122 50932 33134
rect 50876 33070 50878 33122
rect 50930 33070 50932 33122
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 50764 32788 50820 32798
rect 50764 32694 50820 32732
rect 50876 32786 50932 33070
rect 50876 32734 50878 32786
rect 50930 32734 50932 32786
rect 50876 32722 50932 32734
rect 51660 32788 51716 34860
rect 51996 34242 52052 36206
rect 52220 35028 52276 36988
rect 52668 36820 52724 39004
rect 52780 38668 52836 40350
rect 53228 40404 53284 40414
rect 53228 40310 53284 40348
rect 54460 40404 54516 43262
rect 55132 42756 55188 43708
rect 55020 42700 55188 42756
rect 55020 41858 55076 42700
rect 55356 42644 55412 42654
rect 55244 42642 55412 42644
rect 55244 42590 55358 42642
rect 55410 42590 55412 42642
rect 55244 42588 55412 42590
rect 55132 42530 55188 42542
rect 55132 42478 55134 42530
rect 55186 42478 55188 42530
rect 55132 41972 55188 42478
rect 55132 41906 55188 41916
rect 55020 41806 55022 41858
rect 55074 41806 55076 41858
rect 55020 41794 55076 41806
rect 55244 41412 55300 42588
rect 55356 42578 55412 42588
rect 54908 41356 55300 41412
rect 54908 40626 54964 41356
rect 55468 41300 55524 43820
rect 55692 43764 55748 45838
rect 55692 43698 55748 43708
rect 55804 43708 55860 46620
rect 56140 45892 56196 52220
rect 56252 48356 56308 53454
rect 56812 53508 56868 53518
rect 56588 52948 56644 52958
rect 56588 49924 56644 52892
rect 56812 52946 56868 53452
rect 56812 52894 56814 52946
rect 56866 52894 56868 52946
rect 56812 52882 56868 52894
rect 57036 52722 57092 52734
rect 57036 52670 57038 52722
rect 57090 52670 57092 52722
rect 57036 51940 57092 52670
rect 57148 52724 57204 52734
rect 57148 52722 57428 52724
rect 57148 52670 57150 52722
rect 57202 52670 57428 52722
rect 57148 52668 57428 52670
rect 57148 52658 57204 52668
rect 57372 52274 57428 52668
rect 57372 52222 57374 52274
rect 57426 52222 57428 52274
rect 57372 52210 57428 52222
rect 57036 51874 57092 51884
rect 57372 50260 57428 50270
rect 57372 50034 57428 50204
rect 57372 49982 57374 50034
rect 57426 49982 57428 50034
rect 57372 49970 57428 49982
rect 57484 50036 57540 55022
rect 58044 52162 58100 52174
rect 58044 52110 58046 52162
rect 58098 52110 58100 52162
rect 57484 49970 57540 49980
rect 57932 50484 57988 50494
rect 58044 50484 58100 52110
rect 57988 50428 58100 50484
rect 56588 49830 56644 49868
rect 56700 49922 56756 49934
rect 56700 49870 56702 49922
rect 56754 49870 56756 49922
rect 56700 49252 56756 49870
rect 56588 48356 56644 48366
rect 56252 48354 56644 48356
rect 56252 48302 56590 48354
rect 56642 48302 56644 48354
rect 56252 48300 56644 48302
rect 56588 48290 56644 48300
rect 56364 47348 56420 47358
rect 56420 47292 56644 47348
rect 56364 47282 56420 47292
rect 56588 46898 56644 47292
rect 56588 46846 56590 46898
rect 56642 46846 56644 46898
rect 56588 46452 56644 46846
rect 56700 46786 56756 49196
rect 56924 49810 56980 49822
rect 56924 49758 56926 49810
rect 56978 49758 56980 49810
rect 56924 48356 56980 49758
rect 57596 49812 57652 49822
rect 57596 49718 57652 49756
rect 57148 48356 57204 48366
rect 56924 48354 57204 48356
rect 56924 48302 57150 48354
rect 57202 48302 57204 48354
rect 56924 48300 57204 48302
rect 57148 48290 57204 48300
rect 56812 48242 56868 48254
rect 56812 48190 56814 48242
rect 56866 48190 56868 48242
rect 56812 47012 56868 48190
rect 57036 48130 57092 48142
rect 57036 48078 57038 48130
rect 57090 48078 57092 48130
rect 57036 47796 57092 48078
rect 57036 47740 57428 47796
rect 57372 47570 57428 47740
rect 57372 47518 57374 47570
rect 57426 47518 57428 47570
rect 57372 47506 57428 47518
rect 57932 47460 57988 50428
rect 58156 50260 58212 50270
rect 58156 50034 58212 50204
rect 58156 49982 58158 50034
rect 58210 49982 58212 50034
rect 58156 49970 58212 49982
rect 58156 49252 58212 49262
rect 58156 49138 58212 49196
rect 58156 49086 58158 49138
rect 58210 49086 58212 49138
rect 58156 49074 58212 49086
rect 58044 47460 58100 47470
rect 57932 47458 58100 47460
rect 57932 47406 58046 47458
rect 58098 47406 58100 47458
rect 57932 47404 58100 47406
rect 58044 47394 58100 47404
rect 56812 46956 57204 47012
rect 57148 46900 57204 46956
rect 57148 46898 57428 46900
rect 57148 46846 57150 46898
rect 57202 46846 57428 46898
rect 57148 46844 57428 46846
rect 57148 46834 57204 46844
rect 56700 46734 56702 46786
rect 56754 46734 56756 46786
rect 56700 46676 56756 46734
rect 57036 46788 57092 46798
rect 57036 46694 57092 46732
rect 56700 46610 56756 46620
rect 57260 46676 57316 46686
rect 56588 46396 56756 46452
rect 56252 45892 56308 45902
rect 56140 45890 56308 45892
rect 56140 45838 56254 45890
rect 56306 45838 56308 45890
rect 56140 45836 56308 45838
rect 56140 45108 56196 45836
rect 56252 45826 56308 45836
rect 56140 45042 56196 45052
rect 56364 45666 56420 45678
rect 56364 45614 56366 45666
rect 56418 45614 56420 45666
rect 56028 44210 56084 44222
rect 56028 44158 56030 44210
rect 56082 44158 56084 44210
rect 56028 43708 56084 44158
rect 56364 43988 56420 45614
rect 56588 45668 56644 45678
rect 56588 45574 56644 45612
rect 56700 45106 56756 46396
rect 57148 45890 57204 45902
rect 57148 45838 57150 45890
rect 57202 45838 57204 45890
rect 56700 45054 56702 45106
rect 56754 45054 56756 45106
rect 56700 45042 56756 45054
rect 56812 45218 56868 45230
rect 56812 45166 56814 45218
rect 56866 45166 56868 45218
rect 56364 43922 56420 43932
rect 56812 43708 56868 45166
rect 57148 44436 57204 45838
rect 57260 45778 57316 46620
rect 57372 46452 57428 46844
rect 58156 46674 58212 46686
rect 58156 46622 58158 46674
rect 58210 46622 58212 46674
rect 57708 46562 57764 46574
rect 57708 46510 57710 46562
rect 57762 46510 57764 46562
rect 57372 46396 57652 46452
rect 57260 45726 57262 45778
rect 57314 45726 57316 45778
rect 57260 45714 57316 45726
rect 57484 46116 57540 46126
rect 57484 45330 57540 46060
rect 57484 45278 57486 45330
rect 57538 45278 57540 45330
rect 57484 45266 57540 45278
rect 57596 45218 57652 46396
rect 57596 45166 57598 45218
rect 57650 45166 57652 45218
rect 57596 45154 57652 45166
rect 55804 43652 55972 43708
rect 56028 43652 56308 43708
rect 55916 43316 55972 43652
rect 56140 43316 56196 43326
rect 55916 43260 56140 43316
rect 55916 42978 55972 43260
rect 56140 43250 56196 43260
rect 55916 42926 55918 42978
rect 55970 42926 55972 42978
rect 55916 42914 55972 42926
rect 56140 42754 56196 42766
rect 56140 42702 56142 42754
rect 56194 42702 56196 42754
rect 55580 42642 55636 42654
rect 55580 42590 55582 42642
rect 55634 42590 55636 42642
rect 55580 41972 55636 42590
rect 55636 41916 55748 41972
rect 55580 41906 55636 41916
rect 55468 41244 55636 41300
rect 54908 40574 54910 40626
rect 54962 40574 54964 40626
rect 54908 40562 54964 40574
rect 55468 41074 55524 41086
rect 55468 41022 55470 41074
rect 55522 41022 55524 41074
rect 54684 40516 54740 40526
rect 54684 40514 54852 40516
rect 54684 40462 54686 40514
rect 54738 40462 54852 40514
rect 54684 40460 54852 40462
rect 54684 40450 54740 40460
rect 54460 40338 54516 40348
rect 54572 40402 54628 40414
rect 54572 40350 54574 40402
rect 54626 40350 54628 40402
rect 53452 40292 53508 40302
rect 53452 40198 53508 40236
rect 52892 40180 52948 40190
rect 52892 39620 52948 40124
rect 54348 40068 54404 40078
rect 52892 38834 52948 39564
rect 53116 39730 53172 39742
rect 53116 39678 53118 39730
rect 53170 39678 53172 39730
rect 53116 39060 53172 39678
rect 53676 39732 53732 39742
rect 54348 39732 54404 40012
rect 53676 39638 53732 39676
rect 54236 39730 54404 39732
rect 54236 39678 54350 39730
rect 54402 39678 54404 39730
rect 54236 39676 54404 39678
rect 53116 38994 53172 39004
rect 52892 38782 52894 38834
rect 52946 38782 52948 38834
rect 52892 38770 52948 38782
rect 52780 38612 53060 38668
rect 52668 36764 52948 36820
rect 52780 36596 52836 36606
rect 52780 36502 52836 36540
rect 52780 36372 52836 36382
rect 52668 36370 52836 36372
rect 52668 36318 52782 36370
rect 52834 36318 52836 36370
rect 52668 36316 52836 36318
rect 52668 36260 52724 36316
rect 52780 36306 52836 36316
rect 52892 36372 52948 36764
rect 52668 36194 52724 36204
rect 52892 36258 52948 36316
rect 52892 36206 52894 36258
rect 52946 36206 52948 36258
rect 52892 35924 52948 36206
rect 52108 34972 52220 35028
rect 52108 34914 52164 34972
rect 52220 34962 52276 34972
rect 52332 35868 52948 35924
rect 52108 34862 52110 34914
rect 52162 34862 52164 34914
rect 52108 34850 52164 34862
rect 51996 34190 51998 34242
rect 52050 34190 52052 34242
rect 51996 34178 52052 34190
rect 52220 34020 52276 34030
rect 51884 33348 51940 33358
rect 51772 32788 51828 32798
rect 51660 32786 51828 32788
rect 51660 32734 51774 32786
rect 51826 32734 51828 32786
rect 51660 32732 51828 32734
rect 51772 32722 51828 32732
rect 51884 32788 51940 33292
rect 52108 33124 52164 33134
rect 52108 33030 52164 33068
rect 51884 32722 51940 32732
rect 50316 32622 50318 32674
rect 50370 32622 50372 32674
rect 49196 32610 49252 32620
rect 50316 32610 50372 32622
rect 51996 32676 52052 32686
rect 51996 32582 52052 32620
rect 49084 32564 49140 32574
rect 49084 32470 49140 32508
rect 49756 32564 49812 32574
rect 49756 32470 49812 32508
rect 50540 32564 50596 32574
rect 50540 32470 50596 32508
rect 51660 32564 51716 32574
rect 51660 32470 51716 32508
rect 52220 32562 52276 33964
rect 52220 32510 52222 32562
rect 52274 32510 52276 32562
rect 52220 32498 52276 32510
rect 49644 32452 49700 32462
rect 49644 32358 49700 32396
rect 50876 32450 50932 32462
rect 50876 32398 50878 32450
rect 50930 32398 50932 32450
rect 49532 31892 49588 31902
rect 49532 31666 49588 31836
rect 49532 31614 49534 31666
rect 49586 31614 49588 31666
rect 49532 31602 49588 31614
rect 49196 31556 49252 31566
rect 49196 31462 49252 31500
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 48972 31276 49252 31332
rect 50556 31322 50820 31332
rect 48748 31220 48804 31230
rect 48748 31106 48804 31164
rect 48748 31054 48750 31106
rect 48802 31054 48804 31106
rect 48748 31042 48804 31054
rect 48972 30996 49028 31006
rect 48972 30902 49028 30940
rect 48524 30146 48580 30156
rect 48524 29428 48580 29438
rect 48524 28754 48580 29372
rect 48524 28702 48526 28754
rect 48578 28702 48580 28754
rect 48524 28690 48580 28702
rect 48412 28420 48468 28430
rect 48412 28326 48468 28364
rect 48636 28418 48692 28430
rect 48636 28366 48638 28418
rect 48690 28366 48692 28418
rect 48636 28308 48692 28366
rect 48636 26964 48692 28252
rect 48636 26898 48692 26908
rect 49196 25956 49252 31276
rect 49308 30772 49364 30782
rect 49308 30678 49364 30716
rect 49532 30212 49588 30222
rect 49532 29540 49588 30156
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 49644 29652 49700 29662
rect 49644 29558 49700 29596
rect 49308 29428 49364 29438
rect 49532 29428 49588 29484
rect 50764 29540 50820 29550
rect 50764 29446 50820 29484
rect 50876 29540 50932 32398
rect 51884 32450 51940 32462
rect 51884 32398 51886 32450
rect 51938 32398 51940 32450
rect 51884 30660 51940 32398
rect 52332 32452 52388 35868
rect 52892 35698 52948 35710
rect 52892 35646 52894 35698
rect 52946 35646 52948 35698
rect 52892 35028 52948 35646
rect 52892 34914 52948 34972
rect 52892 34862 52894 34914
rect 52946 34862 52948 34914
rect 52892 34850 52948 34862
rect 53004 33572 53060 38612
rect 53116 37154 53172 37166
rect 53116 37102 53118 37154
rect 53170 37102 53172 37154
rect 53116 37044 53172 37102
rect 53116 36978 53172 36988
rect 53900 37044 53956 37054
rect 53900 36482 53956 36988
rect 53900 36430 53902 36482
rect 53954 36430 53956 36482
rect 53340 36370 53396 36382
rect 53340 36318 53342 36370
rect 53394 36318 53396 36370
rect 53116 36258 53172 36270
rect 53116 36206 53118 36258
rect 53170 36206 53172 36258
rect 53116 36148 53172 36206
rect 53116 35364 53172 36092
rect 53116 35298 53172 35308
rect 53340 34020 53396 36318
rect 53396 33964 53508 34020
rect 53340 33954 53396 33964
rect 53004 33506 53060 33516
rect 53004 33348 53060 33358
rect 53340 33348 53396 33358
rect 53004 33346 53396 33348
rect 53004 33294 53006 33346
rect 53058 33294 53342 33346
rect 53394 33294 53396 33346
rect 53004 33292 53396 33294
rect 53004 33282 53060 33292
rect 53340 33282 53396 33292
rect 52668 33234 52724 33246
rect 52668 33182 52670 33234
rect 52722 33182 52724 33234
rect 52556 33124 52612 33134
rect 52556 32788 52612 33068
rect 52668 32900 52724 33182
rect 52780 33236 52836 33246
rect 52780 33012 52836 33180
rect 52780 32956 53060 33012
rect 52668 32844 52948 32900
rect 52556 32732 52724 32788
rect 52668 32676 52724 32732
rect 52668 32674 52836 32676
rect 52668 32622 52670 32674
rect 52722 32622 52836 32674
rect 52668 32620 52836 32622
rect 52668 32610 52724 32620
rect 52556 32564 52612 32574
rect 52556 32470 52612 32508
rect 52332 32386 52388 32396
rect 52668 31892 52724 31902
rect 52668 30996 52724 31836
rect 52780 31666 52836 32620
rect 52892 32564 52948 32844
rect 52892 32340 52948 32508
rect 52892 32274 52948 32284
rect 53004 32788 53060 32956
rect 53004 31778 53060 32732
rect 53004 31726 53006 31778
rect 53058 31726 53060 31778
rect 53004 31714 53060 31726
rect 53116 32676 53172 32686
rect 53116 32562 53172 32620
rect 53116 32510 53118 32562
rect 53170 32510 53172 32562
rect 52780 31614 52782 31666
rect 52834 31614 52836 31666
rect 52780 31602 52836 31614
rect 52892 31220 52948 31230
rect 53116 31220 53172 32510
rect 53340 32340 53396 32350
rect 53340 32246 53396 32284
rect 53228 31780 53284 31790
rect 53228 31686 53284 31724
rect 52892 31218 53172 31220
rect 52892 31166 52894 31218
rect 52946 31166 53172 31218
rect 52892 31164 53172 31166
rect 52892 31154 52948 31164
rect 53340 31108 53396 31118
rect 53452 31108 53508 33964
rect 53564 33346 53620 33358
rect 53564 33294 53566 33346
rect 53618 33294 53620 33346
rect 53564 33124 53620 33294
rect 53900 33236 53956 36430
rect 54012 36258 54068 36270
rect 54012 36206 54014 36258
rect 54066 36206 54068 36258
rect 54012 36148 54068 36206
rect 54012 36082 54068 36092
rect 54236 36258 54292 39676
rect 54348 39666 54404 39676
rect 54572 39396 54628 40350
rect 54796 40180 54852 40460
rect 55468 40404 55524 41022
rect 55356 40348 55524 40404
rect 55244 40292 55300 40302
rect 55244 40198 55300 40236
rect 54796 39618 54852 40124
rect 54908 39732 54964 39742
rect 54964 39676 55076 39732
rect 54908 39666 54964 39676
rect 54796 39566 54798 39618
rect 54850 39566 54852 39618
rect 54796 39554 54852 39566
rect 54572 39172 54628 39340
rect 54572 39106 54628 39116
rect 54908 39508 54964 39518
rect 54908 38836 54964 39452
rect 54684 38834 54964 38836
rect 54684 38782 54910 38834
rect 54962 38782 54964 38834
rect 54684 38780 54964 38782
rect 54460 38276 54516 38286
rect 54460 37826 54516 38220
rect 54460 37774 54462 37826
rect 54514 37774 54516 37826
rect 54460 37762 54516 37774
rect 54348 37044 54404 37054
rect 54348 36594 54404 36988
rect 54348 36542 54350 36594
rect 54402 36542 54404 36594
rect 54348 36530 54404 36542
rect 54236 36206 54238 36258
rect 54290 36206 54292 36258
rect 54236 35364 54292 36206
rect 54348 36260 54404 36270
rect 54404 36204 54516 36260
rect 54348 36166 54404 36204
rect 54460 35698 54516 36204
rect 54460 35646 54462 35698
rect 54514 35646 54516 35698
rect 54460 35634 54516 35646
rect 54684 35700 54740 38780
rect 54908 38770 54964 38780
rect 55020 38668 55076 39676
rect 55244 39620 55300 39630
rect 55356 39620 55412 40348
rect 55468 40180 55524 40190
rect 55580 40180 55636 41244
rect 55692 40628 55748 41916
rect 55692 40516 55748 40572
rect 55804 40516 55860 40526
rect 55692 40514 55860 40516
rect 55692 40462 55806 40514
rect 55858 40462 55860 40514
rect 55692 40460 55860 40462
rect 55804 40450 55860 40460
rect 56140 40404 56196 42702
rect 56252 42530 56308 43652
rect 56700 43652 56868 43708
rect 56924 44380 57204 44436
rect 57484 45106 57540 45118
rect 57484 45054 57486 45106
rect 57538 45054 57540 45106
rect 57484 44436 57540 45054
rect 56924 43876 56980 44380
rect 56700 42644 56756 43652
rect 56924 43540 56980 43820
rect 57484 43708 57540 44380
rect 57036 43652 57540 43708
rect 57036 43650 57092 43652
rect 57036 43598 57038 43650
rect 57090 43598 57092 43650
rect 57036 43586 57092 43598
rect 56812 43484 56980 43540
rect 56812 42980 56868 43484
rect 56924 43316 56980 43326
rect 56924 43222 56980 43260
rect 56924 42980 56980 42990
rect 56812 42978 56980 42980
rect 56812 42926 56926 42978
rect 56978 42926 56980 42978
rect 56812 42924 56980 42926
rect 56924 42914 56980 42924
rect 56812 42644 56868 42654
rect 56700 42642 56868 42644
rect 56700 42590 56814 42642
rect 56866 42590 56868 42642
rect 56700 42588 56868 42590
rect 56252 42478 56254 42530
rect 56306 42478 56308 42530
rect 56252 42466 56308 42478
rect 56812 41972 56868 42588
rect 56812 41906 56868 41916
rect 57708 40628 57764 46510
rect 58156 45668 58212 46622
rect 58156 45666 58324 45668
rect 58156 45614 58158 45666
rect 58210 45614 58324 45666
rect 58156 45612 58324 45614
rect 58156 45602 58212 45612
rect 58268 44548 58324 45612
rect 58268 44482 58324 44492
rect 58156 44436 58212 44446
rect 58156 44342 58212 44380
rect 56140 40338 56196 40348
rect 57484 40572 57764 40628
rect 58156 41972 58212 41982
rect 55468 40178 55636 40180
rect 55468 40126 55470 40178
rect 55522 40126 55636 40178
rect 55468 40124 55636 40126
rect 55916 40178 55972 40190
rect 55916 40126 55918 40178
rect 55970 40126 55972 40178
rect 55468 40114 55524 40124
rect 55916 39732 55972 40126
rect 56028 40180 56084 40190
rect 57484 40180 57540 40572
rect 57820 40514 57876 40526
rect 57820 40462 57822 40514
rect 57874 40462 57876 40514
rect 57596 40402 57652 40414
rect 57596 40350 57598 40402
rect 57650 40350 57652 40402
rect 57596 40292 57652 40350
rect 57596 40226 57652 40236
rect 56028 40178 56196 40180
rect 56028 40126 56030 40178
rect 56082 40126 56196 40178
rect 56028 40124 56196 40126
rect 56028 40114 56084 40124
rect 56028 39732 56084 39742
rect 55916 39730 56084 39732
rect 55916 39678 56030 39730
rect 56082 39678 56084 39730
rect 55916 39676 56084 39678
rect 56028 39666 56084 39676
rect 55300 39564 55412 39620
rect 55244 39526 55300 39564
rect 55804 39172 55860 39182
rect 55468 39060 55524 39070
rect 55468 38966 55524 39004
rect 55804 38946 55860 39116
rect 55804 38894 55806 38946
rect 55858 38894 55860 38946
rect 55804 38882 55860 38894
rect 55916 39060 55972 39070
rect 54908 38612 55076 38668
rect 54908 37938 54964 38612
rect 55916 38050 55972 39004
rect 56140 39058 56196 40124
rect 57484 40114 57540 40124
rect 56140 39006 56142 39058
rect 56194 39006 56196 39058
rect 56140 38994 56196 39006
rect 57820 39060 57876 40462
rect 57820 38994 57876 39004
rect 58044 40402 58100 40414
rect 58044 40350 58046 40402
rect 58098 40350 58100 40402
rect 58044 40292 58100 40350
rect 57708 38834 57764 38846
rect 57708 38782 57710 38834
rect 57762 38782 57764 38834
rect 57148 38722 57204 38734
rect 57148 38670 57150 38722
rect 57202 38670 57204 38722
rect 57148 38164 57204 38670
rect 57148 38098 57204 38108
rect 55916 37998 55918 38050
rect 55970 37998 55972 38050
rect 55916 37986 55972 37998
rect 54908 37886 54910 37938
rect 54962 37886 54964 37938
rect 54908 37268 54964 37886
rect 57708 37940 57764 38782
rect 58044 38724 58100 40236
rect 58156 39730 58212 41916
rect 58156 39678 58158 39730
rect 58210 39678 58212 39730
rect 58156 39666 58212 39678
rect 58268 40180 58324 40190
rect 58156 38724 58212 38734
rect 58044 38668 58156 38724
rect 58156 38658 58212 38668
rect 58156 38052 58212 38062
rect 58268 38052 58324 40124
rect 58156 38050 58324 38052
rect 58156 37998 58158 38050
rect 58210 37998 58324 38050
rect 58156 37996 58324 37998
rect 58156 37986 58212 37996
rect 58044 37940 58100 37950
rect 57708 37938 58100 37940
rect 57708 37886 58046 37938
rect 58098 37886 58100 37938
rect 57708 37884 58100 37886
rect 54908 37202 54964 37212
rect 56028 37266 56084 37278
rect 56028 37214 56030 37266
rect 56082 37214 56084 37266
rect 55244 37156 55300 37166
rect 55244 37062 55300 37100
rect 55356 36596 55412 36606
rect 55356 36482 55412 36540
rect 56028 36596 56084 37214
rect 57820 37268 57876 37278
rect 56588 37156 56644 37166
rect 56588 37062 56644 37100
rect 56700 37154 56756 37166
rect 56700 37102 56702 37154
rect 56754 37102 56756 37154
rect 56700 37044 56756 37102
rect 56700 36978 56756 36988
rect 57820 37042 57876 37212
rect 57820 36990 57822 37042
rect 57874 36990 57876 37042
rect 56028 36530 56084 36540
rect 55356 36430 55358 36482
rect 55410 36430 55412 36482
rect 54908 36372 54964 36382
rect 54908 36278 54964 36316
rect 54796 36148 54852 36158
rect 54796 35924 54852 36092
rect 54908 35924 54964 35934
rect 54796 35922 54964 35924
rect 54796 35870 54910 35922
rect 54962 35870 54964 35922
rect 54796 35868 54964 35870
rect 54908 35858 54964 35868
rect 55132 35812 55188 35822
rect 54236 35298 54292 35308
rect 54124 34020 54180 34030
rect 54124 33926 54180 33964
rect 54572 34018 54628 34030
rect 54572 33966 54574 34018
rect 54626 33966 54628 34018
rect 54572 33796 54628 33966
rect 54572 33730 54628 33740
rect 54236 33236 54292 33246
rect 54572 33236 54628 33246
rect 53900 33180 54180 33236
rect 53620 33068 54068 33124
rect 53564 33058 53620 33068
rect 54012 32786 54068 33068
rect 54012 32734 54014 32786
rect 54066 32734 54068 32786
rect 54012 32722 54068 32734
rect 53676 32338 53732 32350
rect 53676 32286 53678 32338
rect 53730 32286 53732 32338
rect 53676 31892 53732 32286
rect 53900 32340 53956 32350
rect 53900 32246 53956 32284
rect 54124 32116 54180 33180
rect 54236 33234 54628 33236
rect 54236 33182 54238 33234
rect 54290 33182 54574 33234
rect 54626 33182 54628 33234
rect 54236 33180 54628 33182
rect 54236 33170 54292 33180
rect 54572 33170 54628 33180
rect 54236 32788 54292 32798
rect 54236 32694 54292 32732
rect 54460 32564 54516 32574
rect 54460 32470 54516 32508
rect 54684 32116 54740 35644
rect 55020 35756 55132 35812
rect 54796 35588 54852 35598
rect 54796 35494 54852 35532
rect 54796 33796 54852 33806
rect 54852 33740 54964 33796
rect 54796 33730 54852 33740
rect 54796 33460 54852 33470
rect 54796 33366 54852 33404
rect 54908 33346 54964 33740
rect 54908 33294 54910 33346
rect 54962 33294 54964 33346
rect 54908 33282 54964 33294
rect 53676 31826 53732 31836
rect 53900 32060 54180 32116
rect 54236 32060 54740 32116
rect 53676 31668 53732 31678
rect 53676 31574 53732 31612
rect 53340 31106 53508 31108
rect 53340 31054 53342 31106
rect 53394 31054 53508 31106
rect 53340 31052 53508 31054
rect 53340 31042 53396 31052
rect 53004 30996 53060 31006
rect 52668 30994 53284 30996
rect 52668 30942 53006 30994
rect 53058 30942 53284 30994
rect 52668 30940 53284 30942
rect 53004 30930 53060 30940
rect 50988 30604 51940 30660
rect 50988 30210 51044 30604
rect 50988 30158 50990 30210
rect 51042 30158 51044 30210
rect 50988 29764 51044 30158
rect 52220 30324 52276 30334
rect 51100 29988 51156 29998
rect 51100 29986 51828 29988
rect 51100 29934 51102 29986
rect 51154 29934 51828 29986
rect 51100 29932 51828 29934
rect 51100 29922 51156 29932
rect 50988 29708 51156 29764
rect 50988 29540 51044 29550
rect 50876 29538 51044 29540
rect 50876 29486 50990 29538
rect 51042 29486 51044 29538
rect 50876 29484 51044 29486
rect 49644 29428 49700 29438
rect 49532 29426 49700 29428
rect 49532 29374 49646 29426
rect 49698 29374 49700 29426
rect 49532 29372 49700 29374
rect 49308 29334 49364 29372
rect 49644 29362 49700 29372
rect 49980 29428 50036 29438
rect 50652 29428 50708 29438
rect 49980 29426 50372 29428
rect 49980 29374 49982 29426
rect 50034 29374 50372 29426
rect 49980 29372 50372 29374
rect 49980 29362 50036 29372
rect 50204 29202 50260 29214
rect 50204 29150 50206 29202
rect 50258 29150 50260 29202
rect 49756 27132 50036 27188
rect 49756 27074 49812 27132
rect 49756 27022 49758 27074
rect 49810 27022 49812 27074
rect 49756 26908 49812 27022
rect 49196 25890 49252 25900
rect 49308 26852 49812 26908
rect 49868 26964 49924 27002
rect 49868 26898 49924 26908
rect 49308 25730 49364 26852
rect 49980 26290 50036 27132
rect 50204 27074 50260 29150
rect 50316 28866 50372 29372
rect 50652 29334 50708 29372
rect 50876 29204 50932 29484
rect 50988 29474 51044 29484
rect 51100 29426 51156 29708
rect 51548 29652 51604 29662
rect 51548 29558 51604 29596
rect 51772 29650 51828 29932
rect 51772 29598 51774 29650
rect 51826 29598 51828 29650
rect 51772 29586 51828 29598
rect 52220 29428 52276 30268
rect 53228 30212 53284 30940
rect 53452 30772 53508 30782
rect 53452 30770 53620 30772
rect 53452 30718 53454 30770
rect 53506 30718 53620 30770
rect 53452 30716 53620 30718
rect 53452 30706 53508 30716
rect 53340 30212 53396 30222
rect 53228 30210 53396 30212
rect 53228 30158 53342 30210
rect 53394 30158 53396 30210
rect 53228 30156 53396 30158
rect 53340 30146 53396 30156
rect 53564 30210 53620 30716
rect 53676 30324 53732 30334
rect 53676 30230 53732 30268
rect 53564 30158 53566 30210
rect 53618 30158 53620 30210
rect 53564 30146 53620 30158
rect 53788 29988 53844 29998
rect 53788 29894 53844 29932
rect 53900 29764 53956 32060
rect 54236 32004 54292 32060
rect 54124 31948 54292 32004
rect 54012 30212 54068 30222
rect 54012 30118 54068 30156
rect 53788 29708 53956 29764
rect 51100 29374 51102 29426
rect 51154 29374 51156 29426
rect 51100 29362 51156 29374
rect 52108 29426 52276 29428
rect 52108 29374 52222 29426
rect 52274 29374 52276 29426
rect 52108 29372 52276 29374
rect 50316 28814 50318 28866
rect 50370 28814 50372 28866
rect 50316 28802 50372 28814
rect 50428 29148 50932 29204
rect 51660 29314 51716 29326
rect 51660 29262 51662 29314
rect 51714 29262 51716 29314
rect 50428 28754 50484 29148
rect 51660 28868 51716 29262
rect 50428 28702 50430 28754
rect 50482 28702 50484 28754
rect 50428 28690 50484 28702
rect 50988 28812 51716 28868
rect 50988 28642 51044 28812
rect 51996 28756 52052 28766
rect 50988 28590 50990 28642
rect 51042 28590 51044 28642
rect 50988 28578 51044 28590
rect 51324 28644 51380 28654
rect 51324 28550 51380 28588
rect 51548 28644 51604 28654
rect 51548 28550 51604 28588
rect 51996 28530 52052 28700
rect 52108 28642 52164 29372
rect 52220 29362 52276 29372
rect 52780 29428 52836 29438
rect 52780 28756 52836 29372
rect 52780 28754 53060 28756
rect 52780 28702 52782 28754
rect 52834 28702 53060 28754
rect 52780 28700 53060 28702
rect 52780 28690 52836 28700
rect 52108 28590 52110 28642
rect 52162 28590 52164 28642
rect 52108 28578 52164 28590
rect 52668 28644 52724 28654
rect 52668 28550 52724 28588
rect 51996 28478 51998 28530
rect 52050 28478 52052 28530
rect 51996 28466 52052 28478
rect 51100 28418 51156 28430
rect 51100 28366 51102 28418
rect 51154 28366 51156 28418
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 50988 27076 51044 27086
rect 50204 27022 50206 27074
rect 50258 27022 50260 27074
rect 50204 27010 50260 27022
rect 50428 27074 51044 27076
rect 50428 27022 50990 27074
rect 51042 27022 51044 27074
rect 50428 27020 51044 27022
rect 50092 26964 50148 27002
rect 50428 26908 50484 27020
rect 50988 27010 51044 27020
rect 50092 26898 50148 26908
rect 50372 26852 50484 26908
rect 50652 26852 50708 26890
rect 50372 26740 50428 26852
rect 50652 26786 50708 26796
rect 50372 26684 50484 26740
rect 49980 26238 49982 26290
rect 50034 26238 50036 26290
rect 49980 26226 50036 26238
rect 50316 26516 50372 26526
rect 49868 25956 49924 25966
rect 49924 25900 50036 25956
rect 49868 25890 49924 25900
rect 49308 25678 49310 25730
rect 49362 25678 49364 25730
rect 49308 25666 49364 25678
rect 48300 25554 48356 25564
rect 49756 25618 49812 25630
rect 49756 25566 49758 25618
rect 49810 25566 49812 25618
rect 49196 25506 49252 25518
rect 49644 25508 49700 25518
rect 49196 25454 49198 25506
rect 49250 25454 49252 25506
rect 49084 24948 49140 24958
rect 49084 24722 49140 24892
rect 49196 24946 49252 25454
rect 49196 24894 49198 24946
rect 49250 24894 49252 24946
rect 49196 24882 49252 24894
rect 49532 25506 49700 25508
rect 49532 25454 49646 25506
rect 49698 25454 49700 25506
rect 49532 25452 49700 25454
rect 49308 24836 49364 24846
rect 49308 24742 49364 24780
rect 49420 24834 49476 24846
rect 49420 24782 49422 24834
rect 49474 24782 49476 24834
rect 49084 24670 49086 24722
rect 49138 24670 49140 24722
rect 48748 24500 48804 24510
rect 49084 24500 49140 24670
rect 48804 24444 49140 24500
rect 48748 24434 48804 24444
rect 49420 24388 49476 24782
rect 48860 24332 49476 24388
rect 46732 24220 47460 24276
rect 46732 23826 46788 24220
rect 46732 23774 46734 23826
rect 46786 23774 46788 23826
rect 46732 23762 46788 23774
rect 47404 23380 47460 24220
rect 48860 24050 48916 24332
rect 48860 23998 48862 24050
rect 48914 23998 48916 24050
rect 48860 23986 48916 23998
rect 48972 23380 49028 24332
rect 49420 24164 49476 24174
rect 49532 24164 49588 25452
rect 49644 25442 49700 25452
rect 49756 25172 49812 25566
rect 49756 25106 49812 25116
rect 49420 24162 49588 24164
rect 49420 24110 49422 24162
rect 49474 24110 49588 24162
rect 49420 24108 49588 24110
rect 49868 24722 49924 24734
rect 49868 24670 49870 24722
rect 49922 24670 49924 24722
rect 49420 24098 49476 24108
rect 49868 24050 49924 24670
rect 49980 24164 50036 25900
rect 50092 25732 50148 25742
rect 50092 25394 50148 25676
rect 50092 25342 50094 25394
rect 50146 25342 50148 25394
rect 50092 25330 50148 25342
rect 49980 24108 50148 24164
rect 49868 23998 49870 24050
rect 49922 23998 49924 24050
rect 49868 23986 49924 23998
rect 49084 23940 49140 23950
rect 49084 23846 49140 23884
rect 49980 23940 50036 23950
rect 49756 23826 49812 23838
rect 49980 23828 50036 23884
rect 49756 23774 49758 23826
rect 49810 23774 49812 23826
rect 49084 23380 49140 23390
rect 49756 23380 49812 23774
rect 47404 23378 47684 23380
rect 47404 23326 47406 23378
rect 47458 23326 47684 23378
rect 47404 23324 47684 23326
rect 48972 23378 49140 23380
rect 48972 23326 49086 23378
rect 49138 23326 49140 23378
rect 48972 23324 49140 23326
rect 47404 23314 47460 23324
rect 47628 23266 47684 23324
rect 49084 23314 49140 23324
rect 49308 23324 49812 23380
rect 49868 23826 50036 23828
rect 49868 23774 49982 23826
rect 50034 23774 50036 23826
rect 49868 23772 50036 23774
rect 49868 23378 49924 23772
rect 49980 23762 50036 23772
rect 49868 23326 49870 23378
rect 49922 23326 49924 23378
rect 47628 23214 47630 23266
rect 47682 23214 47684 23266
rect 47628 23202 47684 23214
rect 47964 23154 48020 23166
rect 47964 23102 47966 23154
rect 48018 23102 48020 23154
rect 47964 22708 48020 23102
rect 48300 23154 48356 23166
rect 48300 23102 48302 23154
rect 48354 23102 48356 23154
rect 48076 23044 48132 23054
rect 48076 22950 48132 22988
rect 47964 22642 48020 22652
rect 48300 22596 48356 23102
rect 48300 22530 48356 22540
rect 48748 23156 48804 23166
rect 48748 22484 48804 23100
rect 48860 23154 48916 23166
rect 48860 23102 48862 23154
rect 48914 23102 48916 23154
rect 48860 22820 48916 23102
rect 48860 22754 48916 22764
rect 48972 23154 49028 23166
rect 48972 23102 48974 23154
rect 49026 23102 49028 23154
rect 48972 22708 49028 23102
rect 49196 23156 49252 23166
rect 49196 23062 49252 23100
rect 48972 22642 49028 22652
rect 49308 22596 49364 23324
rect 49868 23314 49924 23326
rect 49980 23266 50036 23278
rect 49980 23214 49982 23266
rect 50034 23214 50036 23266
rect 48748 21698 48804 22428
rect 49084 22540 49364 22596
rect 49420 23156 49476 23166
rect 48972 22372 49028 22382
rect 48972 21810 49028 22316
rect 48972 21758 48974 21810
rect 49026 21758 49028 21810
rect 48972 21746 49028 21758
rect 48748 21646 48750 21698
rect 48802 21646 48804 21698
rect 48748 21634 48804 21646
rect 48188 21476 48244 21486
rect 48188 21382 48244 21420
rect 49084 21474 49140 22540
rect 49308 22372 49364 22382
rect 49420 22372 49476 23100
rect 49756 22930 49812 22942
rect 49756 22878 49758 22930
rect 49810 22878 49812 22930
rect 49756 22820 49812 22878
rect 49756 22754 49812 22764
rect 49364 22316 49476 22372
rect 49532 22708 49588 22718
rect 49308 22306 49364 22316
rect 49532 21810 49588 22652
rect 49980 22708 50036 23214
rect 49980 22642 50036 22652
rect 49532 21758 49534 21810
rect 49586 21758 49588 21810
rect 49532 21746 49588 21758
rect 49084 21422 49086 21474
rect 49138 21422 49140 21474
rect 49084 21410 49140 21422
rect 49420 21476 49476 21486
rect 49420 21382 49476 21420
rect 50092 20356 50148 24108
rect 50316 23548 50372 26460
rect 50428 26290 50484 26684
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 50652 26404 50708 26442
rect 50652 26338 50708 26348
rect 51100 26404 51156 28366
rect 51772 28418 51828 28430
rect 51772 28366 51774 28418
rect 51826 28366 51828 28418
rect 51212 27748 51268 27758
rect 51212 27298 51268 27692
rect 51212 27246 51214 27298
rect 51266 27246 51268 27298
rect 51212 27234 51268 27246
rect 51436 27076 51492 27086
rect 51772 27076 51828 28366
rect 51436 27074 51828 27076
rect 51436 27022 51438 27074
rect 51490 27022 51828 27074
rect 51436 27020 51828 27022
rect 52108 27076 52164 27086
rect 51436 27010 51492 27020
rect 51324 26964 51380 26974
rect 51324 26850 51380 26908
rect 51324 26798 51326 26850
rect 51378 26798 51380 26850
rect 51324 26786 51380 26798
rect 52108 26516 52164 27020
rect 52892 27076 52948 27086
rect 52892 26982 52948 27020
rect 52108 26450 52164 26460
rect 53004 26514 53060 28700
rect 53788 28642 53844 29708
rect 53900 28756 53956 28766
rect 53900 28662 53956 28700
rect 53788 28590 53790 28642
rect 53842 28590 53844 28642
rect 53788 26908 53844 28590
rect 54012 28418 54068 28430
rect 54012 28366 54014 28418
rect 54066 28366 54068 28418
rect 54012 28082 54068 28366
rect 54124 28308 54180 31948
rect 54460 31892 54516 31902
rect 54460 31798 54516 31836
rect 54236 31778 54292 31790
rect 54236 31726 54238 31778
rect 54290 31726 54292 31778
rect 54236 31668 54292 31726
rect 54236 29540 54292 31612
rect 54684 31778 54740 31790
rect 54684 31726 54686 31778
rect 54738 31726 54740 31778
rect 54684 30884 54740 31726
rect 54796 31668 54852 31678
rect 54796 31574 54852 31612
rect 54684 30818 54740 30828
rect 54460 30324 54516 30334
rect 55020 30324 55076 35756
rect 55132 35718 55188 35756
rect 54460 30322 55076 30324
rect 54460 30270 54462 30322
rect 54514 30270 55076 30322
rect 54460 30268 55076 30270
rect 55132 35364 55188 35374
rect 54460 30258 54516 30268
rect 54348 30212 54404 30222
rect 54348 30118 54404 30156
rect 54236 29474 54292 29484
rect 54572 29204 54628 30268
rect 54908 29988 54964 29998
rect 54236 29148 54628 29204
rect 54796 29426 54852 29438
rect 54796 29374 54798 29426
rect 54850 29374 54852 29426
rect 54236 28642 54292 29148
rect 54796 28868 54852 29374
rect 54236 28590 54238 28642
rect 54290 28590 54292 28642
rect 54236 28578 54292 28590
rect 54460 28866 54852 28868
rect 54460 28814 54798 28866
rect 54850 28814 54852 28866
rect 54460 28812 54852 28814
rect 54460 28642 54516 28812
rect 54796 28802 54852 28812
rect 54460 28590 54462 28642
rect 54514 28590 54516 28642
rect 54460 28578 54516 28590
rect 54908 28756 54964 29932
rect 54908 28642 54964 28700
rect 54908 28590 54910 28642
rect 54962 28590 54964 28642
rect 54124 28252 54292 28308
rect 54012 28030 54014 28082
rect 54066 28030 54068 28082
rect 54012 28018 54068 28030
rect 54124 27748 54180 27758
rect 54124 27654 54180 27692
rect 54236 27524 54292 28252
rect 53004 26462 53006 26514
rect 53058 26462 53060 26514
rect 53004 26450 53060 26462
rect 53452 26852 53844 26908
rect 54012 27468 54292 27524
rect 51100 26338 51156 26348
rect 52332 26404 52388 26414
rect 52332 26402 52724 26404
rect 52332 26350 52334 26402
rect 52386 26350 52724 26402
rect 52332 26348 52724 26350
rect 52332 26338 52388 26348
rect 50428 26238 50430 26290
rect 50482 26238 50484 26290
rect 50428 24948 50484 26238
rect 52668 26290 52724 26348
rect 52668 26238 52670 26290
rect 52722 26238 52724 26290
rect 52668 26226 52724 26238
rect 52892 26292 52948 26302
rect 53116 26292 53172 26302
rect 53340 26292 53396 26302
rect 52892 26290 53060 26292
rect 52892 26238 52894 26290
rect 52946 26238 53060 26290
rect 52892 26236 53060 26238
rect 52892 26226 52948 26236
rect 50540 26178 50596 26190
rect 50540 26126 50542 26178
rect 50594 26126 50596 26178
rect 50540 25732 50596 26126
rect 50540 25666 50596 25676
rect 52108 26180 52164 26190
rect 51212 25620 51268 25630
rect 51100 25618 51268 25620
rect 51100 25566 51214 25618
rect 51266 25566 51268 25618
rect 51100 25564 51268 25566
rect 50764 25508 50820 25518
rect 50764 25414 50820 25452
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 50988 24948 51044 24958
rect 50428 24946 51044 24948
rect 50428 24894 50990 24946
rect 51042 24894 51044 24946
rect 50428 24892 51044 24894
rect 50988 24882 51044 24892
rect 51100 24834 51156 25564
rect 51212 25554 51268 25564
rect 51772 25396 51828 25406
rect 51772 25302 51828 25340
rect 51212 25282 51268 25294
rect 51212 25230 51214 25282
rect 51266 25230 51268 25282
rect 51212 24948 51268 25230
rect 51212 24882 51268 24892
rect 51324 25282 51380 25294
rect 51324 25230 51326 25282
rect 51378 25230 51380 25282
rect 51100 24782 51102 24834
rect 51154 24782 51156 24834
rect 51100 24770 51156 24782
rect 51324 24724 51380 25230
rect 51548 25284 51604 25294
rect 51548 25190 51604 25228
rect 51324 24164 51380 24668
rect 51324 24098 51380 24108
rect 50556 23548 50820 23558
rect 50316 23492 50484 23548
rect 50428 22370 50484 23492
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 52108 23548 52164 26124
rect 52220 26178 52276 26190
rect 52220 26126 52222 26178
rect 52274 26126 52276 26178
rect 52220 25284 52276 26126
rect 52892 26068 52948 26078
rect 52668 25396 52724 25406
rect 52668 25302 52724 25340
rect 52780 25394 52836 25406
rect 52780 25342 52782 25394
rect 52834 25342 52836 25394
rect 52220 25218 52276 25228
rect 52780 24724 52836 25342
rect 52780 24658 52836 24668
rect 52108 23492 52276 23548
rect 50556 23482 50820 23492
rect 51772 23156 51828 23166
rect 51828 23100 52052 23156
rect 51772 23062 51828 23100
rect 51996 22594 52052 23100
rect 51996 22542 51998 22594
rect 52050 22542 52052 22594
rect 51996 22530 52052 22542
rect 52108 22482 52164 22494
rect 52108 22430 52110 22482
rect 52162 22430 52164 22482
rect 50428 22318 50430 22370
rect 50482 22318 50484 22370
rect 50428 22148 50484 22318
rect 51212 22372 51268 22382
rect 50876 22148 50932 22158
rect 50428 22146 50932 22148
rect 50428 22094 50878 22146
rect 50930 22094 50932 22146
rect 50428 22092 50932 22094
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 50876 20580 50932 22092
rect 50988 21476 51044 21486
rect 51212 21476 51268 22316
rect 52108 22372 52164 22430
rect 52108 22306 52164 22316
rect 50988 21474 51268 21476
rect 50988 21422 50990 21474
rect 51042 21422 51268 21474
rect 50988 21420 51268 21422
rect 50988 21410 51044 21420
rect 52220 20804 52276 23492
rect 52332 23154 52388 23166
rect 52332 23102 52334 23154
rect 52386 23102 52388 23154
rect 52332 22820 52388 23102
rect 52444 23044 52500 23054
rect 52780 23044 52836 23054
rect 52444 23042 52836 23044
rect 52444 22990 52446 23042
rect 52498 22990 52782 23042
rect 52834 22990 52836 23042
rect 52444 22988 52836 22990
rect 52892 23044 52948 26012
rect 53004 24724 53060 26236
rect 53116 26290 53284 26292
rect 53116 26238 53118 26290
rect 53170 26238 53284 26290
rect 53116 26236 53284 26238
rect 53116 26226 53172 26236
rect 53228 25732 53284 26236
rect 53340 26198 53396 26236
rect 53340 25732 53396 25742
rect 53228 25730 53396 25732
rect 53228 25678 53342 25730
rect 53394 25678 53396 25730
rect 53228 25676 53396 25678
rect 53340 25666 53396 25676
rect 53452 25618 53508 26852
rect 53452 25566 53454 25618
rect 53506 25566 53508 25618
rect 53452 25554 53508 25566
rect 53004 24658 53060 24668
rect 53788 24164 53844 24174
rect 53788 24070 53844 24108
rect 53004 23828 53060 23838
rect 53004 23378 53060 23772
rect 53004 23326 53006 23378
rect 53058 23326 53060 23378
rect 53004 23314 53060 23326
rect 53900 23826 53956 23838
rect 53900 23774 53902 23826
rect 53954 23774 53956 23826
rect 53900 23156 53956 23774
rect 53900 23090 53956 23100
rect 52892 22988 53060 23044
rect 52444 22978 52500 22988
rect 52780 22978 52836 22988
rect 52892 22820 52948 22830
rect 52332 22764 52892 22820
rect 52780 22596 52836 22606
rect 52780 22502 52836 22540
rect 52780 22372 52836 22382
rect 52780 22258 52836 22316
rect 52892 22370 52948 22764
rect 52892 22318 52894 22370
rect 52946 22318 52948 22370
rect 52892 22306 52948 22318
rect 52780 22206 52782 22258
rect 52834 22206 52836 22258
rect 52780 22194 52836 22206
rect 52220 20748 52500 20804
rect 50876 20514 50932 20524
rect 52108 20580 52164 20590
rect 52220 20580 52276 20590
rect 52108 20578 52220 20580
rect 52108 20526 52110 20578
rect 52162 20526 52220 20578
rect 52108 20524 52220 20526
rect 52108 20514 52164 20524
rect 49756 20300 50148 20356
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 49756 20244 49812 20300
rect 49084 20188 49812 20244
rect 49084 20130 49140 20188
rect 49084 20078 49086 20130
rect 49138 20078 49140 20130
rect 49084 20066 49140 20078
rect 49756 20130 49812 20188
rect 49756 20078 49758 20130
rect 49810 20078 49812 20130
rect 49756 20066 49812 20078
rect 49196 20020 49252 20030
rect 47516 19908 47572 19918
rect 46956 19906 47684 19908
rect 46956 19854 47518 19906
rect 47570 19854 47684 19906
rect 46956 19852 47684 19854
rect 46620 19404 46900 19460
rect 45388 18622 45390 18674
rect 45442 18622 45444 18674
rect 45388 18610 45444 18622
rect 45500 19236 45556 19246
rect 45052 18450 45444 18452
rect 45052 18398 45054 18450
rect 45106 18398 45444 18450
rect 45052 18396 45444 18398
rect 45052 18386 45108 18396
rect 45388 18340 45444 18396
rect 45388 18274 45444 18284
rect 45276 17556 45332 17566
rect 45276 17108 45332 17500
rect 44492 17054 44494 17106
rect 44546 17054 44548 17106
rect 44492 17042 44548 17054
rect 44604 17106 45332 17108
rect 44604 17054 45278 17106
rect 45330 17054 45332 17106
rect 44604 17052 45332 17054
rect 44380 16770 44436 16782
rect 44380 16718 44382 16770
rect 44434 16718 44436 16770
rect 44380 16324 44436 16718
rect 43932 16268 44436 16324
rect 43932 16098 43988 16268
rect 44604 16212 44660 17052
rect 45276 17042 45332 17052
rect 44940 16884 44996 16894
rect 44940 16882 45220 16884
rect 44940 16830 44942 16882
rect 44994 16830 45220 16882
rect 44940 16828 45220 16830
rect 44940 16818 44996 16828
rect 43932 16046 43934 16098
rect 43986 16046 43988 16098
rect 43932 16034 43988 16046
rect 44268 16156 44660 16212
rect 44268 16098 44324 16156
rect 44268 16046 44270 16098
rect 44322 16046 44324 16098
rect 44268 16034 44324 16046
rect 44044 15988 44100 15998
rect 44044 15894 44100 15932
rect 43820 14642 43876 14654
rect 43820 14590 43822 14642
rect 43874 14590 43876 14642
rect 43820 13860 43876 14590
rect 43820 13794 43876 13804
rect 44268 14644 44324 14654
rect 44268 12962 44324 14588
rect 44268 12910 44270 12962
rect 44322 12910 44324 12962
rect 44268 12898 44324 12910
rect 43596 9986 43652 9996
rect 43372 9202 43428 9212
rect 44268 9716 44324 9726
rect 43708 9156 43764 9166
rect 43708 9062 43764 9100
rect 44268 9044 44324 9660
rect 43260 8988 43652 9044
rect 42476 8652 42756 8708
rect 42140 8372 42196 8382
rect 42140 8278 42196 8316
rect 41468 7980 41972 8036
rect 41356 7700 41412 7710
rect 41244 7698 41412 7700
rect 41244 7646 41358 7698
rect 41410 7646 41412 7698
rect 41244 7644 41412 7646
rect 41356 7634 41412 7644
rect 41132 7588 41188 7598
rect 41132 7586 41300 7588
rect 41132 7534 41134 7586
rect 41186 7534 41300 7586
rect 41132 7532 41300 7534
rect 41132 7522 41188 7532
rect 41244 7476 41300 7532
rect 41468 7476 41524 7980
rect 42252 7812 42308 7822
rect 41244 7420 41524 7476
rect 41580 7476 41636 7486
rect 40908 7382 40964 7420
rect 41580 7382 41636 7420
rect 41132 7362 41188 7374
rect 41132 7310 41134 7362
rect 41186 7310 41188 7362
rect 41132 6692 41188 7310
rect 42252 7362 42308 7756
rect 42700 7700 42756 8652
rect 42700 7698 43316 7700
rect 42700 7646 42702 7698
rect 42754 7646 43316 7698
rect 42700 7644 43316 7646
rect 42700 7634 42756 7644
rect 42252 7310 42254 7362
rect 42306 7310 42308 7362
rect 42252 7028 42308 7310
rect 43148 7362 43204 7374
rect 43148 7310 43150 7362
rect 43202 7310 43204 7362
rect 42252 6962 42308 6972
rect 43036 7250 43092 7262
rect 43036 7198 43038 7250
rect 43090 7198 43092 7250
rect 41132 6626 41188 6636
rect 42252 6804 42308 6814
rect 42252 6690 42308 6748
rect 42252 6638 42254 6690
rect 42306 6638 42308 6690
rect 42252 6626 42308 6638
rect 42700 6692 42756 6702
rect 42700 6598 42756 6636
rect 43036 6690 43092 7198
rect 43148 6804 43204 7310
rect 43148 6738 43204 6748
rect 43260 6802 43316 7644
rect 43596 7698 43652 8988
rect 44268 8370 44324 8988
rect 44268 8318 44270 8370
rect 44322 8318 44324 8370
rect 44268 8306 44324 8318
rect 43596 7646 43598 7698
rect 43650 7646 43652 7698
rect 43596 7250 43652 7646
rect 43596 7198 43598 7250
rect 43650 7198 43652 7250
rect 43596 7186 43652 7198
rect 44156 7476 44212 7486
rect 43484 7028 43540 7038
rect 43484 6914 43540 6972
rect 43484 6862 43486 6914
rect 43538 6862 43540 6914
rect 43484 6850 43540 6862
rect 43708 6916 43764 6926
rect 43260 6750 43262 6802
rect 43314 6750 43316 6802
rect 43260 6738 43316 6750
rect 43036 6638 43038 6690
rect 43090 6638 43092 6690
rect 43036 6626 43092 6638
rect 43708 6690 43764 6860
rect 43708 6638 43710 6690
rect 43762 6638 43764 6690
rect 43708 6626 43764 6638
rect 44044 6690 44100 6702
rect 44044 6638 44046 6690
rect 44098 6638 44100 6690
rect 40236 5796 40292 6524
rect 42588 6468 42644 6478
rect 41916 6466 42644 6468
rect 41916 6414 42590 6466
rect 42642 6414 42644 6466
rect 41916 6412 42644 6414
rect 41132 5908 41188 5918
rect 40348 5796 40404 5806
rect 40236 5794 40404 5796
rect 40236 5742 40350 5794
rect 40402 5742 40404 5794
rect 40236 5740 40404 5742
rect 40348 5730 40404 5740
rect 41132 5794 41188 5852
rect 41132 5742 41134 5794
rect 41186 5742 41188 5794
rect 39564 4386 39620 4396
rect 41020 5236 41076 5246
rect 36204 4338 36372 4340
rect 36204 4286 36206 4338
rect 36258 4286 36372 4338
rect 36204 4284 36372 4286
rect 36204 4274 36260 4284
rect 32172 4174 32174 4226
rect 32226 4174 32228 4226
rect 32172 4162 32228 4174
rect 39004 4226 39060 4238
rect 39004 4174 39006 4226
rect 39058 4174 39060 4226
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 28588 3602 28644 3612
rect 38892 3668 38948 3678
rect 28140 3490 28196 3500
rect 36652 3556 36708 3566
rect 36652 3462 36708 3500
rect 28364 3330 28420 3342
rect 29148 3332 29204 3342
rect 31164 3332 31220 3342
rect 33180 3332 33236 3342
rect 35196 3332 35252 3342
rect 28364 3278 28366 3330
rect 28418 3278 28420 3330
rect 26908 1762 26964 1774
rect 26908 1710 26910 1762
rect 26962 1710 26964 1762
rect 26908 800 26964 1710
rect 28364 1762 28420 3278
rect 28364 1710 28366 1762
rect 28418 1710 28420 1762
rect 28364 1698 28420 1710
rect 28924 3330 29204 3332
rect 28924 3278 29150 3330
rect 29202 3278 29204 3330
rect 28924 3276 29204 3278
rect 28924 800 28980 3276
rect 29148 3266 29204 3276
rect 30940 3330 31220 3332
rect 30940 3278 31166 3330
rect 31218 3278 31220 3330
rect 30940 3276 31220 3278
rect 30940 800 30996 3276
rect 31164 3266 31220 3276
rect 32956 3330 33236 3332
rect 32956 3278 33182 3330
rect 33234 3278 33236 3330
rect 32956 3276 33236 3278
rect 32956 800 33012 3276
rect 33180 3266 33236 3276
rect 34972 3330 35252 3332
rect 34972 3278 35198 3330
rect 35250 3278 35252 3330
rect 34972 3276 35252 3278
rect 34972 800 35028 3276
rect 35196 3266 35252 3276
rect 37660 3330 37716 3342
rect 37660 3278 37662 3330
rect 37714 3278 37716 3330
rect 36988 924 37380 980
rect 36988 800 37044 924
rect 8988 700 9380 756
rect 10752 0 10864 800
rect 12768 0 12880 800
rect 14784 0 14896 800
rect 16800 0 16912 800
rect 18816 0 18928 800
rect 20832 0 20944 800
rect 22848 0 22960 800
rect 24864 0 24976 800
rect 26880 0 26992 800
rect 28896 0 29008 800
rect 30912 0 31024 800
rect 32928 0 33040 800
rect 34944 0 35056 800
rect 36960 0 37072 800
rect 37324 756 37380 924
rect 37660 756 37716 3278
rect 38892 1652 38948 3612
rect 39004 3556 39060 4174
rect 40796 3668 40852 3678
rect 40796 3574 40852 3612
rect 39788 3556 39844 3566
rect 39004 3554 39844 3556
rect 39004 3502 39790 3554
rect 39842 3502 39844 3554
rect 39004 3500 39844 3502
rect 39788 3490 39844 3500
rect 38892 1596 39060 1652
rect 39004 800 39060 1596
rect 41020 800 41076 5180
rect 41132 5124 41188 5742
rect 41356 5234 41412 5246
rect 41356 5182 41358 5234
rect 41410 5182 41412 5234
rect 41356 5124 41412 5182
rect 41692 5124 41748 5134
rect 41356 5122 41748 5124
rect 41356 5070 41694 5122
rect 41746 5070 41748 5122
rect 41356 5068 41748 5070
rect 41132 4338 41188 5068
rect 41692 5058 41748 5068
rect 41916 4450 41972 6412
rect 42588 6402 42644 6412
rect 43484 6466 43540 6478
rect 43484 6414 43486 6466
rect 43538 6414 43540 6466
rect 42700 5236 42756 5246
rect 42700 5142 42756 5180
rect 41916 4398 41918 4450
rect 41970 4398 41972 4450
rect 41916 4386 41972 4398
rect 41132 4286 41134 4338
rect 41186 4286 41188 4338
rect 41132 4274 41188 4286
rect 43036 4116 43092 4126
rect 43036 800 43092 4060
rect 43148 3780 43204 3790
rect 43148 3666 43204 3724
rect 43148 3614 43150 3666
rect 43202 3614 43204 3666
rect 43148 3602 43204 3614
rect 43484 3668 43540 6414
rect 44044 6468 44100 6638
rect 44044 6402 44100 6412
rect 43596 5124 43652 5134
rect 43652 5068 43764 5124
rect 43596 5058 43652 5068
rect 43484 3602 43540 3612
rect 43708 3554 43764 5068
rect 44044 4228 44100 4238
rect 44156 4228 44212 7420
rect 44380 6692 44436 16156
rect 44940 16098 44996 16110
rect 44940 16046 44942 16098
rect 44994 16046 44996 16098
rect 44940 15148 44996 16046
rect 45164 15148 45220 16828
rect 45500 15148 45556 19180
rect 46620 19236 46676 19246
rect 46620 19142 46676 19180
rect 45724 18340 45780 18350
rect 45724 16996 45780 18284
rect 46844 17780 46900 19404
rect 46956 19346 47012 19852
rect 47516 19842 47572 19852
rect 46956 19294 46958 19346
rect 47010 19294 47012 19346
rect 46956 19282 47012 19294
rect 46956 17780 47012 17790
rect 46844 17724 46956 17780
rect 46956 17686 47012 17724
rect 47628 17220 47684 19852
rect 48636 19348 48692 19358
rect 48636 19254 48692 19292
rect 48300 19124 48356 19134
rect 48300 19030 48356 19068
rect 47964 19010 48020 19022
rect 47964 18958 47966 19010
rect 48018 18958 48020 19010
rect 47964 18676 48020 18958
rect 49196 19012 49252 19964
rect 47964 18610 48020 18620
rect 49084 18676 49140 18686
rect 49196 18676 49252 18956
rect 49084 18674 49252 18676
rect 49084 18622 49086 18674
rect 49138 18622 49252 18674
rect 49084 18620 49252 18622
rect 49420 20018 49476 20030
rect 49420 19966 49422 20018
rect 49474 19966 49476 20018
rect 49420 19348 49476 19966
rect 49084 18610 49140 18620
rect 49420 18564 49476 19292
rect 49532 20018 49588 20030
rect 49532 19966 49534 20018
rect 49586 19966 49588 20018
rect 49532 19124 49588 19966
rect 49868 20020 49924 20030
rect 49868 19926 49924 19964
rect 49644 19906 49700 19918
rect 49644 19854 49646 19906
rect 49698 19854 49700 19906
rect 49644 19796 49700 19854
rect 50316 19906 50372 19918
rect 50316 19854 50318 19906
rect 50370 19854 50372 19906
rect 50316 19796 50372 19854
rect 49644 19740 50372 19796
rect 50428 19796 50484 19806
rect 50428 19794 50820 19796
rect 50428 19742 50430 19794
rect 50482 19742 50820 19794
rect 50428 19740 50820 19742
rect 50428 19730 50484 19740
rect 50764 19346 50820 19740
rect 50764 19294 50766 19346
rect 50818 19294 50820 19346
rect 50764 19282 50820 19294
rect 49532 19058 49588 19068
rect 51436 19234 51492 19246
rect 51436 19182 51438 19234
rect 51490 19182 51492 19234
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 49420 18498 49476 18508
rect 50428 18564 50484 18574
rect 48748 18450 48804 18462
rect 48748 18398 48750 18450
rect 48802 18398 48804 18450
rect 48188 18338 48244 18350
rect 48188 18286 48190 18338
rect 48242 18286 48244 18338
rect 48188 18228 48244 18286
rect 48188 18162 48244 18172
rect 48748 18228 48804 18398
rect 48748 18162 48804 18172
rect 46508 17164 47684 17220
rect 46508 17106 46564 17164
rect 46508 17054 46510 17106
rect 46562 17054 46564 17106
rect 46508 17042 46564 17054
rect 45724 16930 45780 16940
rect 46732 16994 46788 17006
rect 46732 16942 46734 16994
rect 46786 16942 46788 16994
rect 46172 16884 46228 16894
rect 46172 16790 46228 16828
rect 46732 16884 46788 16942
rect 47628 16994 47684 17164
rect 47628 16942 47630 16994
rect 47682 16942 47684 16994
rect 47628 16930 47684 16942
rect 47852 17780 47908 17790
rect 46732 16818 46788 16828
rect 47516 16884 47572 16894
rect 47292 16772 47348 16782
rect 47292 16678 47348 16716
rect 46844 16658 46900 16670
rect 46844 16606 46846 16658
rect 46898 16606 46900 16658
rect 45612 15988 45668 15998
rect 46844 15988 46900 16606
rect 47516 16212 47572 16828
rect 47852 16882 47908 17724
rect 47852 16830 47854 16882
rect 47906 16830 47908 16882
rect 47852 16818 47908 16830
rect 48748 16996 48804 17006
rect 48188 16772 48244 16782
rect 47740 16212 47796 16222
rect 47516 16210 47796 16212
rect 47516 16158 47742 16210
rect 47794 16158 47796 16210
rect 47516 16156 47796 16158
rect 45612 15986 46564 15988
rect 45612 15934 45614 15986
rect 45666 15934 46564 15986
rect 45612 15932 46564 15934
rect 45612 15922 45668 15932
rect 46508 15538 46564 15932
rect 46508 15486 46510 15538
rect 46562 15486 46564 15538
rect 46508 15474 46564 15486
rect 46732 15876 46788 15886
rect 46172 15314 46228 15326
rect 46172 15262 46174 15314
rect 46226 15262 46228 15314
rect 44940 15092 45108 15148
rect 45164 15092 45332 15148
rect 45500 15092 45892 15148
rect 45052 14644 45108 15092
rect 45052 14550 45108 14588
rect 44828 13860 44884 13870
rect 44884 13804 44996 13860
rect 44828 13794 44884 13804
rect 44940 12292 44996 13804
rect 45276 13188 45332 15092
rect 45724 13748 45780 13758
rect 45500 13692 45724 13748
rect 45388 13188 45444 13198
rect 45276 13132 45388 13188
rect 45276 12962 45332 12974
rect 45276 12910 45278 12962
rect 45330 12910 45332 12962
rect 45052 12740 45108 12750
rect 45276 12740 45332 12910
rect 45108 12684 45332 12740
rect 45052 12646 45108 12684
rect 45276 12404 45332 12414
rect 45388 12404 45444 13132
rect 45276 12402 45444 12404
rect 45276 12350 45278 12402
rect 45330 12350 45444 12402
rect 45276 12348 45444 12350
rect 45276 12338 45332 12348
rect 45164 12292 45220 12302
rect 44940 12236 45164 12292
rect 45164 12198 45220 12236
rect 45388 11620 45444 12348
rect 45500 12402 45556 13692
rect 45724 13682 45780 13692
rect 45836 12516 45892 15092
rect 45948 13636 46004 13646
rect 46172 13636 46228 15262
rect 46732 15314 46788 15820
rect 46732 15262 46734 15314
rect 46786 15262 46788 15314
rect 46732 15250 46788 15262
rect 46844 15316 46900 15932
rect 47292 15316 47348 15326
rect 46844 15314 47348 15316
rect 46844 15262 47294 15314
rect 47346 15262 47348 15314
rect 46844 15260 47348 15262
rect 47292 15250 47348 15260
rect 46956 14532 47012 14542
rect 46284 13748 46340 13758
rect 46284 13654 46340 13692
rect 46508 13746 46564 13758
rect 46508 13694 46510 13746
rect 46562 13694 46564 13746
rect 45948 13634 46228 13636
rect 45948 13582 45950 13634
rect 46002 13582 46228 13634
rect 45948 13580 46228 13582
rect 46396 13634 46452 13646
rect 46396 13582 46398 13634
rect 46450 13582 46452 13634
rect 45948 13412 46004 13580
rect 45948 12740 46004 13356
rect 46396 12852 46452 13582
rect 46396 12786 46452 12796
rect 45948 12674 46004 12684
rect 45836 12460 46004 12516
rect 45500 12350 45502 12402
rect 45554 12350 45556 12402
rect 45500 12338 45556 12350
rect 45724 12292 45780 12302
rect 45500 11620 45556 11630
rect 45388 11618 45556 11620
rect 45388 11566 45502 11618
rect 45554 11566 45556 11618
rect 45388 11564 45556 11566
rect 45500 11554 45556 11564
rect 45724 11506 45780 12236
rect 45724 11454 45726 11506
rect 45778 11454 45780 11506
rect 45724 11442 45780 11454
rect 45836 12290 45892 12302
rect 45836 12238 45838 12290
rect 45890 12238 45892 12290
rect 45836 12068 45892 12238
rect 45836 11172 45892 12012
rect 45948 12178 46004 12460
rect 45948 12126 45950 12178
rect 46002 12126 46004 12178
rect 45948 11394 46004 12126
rect 46508 11844 46564 13694
rect 46732 13746 46788 13758
rect 46732 13694 46734 13746
rect 46786 13694 46788 13746
rect 46732 12292 46788 13694
rect 46956 12852 47012 14476
rect 47516 13860 47572 13870
rect 47628 13860 47684 16156
rect 47740 16146 47796 16156
rect 48188 16212 48244 16716
rect 48300 16660 48356 16670
rect 48300 16566 48356 16604
rect 48188 16118 48244 16156
rect 48076 15876 48132 15886
rect 47516 13858 47684 13860
rect 47516 13806 47518 13858
rect 47570 13806 47684 13858
rect 47516 13804 47684 13806
rect 47740 15874 48132 15876
rect 47740 15822 48078 15874
rect 48130 15822 48132 15874
rect 47740 15820 48132 15822
rect 47740 15314 47796 15820
rect 48076 15810 48132 15820
rect 47740 15262 47742 15314
rect 47794 15262 47796 15314
rect 47516 13794 47572 13804
rect 47180 13634 47236 13646
rect 47180 13582 47182 13634
rect 47234 13582 47236 13634
rect 47180 13188 47236 13582
rect 47236 13132 47572 13188
rect 47180 13122 47236 13132
rect 47292 12852 47348 12862
rect 46956 12850 47348 12852
rect 46956 12798 47294 12850
rect 47346 12798 47348 12850
rect 46956 12796 47348 12798
rect 46732 12198 46788 12236
rect 46844 12740 46900 12750
rect 46956 12740 47012 12796
rect 47292 12786 47348 12796
rect 46900 12684 47012 12740
rect 46620 12180 46676 12190
rect 46620 12086 46676 12124
rect 46060 11788 46564 11844
rect 46060 11506 46116 11788
rect 46060 11454 46062 11506
rect 46114 11454 46116 11506
rect 46060 11442 46116 11454
rect 45948 11342 45950 11394
rect 46002 11342 46004 11394
rect 45948 11330 46004 11342
rect 46172 11172 46228 11182
rect 45836 11170 46228 11172
rect 45836 11118 46174 11170
rect 46226 11118 46228 11170
rect 45836 11116 46228 11118
rect 46172 11106 46228 11116
rect 46508 10948 46564 11788
rect 46508 10882 46564 10892
rect 45836 10836 45892 10846
rect 45612 10610 45668 10622
rect 45612 10558 45614 10610
rect 45666 10558 45668 10610
rect 45612 10500 45668 10558
rect 45612 6804 45668 10444
rect 45836 8930 45892 10780
rect 46844 10610 46900 12684
rect 47292 12404 47348 12414
rect 47068 12292 47124 12302
rect 46956 11620 47012 11630
rect 46956 10836 47012 11564
rect 47068 11506 47124 12236
rect 47068 11454 47070 11506
rect 47122 11454 47124 11506
rect 47068 11442 47124 11454
rect 47292 11394 47348 12348
rect 47516 12178 47572 13132
rect 47740 12404 47796 15262
rect 48748 15316 48804 16940
rect 49644 16994 49700 17006
rect 49644 16942 49646 16994
rect 49698 16942 49700 16994
rect 49308 16882 49364 16894
rect 49308 16830 49310 16882
rect 49362 16830 49364 16882
rect 48860 16212 48916 16222
rect 48860 16118 48916 16156
rect 49308 15538 49364 16830
rect 49644 16212 49700 16942
rect 49644 16146 49700 16156
rect 49308 15486 49310 15538
rect 49362 15486 49364 15538
rect 49308 15474 49364 15486
rect 48188 15204 48244 15242
rect 48748 15222 48804 15260
rect 48188 15138 48244 15148
rect 48972 15204 49028 15242
rect 48972 15138 49028 15148
rect 49756 15204 49812 15242
rect 49756 15138 49812 15148
rect 49308 14756 49364 14766
rect 48636 14532 48692 14542
rect 48636 14438 48692 14476
rect 48076 13748 48132 13758
rect 48076 13654 48132 13692
rect 49196 13746 49252 13758
rect 49196 13694 49198 13746
rect 49250 13694 49252 13746
rect 48188 13522 48244 13534
rect 48188 13470 48190 13522
rect 48242 13470 48244 13522
rect 47740 12338 47796 12348
rect 48076 12402 48132 12414
rect 48076 12350 48078 12402
rect 48130 12350 48132 12402
rect 47516 12126 47518 12178
rect 47570 12126 47572 12178
rect 47516 12114 47572 12126
rect 47964 12180 48020 12190
rect 47292 11342 47294 11394
rect 47346 11342 47348 11394
rect 47292 11330 47348 11342
rect 47964 11284 48020 12124
rect 48076 11732 48132 12350
rect 48188 12292 48244 13470
rect 49196 13524 49252 13694
rect 49308 13748 49364 14700
rect 50428 13972 50484 18508
rect 51212 18452 51268 18462
rect 51436 18452 51492 19182
rect 52108 19236 52164 19274
rect 52108 19170 52164 19180
rect 51996 19012 52052 19022
rect 51884 19010 52052 19012
rect 51884 18958 51998 19010
rect 52050 18958 52052 19010
rect 51884 18956 52052 18958
rect 51884 18562 51940 18956
rect 51996 18946 52052 18956
rect 51884 18510 51886 18562
rect 51938 18510 51940 18562
rect 51884 18498 51940 18510
rect 51212 18450 51492 18452
rect 51212 18398 51214 18450
rect 51266 18398 51492 18450
rect 51212 18396 51492 18398
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 51212 16884 51268 18396
rect 51436 17892 51492 17902
rect 51436 17108 51492 17836
rect 52108 17668 52164 17678
rect 52220 17668 52276 20524
rect 52164 17612 52276 17668
rect 51884 17444 51940 17454
rect 52108 17444 52164 17612
rect 51772 17108 51828 17118
rect 51436 17106 51828 17108
rect 51436 17054 51438 17106
rect 51490 17054 51774 17106
rect 51826 17054 51828 17106
rect 51436 17052 51828 17054
rect 51436 17042 51492 17052
rect 51772 17042 51828 17052
rect 51212 16818 51268 16828
rect 51660 16884 51716 16894
rect 51884 16884 51940 17388
rect 50988 16212 51044 16222
rect 50988 16118 51044 16156
rect 51660 16098 51716 16828
rect 51660 16046 51662 16098
rect 51714 16046 51716 16098
rect 51660 16034 51716 16046
rect 51772 16828 51940 16884
rect 51996 17442 52164 17444
rect 51996 17390 52110 17442
rect 52162 17390 52164 17442
rect 51996 17388 52164 17390
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 50540 14532 50596 14542
rect 50540 14438 50596 14476
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 51212 13972 51268 13982
rect 50428 13916 50708 13972
rect 49308 13654 49364 13692
rect 49532 13748 49588 13758
rect 49532 13654 49588 13692
rect 49756 13746 49812 13758
rect 49756 13694 49758 13746
rect 49810 13694 49812 13746
rect 49196 13458 49252 13468
rect 49420 13634 49476 13646
rect 49420 13582 49422 13634
rect 49474 13582 49476 13634
rect 49084 12964 49140 12974
rect 48972 12404 49028 12414
rect 48972 12310 49028 12348
rect 49084 12402 49140 12908
rect 49084 12350 49086 12402
rect 49138 12350 49140 12402
rect 48188 12226 48244 12236
rect 48748 12178 48804 12190
rect 48748 12126 48750 12178
rect 48802 12126 48804 12178
rect 48076 11666 48132 11676
rect 48188 12068 48244 12078
rect 48188 11394 48244 12012
rect 48748 11620 48804 12126
rect 49084 12068 49140 12350
rect 49196 12628 49252 12638
rect 49196 12402 49252 12572
rect 49196 12350 49198 12402
rect 49250 12350 49252 12402
rect 49196 12338 49252 12350
rect 49308 12292 49364 12302
rect 49308 12178 49364 12236
rect 49308 12126 49310 12178
rect 49362 12126 49364 12178
rect 49308 12114 49364 12126
rect 49420 12180 49476 13582
rect 49756 13636 49812 13694
rect 49756 13570 49812 13580
rect 50204 13634 50260 13646
rect 50204 13582 50206 13634
rect 50258 13582 50260 13634
rect 50092 13524 50148 13534
rect 50092 13430 50148 13468
rect 49756 12852 49812 12862
rect 49756 12402 49812 12796
rect 49756 12350 49758 12402
rect 49810 12350 49812 12402
rect 49756 12338 49812 12350
rect 49980 12740 50036 12750
rect 49980 12402 50036 12684
rect 50204 12628 50260 13582
rect 50204 12562 50260 12572
rect 49980 12350 49982 12402
rect 50034 12350 50036 12402
rect 49980 12338 50036 12350
rect 50428 12404 50484 13916
rect 50652 13858 50708 13916
rect 50652 13806 50654 13858
rect 50706 13806 50708 13858
rect 50652 13794 50708 13806
rect 50540 13748 50596 13758
rect 50540 13654 50596 13692
rect 50988 12964 51044 12974
rect 50988 12870 51044 12908
rect 50876 12740 50932 12750
rect 50876 12646 50932 12684
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 50764 12404 50820 12414
rect 50428 12402 50820 12404
rect 50428 12350 50766 12402
rect 50818 12350 50820 12402
rect 50428 12348 50820 12350
rect 50764 12338 50820 12348
rect 50988 12402 51044 12414
rect 50988 12350 50990 12402
rect 51042 12350 51044 12402
rect 49420 12114 49476 12124
rect 50204 12290 50260 12302
rect 50204 12238 50206 12290
rect 50258 12238 50260 12290
rect 50204 12180 50260 12238
rect 50204 12114 50260 12124
rect 49084 12002 49140 12012
rect 49868 12066 49924 12078
rect 49868 12014 49870 12066
rect 49922 12014 49924 12066
rect 48748 11554 48804 11564
rect 48188 11342 48190 11394
rect 48242 11342 48244 11394
rect 48188 11330 48244 11342
rect 49644 11394 49700 11406
rect 49644 11342 49646 11394
rect 49698 11342 49700 11394
rect 48076 11284 48132 11294
rect 47964 11282 48132 11284
rect 47964 11230 48078 11282
rect 48130 11230 48132 11282
rect 47964 11228 48132 11230
rect 48076 11218 48132 11228
rect 49420 11282 49476 11294
rect 49420 11230 49422 11282
rect 49474 11230 49476 11282
rect 47852 11172 47908 11182
rect 47628 11170 47908 11172
rect 47628 11118 47854 11170
rect 47906 11118 47908 11170
rect 47628 11116 47908 11118
rect 46956 10770 47012 10780
rect 47180 10948 47236 10958
rect 46844 10558 46846 10610
rect 46898 10558 46900 10610
rect 46732 10500 46788 10510
rect 46844 10500 46900 10558
rect 47180 10610 47236 10892
rect 47180 10558 47182 10610
rect 47234 10558 47236 10610
rect 47180 10546 47236 10558
rect 47628 10610 47684 11116
rect 47852 11106 47908 11116
rect 47628 10558 47630 10610
rect 47682 10558 47684 10610
rect 47628 10546 47684 10558
rect 46788 10444 46900 10500
rect 48860 10498 48916 10510
rect 48860 10446 48862 10498
rect 48914 10446 48916 10498
rect 46732 10434 46788 10444
rect 47404 10388 47460 10398
rect 47404 10294 47460 10332
rect 48076 10386 48132 10398
rect 48076 10334 48078 10386
rect 48130 10334 48132 10386
rect 48076 10164 48132 10334
rect 48748 10388 48804 10398
rect 48748 10294 48804 10332
rect 48076 10108 48580 10164
rect 47740 10052 47796 10062
rect 47740 9958 47796 9996
rect 47404 9828 47460 9838
rect 47180 9826 47460 9828
rect 47180 9774 47406 9826
rect 47458 9774 47460 9826
rect 47180 9772 47460 9774
rect 46172 9044 46228 9054
rect 46172 8950 46228 8988
rect 45836 8878 45838 8930
rect 45890 8878 45892 8930
rect 45836 8866 45892 8878
rect 46284 8818 46340 8830
rect 46284 8766 46286 8818
rect 46338 8766 46340 8818
rect 45612 6738 45668 6748
rect 45724 8036 45780 8046
rect 45724 6802 45780 7980
rect 46284 7924 46340 8766
rect 47180 8482 47236 9772
rect 47404 9762 47460 9772
rect 47964 9828 48020 9838
rect 47964 9734 48020 9772
rect 48524 9826 48580 10108
rect 48860 10052 48916 10446
rect 48860 9986 48916 9996
rect 49420 9938 49476 11230
rect 49420 9886 49422 9938
rect 49474 9886 49476 9938
rect 49420 9874 49476 9886
rect 48524 9774 48526 9826
rect 48578 9774 48580 9826
rect 48524 9762 48580 9774
rect 48860 9826 48916 9838
rect 48860 9774 48862 9826
rect 48914 9774 48916 9826
rect 48076 9156 48132 9166
rect 48076 9062 48132 9100
rect 48188 9044 48244 9054
rect 48188 8950 48244 8988
rect 48748 9044 48804 9054
rect 48860 9044 48916 9774
rect 49084 9828 49140 9838
rect 49084 9266 49140 9772
rect 49644 9716 49700 11342
rect 49756 10724 49812 10734
rect 49868 10724 49924 12014
rect 50876 11732 50932 11742
rect 50204 11396 50260 11406
rect 50204 11302 50260 11340
rect 50876 11282 50932 11676
rect 50876 11230 50878 11282
rect 50930 11230 50932 11282
rect 50876 11218 50932 11230
rect 50988 11394 51044 12350
rect 51212 12178 51268 13916
rect 51212 12126 51214 12178
rect 51266 12126 51268 12178
rect 51212 12114 51268 12126
rect 51772 12180 51828 16828
rect 51884 15314 51940 15326
rect 51884 15262 51886 15314
rect 51938 15262 51940 15314
rect 51884 14868 51940 15262
rect 51884 14802 51940 14812
rect 51996 14700 52052 17388
rect 52108 17378 52164 17388
rect 52444 16996 52500 20748
rect 52892 20802 52948 20814
rect 52892 20750 52894 20802
rect 52946 20750 52948 20802
rect 52892 20580 52948 20750
rect 52892 20514 52948 20524
rect 52780 19348 52836 19358
rect 52668 19346 52836 19348
rect 52668 19294 52782 19346
rect 52834 19294 52836 19346
rect 52668 19292 52836 19294
rect 52556 19236 52612 19246
rect 52668 19236 52724 19292
rect 52780 19282 52836 19292
rect 53004 19348 53060 22988
rect 53116 22930 53172 22942
rect 53116 22878 53118 22930
rect 53170 22878 53172 22930
rect 53116 21698 53172 22878
rect 53116 21646 53118 21698
rect 53170 21646 53172 21698
rect 53116 21634 53172 21646
rect 53900 21588 53956 21598
rect 53900 21494 53956 21532
rect 52612 19180 52724 19236
rect 52892 19236 52948 19246
rect 53004 19236 53060 19292
rect 53788 19348 53844 19358
rect 53788 19254 53844 19292
rect 52892 19234 53060 19236
rect 52892 19182 52894 19234
rect 52946 19182 53060 19234
rect 52892 19180 53060 19182
rect 53228 19234 53284 19246
rect 53228 19182 53230 19234
rect 53282 19182 53284 19234
rect 52556 19170 52612 19180
rect 52892 19170 52948 19180
rect 52780 19124 52836 19134
rect 52668 19122 52836 19124
rect 52668 19070 52782 19122
rect 52834 19070 52836 19122
rect 52668 19068 52836 19070
rect 52668 19012 52724 19068
rect 52780 19058 52836 19068
rect 53116 19124 53172 19134
rect 53116 19030 53172 19068
rect 52668 18946 52724 18956
rect 52892 17668 52948 17678
rect 52892 17574 52948 17612
rect 52780 17556 52836 17566
rect 52780 17108 52836 17500
rect 53228 17444 53284 19182
rect 54012 19236 54068 27468
rect 54236 26852 54292 26862
rect 54236 26402 54292 26796
rect 54908 26852 54964 28590
rect 54908 26786 54964 26796
rect 55020 29540 55076 29550
rect 55020 29426 55076 29484
rect 55020 29374 55022 29426
rect 55074 29374 55076 29426
rect 54236 26350 54238 26402
rect 54290 26350 54292 26402
rect 54236 26338 54292 26350
rect 54348 26404 54404 26414
rect 54348 26310 54404 26348
rect 55020 26404 55076 29374
rect 54124 26292 54180 26302
rect 54124 26198 54180 26236
rect 55020 26290 55076 26348
rect 55020 26238 55022 26290
rect 55074 26238 55076 26290
rect 55020 26226 55076 26238
rect 54796 26066 54852 26078
rect 54796 26014 54798 26066
rect 54850 26014 54852 26066
rect 54460 25506 54516 25518
rect 54460 25454 54462 25506
rect 54514 25454 54516 25506
rect 54460 24612 54516 25454
rect 54684 25508 54740 25518
rect 54796 25508 54852 26014
rect 54684 25506 54852 25508
rect 54684 25454 54686 25506
rect 54738 25454 54852 25506
rect 54684 25452 54852 25454
rect 54908 25732 54964 25742
rect 54908 25506 54964 25676
rect 54908 25454 54910 25506
rect 54962 25454 54964 25506
rect 54572 24724 54628 24734
rect 54572 24630 54628 24668
rect 54460 24546 54516 24556
rect 54684 24500 54740 25452
rect 54908 25442 54964 25454
rect 54796 25284 54852 25294
rect 55132 25284 55188 35308
rect 55356 34804 55412 36430
rect 56028 36372 56084 36382
rect 55580 36370 56084 36372
rect 55580 36318 56030 36370
rect 56082 36318 56084 36370
rect 55580 36316 56084 36318
rect 55580 35922 55636 36316
rect 56028 36306 56084 36316
rect 55580 35870 55582 35922
rect 55634 35870 55636 35922
rect 55580 35858 55636 35870
rect 56028 35700 56084 35710
rect 56028 35606 56084 35644
rect 55468 35588 55524 35598
rect 55468 35494 55524 35532
rect 56700 35586 56756 35598
rect 56700 35534 56702 35586
rect 56754 35534 56756 35586
rect 56700 35364 56756 35534
rect 56700 35298 56756 35308
rect 55468 34804 55524 34814
rect 55356 34802 55524 34804
rect 55356 34750 55470 34802
rect 55522 34750 55524 34802
rect 55356 34748 55524 34750
rect 55244 33796 55300 33806
rect 55244 30212 55300 33740
rect 55356 33346 55412 34748
rect 55468 34738 55524 34748
rect 56028 33460 56084 33470
rect 56028 33366 56084 33404
rect 55356 33294 55358 33346
rect 55410 33294 55412 33346
rect 55356 31778 55412 33294
rect 57372 32788 57428 32798
rect 57372 32694 57428 32732
rect 57708 32452 57764 32462
rect 57820 32452 57876 36990
rect 57708 32450 57876 32452
rect 57708 32398 57710 32450
rect 57762 32398 57876 32450
rect 57708 32396 57876 32398
rect 57708 32386 57764 32396
rect 55356 31726 55358 31778
rect 55410 31726 55412 31778
rect 55356 31714 55412 31726
rect 56028 31668 56084 31678
rect 56028 31574 56084 31612
rect 55244 30210 55860 30212
rect 55244 30158 55246 30210
rect 55298 30158 55860 30210
rect 55244 30156 55860 30158
rect 55244 30146 55300 30156
rect 55804 29650 55860 30156
rect 55804 29598 55806 29650
rect 55858 29598 55860 29650
rect 55804 29586 55860 29598
rect 55244 29316 55300 29326
rect 55580 29316 55636 29326
rect 55244 29314 55636 29316
rect 55244 29262 55246 29314
rect 55298 29262 55582 29314
rect 55634 29262 55636 29314
rect 55244 29260 55636 29262
rect 55244 29250 55300 29260
rect 55580 29250 55636 29260
rect 55916 29202 55972 29214
rect 55916 29150 55918 29202
rect 55970 29150 55972 29202
rect 55916 28756 55972 29150
rect 56028 28756 56084 28766
rect 55916 28754 56084 28756
rect 55916 28702 56030 28754
rect 56082 28702 56084 28754
rect 55916 28700 56084 28702
rect 56028 28690 56084 28700
rect 55356 28642 55412 28654
rect 55356 28590 55358 28642
rect 55410 28590 55412 28642
rect 55356 26962 55412 28590
rect 55356 26910 55358 26962
rect 55410 26910 55412 26962
rect 55244 26178 55300 26190
rect 55244 26126 55246 26178
rect 55298 26126 55300 26178
rect 55244 25732 55300 26126
rect 55244 25666 55300 25676
rect 54796 25190 54852 25228
rect 54908 25228 55188 25284
rect 55356 25506 55412 26910
rect 58044 26908 58100 37884
rect 58156 37154 58212 37166
rect 58156 37102 58158 37154
rect 58210 37102 58212 37154
rect 58156 37042 58212 37102
rect 58156 36990 58158 37042
rect 58210 36990 58212 37042
rect 58156 36978 58212 36990
rect 58156 36594 58212 36606
rect 58156 36542 58158 36594
rect 58210 36542 58212 36594
rect 58156 35812 58212 36542
rect 58156 35746 58212 35756
rect 58156 33458 58212 33470
rect 58156 33406 58158 33458
rect 58210 33406 58212 33458
rect 58156 33348 58212 33406
rect 58156 33282 58212 33292
rect 58156 32788 58212 32798
rect 58156 32694 58212 32732
rect 58156 31890 58212 31902
rect 58156 31838 58158 31890
rect 58210 31838 58212 31890
rect 58156 31780 58212 31838
rect 58156 31714 58212 31724
rect 58156 28756 58212 28766
rect 58156 28662 58212 28700
rect 55468 26852 55524 26862
rect 55468 26402 55524 26796
rect 57596 26852 57652 26862
rect 57596 26514 57652 26796
rect 57596 26462 57598 26514
rect 57650 26462 57652 26514
rect 57596 26450 57652 26462
rect 57820 26852 58100 26908
rect 58156 26852 58212 26862
rect 57820 26514 57876 26852
rect 57820 26462 57822 26514
rect 57874 26462 57876 26514
rect 57820 26450 57876 26462
rect 58156 26514 58212 26796
rect 58156 26462 58158 26514
rect 58210 26462 58212 26514
rect 58156 26450 58212 26462
rect 55468 26350 55470 26402
rect 55522 26350 55524 26402
rect 55468 26338 55524 26350
rect 55692 26292 55748 26302
rect 55692 25620 55748 26236
rect 55692 25554 55748 25564
rect 58156 25620 58212 25630
rect 58156 25526 58212 25564
rect 55356 25454 55358 25506
rect 55410 25454 55412 25506
rect 54796 24500 54852 24510
rect 54684 24498 54852 24500
rect 54684 24446 54798 24498
rect 54850 24446 54852 24498
rect 54684 24444 54852 24446
rect 54796 24388 54852 24444
rect 54796 24322 54852 24332
rect 54684 22930 54740 22942
rect 54684 22878 54686 22930
rect 54738 22878 54740 22930
rect 54684 22820 54740 22878
rect 54684 22754 54740 22764
rect 54796 20132 54852 20142
rect 54908 20132 54964 25228
rect 55132 24500 55188 24510
rect 55020 24444 55132 24500
rect 55020 23154 55076 24444
rect 55132 24406 55188 24444
rect 55356 23938 55412 25454
rect 56028 25394 56084 25406
rect 56028 25342 56030 25394
rect 56082 25342 56084 25394
rect 56028 25284 56084 25342
rect 56028 25218 56084 25228
rect 55916 24946 55972 24958
rect 55916 24894 55918 24946
rect 55970 24894 55972 24946
rect 55580 24612 55636 24622
rect 55580 24518 55636 24556
rect 55356 23886 55358 23938
rect 55410 23886 55412 23938
rect 55356 23874 55412 23886
rect 55804 24500 55860 24510
rect 55692 23266 55748 23278
rect 55692 23214 55694 23266
rect 55746 23214 55748 23266
rect 55020 23102 55022 23154
rect 55074 23102 55076 23154
rect 55020 23090 55076 23102
rect 55244 23156 55300 23166
rect 55692 23156 55748 23214
rect 55804 23268 55860 24444
rect 55916 24052 55972 24894
rect 56028 24724 56084 24734
rect 56700 24724 56756 24734
rect 56028 24722 56756 24724
rect 56028 24670 56030 24722
rect 56082 24670 56702 24722
rect 56754 24670 56756 24722
rect 56028 24668 56756 24670
rect 56028 24658 56084 24668
rect 56700 24658 56756 24668
rect 56924 24724 56980 24734
rect 56028 24500 56084 24510
rect 56084 24444 56196 24500
rect 56028 24434 56084 24444
rect 56028 24052 56084 24062
rect 55916 24050 56084 24052
rect 55916 23998 56030 24050
rect 56082 23998 56084 24050
rect 55916 23996 56084 23998
rect 56028 23986 56084 23996
rect 55916 23268 55972 23278
rect 55804 23266 55972 23268
rect 55804 23214 55918 23266
rect 55970 23214 55972 23266
rect 55804 23212 55972 23214
rect 55916 23202 55972 23212
rect 55300 23100 55748 23156
rect 55244 23062 55300 23100
rect 55580 22930 55636 22942
rect 55580 22878 55582 22930
rect 55634 22878 55636 22930
rect 55244 22820 55300 22830
rect 55300 22764 55412 22820
rect 55244 22754 55300 22764
rect 55244 22370 55300 22382
rect 55244 22318 55246 22370
rect 55298 22318 55300 22370
rect 55244 21588 55300 22318
rect 55244 20692 55300 21532
rect 55356 21586 55412 22764
rect 55356 21534 55358 21586
rect 55410 21534 55412 21586
rect 55356 21522 55412 21534
rect 55468 21588 55524 21598
rect 55580 21588 55636 22878
rect 55692 22484 55748 23100
rect 55692 22418 55748 22428
rect 56028 22260 56084 22270
rect 55804 22258 56084 22260
rect 55804 22206 56030 22258
rect 56082 22206 56084 22258
rect 55804 22204 56084 22206
rect 55804 21698 55860 22204
rect 56028 22194 56084 22204
rect 55804 21646 55806 21698
rect 55858 21646 55860 21698
rect 55804 21634 55860 21646
rect 55468 21586 55636 21588
rect 55468 21534 55470 21586
rect 55522 21534 55636 21586
rect 55468 21532 55636 21534
rect 55468 21522 55524 21532
rect 55692 21476 55748 21486
rect 56140 21476 56196 24444
rect 56588 24498 56644 24510
rect 56588 24446 56590 24498
rect 56642 24446 56644 24498
rect 56588 24388 56644 24446
rect 56588 24322 56644 24332
rect 56924 24052 56980 24668
rect 56924 23986 56980 23996
rect 58156 24052 58212 24062
rect 58156 23958 58212 23996
rect 58156 22484 58212 22494
rect 58156 22390 58212 22428
rect 57820 21700 57876 21710
rect 57820 21606 57876 21644
rect 58156 21586 58212 21598
rect 58156 21534 58158 21586
rect 58210 21534 58212 21586
rect 55692 21474 56196 21476
rect 55692 21422 55694 21474
rect 55746 21422 56196 21474
rect 55692 21420 56196 21422
rect 57596 21476 57652 21486
rect 58156 21476 58212 21534
rect 57596 21474 58212 21476
rect 57596 21422 57598 21474
rect 57650 21422 58212 21474
rect 57596 21420 58212 21422
rect 55692 21410 55748 21420
rect 57596 21410 57652 21420
rect 58156 21140 58212 21420
rect 58156 21074 58212 21084
rect 55356 20692 55412 20702
rect 55244 20690 55412 20692
rect 55244 20638 55358 20690
rect 55410 20638 55412 20690
rect 55244 20636 55412 20638
rect 54796 20130 54908 20132
rect 54796 20078 54798 20130
rect 54850 20078 54908 20130
rect 54796 20076 54908 20078
rect 54796 20066 54852 20076
rect 54908 20038 54964 20076
rect 54460 20018 54516 20030
rect 54460 19966 54462 20018
rect 54514 19966 54516 20018
rect 54460 19348 54516 19966
rect 54012 19170 54068 19180
rect 54348 19292 54460 19348
rect 54236 19122 54292 19134
rect 54236 19070 54238 19122
rect 54290 19070 54292 19122
rect 53228 17378 53284 17388
rect 54012 18338 54068 18350
rect 54012 18286 54014 18338
rect 54066 18286 54068 18338
rect 54012 17444 54068 18286
rect 54012 17378 54068 17388
rect 52780 17106 53060 17108
rect 52780 17054 52782 17106
rect 52834 17054 53060 17106
rect 52780 17052 53060 17054
rect 52780 17042 52836 17052
rect 52332 16884 52388 16894
rect 52444 16884 52500 16940
rect 52332 16882 52500 16884
rect 52332 16830 52334 16882
rect 52386 16830 52500 16882
rect 52332 16828 52500 16830
rect 52332 16818 52388 16828
rect 52668 16660 52724 16670
rect 52108 15426 52164 15438
rect 52108 15374 52110 15426
rect 52162 15374 52164 15426
rect 52108 15204 52164 15374
rect 52668 15314 52724 16604
rect 53004 16098 53060 17052
rect 54012 16884 54068 16894
rect 54236 16884 54292 19070
rect 54348 18564 54404 19292
rect 54460 19282 54516 19292
rect 54572 20018 54628 20030
rect 54572 19966 54574 20018
rect 54626 19966 54628 20018
rect 54460 19124 54516 19134
rect 54572 19124 54628 19966
rect 55020 20020 55076 20030
rect 55020 20018 55188 20020
rect 55020 19966 55022 20018
rect 55074 19966 55188 20018
rect 55020 19964 55188 19966
rect 55020 19954 55076 19964
rect 54684 19908 54740 19918
rect 54684 19814 54740 19852
rect 54796 19348 54852 19358
rect 54796 19346 55076 19348
rect 54796 19294 54798 19346
rect 54850 19294 55076 19346
rect 54796 19292 55076 19294
rect 54796 19282 54852 19292
rect 54684 19236 54740 19246
rect 54684 19142 54740 19180
rect 54516 19068 54628 19124
rect 54460 19030 54516 19068
rect 54796 19012 54852 19022
rect 54796 18918 54852 18956
rect 55020 18788 55076 19292
rect 55132 19012 55188 19964
rect 55356 19236 55412 20636
rect 56140 20132 56196 20142
rect 56140 20038 56196 20076
rect 55468 19908 55524 19918
rect 55468 19814 55524 19852
rect 55580 19796 55636 19806
rect 55580 19794 56084 19796
rect 55580 19742 55582 19794
rect 55634 19742 56084 19794
rect 55580 19740 56084 19742
rect 55580 19730 55636 19740
rect 56028 19346 56084 19740
rect 56028 19294 56030 19346
rect 56082 19294 56084 19346
rect 56028 19282 56084 19294
rect 58156 19348 58212 19358
rect 58156 19254 58212 19292
rect 55916 19236 55972 19246
rect 55356 19234 55524 19236
rect 55356 19182 55358 19234
rect 55410 19182 55524 19234
rect 55356 19180 55524 19182
rect 55356 19170 55412 19180
rect 55132 18946 55188 18956
rect 55020 18732 55300 18788
rect 54460 18564 54516 18574
rect 54348 18562 54516 18564
rect 54348 18510 54462 18562
rect 54514 18510 54516 18562
rect 54348 18508 54516 18510
rect 55244 18564 55300 18732
rect 55356 18564 55412 18574
rect 55244 18562 55412 18564
rect 55244 18510 55358 18562
rect 55410 18510 55412 18562
rect 55244 18508 55412 18510
rect 54460 18498 54516 18508
rect 55356 18498 55412 18508
rect 55468 18452 55524 19180
rect 55916 18452 55972 19180
rect 56028 18452 56084 18462
rect 55916 18450 56084 18452
rect 55916 18398 56030 18450
rect 56082 18398 56084 18450
rect 55916 18396 56084 18398
rect 55468 18386 55524 18396
rect 56028 18386 56084 18396
rect 55244 18340 55300 18350
rect 54348 18228 54404 18238
rect 54348 18226 54740 18228
rect 54348 18174 54350 18226
rect 54402 18174 54740 18226
rect 54348 18172 54740 18174
rect 54348 18162 54404 18172
rect 54012 16882 54292 16884
rect 54012 16830 54014 16882
rect 54066 16830 54292 16882
rect 54012 16828 54292 16830
rect 53004 16046 53006 16098
rect 53058 16046 53060 16098
rect 53004 16034 53060 16046
rect 53900 16658 53956 16670
rect 53900 16606 53902 16658
rect 53954 16606 53956 16658
rect 53228 15986 53284 15998
rect 53228 15934 53230 15986
rect 53282 15934 53284 15986
rect 53004 15540 53060 15550
rect 53228 15540 53284 15934
rect 53340 15988 53396 15998
rect 53788 15988 53844 15998
rect 53340 15986 53732 15988
rect 53340 15934 53342 15986
rect 53394 15934 53732 15986
rect 53340 15932 53732 15934
rect 53340 15922 53396 15932
rect 53004 15538 53284 15540
rect 53004 15486 53006 15538
rect 53058 15486 53284 15538
rect 53004 15484 53284 15486
rect 53676 15538 53732 15932
rect 53788 15894 53844 15932
rect 53676 15486 53678 15538
rect 53730 15486 53732 15538
rect 53004 15474 53060 15484
rect 53452 15426 53508 15438
rect 53452 15374 53454 15426
rect 53506 15374 53508 15426
rect 52668 15262 52670 15314
rect 52722 15262 52724 15314
rect 52444 15204 52500 15214
rect 52108 15202 52500 15204
rect 52108 15150 52446 15202
rect 52498 15150 52500 15202
rect 52108 15148 52500 15150
rect 52444 15092 52500 15148
rect 52444 15026 52500 15036
rect 52668 14756 52724 15262
rect 53340 15314 53396 15326
rect 53340 15262 53342 15314
rect 53394 15262 53396 15314
rect 53340 15148 53396 15262
rect 51884 14644 52052 14700
rect 52444 14700 52724 14756
rect 52780 15092 52836 15102
rect 51884 14578 51940 14588
rect 51996 14532 52052 14542
rect 51996 13972 52052 14476
rect 51996 13878 52052 13916
rect 52444 13748 52500 14700
rect 52444 13654 52500 13692
rect 52668 13748 52724 13758
rect 52780 13748 52836 15036
rect 53228 15092 53396 15148
rect 53452 15092 53508 15374
rect 52668 13746 52836 13748
rect 52668 13694 52670 13746
rect 52722 13694 52836 13746
rect 52668 13692 52836 13694
rect 52668 13682 52724 13692
rect 51884 13636 51940 13646
rect 51884 13542 51940 13580
rect 52780 13188 52836 13692
rect 52892 13858 52948 13870
rect 52892 13806 52894 13858
rect 52946 13806 52948 13858
rect 52892 13636 52948 13806
rect 52892 13412 52948 13580
rect 53228 13748 53284 15092
rect 53452 15026 53508 15036
rect 53676 14642 53732 15486
rect 53900 15148 53956 16606
rect 54012 16212 54068 16828
rect 54012 16146 54068 16156
rect 54572 15988 54628 15998
rect 54572 15894 54628 15932
rect 53676 14590 53678 14642
rect 53730 14590 53732 14642
rect 53676 14578 53732 14590
rect 53788 15092 53956 15148
rect 54348 15204 54404 15214
rect 53340 14532 53396 14542
rect 53340 14438 53396 14476
rect 53004 13524 53060 13534
rect 53004 13522 53172 13524
rect 53004 13470 53006 13522
rect 53058 13470 53172 13522
rect 53004 13468 53172 13470
rect 53004 13458 53060 13468
rect 52892 13346 52948 13356
rect 52780 13132 53060 13188
rect 52668 12962 52724 12974
rect 52668 12910 52670 12962
rect 52722 12910 52724 12962
rect 52108 12292 52164 12302
rect 52108 12198 52164 12236
rect 51772 12178 52052 12180
rect 51772 12126 51774 12178
rect 51826 12126 52052 12178
rect 51772 12124 52052 12126
rect 51772 12114 51828 12124
rect 51996 11506 52052 12124
rect 51996 11454 51998 11506
rect 52050 11454 52052 11506
rect 51996 11442 52052 11454
rect 52668 11508 52724 12910
rect 53004 12962 53060 13132
rect 53004 12910 53006 12962
rect 53058 12910 53060 12962
rect 53004 12898 53060 12910
rect 52892 12852 52948 12862
rect 52892 12758 52948 12796
rect 52780 12740 52836 12750
rect 52780 12292 52836 12684
rect 52780 12178 52836 12236
rect 52780 12126 52782 12178
rect 52834 12126 52836 12178
rect 52780 12114 52836 12126
rect 53004 12180 53060 12190
rect 53116 12180 53172 13468
rect 53228 12962 53284 13692
rect 53228 12910 53230 12962
rect 53282 12910 53284 12962
rect 53228 12898 53284 12910
rect 53340 13412 53396 13422
rect 53340 12852 53396 13356
rect 53788 12964 53844 15092
rect 54348 14756 54404 15148
rect 53900 14700 54404 14756
rect 53900 13636 53956 14700
rect 54348 14698 54404 14700
rect 54348 14646 54350 14698
rect 54402 14646 54404 14698
rect 54348 14624 54404 14646
rect 54572 14530 54628 14542
rect 54572 14478 54574 14530
rect 54626 14478 54628 14530
rect 54012 14420 54068 14430
rect 54572 14420 54628 14478
rect 54012 14418 54628 14420
rect 54012 14366 54014 14418
rect 54066 14366 54628 14418
rect 54012 14364 54628 14366
rect 54012 14354 54068 14364
rect 54012 13636 54068 13646
rect 53900 13634 54068 13636
rect 53900 13582 54014 13634
rect 54066 13582 54068 13634
rect 53900 13580 54068 13582
rect 54012 13188 54068 13580
rect 54012 13132 54404 13188
rect 53340 12786 53396 12796
rect 53564 12908 53844 12964
rect 53004 12178 53172 12180
rect 53004 12126 53006 12178
rect 53058 12126 53172 12178
rect 53004 12124 53172 12126
rect 53004 12114 53060 12124
rect 53340 11956 53396 11966
rect 53340 11862 53396 11900
rect 53116 11508 53172 11518
rect 52668 11452 53116 11508
rect 50988 11342 50990 11394
rect 51042 11342 51044 11394
rect 50316 11172 50372 11182
rect 49756 10722 49924 10724
rect 49756 10670 49758 10722
rect 49810 10670 49924 10722
rect 49756 10668 49924 10670
rect 50092 10724 50148 10734
rect 49756 10658 49812 10668
rect 50092 10630 50148 10668
rect 50316 10722 50372 11116
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 50316 10670 50318 10722
rect 50370 10670 50372 10722
rect 50316 10658 50372 10670
rect 50988 10724 51044 11342
rect 53116 11394 53172 11452
rect 53564 11396 53620 12908
rect 54012 12852 54068 12862
rect 54012 12850 54180 12852
rect 54012 12798 54014 12850
rect 54066 12798 54180 12850
rect 54012 12796 54180 12798
rect 54012 12786 54068 12796
rect 53676 12738 53732 12750
rect 53676 12686 53678 12738
rect 53730 12686 53732 12738
rect 53676 12180 53732 12686
rect 53900 12740 53956 12750
rect 53900 12646 53956 12684
rect 53676 12124 53956 12180
rect 53116 11342 53118 11394
rect 53170 11342 53172 11394
rect 53116 11330 53172 11342
rect 53228 11394 53620 11396
rect 53228 11342 53566 11394
rect 53618 11342 53620 11394
rect 53228 11340 53620 11342
rect 51436 11284 51492 11294
rect 51436 11190 51492 11228
rect 53004 11284 53060 11294
rect 51324 11172 51380 11182
rect 51324 11078 51380 11116
rect 52108 11172 52164 11182
rect 52780 11172 52836 11182
rect 52108 11170 52836 11172
rect 52108 11118 52110 11170
rect 52162 11118 52782 11170
rect 52834 11118 52836 11170
rect 52108 11116 52836 11118
rect 52108 11106 52164 11116
rect 52780 11106 52836 11116
rect 53004 11170 53060 11228
rect 53004 11118 53006 11170
rect 53058 11118 53060 11170
rect 53004 11106 53060 11118
rect 50988 10658 51044 10668
rect 49868 10498 49924 10510
rect 49868 10446 49870 10498
rect 49922 10446 49924 10498
rect 49868 9826 49924 10446
rect 49868 9774 49870 9826
rect 49922 9774 49924 9826
rect 49868 9762 49924 9774
rect 50540 9828 50596 9838
rect 50540 9734 50596 9772
rect 51324 9828 51380 9838
rect 49644 9660 49812 9716
rect 49644 9492 49700 9502
rect 49084 9214 49086 9266
rect 49138 9214 49140 9266
rect 49084 9202 49140 9214
rect 49420 9436 49644 9492
rect 49756 9492 49812 9660
rect 49980 9602 50036 9614
rect 49980 9550 49982 9602
rect 50034 9550 50036 9602
rect 49980 9492 50036 9550
rect 49756 9436 49924 9492
rect 48748 9042 48916 9044
rect 48748 8990 48750 9042
rect 48802 8990 48916 9042
rect 48748 8988 48916 8990
rect 48972 9044 49028 9054
rect 47180 8430 47182 8482
rect 47234 8430 47236 8482
rect 47180 8418 47236 8430
rect 47628 8484 47684 8494
rect 47628 8390 47684 8428
rect 48748 8484 48804 8988
rect 48972 8950 49028 8988
rect 49420 9042 49476 9436
rect 49644 9426 49700 9436
rect 49756 9268 49812 9278
rect 49644 9266 49812 9268
rect 49644 9214 49758 9266
rect 49810 9214 49812 9266
rect 49644 9212 49812 9214
rect 49644 9156 49700 9212
rect 49644 9090 49700 9100
rect 49420 8990 49422 9042
rect 49474 8990 49476 9042
rect 49420 8978 49476 8990
rect 48748 8418 48804 8428
rect 49756 8370 49812 9212
rect 49868 9266 49924 9436
rect 49980 9426 50036 9436
rect 50092 9602 50148 9614
rect 50092 9550 50094 9602
rect 50146 9550 50148 9602
rect 49868 9214 49870 9266
rect 49922 9214 49924 9266
rect 49868 9202 49924 9214
rect 49980 9156 50036 9166
rect 50092 9156 50148 9550
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 51324 9266 51380 9772
rect 52108 9828 52164 9838
rect 52892 9828 52948 9838
rect 52108 9826 52948 9828
rect 52108 9774 52110 9826
rect 52162 9774 52894 9826
rect 52946 9774 52948 9826
rect 52108 9772 52948 9774
rect 51324 9214 51326 9266
rect 51378 9214 51380 9266
rect 51324 9202 51380 9214
rect 51660 9604 51716 9614
rect 49980 9154 50092 9156
rect 49980 9102 49982 9154
rect 50034 9102 50092 9154
rect 49980 9100 50092 9102
rect 49980 9090 50036 9100
rect 50092 9062 50148 9100
rect 50988 9042 51044 9054
rect 50988 8990 50990 9042
rect 51042 8990 51044 9042
rect 49756 8318 49758 8370
rect 49810 8318 49812 8370
rect 49756 8306 49812 8318
rect 49980 8820 50036 8830
rect 49980 8258 50036 8764
rect 50988 8428 51044 8990
rect 51212 9044 51268 9054
rect 51212 8950 51268 8988
rect 51436 9042 51492 9054
rect 51436 8990 51438 9042
rect 51490 8990 51492 9042
rect 50316 8372 51044 8428
rect 50316 8370 50372 8372
rect 50316 8318 50318 8370
rect 50370 8318 50372 8370
rect 50316 8306 50372 8318
rect 49980 8206 49982 8258
rect 50034 8206 50036 8258
rect 49980 8194 50036 8206
rect 46284 7858 46340 7868
rect 46844 8146 46900 8158
rect 47516 8148 47572 8158
rect 46844 8094 46846 8146
rect 46898 8094 46900 8146
rect 46060 7700 46116 7710
rect 46060 7698 46676 7700
rect 46060 7646 46062 7698
rect 46114 7646 46676 7698
rect 46060 7644 46676 7646
rect 46060 7634 46116 7644
rect 45948 7476 46004 7486
rect 45724 6750 45726 6802
rect 45778 6750 45780 6802
rect 45724 6738 45780 6750
rect 45836 7420 45948 7476
rect 44380 6626 44436 6636
rect 45052 6692 45108 6702
rect 45052 6598 45108 6636
rect 45388 6690 45444 6702
rect 45388 6638 45390 6690
rect 45442 6638 45444 6690
rect 45388 6580 45444 6638
rect 44828 6468 44884 6478
rect 44828 5346 44884 6412
rect 45388 6356 45444 6524
rect 45388 6290 45444 6300
rect 45500 6692 45556 6702
rect 44828 5294 44830 5346
rect 44882 5294 44884 5346
rect 44828 5282 44884 5294
rect 45500 6132 45556 6636
rect 45836 6690 45892 7420
rect 45948 7382 46004 7420
rect 46396 7476 46452 7486
rect 46396 7474 46564 7476
rect 46396 7422 46398 7474
rect 46450 7422 46564 7474
rect 46396 7420 46564 7422
rect 46396 7410 46452 7420
rect 45836 6638 45838 6690
rect 45890 6638 45892 6690
rect 45836 6626 45892 6638
rect 46172 6692 46228 6702
rect 46060 6580 46116 6590
rect 46060 6486 46116 6524
rect 45612 6468 45668 6478
rect 45612 6374 45668 6412
rect 45500 5234 45556 6076
rect 46172 5906 46228 6636
rect 46396 6578 46452 6590
rect 46396 6526 46398 6578
rect 46450 6526 46452 6578
rect 46396 6356 46452 6526
rect 46396 6290 46452 6300
rect 46508 6020 46564 7420
rect 46620 7474 46676 7644
rect 46620 7422 46622 7474
rect 46674 7422 46676 7474
rect 46620 7410 46676 7422
rect 46844 7474 46900 8094
rect 47180 8146 47572 8148
rect 47180 8094 47518 8146
rect 47570 8094 47572 8146
rect 47180 8092 47572 8094
rect 47068 8036 47124 8046
rect 47068 7942 47124 7980
rect 47180 7812 47236 8092
rect 47516 8082 47572 8092
rect 47628 8036 47684 8046
rect 47628 7942 47684 7980
rect 49644 8034 49700 8046
rect 49644 7982 49646 8034
rect 49698 7982 49700 8034
rect 46956 7756 47236 7812
rect 47292 7924 47348 7934
rect 46956 7698 47012 7756
rect 46956 7646 46958 7698
rect 47010 7646 47012 7698
rect 46956 7634 47012 7646
rect 47068 7588 47124 7598
rect 47292 7588 47348 7868
rect 49644 7924 49700 7982
rect 49644 7858 49700 7868
rect 49868 8034 49924 8046
rect 49868 7982 49870 8034
rect 49922 7982 49924 8034
rect 49868 7700 49924 7982
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 49980 7700 50036 7710
rect 50988 7700 51044 8372
rect 51436 8260 51492 8990
rect 51660 9042 51716 9548
rect 51660 8990 51662 9042
rect 51714 8990 51716 9042
rect 51660 8978 51716 8990
rect 51436 8194 51492 8204
rect 49868 7698 50260 7700
rect 49868 7646 49982 7698
rect 50034 7646 50260 7698
rect 49868 7644 50260 7646
rect 49980 7634 50036 7644
rect 47068 7586 47348 7588
rect 47068 7534 47070 7586
rect 47122 7534 47348 7586
rect 47068 7532 47348 7534
rect 47068 7522 47124 7532
rect 46844 7422 46846 7474
rect 46898 7422 46900 7474
rect 46844 7252 46900 7422
rect 46620 7196 46900 7252
rect 47404 7474 47460 7486
rect 47404 7422 47406 7474
rect 47458 7422 47460 7474
rect 46620 6802 46676 7196
rect 46620 6750 46622 6802
rect 46674 6750 46676 6802
rect 46620 6738 46676 6750
rect 47180 6692 47236 6702
rect 47180 6598 47236 6636
rect 46956 6580 47012 6590
rect 46620 6468 46676 6478
rect 46620 6374 46676 6412
rect 46956 6020 47012 6524
rect 47404 6580 47460 7422
rect 50092 7474 50148 7486
rect 50092 7422 50094 7474
rect 50146 7422 50148 7474
rect 49980 7250 50036 7262
rect 49980 7198 49982 7250
rect 50034 7198 50036 7250
rect 48972 6916 49028 6926
rect 48972 6822 49028 6860
rect 49644 6916 49700 6926
rect 49308 6804 49364 6814
rect 49308 6692 49364 6748
rect 49308 6690 49588 6692
rect 49308 6638 49310 6690
rect 49362 6638 49588 6690
rect 49308 6636 49588 6638
rect 49308 6626 49364 6636
rect 47404 6514 47460 6524
rect 49084 6466 49140 6478
rect 49084 6414 49086 6466
rect 49138 6414 49140 6466
rect 46508 5964 46676 6020
rect 46172 5854 46174 5906
rect 46226 5854 46228 5906
rect 46172 5842 46228 5854
rect 46508 5796 46564 5806
rect 46284 5794 46564 5796
rect 46284 5742 46510 5794
rect 46562 5742 46564 5794
rect 46284 5740 46564 5742
rect 46284 5460 46340 5740
rect 46508 5730 46564 5740
rect 46620 5796 46676 5964
rect 46956 5906 47012 5964
rect 47852 6020 47908 6030
rect 47852 5926 47908 5964
rect 46956 5854 46958 5906
rect 47010 5854 47012 5906
rect 46956 5842 47012 5854
rect 47404 5908 47460 5918
rect 47404 5814 47460 5852
rect 46620 5572 46676 5740
rect 47964 5796 48020 5806
rect 47964 5702 48020 5740
rect 49084 5796 49140 6414
rect 49532 6468 49588 6636
rect 49644 6690 49700 6860
rect 49644 6638 49646 6690
rect 49698 6638 49700 6690
rect 49644 6626 49700 6638
rect 49868 6578 49924 6590
rect 49868 6526 49870 6578
rect 49922 6526 49924 6578
rect 49868 6468 49924 6526
rect 49532 6412 49924 6468
rect 49644 6132 49700 6142
rect 49644 6038 49700 6076
rect 49980 5908 50036 7198
rect 50092 6916 50148 7422
rect 50092 6822 50148 6860
rect 50204 6804 50260 7644
rect 50988 7634 51044 7644
rect 50204 6738 50260 6748
rect 50764 6804 50820 6814
rect 50764 6578 50820 6748
rect 52108 6692 52164 9772
rect 52892 9762 52948 9772
rect 52780 9604 52836 9614
rect 52780 9266 52836 9548
rect 52780 9214 52782 9266
rect 52834 9214 52836 9266
rect 52780 9202 52836 9214
rect 52892 9156 52948 9166
rect 52892 9062 52948 9100
rect 53004 9044 53060 9054
rect 53004 9042 53172 9044
rect 53004 8990 53006 9042
rect 53058 8990 53172 9042
rect 53004 8988 53172 8990
rect 53004 8978 53060 8988
rect 52332 8930 52388 8942
rect 52332 8878 52334 8930
rect 52386 8878 52388 8930
rect 52332 8820 52388 8878
rect 52220 7140 52276 7150
rect 52220 6802 52276 7084
rect 52332 7028 52388 8764
rect 52892 8260 52948 8270
rect 52332 6962 52388 6972
rect 52668 7250 52724 7262
rect 52668 7198 52670 7250
rect 52722 7198 52724 7250
rect 52668 6916 52724 7198
rect 52668 6850 52724 6860
rect 52780 7028 52836 7038
rect 52220 6750 52222 6802
rect 52274 6750 52276 6802
rect 52220 6738 52276 6750
rect 50764 6526 50766 6578
rect 50818 6526 50820 6578
rect 50764 6514 50820 6526
rect 51100 6580 51156 6590
rect 50428 6468 50484 6478
rect 50204 6466 50484 6468
rect 50204 6414 50430 6466
rect 50482 6414 50484 6466
rect 50204 6412 50484 6414
rect 50092 6132 50148 6142
rect 50092 6018 50148 6076
rect 50092 5966 50094 6018
rect 50146 5966 50148 6018
rect 50092 5954 50148 5966
rect 50204 6018 50260 6412
rect 50428 6402 50484 6412
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 50204 5966 50206 6018
rect 50258 5966 50260 6018
rect 50204 5954 50260 5966
rect 49980 5842 50036 5852
rect 50316 5908 50372 5918
rect 50316 5814 50372 5852
rect 49084 5730 49140 5740
rect 45724 5404 46340 5460
rect 46396 5516 46676 5572
rect 50764 5682 50820 5694
rect 50764 5630 50766 5682
rect 50818 5630 50820 5682
rect 45724 5346 45780 5404
rect 45724 5294 45726 5346
rect 45778 5294 45780 5346
rect 45724 5282 45780 5294
rect 45500 5182 45502 5234
rect 45554 5182 45556 5234
rect 45500 5170 45556 5182
rect 46396 5234 46452 5516
rect 46396 5182 46398 5234
rect 46450 5182 46452 5234
rect 46396 5170 46452 5182
rect 49308 5124 49364 5134
rect 50764 5124 50820 5630
rect 50988 5124 51044 5134
rect 50764 5122 51044 5124
rect 50764 5070 50990 5122
rect 51042 5070 51044 5122
rect 50764 5068 51044 5070
rect 49308 5030 49364 5068
rect 50988 5058 51044 5068
rect 44940 5012 44996 5022
rect 44940 4918 44996 4956
rect 46508 5012 46564 5022
rect 48524 5012 48580 5022
rect 46060 4900 46116 4910
rect 46060 4806 46116 4844
rect 44044 4226 44212 4228
rect 44044 4174 44046 4226
rect 44098 4174 44212 4226
rect 44044 4172 44212 4174
rect 44492 4338 44548 4350
rect 44492 4286 44494 4338
rect 44546 4286 44548 4338
rect 44044 4162 44100 4172
rect 44492 3780 44548 4286
rect 45388 4116 45444 4126
rect 45388 4022 45444 4060
rect 44492 3714 44548 3724
rect 44380 3668 44436 3678
rect 44380 3574 44436 3612
rect 46508 3666 46564 4956
rect 47740 5010 48580 5012
rect 47740 4958 48526 5010
rect 48578 4958 48580 5010
rect 47740 4956 48580 4958
rect 47404 4900 47460 4910
rect 47404 4450 47460 4844
rect 47740 4562 47796 4956
rect 48524 4946 48580 4956
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 47740 4510 47742 4562
rect 47794 4510 47796 4562
rect 47740 4498 47796 4510
rect 47404 4398 47406 4450
rect 47458 4398 47460 4450
rect 47404 4386 47460 4398
rect 48076 4450 48132 4462
rect 48076 4398 48078 4450
rect 48130 4398 48132 4450
rect 46508 3614 46510 3666
rect 46562 3614 46564 3666
rect 46508 3602 46564 3614
rect 43708 3502 43710 3554
rect 43762 3502 43764 3554
rect 43708 3490 43764 3502
rect 47404 3556 47460 3566
rect 47404 3462 47460 3500
rect 45052 3444 45108 3454
rect 48076 3388 48132 4398
rect 48860 4226 48916 4238
rect 48860 4174 48862 4226
rect 48914 4174 48916 4226
rect 48860 3556 48916 4174
rect 50540 4228 50596 4238
rect 51100 4228 51156 6524
rect 52108 5236 52164 6636
rect 52780 6580 52836 6972
rect 52892 6804 52948 8204
rect 53116 8260 53172 8988
rect 53228 9042 53284 11340
rect 53564 11330 53620 11340
rect 53900 11954 53956 12124
rect 53900 11902 53902 11954
rect 53954 11902 53956 11954
rect 53676 11282 53732 11294
rect 53676 11230 53678 11282
rect 53730 11230 53732 11282
rect 53564 10836 53620 10846
rect 53676 10836 53732 11230
rect 53564 10834 53732 10836
rect 53564 10782 53566 10834
rect 53618 10782 53732 10834
rect 53564 10780 53732 10782
rect 53564 9156 53620 10780
rect 53228 8990 53230 9042
rect 53282 8990 53284 9042
rect 53228 8978 53284 8990
rect 53452 9044 53508 9054
rect 53564 9044 53620 9100
rect 53452 9042 53620 9044
rect 53452 8990 53454 9042
rect 53506 8990 53620 9042
rect 53452 8988 53620 8990
rect 53676 10498 53732 10510
rect 53676 10446 53678 10498
rect 53730 10446 53732 10498
rect 53676 9044 53732 10446
rect 53788 10386 53844 10398
rect 53788 10334 53790 10386
rect 53842 10334 53844 10386
rect 53788 10276 53844 10334
rect 53900 10276 53956 11902
rect 54012 11956 54068 11966
rect 54012 11862 54068 11900
rect 54012 11508 54068 11518
rect 54124 11508 54180 12796
rect 54068 11452 54180 11508
rect 54236 12740 54292 12750
rect 54236 11954 54292 12684
rect 54236 11902 54238 11954
rect 54290 11902 54292 11954
rect 54236 11844 54292 11902
rect 54012 11442 54068 11452
rect 54012 10276 54068 10286
rect 53788 10220 54012 10276
rect 54012 10210 54068 10220
rect 53788 9044 53844 9054
rect 53676 9042 53844 9044
rect 53676 8990 53790 9042
rect 53842 8990 53844 9042
rect 53676 8988 53844 8990
rect 53452 8978 53508 8988
rect 53788 8978 53844 8988
rect 54236 9042 54292 11788
rect 54236 8990 54238 9042
rect 54290 8990 54292 9042
rect 54012 8818 54068 8830
rect 54012 8766 54014 8818
rect 54066 8766 54068 8818
rect 54012 8372 54068 8766
rect 54012 8278 54068 8316
rect 53116 8148 53172 8204
rect 53900 8260 53956 8270
rect 53116 8146 53284 8148
rect 53116 8094 53118 8146
rect 53170 8094 53284 8146
rect 53116 8092 53284 8094
rect 53116 8082 53172 8092
rect 53116 7588 53172 7598
rect 53116 7494 53172 7532
rect 53228 7586 53284 8092
rect 53228 7534 53230 7586
rect 53282 7534 53284 7586
rect 53228 7522 53284 7534
rect 53340 7700 53396 7710
rect 53340 7588 53396 7644
rect 53788 7588 53844 7598
rect 53340 7586 53844 7588
rect 53340 7534 53342 7586
rect 53394 7534 53790 7586
rect 53842 7534 53844 7586
rect 53340 7532 53844 7534
rect 53900 7588 53956 8204
rect 54236 8148 54292 8990
rect 54348 8596 54404 13132
rect 54460 12740 54516 12750
rect 54460 12646 54516 12684
rect 54684 12628 54740 18172
rect 55244 16098 55300 18284
rect 55468 18228 55524 18238
rect 55468 18226 55972 18228
rect 55468 18174 55470 18226
rect 55522 18174 55972 18226
rect 55468 18172 55972 18174
rect 55468 18162 55524 18172
rect 55244 16046 55246 16098
rect 55298 16046 55300 16098
rect 55244 16034 55300 16046
rect 55356 17554 55412 17566
rect 55356 17502 55358 17554
rect 55410 17502 55412 17554
rect 55356 16884 55412 17502
rect 54908 15874 54964 15886
rect 54908 15822 54910 15874
rect 54962 15822 54964 15874
rect 54908 14644 54964 15822
rect 54908 14578 54964 14588
rect 55356 14530 55412 16828
rect 55916 16212 55972 18172
rect 56028 16212 56084 16222
rect 55916 16210 56084 16212
rect 55916 16158 56030 16210
rect 56082 16158 56084 16210
rect 55916 16156 56084 16158
rect 56028 16146 56084 16156
rect 58156 16212 58212 16222
rect 58156 16118 58212 16156
rect 57820 15428 57876 15438
rect 57820 15334 57876 15372
rect 57596 15316 57652 15326
rect 57596 15222 57652 15260
rect 58156 15316 58212 15326
rect 58156 15222 58212 15260
rect 58156 14868 58212 14878
rect 56028 14644 56084 14654
rect 56028 14550 56084 14588
rect 58156 14642 58212 14812
rect 58156 14590 58158 14642
rect 58210 14590 58212 14642
rect 58156 14578 58212 14590
rect 55356 14478 55358 14530
rect 55410 14478 55412 14530
rect 55356 14466 55412 14478
rect 54908 14308 54964 14318
rect 54908 14214 54964 14252
rect 55692 14308 55748 14318
rect 55692 13858 55748 14252
rect 55692 13806 55694 13858
rect 55746 13806 55748 13858
rect 55692 13794 55748 13806
rect 56028 13858 56084 13870
rect 56028 13806 56030 13858
rect 56082 13806 56084 13858
rect 56028 13074 56084 13806
rect 56028 13022 56030 13074
rect 56082 13022 56084 13074
rect 56028 13010 56084 13022
rect 58156 13074 58212 13086
rect 58156 13022 58158 13074
rect 58210 13022 58212 13074
rect 55244 12962 55300 12974
rect 55244 12910 55246 12962
rect 55298 12910 55300 12962
rect 54684 12562 54740 12572
rect 55132 12628 55188 12638
rect 54460 12516 54516 12526
rect 54460 12178 54516 12460
rect 55020 12516 55076 12526
rect 55020 12402 55076 12460
rect 55020 12350 55022 12402
rect 55074 12350 55076 12402
rect 55020 12338 55076 12350
rect 54460 12126 54462 12178
rect 54514 12126 54516 12178
rect 54460 12114 54516 12126
rect 54572 12180 54628 12190
rect 54572 12086 54628 12124
rect 55132 9604 55188 12572
rect 55244 11732 55300 12910
rect 58156 12852 58212 13022
rect 58156 12786 58212 12796
rect 55692 12290 55748 12302
rect 55692 12238 55694 12290
rect 55746 12238 55748 12290
rect 55356 12180 55412 12190
rect 55356 12086 55412 12124
rect 55244 11676 55524 11732
rect 55244 11508 55300 11518
rect 55244 11414 55300 11452
rect 55468 11396 55524 11676
rect 55692 11508 55748 12238
rect 55692 11442 55748 11452
rect 57372 11508 57428 11518
rect 57372 11414 57428 11452
rect 55132 9538 55188 9548
rect 55244 10276 55300 10286
rect 54572 9044 54628 9054
rect 54572 8950 54628 8988
rect 55244 9042 55300 10220
rect 55468 9938 55524 11340
rect 55468 9886 55470 9938
rect 55522 9886 55524 9938
rect 55468 9874 55524 9886
rect 58044 11396 58100 11406
rect 57596 9492 57652 9502
rect 57596 9266 57652 9436
rect 57596 9214 57598 9266
rect 57650 9214 57652 9266
rect 57596 9202 57652 9214
rect 57820 9268 57876 9278
rect 57820 9174 57876 9212
rect 55468 9156 55524 9166
rect 55468 9044 55524 9100
rect 56924 9156 56980 9166
rect 56924 9154 57092 9156
rect 56924 9102 56926 9154
rect 56978 9102 57092 9154
rect 56924 9100 57092 9102
rect 56924 9090 56980 9100
rect 55244 8990 55246 9042
rect 55298 8990 55300 9042
rect 55244 8978 55300 8990
rect 55356 9042 55524 9044
rect 55356 8990 55470 9042
rect 55522 8990 55524 9042
rect 55356 8988 55524 8990
rect 54460 8820 54516 8830
rect 54460 8726 54516 8764
rect 54908 8818 54964 8830
rect 54908 8766 54910 8818
rect 54962 8766 54964 8818
rect 54348 8530 54404 8540
rect 54124 8092 54236 8148
rect 54012 7588 54068 7598
rect 53900 7586 54068 7588
rect 53900 7534 54014 7586
rect 54066 7534 54068 7586
rect 53900 7532 54068 7534
rect 53340 7522 53396 7532
rect 53116 6916 53172 6926
rect 53116 6804 53172 6860
rect 53340 6916 53396 6926
rect 53340 6822 53396 6860
rect 53228 6804 53284 6814
rect 53116 6802 53284 6804
rect 53116 6750 53230 6802
rect 53282 6750 53284 6802
rect 53116 6748 53284 6750
rect 52892 6738 52948 6748
rect 53228 6738 53284 6748
rect 52892 6580 52948 6590
rect 53452 6580 53508 7532
rect 53788 7522 53844 7532
rect 54012 7522 54068 7532
rect 54124 7140 54180 8092
rect 54236 8082 54292 8092
rect 54348 8372 54404 8382
rect 54348 7588 54404 8316
rect 54908 8372 54964 8766
rect 54908 8306 54964 8316
rect 55244 8372 55300 8382
rect 55356 8372 55412 8988
rect 55468 8978 55524 8988
rect 56588 9044 56644 9054
rect 56588 8950 56644 8988
rect 57036 8428 57092 9100
rect 57036 8372 57428 8428
rect 55244 8370 55412 8372
rect 55244 8318 55246 8370
rect 55298 8318 55412 8370
rect 55244 8316 55412 8318
rect 57372 8370 57428 8372
rect 57372 8318 57374 8370
rect 57426 8318 57428 8370
rect 55244 8306 55300 8316
rect 57372 8306 57428 8318
rect 58044 8258 58100 11340
rect 58156 9492 58212 9502
rect 58156 9266 58212 9436
rect 58156 9214 58158 9266
rect 58210 9214 58212 9266
rect 58156 9202 58212 9214
rect 58044 8206 58046 8258
rect 58098 8206 58100 8258
rect 54460 8148 54516 8158
rect 54908 8148 54964 8158
rect 54460 8146 54852 8148
rect 54460 8094 54462 8146
rect 54514 8094 54852 8146
rect 54460 8092 54852 8094
rect 54460 8082 54516 8092
rect 54796 7700 54852 8092
rect 54908 8054 54964 8092
rect 54796 7644 55076 7700
rect 54348 7494 54404 7532
rect 55020 7474 55076 7644
rect 56924 7588 56980 7598
rect 56924 7586 57092 7588
rect 56924 7534 56926 7586
rect 56978 7534 57092 7586
rect 56924 7532 57092 7534
rect 56924 7522 56980 7532
rect 55020 7422 55022 7474
rect 55074 7422 55076 7474
rect 55020 7410 55076 7422
rect 55356 7476 55412 7486
rect 55356 7382 55412 7420
rect 56588 7476 56644 7486
rect 56588 7382 56644 7420
rect 53564 7028 53620 7038
rect 53620 6972 53844 7028
rect 53564 6962 53620 6972
rect 53788 6914 53844 6972
rect 53788 6862 53790 6914
rect 53842 6862 53844 6914
rect 53788 6850 53844 6862
rect 54124 6804 54180 7084
rect 54236 7362 54292 7374
rect 54236 7310 54238 7362
rect 54290 7310 54292 7362
rect 54236 6916 54292 7310
rect 54796 7362 54852 7374
rect 54796 7310 54798 7362
rect 54850 7310 54852 7362
rect 54796 7252 54852 7310
rect 54236 6850 54292 6860
rect 54572 7196 54796 7252
rect 53900 6748 54180 6804
rect 54572 6802 54628 7196
rect 54796 7186 54852 7196
rect 54572 6750 54574 6802
rect 54626 6750 54628 6802
rect 53564 6692 53620 6702
rect 53900 6692 53956 6748
rect 54572 6738 54628 6750
rect 55244 6804 55300 6814
rect 55244 6710 55300 6748
rect 53564 6690 53956 6692
rect 53564 6638 53566 6690
rect 53618 6638 53956 6690
rect 53564 6636 53956 6638
rect 56028 6692 56084 6702
rect 57036 6692 57092 7532
rect 57372 6692 57428 6702
rect 57036 6690 57428 6692
rect 57036 6638 57374 6690
rect 57426 6638 57428 6690
rect 57036 6636 57428 6638
rect 53564 6626 53620 6636
rect 52780 6578 52948 6580
rect 52780 6526 52894 6578
rect 52946 6526 52948 6578
rect 52780 6524 52948 6526
rect 52892 6514 52948 6524
rect 53116 6524 53508 6580
rect 53116 5794 53172 6524
rect 53116 5742 53118 5794
rect 53170 5742 53172 5794
rect 53116 5730 53172 5742
rect 53676 6466 53732 6478
rect 53676 6414 53678 6466
rect 53730 6414 53732 6466
rect 52220 5236 52276 5246
rect 52108 5234 52276 5236
rect 52108 5182 52222 5234
rect 52274 5182 52276 5234
rect 52108 5180 52276 5182
rect 52220 5124 52276 5180
rect 53452 5236 53508 5246
rect 52668 5124 52724 5134
rect 52220 5122 52724 5124
rect 52220 5070 52670 5122
rect 52722 5070 52724 5122
rect 52220 5068 52724 5070
rect 52668 5058 52724 5068
rect 51324 4900 51380 4910
rect 51324 4806 51380 4844
rect 52668 4900 52724 4910
rect 52668 4450 52724 4844
rect 52668 4398 52670 4450
rect 52722 4398 52724 4450
rect 52668 4386 52724 4398
rect 53452 4338 53508 5180
rect 53676 4452 53732 6414
rect 56028 5906 56084 6636
rect 57372 6626 57428 6636
rect 58044 6692 58100 8206
rect 58044 6598 58100 6636
rect 56028 5854 56030 5906
rect 56082 5854 56084 5906
rect 56028 5842 56084 5854
rect 55244 5796 55300 5806
rect 54124 5794 55300 5796
rect 54124 5742 55246 5794
rect 55298 5742 55300 5794
rect 54124 5740 55300 5742
rect 54124 4562 54180 5740
rect 55244 5730 55300 5740
rect 54684 5236 54740 5246
rect 54684 5142 54740 5180
rect 54124 4510 54126 4562
rect 54178 4510 54180 4562
rect 54124 4498 54180 4510
rect 53788 4452 53844 4462
rect 53676 4450 53844 4452
rect 53676 4398 53790 4450
rect 53842 4398 53844 4450
rect 53676 4396 53844 4398
rect 53788 4386 53844 4396
rect 57820 4452 57876 4462
rect 57820 4358 57876 4396
rect 53452 4286 53454 4338
rect 53506 4286 53508 4338
rect 53452 4274 53508 4286
rect 58156 4338 58212 4350
rect 58156 4286 58158 4338
rect 58210 4286 58212 4338
rect 50540 4226 51156 4228
rect 50540 4174 50542 4226
rect 50594 4174 51156 4226
rect 50540 4172 51156 4174
rect 57596 4228 57652 4238
rect 58156 4228 58212 4286
rect 57596 4226 58212 4228
rect 57596 4174 57598 4226
rect 57650 4174 58212 4226
rect 57596 4172 58212 4174
rect 50540 4162 50596 4172
rect 57596 4162 57652 4172
rect 58156 3668 58212 4172
rect 58156 3602 58212 3612
rect 48860 3490 48916 3500
rect 45052 800 45108 3388
rect 47852 3332 48132 3388
rect 48972 3444 49028 3482
rect 48972 3378 49028 3388
rect 47068 924 47348 980
rect 47068 800 47124 924
rect 37324 700 37716 756
rect 38976 0 39088 800
rect 40992 0 41104 800
rect 43008 0 43120 800
rect 45024 0 45136 800
rect 47040 0 47152 800
rect 47292 756 47348 924
rect 47852 756 47908 3332
rect 50316 3330 50372 3342
rect 51324 3332 51380 3342
rect 53340 3332 53396 3342
rect 55356 3332 55412 3342
rect 57372 3332 57428 3342
rect 50316 3278 50318 3330
rect 50370 3278 50372 3330
rect 49084 1762 49140 1774
rect 49084 1710 49086 1762
rect 49138 1710 49140 1762
rect 49084 800 49140 1710
rect 50316 1762 50372 3278
rect 51100 3330 51380 3332
rect 51100 3278 51326 3330
rect 51378 3278 51380 3330
rect 51100 3276 51380 3278
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 50316 1710 50318 1762
rect 50370 1710 50372 1762
rect 50316 1698 50372 1710
rect 51100 800 51156 3276
rect 51324 3266 51380 3276
rect 53116 3330 53396 3332
rect 53116 3278 53342 3330
rect 53394 3278 53396 3330
rect 53116 3276 53396 3278
rect 53116 800 53172 3276
rect 53340 3266 53396 3276
rect 55132 3330 55412 3332
rect 55132 3278 55358 3330
rect 55410 3278 55412 3330
rect 55132 3276 55412 3278
rect 55132 800 55188 3276
rect 55356 3266 55412 3276
rect 57148 3330 57428 3332
rect 57148 3278 57374 3330
rect 57426 3278 57428 3330
rect 57148 3276 57428 3278
rect 57148 800 57204 3276
rect 57372 3266 57428 3276
rect 47292 700 47908 756
rect 49056 0 49168 800
rect 51072 0 51184 800
rect 53088 0 53200 800
rect 55104 0 55216 800
rect 57120 0 57232 800
<< via2 >>
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 23100 55970 23156 55972
rect 23100 55918 23102 55970
rect 23102 55918 23154 55970
rect 23154 55918 23156 55970
rect 23100 55916 23156 55918
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 6860 48130 6916 48132
rect 6860 48078 6862 48130
rect 6862 48078 6914 48130
rect 6914 48078 6916 48130
rect 6860 48076 6916 48078
rect 6188 47570 6244 47572
rect 6188 47518 6190 47570
rect 6190 47518 6242 47570
rect 6242 47518 6244 47570
rect 6188 47516 6244 47518
rect 6972 47516 7028 47572
rect 6300 46562 6356 46564
rect 6300 46510 6302 46562
rect 6302 46510 6354 46562
rect 6354 46510 6356 46562
rect 6300 46508 6356 46510
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 7196 45948 7252 46004
rect 4172 45836 4228 45892
rect 6748 45890 6804 45892
rect 6748 45838 6750 45890
rect 6750 45838 6802 45890
rect 6802 45838 6804 45890
rect 6748 45836 6804 45838
rect 7420 45500 7476 45556
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4732 43820 4788 43876
rect 18284 55186 18340 55188
rect 18284 55134 18286 55186
rect 18286 55134 18338 55186
rect 18338 55134 18340 55186
rect 18284 55132 18340 55134
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 20300 54402 20356 54404
rect 20300 54350 20302 54402
rect 20302 54350 20354 54402
rect 20354 54350 20356 54402
rect 20300 54348 20356 54350
rect 18172 53676 18228 53732
rect 20188 53730 20244 53732
rect 20188 53678 20190 53730
rect 20190 53678 20242 53730
rect 20242 53678 20244 53730
rect 20188 53676 20244 53678
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 19068 52946 19124 52948
rect 19068 52894 19070 52946
rect 19070 52894 19122 52946
rect 19122 52894 19124 52946
rect 19068 52892 19124 52894
rect 17500 52780 17556 52836
rect 18060 52274 18116 52276
rect 18060 52222 18062 52274
rect 18062 52222 18114 52274
rect 18114 52222 18116 52274
rect 18060 52220 18116 52222
rect 15932 52050 15988 52052
rect 15932 51998 15934 52050
rect 15934 51998 15986 52050
rect 15986 51998 15988 52050
rect 15932 51996 15988 51998
rect 16156 51100 16212 51156
rect 14364 49756 14420 49812
rect 7644 46562 7700 46564
rect 7644 46510 7646 46562
rect 7646 46510 7698 46562
rect 7698 46510 7700 46562
rect 7644 46508 7700 46510
rect 8092 48802 8148 48804
rect 8092 48750 8094 48802
rect 8094 48750 8146 48802
rect 8146 48750 8148 48802
rect 8092 48748 8148 48750
rect 10444 48748 10500 48804
rect 8316 48300 8372 48356
rect 9548 48354 9604 48356
rect 9548 48302 9550 48354
rect 9550 48302 9602 48354
rect 9602 48302 9604 48354
rect 9548 48300 9604 48302
rect 9660 48130 9716 48132
rect 9660 48078 9662 48130
rect 9662 48078 9714 48130
rect 9714 48078 9716 48130
rect 9660 48076 9716 48078
rect 7980 45948 8036 46004
rect 7756 45500 7812 45556
rect 8204 45052 8260 45108
rect 7644 44434 7700 44436
rect 7644 44382 7646 44434
rect 7646 44382 7698 44434
rect 7698 44382 7700 44434
rect 7644 44380 7700 44382
rect 7868 44322 7924 44324
rect 7868 44270 7870 44322
rect 7870 44270 7922 44322
rect 7922 44270 7924 44322
rect 7868 44268 7924 44270
rect 10444 47180 10500 47236
rect 9548 45836 9604 45892
rect 8540 45164 8596 45220
rect 9660 45218 9716 45220
rect 9660 45166 9662 45218
rect 9662 45166 9714 45218
rect 9714 45166 9716 45218
rect 9660 45164 9716 45166
rect 9884 45106 9940 45108
rect 9884 45054 9886 45106
rect 9886 45054 9938 45106
rect 9938 45054 9940 45106
rect 9884 45052 9940 45054
rect 8316 44268 8372 44324
rect 8540 44380 8596 44436
rect 9100 44044 9156 44100
rect 8428 43932 8484 43988
rect 8204 43820 8260 43876
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 4956 40572 5012 40628
rect 1820 40460 1876 40516
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 2492 38892 2548 38948
rect 5292 39004 5348 39060
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 2492 38108 2548 38164
rect 7308 39340 7364 39396
rect 5180 38444 5236 38500
rect 5740 38780 5796 38836
rect 6300 38834 6356 38836
rect 6300 38782 6302 38834
rect 6302 38782 6354 38834
rect 6354 38782 6356 38834
rect 6300 38780 6356 38782
rect 6748 38834 6804 38836
rect 6748 38782 6750 38834
rect 6750 38782 6802 38834
rect 6802 38782 6804 38834
rect 6748 38780 6804 38782
rect 6188 38444 6244 38500
rect 5852 38162 5908 38164
rect 5852 38110 5854 38162
rect 5854 38110 5906 38162
rect 5906 38110 5908 38162
rect 5852 38108 5908 38110
rect 5628 37996 5684 38052
rect 5180 37772 5236 37828
rect 2492 36370 2548 36372
rect 2492 36318 2494 36370
rect 2494 36318 2546 36370
rect 2546 36318 2548 36370
rect 2492 36316 2548 36318
rect 4172 35756 4228 35812
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4508 36316 4564 36372
rect 4732 36204 4788 36260
rect 7196 38834 7252 38836
rect 7196 38782 7198 38834
rect 7198 38782 7250 38834
rect 7250 38782 7252 38834
rect 7196 38780 7252 38782
rect 6860 38050 6916 38052
rect 6860 37998 6862 38050
rect 6862 37998 6914 38050
rect 6914 37998 6916 38050
rect 6860 37996 6916 37998
rect 6748 37826 6804 37828
rect 6748 37774 6750 37826
rect 6750 37774 6802 37826
rect 6802 37774 6804 37826
rect 6748 37772 6804 37774
rect 5516 36258 5572 36260
rect 5516 36206 5518 36258
rect 5518 36206 5570 36258
rect 5570 36206 5572 36258
rect 5516 36204 5572 36206
rect 5068 35756 5124 35812
rect 4844 35644 4900 35700
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4844 35084 4900 35140
rect 2492 34636 2548 34692
rect 1820 33346 1876 33348
rect 1820 33294 1822 33346
rect 1822 33294 1874 33346
rect 1874 33294 1876 33346
rect 1820 33292 1876 33294
rect 2492 32450 2548 32452
rect 2492 32398 2494 32450
rect 2494 32398 2546 32450
rect 2546 32398 2548 32450
rect 2492 32396 2548 32398
rect 4620 34802 4676 34804
rect 4620 34750 4622 34802
rect 4622 34750 4674 34802
rect 4674 34750 4676 34802
rect 4620 34748 4676 34750
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 5068 35308 5124 35364
rect 5516 35698 5572 35700
rect 5516 35646 5518 35698
rect 5518 35646 5570 35698
rect 5570 35646 5572 35698
rect 5516 35644 5572 35646
rect 6076 35810 6132 35812
rect 6076 35758 6078 35810
rect 6078 35758 6130 35810
rect 6130 35758 6132 35810
rect 6076 35756 6132 35758
rect 6076 35196 6132 35252
rect 5964 35084 6020 35140
rect 4956 33292 5012 33348
rect 4620 32732 4676 32788
rect 4172 32508 4228 32564
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 5628 34802 5684 34804
rect 5628 34750 5630 34802
rect 5630 34750 5682 34802
rect 5682 34750 5684 34802
rect 5628 34748 5684 34750
rect 5740 34690 5796 34692
rect 5740 34638 5742 34690
rect 5742 34638 5794 34690
rect 5794 34638 5796 34690
rect 5740 34636 5796 34638
rect 6412 33516 6468 33572
rect 6860 33516 6916 33572
rect 5180 32732 5236 32788
rect 4956 32508 5012 32564
rect 5964 32786 6020 32788
rect 5964 32734 5966 32786
rect 5966 32734 6018 32786
rect 6018 32734 6020 32786
rect 5964 32732 6020 32734
rect 5068 32450 5124 32452
rect 5068 32398 5070 32450
rect 5070 32398 5122 32450
rect 5122 32398 5124 32450
rect 5068 32396 5124 32398
rect 6076 32562 6132 32564
rect 6076 32510 6078 32562
rect 6078 32510 6130 32562
rect 6130 32510 6132 32562
rect 6076 32508 6132 32510
rect 4060 31500 4116 31556
rect 2492 30828 2548 30884
rect 4508 31106 4564 31108
rect 4508 31054 4510 31106
rect 4510 31054 4562 31106
rect 4562 31054 4564 31106
rect 4508 31052 4564 31054
rect 4732 31500 4788 31556
rect 5628 31554 5684 31556
rect 5628 31502 5630 31554
rect 5630 31502 5682 31554
rect 5682 31502 5684 31554
rect 5628 31500 5684 31502
rect 5964 31218 6020 31220
rect 5964 31166 5966 31218
rect 5966 31166 6018 31218
rect 6018 31166 6020 31218
rect 5964 31164 6020 31166
rect 4956 30882 5012 30884
rect 4956 30830 4958 30882
rect 4958 30830 5010 30882
rect 5010 30830 5012 30882
rect 4956 30828 5012 30830
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 6188 31052 6244 31108
rect 4956 29932 5012 29988
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 3836 27804 3892 27860
rect 2492 27746 2548 27748
rect 2492 27694 2494 27746
rect 2494 27694 2546 27746
rect 2546 27694 2548 27746
rect 2492 27692 2548 27694
rect 3948 27692 4004 27748
rect 4508 27580 4564 27636
rect 4844 27858 4900 27860
rect 4844 27806 4846 27858
rect 4846 27806 4898 27858
rect 4898 27806 4900 27858
rect 4844 27804 4900 27806
rect 5740 29986 5796 29988
rect 5740 29934 5742 29986
rect 5742 29934 5794 29986
rect 5794 29934 5796 29986
rect 5740 29932 5796 29934
rect 6524 29820 6580 29876
rect 5852 29650 5908 29652
rect 5852 29598 5854 29650
rect 5854 29598 5906 29650
rect 5906 29598 5908 29650
rect 5852 29596 5908 29598
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4396 26962 4452 26964
rect 4396 26910 4398 26962
rect 4398 26910 4450 26962
rect 4450 26910 4452 26962
rect 4396 26908 4452 26910
rect 4956 27580 5012 27636
rect 4956 27074 5012 27076
rect 4956 27022 4958 27074
rect 4958 27022 5010 27074
rect 5010 27022 5012 27074
rect 4956 27020 5012 27022
rect 3276 26514 3332 26516
rect 3276 26462 3278 26514
rect 3278 26462 3330 26514
rect 3330 26462 3332 26514
rect 3276 26460 3332 26462
rect 3164 26402 3220 26404
rect 3164 26350 3166 26402
rect 3166 26350 3218 26402
rect 3218 26350 3220 26402
rect 3164 26348 3220 26350
rect 4732 26460 4788 26516
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4284 25506 4340 25508
rect 4284 25454 4286 25506
rect 4286 25454 4338 25506
rect 4338 25454 4340 25506
rect 4284 25452 4340 25454
rect 2492 25228 2548 25284
rect 3836 25282 3892 25284
rect 3836 25230 3838 25282
rect 3838 25230 3890 25282
rect 3890 25230 3892 25282
rect 3836 25228 3892 25230
rect 1820 24722 1876 24724
rect 1820 24670 1822 24722
rect 1822 24670 1874 24722
rect 1874 24670 1876 24722
rect 1820 24668 1876 24670
rect 6972 33346 7028 33348
rect 6972 33294 6974 33346
rect 6974 33294 7026 33346
rect 7026 33294 7028 33346
rect 6972 33292 7028 33294
rect 6860 28642 6916 28644
rect 6860 28590 6862 28642
rect 6862 28590 6914 28642
rect 6914 28590 6916 28642
rect 6860 28588 6916 28590
rect 7308 31778 7364 31780
rect 7308 31726 7310 31778
rect 7310 31726 7362 31778
rect 7362 31726 7364 31778
rect 7308 31724 7364 31726
rect 5628 27074 5684 27076
rect 5628 27022 5630 27074
rect 5630 27022 5682 27074
rect 5682 27022 5684 27074
rect 5628 27020 5684 27022
rect 6524 27020 6580 27076
rect 5180 26348 5236 26404
rect 4956 26290 5012 26292
rect 4956 26238 4958 26290
rect 4958 26238 5010 26290
rect 5010 26238 5012 26290
rect 4956 26236 5012 26238
rect 5180 25564 5236 25620
rect 5628 26796 5684 26852
rect 7644 43538 7700 43540
rect 7644 43486 7646 43538
rect 7646 43486 7698 43538
rect 7698 43486 7700 43538
rect 7644 43484 7700 43486
rect 9436 43932 9492 43988
rect 9548 44156 9604 44212
rect 9996 44098 10052 44100
rect 9996 44046 9998 44098
rect 9998 44046 10050 44098
rect 10050 44046 10052 44098
rect 9996 44044 10052 44046
rect 10220 43932 10276 43988
rect 10108 43820 10164 43876
rect 10332 43484 10388 43540
rect 10332 41916 10388 41972
rect 11340 47404 11396 47460
rect 15372 49756 15428 49812
rect 19068 50652 19124 50708
rect 18396 50316 18452 50372
rect 19404 52220 19460 52276
rect 19964 52220 20020 52276
rect 25788 55410 25844 55412
rect 25788 55358 25790 55410
rect 25790 55358 25842 55410
rect 25842 55358 25844 55410
rect 25788 55356 25844 55358
rect 21308 54348 21364 54404
rect 20972 54012 21028 54068
rect 20412 53676 20468 53732
rect 21420 53564 21476 53620
rect 21644 53788 21700 53844
rect 21868 54012 21924 54068
rect 22988 55298 23044 55300
rect 22988 55246 22990 55298
rect 22990 55246 23042 55298
rect 23042 55246 23044 55298
rect 22988 55244 23044 55246
rect 25452 55244 25508 55300
rect 22764 55132 22820 55188
rect 26124 55132 26180 55188
rect 23100 54460 23156 54516
rect 21980 53788 22036 53844
rect 22540 54012 22596 54068
rect 21868 53730 21924 53732
rect 21868 53678 21870 53730
rect 21870 53678 21922 53730
rect 21922 53678 21924 53730
rect 21868 53676 21924 53678
rect 22092 53730 22148 53732
rect 22092 53678 22094 53730
rect 22094 53678 22146 53730
rect 22146 53678 22148 53730
rect 22092 53676 22148 53678
rect 20300 51996 20356 52052
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 20412 51324 20468 51380
rect 19628 51212 19684 51268
rect 21084 51378 21140 51380
rect 21084 51326 21086 51378
rect 21086 51326 21138 51378
rect 21138 51326 21140 51378
rect 21084 51324 21140 51326
rect 20636 51212 20692 51268
rect 20188 50428 20244 50484
rect 21196 51154 21252 51156
rect 21196 51102 21198 51154
rect 21198 51102 21250 51154
rect 21250 51102 21252 51154
rect 21196 51100 21252 51102
rect 21308 50706 21364 50708
rect 21308 50654 21310 50706
rect 21310 50654 21362 50706
rect 21362 50654 21364 50706
rect 21308 50652 21364 50654
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 21980 50428 22036 50484
rect 21532 50370 21588 50372
rect 21532 50318 21534 50370
rect 21534 50318 21586 50370
rect 21586 50318 21588 50370
rect 21532 50316 21588 50318
rect 18956 49084 19012 49140
rect 14700 48130 14756 48132
rect 14700 48078 14702 48130
rect 14702 48078 14754 48130
rect 14754 48078 14756 48130
rect 14700 48076 14756 48078
rect 15932 48076 15988 48132
rect 16044 47628 16100 47684
rect 13468 47292 13524 47348
rect 14588 47404 14644 47460
rect 11004 47180 11060 47236
rect 10556 44994 10612 44996
rect 10556 44942 10558 44994
rect 10558 44942 10610 44994
rect 10610 44942 10612 44994
rect 10556 44940 10612 44942
rect 11676 45778 11732 45780
rect 11676 45726 11678 45778
rect 11678 45726 11730 45778
rect 11730 45726 11732 45778
rect 11676 45724 11732 45726
rect 11340 45500 11396 45556
rect 11228 45106 11284 45108
rect 11228 45054 11230 45106
rect 11230 45054 11282 45106
rect 11282 45054 11284 45106
rect 11228 45052 11284 45054
rect 12572 45778 12628 45780
rect 12572 45726 12574 45778
rect 12574 45726 12626 45778
rect 12626 45726 12628 45778
rect 12572 45724 12628 45726
rect 12684 45666 12740 45668
rect 12684 45614 12686 45666
rect 12686 45614 12738 45666
rect 12738 45614 12740 45666
rect 12684 45612 12740 45614
rect 12460 45276 12516 45332
rect 15260 47346 15316 47348
rect 15260 47294 15262 47346
rect 15262 47294 15314 47346
rect 15314 47294 15316 47346
rect 15260 47292 15316 47294
rect 15820 47346 15876 47348
rect 15820 47294 15822 47346
rect 15822 47294 15874 47346
rect 15874 47294 15876 47346
rect 15820 47292 15876 47294
rect 16268 47180 16324 47236
rect 17612 47682 17668 47684
rect 17612 47630 17614 47682
rect 17614 47630 17666 47682
rect 17666 47630 17668 47682
rect 17612 47628 17668 47630
rect 17052 47458 17108 47460
rect 17052 47406 17054 47458
rect 17054 47406 17106 47458
rect 17106 47406 17108 47458
rect 17052 47404 17108 47406
rect 17500 47404 17556 47460
rect 16940 47234 16996 47236
rect 16940 47182 16942 47234
rect 16942 47182 16994 47234
rect 16994 47182 16996 47234
rect 16940 47180 16996 47182
rect 14252 45778 14308 45780
rect 14252 45726 14254 45778
rect 14254 45726 14306 45778
rect 14306 45726 14308 45778
rect 14252 45724 14308 45726
rect 13020 45276 13076 45332
rect 13244 45612 13300 45668
rect 13916 45500 13972 45556
rect 12236 45052 12292 45108
rect 13020 45106 13076 45108
rect 13020 45054 13022 45106
rect 13022 45054 13074 45106
rect 13074 45054 13076 45106
rect 13020 45052 13076 45054
rect 13356 45106 13412 45108
rect 13356 45054 13358 45106
rect 13358 45054 13410 45106
rect 13410 45054 13412 45106
rect 13356 45052 13412 45054
rect 12012 44940 12068 44996
rect 10668 44380 10724 44436
rect 11116 44044 11172 44100
rect 10444 43372 10500 43428
rect 10108 41692 10164 41748
rect 8316 40514 8372 40516
rect 8316 40462 8318 40514
rect 8318 40462 8370 40514
rect 8370 40462 8372 40514
rect 8316 40460 8372 40462
rect 8428 40460 8484 40516
rect 9660 40572 9716 40628
rect 10668 43932 10724 43988
rect 13580 43372 13636 43428
rect 17388 47180 17444 47236
rect 15036 46396 15092 46452
rect 14700 45666 14756 45668
rect 14700 45614 14702 45666
rect 14702 45614 14754 45666
rect 14754 45614 14756 45666
rect 14700 45612 14756 45614
rect 14364 45330 14420 45332
rect 14364 45278 14366 45330
rect 14366 45278 14418 45330
rect 14418 45278 14420 45330
rect 14364 45276 14420 45278
rect 14700 45276 14756 45332
rect 14588 45218 14644 45220
rect 14588 45166 14590 45218
rect 14590 45166 14642 45218
rect 14642 45166 14644 45218
rect 14588 45164 14644 45166
rect 14700 45106 14756 45108
rect 14700 45054 14702 45106
rect 14702 45054 14754 45106
rect 14754 45054 14756 45106
rect 14700 45052 14756 45054
rect 14252 44380 14308 44436
rect 14140 44268 14196 44324
rect 14364 42754 14420 42756
rect 14364 42702 14366 42754
rect 14366 42702 14418 42754
rect 14418 42702 14420 42754
rect 14364 42700 14420 42702
rect 12684 42476 12740 42532
rect 11340 41916 11396 41972
rect 11340 41692 11396 41748
rect 10444 40572 10500 40628
rect 8540 39116 8596 39172
rect 7532 38668 7588 38724
rect 8876 39004 8932 39060
rect 8204 38668 8260 38724
rect 7756 38556 7812 38612
rect 7644 36988 7700 37044
rect 7756 35810 7812 35812
rect 7756 35758 7758 35810
rect 7758 35758 7810 35810
rect 7810 35758 7812 35810
rect 7756 35756 7812 35758
rect 8092 35868 8148 35924
rect 9324 39394 9380 39396
rect 9324 39342 9326 39394
rect 9326 39342 9378 39394
rect 9378 39342 9380 39394
rect 9324 39340 9380 39342
rect 8876 38722 8932 38724
rect 8876 38670 8878 38722
rect 8878 38670 8930 38722
rect 8930 38670 8932 38722
rect 8876 38668 8932 38670
rect 8876 38050 8932 38052
rect 8876 37998 8878 38050
rect 8878 37998 8930 38050
rect 8930 37998 8932 38050
rect 8876 37996 8932 37998
rect 7532 35644 7588 35700
rect 7532 33516 7588 33572
rect 7868 31666 7924 31668
rect 7868 31614 7870 31666
rect 7870 31614 7922 31666
rect 7922 31614 7924 31666
rect 7868 31612 7924 31614
rect 7532 31164 7588 31220
rect 7420 29932 7476 29988
rect 7084 29820 7140 29876
rect 7756 29820 7812 29876
rect 7532 28588 7588 28644
rect 7868 28700 7924 28756
rect 7980 28530 8036 28532
rect 7980 28478 7982 28530
rect 7982 28478 8034 28530
rect 8034 28478 8036 28530
rect 7980 28476 8036 28478
rect 9660 37996 9716 38052
rect 8652 37042 8708 37044
rect 8652 36990 8654 37042
rect 8654 36990 8706 37042
rect 8706 36990 8708 37042
rect 8652 36988 8708 36990
rect 8876 35810 8932 35812
rect 8876 35758 8878 35810
rect 8878 35758 8930 35810
rect 8930 35758 8932 35810
rect 8876 35756 8932 35758
rect 8764 35698 8820 35700
rect 8764 35646 8766 35698
rect 8766 35646 8818 35698
rect 8818 35646 8820 35698
rect 8764 35644 8820 35646
rect 8204 34130 8260 34132
rect 8204 34078 8206 34130
rect 8206 34078 8258 34130
rect 8258 34078 8260 34130
rect 8204 34076 8260 34078
rect 8204 31778 8260 31780
rect 8204 31726 8206 31778
rect 8206 31726 8258 31778
rect 8258 31726 8260 31778
rect 8204 31724 8260 31726
rect 8204 31218 8260 31220
rect 8204 31166 8206 31218
rect 8206 31166 8258 31218
rect 8258 31166 8260 31218
rect 8204 31164 8260 31166
rect 9324 35644 9380 35700
rect 9660 34972 9716 35028
rect 12012 41970 12068 41972
rect 12012 41918 12014 41970
rect 12014 41918 12066 41970
rect 12066 41918 12068 41970
rect 12012 41916 12068 41918
rect 13916 42530 13972 42532
rect 13916 42478 13918 42530
rect 13918 42478 13970 42530
rect 13970 42478 13972 42530
rect 13916 42476 13972 42478
rect 14812 44098 14868 44100
rect 14812 44046 14814 44098
rect 14814 44046 14866 44098
rect 14866 44046 14868 44098
rect 14812 44044 14868 44046
rect 14700 43596 14756 43652
rect 14476 42028 14532 42084
rect 16156 46450 16212 46452
rect 16156 46398 16158 46450
rect 16158 46398 16210 46450
rect 16210 46398 16212 46450
rect 16156 46396 16212 46398
rect 15260 45724 15316 45780
rect 15484 45276 15540 45332
rect 15372 45106 15428 45108
rect 15372 45054 15374 45106
rect 15374 45054 15426 45106
rect 15426 45054 15428 45106
rect 15372 45052 15428 45054
rect 16604 45106 16660 45108
rect 16604 45054 16606 45106
rect 16606 45054 16658 45106
rect 16658 45054 16660 45106
rect 16604 45052 16660 45054
rect 16268 44322 16324 44324
rect 16268 44270 16270 44322
rect 16270 44270 16322 44322
rect 16322 44270 16324 44322
rect 16268 44268 16324 44270
rect 16044 44044 16100 44100
rect 15372 43650 15428 43652
rect 15372 43598 15374 43650
rect 15374 43598 15426 43650
rect 15426 43598 15428 43650
rect 15372 43596 15428 43598
rect 16380 43650 16436 43652
rect 16380 43598 16382 43650
rect 16382 43598 16434 43650
rect 16434 43598 16436 43650
rect 16380 43596 16436 43598
rect 15820 42700 15876 42756
rect 15820 42028 15876 42084
rect 15372 41970 15428 41972
rect 15372 41918 15374 41970
rect 15374 41918 15426 41970
rect 15426 41918 15428 41970
rect 15372 41916 15428 41918
rect 17948 47458 18004 47460
rect 17948 47406 17950 47458
rect 17950 47406 18002 47458
rect 18002 47406 18004 47458
rect 17948 47404 18004 47406
rect 17948 47180 18004 47236
rect 18620 47404 18676 47460
rect 18620 46732 18676 46788
rect 18732 46674 18788 46676
rect 18732 46622 18734 46674
rect 18734 46622 18786 46674
rect 18786 46622 18788 46674
rect 18732 46620 18788 46622
rect 18620 46060 18676 46116
rect 18284 44380 18340 44436
rect 16604 43708 16660 43764
rect 17948 43762 18004 43764
rect 17948 43710 17950 43762
rect 17950 43710 18002 43762
rect 18002 43710 18004 43762
rect 17948 43708 18004 43710
rect 17388 43596 17444 43652
rect 15260 40572 15316 40628
rect 14252 40348 14308 40404
rect 12796 40236 12852 40292
rect 11004 39116 11060 39172
rect 12572 38780 12628 38836
rect 11676 38722 11732 38724
rect 11676 38670 11678 38722
rect 11678 38670 11730 38722
rect 11730 38670 11732 38722
rect 11676 38668 11732 38670
rect 11676 37436 11732 37492
rect 12348 37436 12404 37492
rect 10556 36876 10612 36932
rect 9884 35698 9940 35700
rect 9884 35646 9886 35698
rect 9886 35646 9938 35698
rect 9938 35646 9940 35698
rect 9884 35644 9940 35646
rect 10556 35026 10612 35028
rect 10556 34974 10558 35026
rect 10558 34974 10610 35026
rect 10610 34974 10612 35026
rect 10556 34972 10612 34974
rect 9660 34130 9716 34132
rect 9660 34078 9662 34130
rect 9662 34078 9714 34130
rect 9714 34078 9716 34130
rect 9660 34076 9716 34078
rect 12124 36988 12180 37044
rect 11340 35196 11396 35252
rect 11788 35196 11844 35252
rect 11340 33516 11396 33572
rect 14812 39340 14868 39396
rect 13468 38780 13524 38836
rect 16380 41186 16436 41188
rect 16380 41134 16382 41186
rect 16382 41134 16434 41186
rect 16434 41134 16436 41186
rect 16380 41132 16436 41134
rect 16604 40572 16660 40628
rect 16156 40402 16212 40404
rect 16156 40350 16158 40402
rect 16158 40350 16210 40402
rect 16210 40350 16212 40402
rect 16156 40348 16212 40350
rect 16604 40402 16660 40404
rect 16604 40350 16606 40402
rect 16606 40350 16658 40402
rect 16658 40350 16660 40402
rect 16604 40348 16660 40350
rect 16492 40290 16548 40292
rect 16492 40238 16494 40290
rect 16494 40238 16546 40290
rect 16546 40238 16548 40290
rect 16492 40236 16548 40238
rect 17276 40236 17332 40292
rect 17164 39618 17220 39620
rect 17164 39566 17166 39618
rect 17166 39566 17218 39618
rect 17218 39566 17220 39618
rect 17164 39564 17220 39566
rect 16940 39506 16996 39508
rect 16940 39454 16942 39506
rect 16942 39454 16994 39506
rect 16994 39454 16996 39506
rect 16940 39452 16996 39454
rect 17052 39394 17108 39396
rect 17052 39342 17054 39394
rect 17054 39342 17106 39394
rect 17106 39342 17108 39394
rect 17052 39340 17108 39342
rect 17052 38556 17108 38612
rect 12572 37266 12628 37268
rect 12572 37214 12574 37266
rect 12574 37214 12626 37266
rect 12626 37214 12628 37266
rect 12572 37212 12628 37214
rect 13244 36204 13300 36260
rect 13356 35922 13412 35924
rect 13356 35870 13358 35922
rect 13358 35870 13410 35922
rect 13410 35870 13412 35922
rect 13356 35868 13412 35870
rect 12572 35196 12628 35252
rect 12684 35644 12740 35700
rect 14140 36316 14196 36372
rect 13804 36258 13860 36260
rect 13804 36206 13806 36258
rect 13806 36206 13858 36258
rect 13858 36206 13860 36258
rect 13804 36204 13860 36206
rect 14252 35922 14308 35924
rect 14252 35870 14254 35922
rect 14254 35870 14306 35922
rect 14306 35870 14308 35922
rect 14252 35868 14308 35870
rect 14924 35868 14980 35924
rect 13580 35698 13636 35700
rect 13580 35646 13582 35698
rect 13582 35646 13634 35698
rect 13634 35646 13636 35698
rect 13580 35644 13636 35646
rect 8652 31666 8708 31668
rect 8652 31614 8654 31666
rect 8654 31614 8706 31666
rect 8706 31614 8708 31666
rect 8652 31612 8708 31614
rect 8428 30268 8484 30324
rect 8092 28140 8148 28196
rect 7308 27020 7364 27076
rect 7196 26962 7252 26964
rect 7196 26910 7198 26962
rect 7198 26910 7250 26962
rect 7250 26910 7252 26962
rect 7196 26908 7252 26910
rect 5740 26460 5796 26516
rect 5628 25506 5684 25508
rect 5628 25454 5630 25506
rect 5630 25454 5682 25506
rect 5682 25454 5684 25506
rect 5628 25452 5684 25454
rect 6524 25506 6580 25508
rect 6524 25454 6526 25506
rect 6526 25454 6578 25506
rect 6578 25454 6580 25506
rect 6524 25452 6580 25454
rect 6636 25394 6692 25396
rect 6636 25342 6638 25394
rect 6638 25342 6690 25394
rect 6690 25342 6692 25394
rect 6636 25340 6692 25342
rect 5068 25116 5124 25172
rect 5068 24722 5124 24724
rect 5068 24670 5070 24722
rect 5070 24670 5122 24722
rect 5122 24670 5124 24722
rect 5068 24668 5124 24670
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 8540 30156 8596 30212
rect 11228 31612 11284 31668
rect 9548 31106 9604 31108
rect 9548 31054 9550 31106
rect 9550 31054 9602 31106
rect 9602 31054 9604 31106
rect 9548 31052 9604 31054
rect 8988 30044 9044 30100
rect 8540 29596 8596 29652
rect 9548 30156 9604 30212
rect 8652 29426 8708 29428
rect 8652 29374 8654 29426
rect 8654 29374 8706 29426
rect 8706 29374 8708 29426
rect 8652 29372 8708 29374
rect 8988 28588 9044 28644
rect 8764 28140 8820 28196
rect 8652 27858 8708 27860
rect 8652 27806 8654 27858
rect 8654 27806 8706 27858
rect 8706 27806 8708 27858
rect 8652 27804 8708 27806
rect 7980 26962 8036 26964
rect 7980 26910 7982 26962
rect 7982 26910 8034 26962
rect 8034 26910 8036 26962
rect 7980 26908 8036 26910
rect 7420 25394 7476 25396
rect 7420 25342 7422 25394
rect 7422 25342 7474 25394
rect 7474 25342 7476 25394
rect 7420 25340 7476 25342
rect 7868 25340 7924 25396
rect 8540 27580 8596 27636
rect 9772 28700 9828 28756
rect 9660 28642 9716 28644
rect 9660 28590 9662 28642
rect 9662 28590 9714 28642
rect 9714 28590 9716 28642
rect 9660 28588 9716 28590
rect 9660 27580 9716 27636
rect 10556 30268 10612 30324
rect 10668 30098 10724 30100
rect 10668 30046 10670 30098
rect 10670 30046 10722 30098
rect 10722 30046 10724 30098
rect 10668 30044 10724 30046
rect 10668 28588 10724 28644
rect 10892 28642 10948 28644
rect 10892 28590 10894 28642
rect 10894 28590 10946 28642
rect 10946 28590 10948 28642
rect 10892 28588 10948 28590
rect 10220 27580 10276 27636
rect 9100 27074 9156 27076
rect 9100 27022 9102 27074
rect 9102 27022 9154 27074
rect 9154 27022 9156 27074
rect 9100 27020 9156 27022
rect 8876 26236 8932 26292
rect 8428 25564 8484 25620
rect 8764 25618 8820 25620
rect 8764 25566 8766 25618
rect 8766 25566 8818 25618
rect 8818 25566 8820 25618
rect 8764 25564 8820 25566
rect 8316 25340 8372 25396
rect 7980 25116 8036 25172
rect 8652 24162 8708 24164
rect 8652 24110 8654 24162
rect 8654 24110 8706 24162
rect 8706 24110 8708 24162
rect 8652 24108 8708 24110
rect 4620 22876 4676 22932
rect 5628 22876 5684 22932
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 2492 22540 2548 22596
rect 4732 22594 4788 22596
rect 4732 22542 4734 22594
rect 4734 22542 4786 22594
rect 4786 22542 4788 22594
rect 4732 22540 4788 22542
rect 3388 22482 3444 22484
rect 3388 22430 3390 22482
rect 3390 22430 3442 22482
rect 3442 22430 3444 22482
rect 3388 22428 3444 22430
rect 3948 22482 4004 22484
rect 3948 22430 3950 22482
rect 3950 22430 4002 22482
rect 4002 22430 4004 22482
rect 3948 22428 4004 22430
rect 1820 21644 1876 21700
rect 4956 22428 5012 22484
rect 4844 22146 4900 22148
rect 4844 22094 4846 22146
rect 4846 22094 4898 22146
rect 4898 22094 4900 22146
rect 4844 22092 4900 22094
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 5964 22316 6020 22372
rect 5068 20636 5124 20692
rect 4508 20018 4564 20020
rect 4508 19966 4510 20018
rect 4510 19966 4562 20018
rect 4562 19966 4564 20018
rect 4508 19964 4564 19966
rect 3164 18338 3220 18340
rect 3164 18286 3166 18338
rect 3166 18286 3218 18338
rect 3218 18286 3220 18338
rect 3164 18284 3220 18286
rect 3612 18338 3668 18340
rect 3612 18286 3614 18338
rect 3614 18286 3666 18338
rect 3666 18286 3668 18338
rect 3612 18284 3668 18286
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4508 18338 4564 18340
rect 4508 18286 4510 18338
rect 4510 18286 4562 18338
rect 4562 18286 4564 18338
rect 4508 18284 4564 18286
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4172 13916 4228 13972
rect 4620 13970 4676 13972
rect 4620 13918 4622 13970
rect 4622 13918 4674 13970
rect 4674 13918 4676 13970
rect 4620 13916 4676 13918
rect 3276 13634 3332 13636
rect 3276 13582 3278 13634
rect 3278 13582 3330 13634
rect 3330 13582 3332 13634
rect 3276 13580 3332 13582
rect 3724 13634 3780 13636
rect 3724 13582 3726 13634
rect 3726 13582 3778 13634
rect 3778 13582 3780 13634
rect 3724 13580 3780 13582
rect 3052 13468 3108 13524
rect 3948 13468 4004 13524
rect 1820 12012 1876 12068
rect 2492 12684 2548 12740
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 3948 11228 4004 11284
rect 4396 12738 4452 12740
rect 4396 12686 4398 12738
rect 4398 12686 4450 12738
rect 4450 12686 4452 12738
rect 4396 12684 4452 12686
rect 6188 22146 6244 22148
rect 6188 22094 6190 22146
rect 6190 22094 6242 22146
rect 6242 22094 6244 22146
rect 6188 22092 6244 22094
rect 6412 21698 6468 21700
rect 6412 21646 6414 21698
rect 6414 21646 6466 21698
rect 6466 21646 6468 21698
rect 6412 21644 6468 21646
rect 6860 22092 6916 22148
rect 6636 20412 6692 20468
rect 6300 19964 6356 20020
rect 6636 18284 6692 18340
rect 7308 20690 7364 20692
rect 7308 20638 7310 20690
rect 7310 20638 7362 20690
rect 7362 20638 7364 20690
rect 7308 20636 7364 20638
rect 8988 25900 9044 25956
rect 6972 20412 7028 20468
rect 12348 33570 12404 33572
rect 12348 33518 12350 33570
rect 12350 33518 12402 33570
rect 12402 33518 12404 33570
rect 12348 33516 12404 33518
rect 14588 35644 14644 35700
rect 13916 35196 13972 35252
rect 16492 37212 16548 37268
rect 16044 36428 16100 36484
rect 15148 36316 15204 36372
rect 15148 35810 15204 35812
rect 15148 35758 15150 35810
rect 15150 35758 15202 35810
rect 15202 35758 15204 35810
rect 15148 35756 15204 35758
rect 14924 35308 14980 35364
rect 14700 33068 14756 33124
rect 11564 30268 11620 30324
rect 11676 30044 11732 30100
rect 11340 28418 11396 28420
rect 11340 28366 11342 28418
rect 11342 28366 11394 28418
rect 11394 28366 11396 28418
rect 11340 28364 11396 28366
rect 10668 27580 10724 27636
rect 10892 27804 10948 27860
rect 10556 27020 10612 27076
rect 9772 26290 9828 26292
rect 9772 26238 9774 26290
rect 9774 26238 9826 26290
rect 9826 26238 9828 26290
rect 9772 26236 9828 26238
rect 12124 31666 12180 31668
rect 12124 31614 12126 31666
rect 12126 31614 12178 31666
rect 12178 31614 12180 31666
rect 12124 31612 12180 31614
rect 12124 28754 12180 28756
rect 12124 28702 12126 28754
rect 12126 28702 12178 28754
rect 12178 28702 12180 28754
rect 12124 28700 12180 28702
rect 12012 28642 12068 28644
rect 12012 28590 12014 28642
rect 12014 28590 12066 28642
rect 12066 28590 12068 28642
rect 12012 28588 12068 28590
rect 11228 27804 11284 27860
rect 11900 27804 11956 27860
rect 11116 27020 11172 27076
rect 13804 29596 13860 29652
rect 15372 35532 15428 35588
rect 15148 28924 15204 28980
rect 15484 35308 15540 35364
rect 13020 28364 13076 28420
rect 10892 25900 10948 25956
rect 10108 24668 10164 24724
rect 9660 23714 9716 23716
rect 9660 23662 9662 23714
rect 9662 23662 9714 23714
rect 9714 23662 9716 23714
rect 9660 23660 9716 23662
rect 8652 20300 8708 20356
rect 7420 18450 7476 18452
rect 7420 18398 7422 18450
rect 7422 18398 7474 18450
rect 7474 18398 7476 18450
rect 7420 18396 7476 18398
rect 7756 18338 7812 18340
rect 7756 18286 7758 18338
rect 7758 18286 7810 18338
rect 7810 18286 7812 18338
rect 7756 18284 7812 18286
rect 6860 18172 6916 18228
rect 7980 18226 8036 18228
rect 7980 18174 7982 18226
rect 7982 18174 8034 18226
rect 8034 18174 8036 18226
rect 7980 18172 8036 18174
rect 6412 17500 6468 17556
rect 6748 17500 6804 17556
rect 7420 17554 7476 17556
rect 7420 17502 7422 17554
rect 7422 17502 7474 17554
rect 7474 17502 7476 17554
rect 7420 17500 7476 17502
rect 5516 15820 5572 15876
rect 6972 15874 7028 15876
rect 6972 15822 6974 15874
rect 6974 15822 7026 15874
rect 7026 15822 7028 15874
rect 6972 15820 7028 15822
rect 6748 15372 6804 15428
rect 7420 15372 7476 15428
rect 7980 16098 8036 16100
rect 7980 16046 7982 16098
rect 7982 16046 8034 16098
rect 8034 16046 8036 16098
rect 7980 16044 8036 16046
rect 8540 16044 8596 16100
rect 7980 15372 8036 15428
rect 8204 15202 8260 15204
rect 8204 15150 8206 15202
rect 8206 15150 8258 15202
rect 8258 15150 8260 15202
rect 8204 15148 8260 15150
rect 8540 15708 8596 15764
rect 9884 23660 9940 23716
rect 10780 24722 10836 24724
rect 10780 24670 10782 24722
rect 10782 24670 10834 24722
rect 10834 24670 10836 24722
rect 10780 24668 10836 24670
rect 11452 24610 11508 24612
rect 11452 24558 11454 24610
rect 11454 24558 11506 24610
rect 11506 24558 11508 24610
rect 11452 24556 11508 24558
rect 10220 23714 10276 23716
rect 10220 23662 10222 23714
rect 10222 23662 10274 23714
rect 10274 23662 10276 23714
rect 10220 23660 10276 23662
rect 10780 21756 10836 21812
rect 8764 19794 8820 19796
rect 8764 19742 8766 19794
rect 8766 19742 8818 19794
rect 8818 19742 8820 19794
rect 8764 19740 8820 19742
rect 10332 19906 10388 19908
rect 10332 19854 10334 19906
rect 10334 19854 10386 19906
rect 10386 19854 10388 19906
rect 10332 19852 10388 19854
rect 9996 19740 10052 19796
rect 9660 18396 9716 18452
rect 9212 16492 9268 16548
rect 8876 16044 8932 16100
rect 10220 18450 10276 18452
rect 10220 18398 10222 18450
rect 10222 18398 10274 18450
rect 10274 18398 10276 18450
rect 10220 18396 10276 18398
rect 11004 18338 11060 18340
rect 11004 18286 11006 18338
rect 11006 18286 11058 18338
rect 11058 18286 11060 18338
rect 11004 18284 11060 18286
rect 10332 16044 10388 16100
rect 9548 15708 9604 15764
rect 5068 13916 5124 13972
rect 6636 13916 6692 13972
rect 4844 12236 4900 12292
rect 6300 12290 6356 12292
rect 6300 12238 6302 12290
rect 6302 12238 6354 12290
rect 6354 12238 6356 12290
rect 6300 12236 6356 12238
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4844 11452 4900 11508
rect 5740 11506 5796 11508
rect 5740 11454 5742 11506
rect 5742 11454 5794 11506
rect 5794 11454 5796 11506
rect 5740 11452 5796 11454
rect 4620 11340 4676 11396
rect 4172 10834 4228 10836
rect 4172 10782 4174 10834
rect 4174 10782 4226 10834
rect 4226 10782 4228 10834
rect 4172 10780 4228 10782
rect 5852 11394 5908 11396
rect 5852 11342 5854 11394
rect 5854 11342 5906 11394
rect 5906 11342 5908 11394
rect 5852 11340 5908 11342
rect 5628 11282 5684 11284
rect 5628 11230 5630 11282
rect 5630 11230 5682 11282
rect 5682 11230 5684 11282
rect 5628 11228 5684 11230
rect 5516 10834 5572 10836
rect 5516 10782 5518 10834
rect 5518 10782 5570 10834
rect 5570 10782 5572 10834
rect 5516 10780 5572 10782
rect 5628 10610 5684 10612
rect 5628 10558 5630 10610
rect 5630 10558 5682 10610
rect 5682 10558 5684 10610
rect 5628 10556 5684 10558
rect 5740 10444 5796 10500
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 5628 10220 5684 10276
rect 5964 10556 6020 10612
rect 2940 9212 2996 9268
rect 8204 12572 8260 12628
rect 7084 11452 7140 11508
rect 8316 12348 8372 12404
rect 8652 12124 8708 12180
rect 8428 11506 8484 11508
rect 8428 11454 8430 11506
rect 8430 11454 8482 11506
rect 8482 11454 8484 11506
rect 8428 11452 8484 11454
rect 10108 15484 10164 15540
rect 9996 15372 10052 15428
rect 9772 15202 9828 15204
rect 9772 15150 9774 15202
rect 9774 15150 9826 15202
rect 9826 15150 9828 15202
rect 9772 15148 9828 15150
rect 11676 16098 11732 16100
rect 11676 16046 11678 16098
rect 11678 16046 11730 16098
rect 11730 16046 11732 16098
rect 11676 16044 11732 16046
rect 11004 15484 11060 15540
rect 10556 15426 10612 15428
rect 10556 15374 10558 15426
rect 10558 15374 10610 15426
rect 10610 15374 10612 15426
rect 10556 15372 10612 15374
rect 11116 15148 11172 15204
rect 9436 12348 9492 12404
rect 9212 12124 9268 12180
rect 9772 12178 9828 12180
rect 9772 12126 9774 12178
rect 9774 12126 9826 12178
rect 9826 12126 9828 12178
rect 9772 12124 9828 12126
rect 8764 11116 8820 11172
rect 9324 11170 9380 11172
rect 9324 11118 9326 11170
rect 9326 11118 9378 11170
rect 9378 11118 9380 11170
rect 9324 11116 9380 11118
rect 6188 9714 6244 9716
rect 6188 9662 6190 9714
rect 6190 9662 6242 9714
rect 6242 9662 6244 9714
rect 6188 9660 6244 9662
rect 6860 9660 6916 9716
rect 6076 9266 6132 9268
rect 6076 9214 6078 9266
rect 6078 9214 6130 9266
rect 6130 9214 6132 9266
rect 6076 9212 6132 9214
rect 6300 9042 6356 9044
rect 6300 8990 6302 9042
rect 6302 8990 6354 9042
rect 6354 8990 6356 9042
rect 6300 8988 6356 8990
rect 7308 9100 7364 9156
rect 8764 9154 8820 9156
rect 8764 9102 8766 9154
rect 8766 9102 8818 9154
rect 8818 9102 8820 9154
rect 8764 9100 8820 9102
rect 6636 8988 6692 9044
rect 8428 9042 8484 9044
rect 8428 8990 8430 9042
rect 8430 8990 8482 9042
rect 8482 8990 8484 9042
rect 8428 8988 8484 8990
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 5964 7420 6020 7476
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 8652 8370 8708 8372
rect 8652 8318 8654 8370
rect 8654 8318 8706 8370
rect 8706 8318 8708 8370
rect 8652 8316 8708 8318
rect 7756 8092 7812 8148
rect 9772 9154 9828 9156
rect 9772 9102 9774 9154
rect 9774 9102 9826 9154
rect 9826 9102 9828 9154
rect 9772 9100 9828 9102
rect 9212 8988 9268 9044
rect 10220 12572 10276 12628
rect 9996 12124 10052 12180
rect 10332 11788 10388 11844
rect 10108 9660 10164 9716
rect 10220 9212 10276 9268
rect 8988 8146 9044 8148
rect 8988 8094 8990 8146
rect 8990 8094 9042 8146
rect 9042 8094 9044 8146
rect 8988 8092 9044 8094
rect 7756 7474 7812 7476
rect 7756 7422 7758 7474
rect 7758 7422 7810 7474
rect 7810 7422 7812 7474
rect 7756 7420 7812 7422
rect 7868 6018 7924 6020
rect 7868 5966 7870 6018
rect 7870 5966 7922 6018
rect 7922 5966 7924 6018
rect 7868 5964 7924 5966
rect 8876 6690 8932 6692
rect 8876 6638 8878 6690
rect 8878 6638 8930 6690
rect 8930 6638 8932 6690
rect 8876 6636 8932 6638
rect 8540 6018 8596 6020
rect 8540 5966 8542 6018
rect 8542 5966 8594 6018
rect 8594 5966 8596 6018
rect 8540 5964 8596 5966
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 10780 12012 10836 12068
rect 10668 9266 10724 9268
rect 10668 9214 10670 9266
rect 10670 9214 10722 9266
rect 10722 9214 10724 9266
rect 10668 9212 10724 9214
rect 14700 27746 14756 27748
rect 14700 27694 14702 27746
rect 14702 27694 14754 27746
rect 14754 27694 14756 27746
rect 14700 27692 14756 27694
rect 13916 24722 13972 24724
rect 13916 24670 13918 24722
rect 13918 24670 13970 24722
rect 13970 24670 13972 24722
rect 13916 24668 13972 24670
rect 15036 24668 15092 24724
rect 12348 24556 12404 24612
rect 14700 24610 14756 24612
rect 14700 24558 14702 24610
rect 14702 24558 14754 24610
rect 14754 24558 14756 24610
rect 14700 24556 14756 24558
rect 12684 23826 12740 23828
rect 12684 23774 12686 23826
rect 12686 23774 12738 23826
rect 12738 23774 12740 23826
rect 12684 23772 12740 23774
rect 14588 23938 14644 23940
rect 14588 23886 14590 23938
rect 14590 23886 14642 23938
rect 14642 23886 14644 23938
rect 14588 23884 14644 23886
rect 15036 23884 15092 23940
rect 14140 23826 14196 23828
rect 14140 23774 14142 23826
rect 14142 23774 14194 23826
rect 14194 23774 14196 23826
rect 14140 23772 14196 23774
rect 12348 22876 12404 22932
rect 13468 22930 13524 22932
rect 13468 22878 13470 22930
rect 13470 22878 13522 22930
rect 13522 22878 13524 22930
rect 13468 22876 13524 22878
rect 13804 22930 13860 22932
rect 13804 22878 13806 22930
rect 13806 22878 13858 22930
rect 13858 22878 13860 22930
rect 13804 22876 13860 22878
rect 14140 22876 14196 22932
rect 12348 22316 12404 22372
rect 12796 21810 12852 21812
rect 12796 21758 12798 21810
rect 12798 21758 12850 21810
rect 12850 21758 12852 21810
rect 12796 21756 12852 21758
rect 13468 21810 13524 21812
rect 13468 21758 13470 21810
rect 13470 21758 13522 21810
rect 13522 21758 13524 21810
rect 13468 21756 13524 21758
rect 14700 21756 14756 21812
rect 13244 21586 13300 21588
rect 13244 21534 13246 21586
rect 13246 21534 13298 21586
rect 13298 21534 13300 21586
rect 13244 21532 13300 21534
rect 12684 20748 12740 20804
rect 13132 20748 13188 20804
rect 12908 20524 12964 20580
rect 13468 20802 13524 20804
rect 13468 20750 13470 20802
rect 13470 20750 13522 20802
rect 13522 20750 13524 20802
rect 13468 20748 13524 20750
rect 13692 20578 13748 20580
rect 13692 20526 13694 20578
rect 13694 20526 13746 20578
rect 13746 20526 13748 20578
rect 13692 20524 13748 20526
rect 13580 20300 13636 20356
rect 13580 20076 13636 20132
rect 14476 21586 14532 21588
rect 14476 21534 14478 21586
rect 14478 21534 14530 21586
rect 14530 21534 14532 21586
rect 14476 21532 14532 21534
rect 14140 20748 14196 20804
rect 14028 20130 14084 20132
rect 14028 20078 14030 20130
rect 14030 20078 14082 20130
rect 14082 20078 14084 20130
rect 14028 20076 14084 20078
rect 13916 19906 13972 19908
rect 13916 19854 13918 19906
rect 13918 19854 13970 19906
rect 13970 19854 13972 19906
rect 13916 19852 13972 19854
rect 13580 19010 13636 19012
rect 13580 18958 13582 19010
rect 13582 18958 13634 19010
rect 13634 18958 13636 19010
rect 13580 18956 13636 18958
rect 13468 18450 13524 18452
rect 13468 18398 13470 18450
rect 13470 18398 13522 18450
rect 13522 18398 13524 18450
rect 13468 18396 13524 18398
rect 13692 18396 13748 18452
rect 14924 19346 14980 19348
rect 14924 19294 14926 19346
rect 14926 19294 14978 19346
rect 14978 19294 14980 19346
rect 14924 19292 14980 19294
rect 14028 18450 14084 18452
rect 14028 18398 14030 18450
rect 14030 18398 14082 18450
rect 14082 18398 14084 18450
rect 14028 18396 14084 18398
rect 14252 18956 14308 19012
rect 14700 18450 14756 18452
rect 14700 18398 14702 18450
rect 14702 18398 14754 18450
rect 14754 18398 14756 18450
rect 14700 18396 14756 18398
rect 14476 18338 14532 18340
rect 14476 18286 14478 18338
rect 14478 18286 14530 18338
rect 14530 18286 14532 18338
rect 14476 18284 14532 18286
rect 14140 18172 14196 18228
rect 15148 20412 15204 20468
rect 13804 16882 13860 16884
rect 13804 16830 13806 16882
rect 13806 16830 13858 16882
rect 13858 16830 13860 16882
rect 13804 16828 13860 16830
rect 15148 17052 15204 17108
rect 15260 16882 15316 16884
rect 15260 16830 15262 16882
rect 15262 16830 15314 16882
rect 15314 16830 15316 16882
rect 15260 16828 15316 16830
rect 14700 16210 14756 16212
rect 14700 16158 14702 16210
rect 14702 16158 14754 16210
rect 14754 16158 14756 16210
rect 14700 16156 14756 16158
rect 14812 16604 14868 16660
rect 14476 16044 14532 16100
rect 13356 15202 13412 15204
rect 13356 15150 13358 15202
rect 13358 15150 13410 15202
rect 13410 15150 13412 15202
rect 13356 15148 13412 15150
rect 13244 14476 13300 14532
rect 15372 16604 15428 16660
rect 15708 35196 15764 35252
rect 16268 35810 16324 35812
rect 16268 35758 16270 35810
rect 16270 35758 16322 35810
rect 16322 35758 16324 35810
rect 16268 35756 16324 35758
rect 16156 35698 16212 35700
rect 16156 35646 16158 35698
rect 16158 35646 16210 35698
rect 16210 35646 16212 35698
rect 16156 35644 16212 35646
rect 16380 35196 16436 35252
rect 16604 36482 16660 36484
rect 16604 36430 16606 36482
rect 16606 36430 16658 36482
rect 16658 36430 16660 36482
rect 16604 36428 16660 36430
rect 16716 35644 16772 35700
rect 16380 34076 16436 34132
rect 17500 41132 17556 41188
rect 17612 41244 17668 41300
rect 17500 40348 17556 40404
rect 19964 49138 20020 49140
rect 19964 49086 19966 49138
rect 19966 49086 20018 49138
rect 20018 49086 20020 49138
rect 19964 49084 20020 49086
rect 19740 48748 19796 48804
rect 20076 48802 20132 48804
rect 20076 48750 20078 48802
rect 20078 48750 20130 48802
rect 20130 48750 20132 48802
rect 20076 48748 20132 48750
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 22876 53730 22932 53732
rect 22876 53678 22878 53730
rect 22878 53678 22930 53730
rect 22930 53678 22932 53730
rect 22876 53676 22932 53678
rect 22988 53506 23044 53508
rect 22988 53454 22990 53506
rect 22990 53454 23042 53506
rect 23042 53454 23044 53506
rect 22988 53452 23044 53454
rect 22652 52834 22708 52836
rect 22652 52782 22654 52834
rect 22654 52782 22706 52834
rect 22706 52782 22708 52834
rect 22652 52780 22708 52782
rect 22988 52162 23044 52164
rect 22988 52110 22990 52162
rect 22990 52110 23042 52162
rect 23042 52110 23044 52162
rect 22988 52108 23044 52110
rect 23548 54514 23604 54516
rect 23548 54462 23550 54514
rect 23550 54462 23602 54514
rect 23602 54462 23604 54514
rect 23548 54460 23604 54462
rect 24780 54402 24836 54404
rect 24780 54350 24782 54402
rect 24782 54350 24834 54402
rect 24834 54350 24836 54402
rect 24780 54348 24836 54350
rect 23884 53676 23940 53732
rect 25228 53730 25284 53732
rect 25228 53678 25230 53730
rect 25230 53678 25282 53730
rect 25282 53678 25284 53730
rect 25228 53676 25284 53678
rect 24668 52946 24724 52948
rect 24668 52894 24670 52946
rect 24670 52894 24722 52946
rect 24722 52894 24724 52946
rect 24668 52892 24724 52894
rect 25452 53452 25508 53508
rect 23996 52162 24052 52164
rect 23996 52110 23998 52162
rect 23998 52110 24050 52162
rect 24050 52110 24052 52162
rect 23996 52108 24052 52110
rect 24556 52162 24612 52164
rect 24556 52110 24558 52162
rect 24558 52110 24610 52162
rect 24610 52110 24612 52162
rect 24556 52108 24612 52110
rect 22764 50652 22820 50708
rect 20748 48860 20804 48916
rect 21644 48914 21700 48916
rect 21644 48862 21646 48914
rect 21646 48862 21698 48914
rect 21698 48862 21700 48914
rect 21644 48860 21700 48862
rect 22092 48914 22148 48916
rect 22092 48862 22094 48914
rect 22094 48862 22146 48914
rect 22146 48862 22148 48914
rect 22092 48860 22148 48862
rect 21420 48748 21476 48804
rect 19964 47458 20020 47460
rect 19964 47406 19966 47458
rect 19966 47406 20018 47458
rect 20018 47406 20020 47458
rect 19964 47404 20020 47406
rect 20188 47180 20244 47236
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 21532 47404 21588 47460
rect 21196 47180 21252 47236
rect 21532 47068 21588 47124
rect 21644 48412 21700 48468
rect 19628 46620 19684 46676
rect 21420 46060 21476 46116
rect 19516 45724 19572 45780
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 22540 48412 22596 48468
rect 21756 47180 21812 47236
rect 21756 45836 21812 45892
rect 22988 51378 23044 51380
rect 22988 51326 22990 51378
rect 22990 51326 23042 51378
rect 23042 51326 23044 51378
rect 22988 51324 23044 51326
rect 23324 51266 23380 51268
rect 23324 51214 23326 51266
rect 23326 51214 23378 51266
rect 23378 51214 23380 51266
rect 23324 51212 23380 51214
rect 23772 51324 23828 51380
rect 23996 51212 24052 51268
rect 22876 48748 22932 48804
rect 23324 50316 23380 50372
rect 24556 49756 24612 49812
rect 25340 49644 25396 49700
rect 26684 55132 26740 55188
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 27132 55356 27188 55412
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 27356 55020 27412 55076
rect 27468 55186 27524 55188
rect 27468 55134 27470 55186
rect 27470 55134 27522 55186
rect 27522 55134 27524 55186
rect 27468 55132 27524 55134
rect 26908 54012 26964 54068
rect 26348 53564 26404 53620
rect 25788 52108 25844 52164
rect 25900 50428 25956 50484
rect 25676 49810 25732 49812
rect 25676 49758 25678 49810
rect 25678 49758 25730 49810
rect 25730 49758 25732 49810
rect 25676 49756 25732 49758
rect 25900 49308 25956 49364
rect 23100 47292 23156 47348
rect 22652 46844 22708 46900
rect 22876 47180 22932 47236
rect 19852 44882 19908 44884
rect 19852 44830 19854 44882
rect 19854 44830 19906 44882
rect 19906 44830 19908 44882
rect 19852 44828 19908 44830
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 18732 43596 18788 43652
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 18508 41132 18564 41188
rect 19852 41356 19908 41412
rect 18956 40626 19012 40628
rect 18956 40574 18958 40626
rect 18958 40574 19010 40626
rect 19010 40574 19012 40626
rect 18956 40572 19012 40574
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19628 40626 19684 40628
rect 19628 40574 19630 40626
rect 19630 40574 19682 40626
rect 19682 40574 19684 40626
rect 19628 40572 19684 40574
rect 18172 40236 18228 40292
rect 18620 40236 18676 40292
rect 17836 39618 17892 39620
rect 17836 39566 17838 39618
rect 17838 39566 17890 39618
rect 17890 39566 17892 39618
rect 17836 39564 17892 39566
rect 19068 40236 19124 40292
rect 18844 39452 18900 39508
rect 18508 38780 18564 38836
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 18060 38722 18116 38724
rect 18060 38670 18062 38722
rect 18062 38670 18114 38722
rect 18114 38670 18116 38722
rect 18060 38668 18116 38670
rect 17948 38610 18004 38612
rect 17948 38558 17950 38610
rect 17950 38558 18002 38610
rect 18002 38558 18004 38610
rect 17948 38556 18004 38558
rect 18844 38722 18900 38724
rect 18844 38670 18846 38722
rect 18846 38670 18898 38722
rect 18898 38670 18900 38722
rect 18844 38668 18900 38670
rect 19180 38780 19236 38836
rect 19068 38668 19124 38724
rect 19516 37266 19572 37268
rect 19516 37214 19518 37266
rect 19518 37214 19570 37266
rect 19570 37214 19572 37266
rect 19516 37212 19572 37214
rect 20076 38722 20132 38724
rect 20076 38670 20078 38722
rect 20078 38670 20130 38722
rect 20130 38670 20132 38722
rect 20076 38668 20132 38670
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 20412 44882 20468 44884
rect 20412 44830 20414 44882
rect 20414 44830 20466 44882
rect 20466 44830 20468 44882
rect 20412 44828 20468 44830
rect 21420 43372 21476 43428
rect 20748 42754 20804 42756
rect 20748 42702 20750 42754
rect 20750 42702 20802 42754
rect 20802 42702 20804 42754
rect 20748 42700 20804 42702
rect 21420 42700 21476 42756
rect 21196 42476 21252 42532
rect 20412 40124 20468 40180
rect 20860 40124 20916 40180
rect 21532 39788 21588 39844
rect 23212 47068 23268 47124
rect 23436 45724 23492 45780
rect 23436 45500 23492 45556
rect 22652 45052 22708 45108
rect 21980 42530 22036 42532
rect 21980 42478 21982 42530
rect 21982 42478 22034 42530
rect 22034 42478 22036 42530
rect 21980 42476 22036 42478
rect 22092 41916 22148 41972
rect 22316 39842 22372 39844
rect 22316 39790 22318 39842
rect 22318 39790 22370 39842
rect 22370 39790 22372 39842
rect 22316 39788 22372 39790
rect 22428 39730 22484 39732
rect 22428 39678 22430 39730
rect 22430 39678 22482 39730
rect 22482 39678 22484 39730
rect 22428 39676 22484 39678
rect 21980 39340 22036 39396
rect 21196 38108 21252 38164
rect 19740 37100 19796 37156
rect 22876 44268 22932 44324
rect 24108 47234 24164 47236
rect 24108 47182 24110 47234
rect 24110 47182 24162 47234
rect 24162 47182 24164 47234
rect 24108 47180 24164 47182
rect 24332 46674 24388 46676
rect 24332 46622 24334 46674
rect 24334 46622 24386 46674
rect 24386 46622 24388 46674
rect 24332 46620 24388 46622
rect 24108 45890 24164 45892
rect 24108 45838 24110 45890
rect 24110 45838 24162 45890
rect 24162 45838 24164 45890
rect 24108 45836 24164 45838
rect 23660 45164 23716 45220
rect 23772 45106 23828 45108
rect 23772 45054 23774 45106
rect 23774 45054 23826 45106
rect 23826 45054 23828 45106
rect 23772 45052 23828 45054
rect 23772 43596 23828 43652
rect 25228 46620 25284 46676
rect 25116 43260 25172 43316
rect 23324 41858 23380 41860
rect 23324 41806 23326 41858
rect 23326 41806 23378 41858
rect 23378 41806 23380 41858
rect 23324 41804 23380 41806
rect 23772 41804 23828 41860
rect 23996 41970 24052 41972
rect 23996 41918 23998 41970
rect 23998 41918 24050 41970
rect 24050 41918 24052 41970
rect 23996 41916 24052 41918
rect 23884 41692 23940 41748
rect 24220 41970 24276 41972
rect 24220 41918 24222 41970
rect 24222 41918 24274 41970
rect 24274 41918 24276 41970
rect 24220 41916 24276 41918
rect 24108 41356 24164 41412
rect 24444 41692 24500 41748
rect 24332 39676 24388 39732
rect 24444 40236 24500 40292
rect 23100 38892 23156 38948
rect 23884 39564 23940 39620
rect 23436 38668 23492 38724
rect 23660 38162 23716 38164
rect 23660 38110 23662 38162
rect 23662 38110 23714 38162
rect 23714 38110 23716 38162
rect 23660 38108 23716 38110
rect 20524 37212 20580 37268
rect 20188 37154 20244 37156
rect 20188 37102 20190 37154
rect 20190 37102 20242 37154
rect 20242 37102 20244 37154
rect 20188 37100 20244 37102
rect 20076 36204 20132 36260
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 17500 35756 17556 35812
rect 17388 34914 17444 34916
rect 17388 34862 17390 34914
rect 17390 34862 17442 34914
rect 17442 34862 17444 34914
rect 17388 34860 17444 34862
rect 19180 34914 19236 34916
rect 19180 34862 19182 34914
rect 19182 34862 19234 34914
rect 19234 34862 19236 34914
rect 19180 34860 19236 34862
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 16492 33964 16548 34020
rect 16044 33906 16100 33908
rect 16044 33854 16046 33906
rect 16046 33854 16098 33906
rect 16098 33854 16100 33906
rect 16044 33852 16100 33854
rect 16492 33122 16548 33124
rect 16492 33070 16494 33122
rect 16494 33070 16546 33122
rect 16546 33070 16548 33122
rect 16492 33068 16548 33070
rect 16380 32732 16436 32788
rect 19516 34130 19572 34132
rect 19516 34078 19518 34130
rect 19518 34078 19570 34130
rect 19570 34078 19572 34130
rect 19516 34076 19572 34078
rect 22540 37266 22596 37268
rect 22540 37214 22542 37266
rect 22542 37214 22594 37266
rect 22594 37214 22596 37266
rect 22540 37212 22596 37214
rect 20636 37100 20692 37156
rect 21196 36204 21252 36260
rect 20860 34860 20916 34916
rect 20524 34188 20580 34244
rect 20300 34130 20356 34132
rect 20300 34078 20302 34130
rect 20302 34078 20354 34130
rect 20354 34078 20356 34130
rect 20300 34076 20356 34078
rect 17388 34018 17444 34020
rect 17388 33966 17390 34018
rect 17390 33966 17442 34018
rect 17442 33966 17444 34018
rect 17388 33964 17444 33966
rect 19516 33852 19572 33908
rect 16492 31836 16548 31892
rect 17388 32786 17444 32788
rect 17388 32734 17390 32786
rect 17390 32734 17442 32786
rect 17442 32734 17444 32786
rect 17388 32732 17444 32734
rect 16828 31890 16884 31892
rect 16828 31838 16830 31890
rect 16830 31838 16882 31890
rect 16882 31838 16884 31890
rect 16828 31836 16884 31838
rect 16492 30828 16548 30884
rect 15932 30156 15988 30212
rect 16380 30210 16436 30212
rect 16380 30158 16382 30210
rect 16382 30158 16434 30210
rect 16434 30158 16436 30210
rect 16380 30156 16436 30158
rect 16268 29650 16324 29652
rect 16268 29598 16270 29650
rect 16270 29598 16322 29650
rect 16322 29598 16324 29650
rect 16268 29596 16324 29598
rect 16716 30210 16772 30212
rect 16716 30158 16718 30210
rect 16718 30158 16770 30210
rect 16770 30158 16772 30210
rect 16716 30156 16772 30158
rect 16380 28476 16436 28532
rect 16716 28530 16772 28532
rect 16716 28478 16718 28530
rect 16718 28478 16770 28530
rect 16770 28478 16772 28530
rect 16716 28476 16772 28478
rect 16268 27692 16324 27748
rect 16940 30044 16996 30100
rect 17164 31164 17220 31220
rect 17836 31218 17892 31220
rect 17836 31166 17838 31218
rect 17838 31166 17890 31218
rect 17890 31166 17892 31218
rect 17836 31164 17892 31166
rect 17500 30882 17556 30884
rect 17500 30830 17502 30882
rect 17502 30830 17554 30882
rect 17554 30830 17556 30882
rect 17500 30828 17556 30830
rect 17612 30156 17668 30212
rect 18956 32172 19012 32228
rect 17948 30044 18004 30100
rect 18508 29820 18564 29876
rect 18396 28754 18452 28756
rect 18396 28702 18398 28754
rect 18398 28702 18450 28754
rect 18450 28702 18452 28754
rect 18396 28700 18452 28702
rect 15932 24556 15988 24612
rect 15820 20412 15876 20468
rect 16716 23100 16772 23156
rect 16156 21980 16212 22036
rect 17724 27692 17780 27748
rect 18060 25228 18116 25284
rect 17836 24556 17892 24612
rect 17164 23100 17220 23156
rect 17612 22540 17668 22596
rect 16716 21980 16772 22036
rect 17724 22316 17780 22372
rect 16604 21532 16660 21588
rect 17388 21586 17444 21588
rect 17388 21534 17390 21586
rect 17390 21534 17442 21586
rect 17442 21534 17444 21586
rect 17388 21532 17444 21534
rect 17948 23154 18004 23156
rect 17948 23102 17950 23154
rect 17950 23102 18002 23154
rect 18002 23102 18004 23154
rect 17948 23100 18004 23102
rect 17948 22540 18004 22596
rect 17948 20972 18004 21028
rect 17612 20130 17668 20132
rect 17612 20078 17614 20130
rect 17614 20078 17666 20130
rect 17666 20078 17668 20130
rect 17612 20076 17668 20078
rect 16604 19740 16660 19796
rect 16492 19292 16548 19348
rect 16492 18674 16548 18676
rect 16492 18622 16494 18674
rect 16494 18622 16546 18674
rect 16546 18622 16548 18674
rect 16492 18620 16548 18622
rect 17388 19794 17444 19796
rect 17388 19742 17390 19794
rect 17390 19742 17442 19794
rect 17442 19742 17444 19794
rect 17388 19740 17444 19742
rect 17388 18620 17444 18676
rect 16716 18396 16772 18452
rect 17612 18450 17668 18452
rect 17612 18398 17614 18450
rect 17614 18398 17666 18450
rect 17666 18398 17668 18450
rect 17612 18396 17668 18398
rect 16044 18172 16100 18228
rect 18172 18956 18228 19012
rect 18284 20972 18340 21028
rect 19292 30098 19348 30100
rect 19292 30046 19294 30098
rect 19294 30046 19346 30098
rect 19346 30046 19348 30098
rect 19292 30044 19348 30046
rect 19068 29820 19124 29876
rect 19404 29650 19460 29652
rect 19404 29598 19406 29650
rect 19406 29598 19458 29650
rect 19458 29598 19460 29650
rect 19404 29596 19460 29598
rect 18732 28476 18788 28532
rect 19292 27692 19348 27748
rect 19180 25282 19236 25284
rect 19180 25230 19182 25282
rect 19182 25230 19234 25282
rect 19234 25230 19236 25282
rect 19180 25228 19236 25230
rect 18620 24610 18676 24612
rect 18620 24558 18622 24610
rect 18622 24558 18674 24610
rect 18674 24558 18676 24610
rect 18620 24556 18676 24558
rect 19292 24556 19348 24612
rect 20300 33234 20356 33236
rect 20300 33182 20302 33234
rect 20302 33182 20354 33234
rect 20354 33182 20356 33234
rect 20300 33180 20356 33182
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 20412 31666 20468 31668
rect 20412 31614 20414 31666
rect 20414 31614 20466 31666
rect 20466 31614 20468 31666
rect 20412 31612 20468 31614
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20412 29820 20468 29876
rect 20044 29764 20100 29766
rect 19852 29650 19908 29652
rect 19852 29598 19854 29650
rect 19854 29598 19906 29650
rect 19906 29598 19908 29650
rect 19852 29596 19908 29598
rect 20860 33458 20916 33460
rect 20860 33406 20862 33458
rect 20862 33406 20914 33458
rect 20914 33406 20916 33458
rect 20860 33404 20916 33406
rect 20524 29596 20580 29652
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 20972 28028 21028 28084
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 20076 26402 20132 26404
rect 20076 26350 20078 26402
rect 20078 26350 20130 26402
rect 20130 26350 20132 26402
rect 20076 26348 20132 26350
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19516 23100 19572 23156
rect 19628 24108 19684 24164
rect 20748 24050 20804 24052
rect 20748 23998 20750 24050
rect 20750 23998 20802 24050
rect 20802 23998 20804 24050
rect 20748 23996 20804 23998
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19852 23100 19908 23156
rect 19628 22930 19684 22932
rect 19628 22878 19630 22930
rect 19630 22878 19682 22930
rect 19682 22878 19684 22930
rect 19628 22876 19684 22878
rect 20300 22876 20356 22932
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19180 20972 19236 21028
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 18844 20076 18900 20132
rect 19404 20130 19460 20132
rect 19404 20078 19406 20130
rect 19406 20078 19458 20130
rect 19458 20078 19460 20130
rect 19404 20076 19460 20078
rect 18284 18620 18340 18676
rect 17948 18508 18004 18564
rect 17836 17666 17892 17668
rect 17836 17614 17838 17666
rect 17838 17614 17890 17666
rect 17890 17614 17892 17666
rect 17836 17612 17892 17614
rect 18060 17554 18116 17556
rect 18060 17502 18062 17554
rect 18062 17502 18114 17554
rect 18114 17502 18116 17554
rect 18060 17500 18116 17502
rect 18396 18508 18452 18564
rect 15932 17388 15988 17444
rect 15708 17106 15764 17108
rect 15708 17054 15710 17106
rect 15710 17054 15762 17106
rect 15762 17054 15764 17106
rect 15708 17052 15764 17054
rect 15036 16098 15092 16100
rect 15036 16046 15038 16098
rect 15038 16046 15090 16098
rect 15090 16046 15092 16098
rect 15036 16044 15092 16046
rect 13244 13634 13300 13636
rect 13244 13582 13246 13634
rect 13246 13582 13298 13634
rect 13298 13582 13300 13634
rect 13244 13580 13300 13582
rect 16044 16716 16100 16772
rect 16828 16828 16884 16884
rect 14028 14530 14084 14532
rect 14028 14478 14030 14530
rect 14030 14478 14082 14530
rect 14082 14478 14084 14530
rect 14028 14476 14084 14478
rect 15260 14252 15316 14308
rect 13692 13746 13748 13748
rect 13692 13694 13694 13746
rect 13694 13694 13746 13746
rect 13746 13694 13748 13746
rect 13692 13692 13748 13694
rect 13580 13580 13636 13636
rect 13468 12572 13524 12628
rect 13916 12572 13972 12628
rect 12236 12178 12292 12180
rect 12236 12126 12238 12178
rect 12238 12126 12290 12178
rect 12290 12126 12292 12178
rect 12236 12124 12292 12126
rect 12348 12066 12404 12068
rect 12348 12014 12350 12066
rect 12350 12014 12402 12066
rect 12402 12014 12404 12066
rect 12348 12012 12404 12014
rect 12796 11452 12852 11508
rect 12908 11340 12964 11396
rect 13468 12124 13524 12180
rect 13580 11506 13636 11508
rect 13580 11454 13582 11506
rect 13582 11454 13634 11506
rect 13634 11454 13636 11506
rect 13580 11452 13636 11454
rect 13692 11394 13748 11396
rect 13692 11342 13694 11394
rect 13694 11342 13746 11394
rect 13746 11342 13748 11394
rect 13692 11340 13748 11342
rect 14924 12236 14980 12292
rect 14252 12124 14308 12180
rect 14588 12178 14644 12180
rect 14588 12126 14590 12178
rect 14590 12126 14642 12178
rect 14642 12126 14644 12178
rect 14588 12124 14644 12126
rect 14028 11788 14084 11844
rect 14476 11340 14532 11396
rect 14700 11788 14756 11844
rect 13580 9660 13636 9716
rect 10332 8316 10388 8372
rect 12684 8092 12740 8148
rect 11228 6636 11284 6692
rect 9548 4898 9604 4900
rect 9548 4846 9550 4898
rect 9550 4846 9602 4898
rect 9602 4846 9604 4898
rect 9548 4844 9604 4846
rect 10892 4844 10948 4900
rect 10220 4338 10276 4340
rect 10220 4286 10222 4338
rect 10222 4286 10274 4338
rect 10274 4286 10276 4338
rect 10220 4284 10276 4286
rect 14924 11452 14980 11508
rect 14924 11116 14980 11172
rect 14252 6578 14308 6580
rect 14252 6526 14254 6578
rect 14254 6526 14306 6578
rect 14306 6526 14308 6578
rect 14252 6524 14308 6526
rect 15484 14476 15540 14532
rect 15484 13970 15540 13972
rect 15484 13918 15486 13970
rect 15486 13918 15538 13970
rect 15538 13918 15540 13970
rect 15484 13916 15540 13918
rect 16716 14588 16772 14644
rect 15708 13746 15764 13748
rect 15708 13694 15710 13746
rect 15710 13694 15762 13746
rect 15762 13694 15764 13746
rect 15708 13692 15764 13694
rect 15596 12178 15652 12180
rect 15596 12126 15598 12178
rect 15598 12126 15650 12178
rect 15650 12126 15652 12178
rect 15596 12124 15652 12126
rect 16492 14306 16548 14308
rect 16492 14254 16494 14306
rect 16494 14254 16546 14306
rect 16546 14254 16548 14306
rect 16492 14252 16548 14254
rect 16380 13970 16436 13972
rect 16380 13918 16382 13970
rect 16382 13918 16434 13970
rect 16434 13918 16436 13970
rect 16380 13916 16436 13918
rect 16268 13804 16324 13860
rect 17052 16156 17108 16212
rect 18620 17612 18676 17668
rect 18284 16716 18340 16772
rect 20076 20018 20132 20020
rect 20076 19966 20078 20018
rect 20078 19966 20130 20018
rect 20130 19966 20132 20018
rect 20076 19964 20132 19966
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19068 18674 19124 18676
rect 19068 18622 19070 18674
rect 19070 18622 19122 18674
rect 19122 18622 19124 18674
rect 19068 18620 19124 18622
rect 18956 18562 19012 18564
rect 18956 18510 18958 18562
rect 18958 18510 19010 18562
rect 19010 18510 19012 18562
rect 18956 18508 19012 18510
rect 20524 20130 20580 20132
rect 20524 20078 20526 20130
rect 20526 20078 20578 20130
rect 20578 20078 20580 20130
rect 20524 20076 20580 20078
rect 21868 34130 21924 34132
rect 21868 34078 21870 34130
rect 21870 34078 21922 34130
rect 21922 34078 21924 34130
rect 21868 34076 21924 34078
rect 21756 32450 21812 32452
rect 21756 32398 21758 32450
rect 21758 32398 21810 32450
rect 21810 32398 21812 32450
rect 21756 32396 21812 32398
rect 21308 32172 21364 32228
rect 21868 32172 21924 32228
rect 22988 37212 23044 37268
rect 22428 33180 22484 33236
rect 22540 32732 22596 32788
rect 22764 32844 22820 32900
rect 23548 37154 23604 37156
rect 23548 37102 23550 37154
rect 23550 37102 23602 37154
rect 23602 37102 23604 37154
rect 23548 37100 23604 37102
rect 23660 35420 23716 35476
rect 24220 39564 24276 39620
rect 23996 37826 24052 37828
rect 23996 37774 23998 37826
rect 23998 37774 24050 37826
rect 24050 37774 24052 37826
rect 23996 37772 24052 37774
rect 24108 37266 24164 37268
rect 24108 37214 24110 37266
rect 24110 37214 24162 37266
rect 24162 37214 24164 37266
rect 24108 37212 24164 37214
rect 24668 41916 24724 41972
rect 24780 40460 24836 40516
rect 24556 40124 24612 40180
rect 25340 45500 25396 45556
rect 25788 46674 25844 46676
rect 25788 46622 25790 46674
rect 25790 46622 25842 46674
rect 25842 46622 25844 46674
rect 25788 46620 25844 46622
rect 25564 45778 25620 45780
rect 25564 45726 25566 45778
rect 25566 45726 25618 45778
rect 25618 45726 25620 45778
rect 25564 45724 25620 45726
rect 26460 53452 26516 53508
rect 27468 54684 27524 54740
rect 28252 54684 28308 54740
rect 28140 53788 28196 53844
rect 27244 53506 27300 53508
rect 27244 53454 27246 53506
rect 27246 53454 27298 53506
rect 27298 53454 27300 53506
rect 27244 53452 27300 53454
rect 27580 53730 27636 53732
rect 27580 53678 27582 53730
rect 27582 53678 27634 53730
rect 27634 53678 27636 53730
rect 27580 53676 27636 53678
rect 27916 53452 27972 53508
rect 28252 53730 28308 53732
rect 28252 53678 28254 53730
rect 28254 53678 28306 53730
rect 28306 53678 28308 53730
rect 28252 53676 28308 53678
rect 29036 54514 29092 54516
rect 29036 54462 29038 54514
rect 29038 54462 29090 54514
rect 29090 54462 29092 54514
rect 29036 54460 29092 54462
rect 28364 52946 28420 52948
rect 28364 52894 28366 52946
rect 28366 52894 28418 52946
rect 28418 52894 28420 52946
rect 28364 52892 28420 52894
rect 32060 55298 32116 55300
rect 32060 55246 32062 55298
rect 32062 55246 32114 55298
rect 32114 55246 32116 55298
rect 32060 55244 32116 55246
rect 33516 55298 33572 55300
rect 33516 55246 33518 55298
rect 33518 55246 33570 55298
rect 33570 55246 33572 55298
rect 33516 55244 33572 55246
rect 34076 55244 34132 55300
rect 29820 55132 29876 55188
rect 29484 53954 29540 53956
rect 29484 53902 29486 53954
rect 29486 53902 29538 53954
rect 29538 53902 29540 53954
rect 29484 53900 29540 53902
rect 29372 53842 29428 53844
rect 29372 53790 29374 53842
rect 29374 53790 29426 53842
rect 29426 53790 29428 53842
rect 29372 53788 29428 53790
rect 29708 53842 29764 53844
rect 29708 53790 29710 53842
rect 29710 53790 29762 53842
rect 29762 53790 29764 53842
rect 29708 53788 29764 53790
rect 31276 55186 31332 55188
rect 31276 55134 31278 55186
rect 31278 55134 31330 55186
rect 31330 55134 31332 55186
rect 31276 55132 31332 55134
rect 31388 55020 31444 55076
rect 30604 53506 30660 53508
rect 30604 53454 30606 53506
rect 30606 53454 30658 53506
rect 30658 53454 30660 53506
rect 30604 53452 30660 53454
rect 29260 52892 29316 52948
rect 27132 50876 27188 50932
rect 26908 50594 26964 50596
rect 26908 50542 26910 50594
rect 26910 50542 26962 50594
rect 26962 50542 26964 50594
rect 26908 50540 26964 50542
rect 26236 50092 26292 50148
rect 26908 50092 26964 50148
rect 26124 49698 26180 49700
rect 26124 49646 26126 49698
rect 26126 49646 26178 49698
rect 26178 49646 26180 49698
rect 26124 49644 26180 49646
rect 26572 49644 26628 49700
rect 26348 49586 26404 49588
rect 26348 49534 26350 49586
rect 26350 49534 26402 49586
rect 26402 49534 26404 49586
rect 26348 49532 26404 49534
rect 26348 49308 26404 49364
rect 26796 48188 26852 48244
rect 26460 46844 26516 46900
rect 26124 46562 26180 46564
rect 26124 46510 26126 46562
rect 26126 46510 26178 46562
rect 26178 46510 26180 46562
rect 26124 46508 26180 46510
rect 26348 45164 26404 45220
rect 26460 45052 26516 45108
rect 25788 44268 25844 44324
rect 25452 43596 25508 43652
rect 25564 43314 25620 43316
rect 25564 43262 25566 43314
rect 25566 43262 25618 43314
rect 25618 43262 25620 43314
rect 25564 43260 25620 43262
rect 25340 42140 25396 42196
rect 25676 42140 25732 42196
rect 25340 41356 25396 41412
rect 25340 40348 25396 40404
rect 25004 40236 25060 40292
rect 24556 39564 24612 39620
rect 25340 39618 25396 39620
rect 25340 39566 25342 39618
rect 25342 39566 25394 39618
rect 25394 39566 25396 39618
rect 25340 39564 25396 39566
rect 24444 39452 24500 39508
rect 24892 39506 24948 39508
rect 24892 39454 24894 39506
rect 24894 39454 24946 39506
rect 24946 39454 24948 39506
rect 24892 39452 24948 39454
rect 24444 39116 24500 39172
rect 25452 36428 25508 36484
rect 25004 36370 25060 36372
rect 25004 36318 25006 36370
rect 25006 36318 25058 36370
rect 25058 36318 25060 36370
rect 25004 36316 25060 36318
rect 25788 41970 25844 41972
rect 25788 41918 25790 41970
rect 25790 41918 25842 41970
rect 25842 41918 25844 41970
rect 25788 41916 25844 41918
rect 26012 42082 26068 42084
rect 26012 42030 26014 42082
rect 26014 42030 26066 42082
rect 26066 42030 26068 42082
rect 26012 42028 26068 42030
rect 26012 41244 26068 41300
rect 26236 41970 26292 41972
rect 26236 41918 26238 41970
rect 26238 41918 26290 41970
rect 26290 41918 26292 41970
rect 26236 41916 26292 41918
rect 26460 44156 26516 44212
rect 26460 42812 26516 42868
rect 26124 41692 26180 41748
rect 25788 41186 25844 41188
rect 25788 41134 25790 41186
rect 25790 41134 25842 41186
rect 25842 41134 25844 41186
rect 25788 41132 25844 41134
rect 25900 40962 25956 40964
rect 25900 40910 25902 40962
rect 25902 40910 25954 40962
rect 25954 40910 25956 40962
rect 25900 40908 25956 40910
rect 26012 40460 26068 40516
rect 26012 39506 26068 39508
rect 26012 39454 26014 39506
rect 26014 39454 26066 39506
rect 26066 39454 26068 39506
rect 26012 39452 26068 39454
rect 26124 36316 26180 36372
rect 26012 35420 26068 35476
rect 24108 32844 24164 32900
rect 22316 32674 22372 32676
rect 22316 32622 22318 32674
rect 22318 32622 22370 32674
rect 22370 32622 22372 32674
rect 22316 32620 22372 32622
rect 22092 32396 22148 32452
rect 22428 32508 22484 32564
rect 23548 32786 23604 32788
rect 23548 32734 23550 32786
rect 23550 32734 23602 32786
rect 23602 32734 23604 32786
rect 23548 32732 23604 32734
rect 24108 32562 24164 32564
rect 24108 32510 24110 32562
rect 24110 32510 24162 32562
rect 24162 32510 24164 32562
rect 24108 32508 24164 32510
rect 24444 32674 24500 32676
rect 24444 32622 24446 32674
rect 24446 32622 24498 32674
rect 24498 32622 24500 32674
rect 24444 32620 24500 32622
rect 22428 31778 22484 31780
rect 22428 31726 22430 31778
rect 22430 31726 22482 31778
rect 22482 31726 22484 31778
rect 22428 31724 22484 31726
rect 23324 32172 23380 32228
rect 25228 33404 25284 33460
rect 24220 32396 24276 32452
rect 22988 31724 23044 31780
rect 22316 31666 22372 31668
rect 22316 31614 22318 31666
rect 22318 31614 22370 31666
rect 22370 31614 22372 31666
rect 22316 31612 22372 31614
rect 24108 31948 24164 32004
rect 21308 27580 21364 27636
rect 21644 27186 21700 27188
rect 21644 27134 21646 27186
rect 21646 27134 21698 27186
rect 21698 27134 21700 27186
rect 21644 27132 21700 27134
rect 22092 28812 22148 28868
rect 22316 28924 22372 28980
rect 26348 41074 26404 41076
rect 26348 41022 26350 41074
rect 26350 41022 26402 41074
rect 26402 41022 26404 41074
rect 26348 41020 26404 41022
rect 28364 51100 28420 51156
rect 28700 50764 28756 50820
rect 28252 50482 28308 50484
rect 28252 50430 28254 50482
rect 28254 50430 28306 50482
rect 28306 50430 28308 50482
rect 28252 50428 28308 50430
rect 28588 50482 28644 50484
rect 28588 50430 28590 50482
rect 28590 50430 28642 50482
rect 28642 50430 28644 50482
rect 28588 50428 28644 50430
rect 28028 48972 28084 49028
rect 27804 48914 27860 48916
rect 27804 48862 27806 48914
rect 27806 48862 27858 48914
rect 27858 48862 27860 48914
rect 27804 48860 27860 48862
rect 28588 47570 28644 47572
rect 28588 47518 28590 47570
rect 28590 47518 28642 47570
rect 28642 47518 28644 47570
rect 28588 47516 28644 47518
rect 26908 46674 26964 46676
rect 26908 46622 26910 46674
rect 26910 46622 26962 46674
rect 26962 46622 26964 46674
rect 26908 46620 26964 46622
rect 26796 46508 26852 46564
rect 26908 46396 26964 46452
rect 26908 45276 26964 45332
rect 27020 45164 27076 45220
rect 28364 46674 28420 46676
rect 28364 46622 28366 46674
rect 28366 46622 28418 46674
rect 28418 46622 28420 46674
rect 28364 46620 28420 46622
rect 28364 45388 28420 45444
rect 27692 45276 27748 45332
rect 27692 44268 27748 44324
rect 27244 42866 27300 42868
rect 27244 42814 27246 42866
rect 27246 42814 27298 42866
rect 27298 42814 27300 42866
rect 27244 42812 27300 42814
rect 26908 41916 26964 41972
rect 27244 41970 27300 41972
rect 27244 41918 27246 41970
rect 27246 41918 27298 41970
rect 27298 41918 27300 41970
rect 27244 41916 27300 41918
rect 26684 41020 26740 41076
rect 26908 40962 26964 40964
rect 26908 40910 26910 40962
rect 26910 40910 26962 40962
rect 26962 40910 26964 40962
rect 26908 40908 26964 40910
rect 26908 39564 26964 39620
rect 26796 38892 26852 38948
rect 26796 36316 26852 36372
rect 27020 38556 27076 38612
rect 27020 37660 27076 37716
rect 27804 44210 27860 44212
rect 27804 44158 27806 44210
rect 27806 44158 27858 44210
rect 27858 44158 27860 44210
rect 27804 44156 27860 44158
rect 27692 42028 27748 42084
rect 27468 41132 27524 41188
rect 27580 38722 27636 38724
rect 27580 38670 27582 38722
rect 27582 38670 27634 38722
rect 27634 38670 27636 38722
rect 27580 38668 27636 38670
rect 27804 40962 27860 40964
rect 27804 40910 27806 40962
rect 27806 40910 27858 40962
rect 27858 40910 27860 40962
rect 27804 40908 27860 40910
rect 28588 46844 28644 46900
rect 28588 45106 28644 45108
rect 28588 45054 28590 45106
rect 28590 45054 28642 45106
rect 28642 45054 28644 45106
rect 28588 45052 28644 45054
rect 29036 48242 29092 48244
rect 29036 48190 29038 48242
rect 29038 48190 29090 48242
rect 29090 48190 29092 48242
rect 29036 48188 29092 48190
rect 30380 51436 30436 51492
rect 30156 50764 30212 50820
rect 29484 50706 29540 50708
rect 29484 50654 29486 50706
rect 29486 50654 29538 50706
rect 29538 50654 29540 50706
rect 29484 50652 29540 50654
rect 30492 50876 30548 50932
rect 29932 50428 29988 50484
rect 31836 53788 31892 53844
rect 31388 52386 31444 52388
rect 31388 52334 31390 52386
rect 31390 52334 31442 52386
rect 31442 52334 31444 52386
rect 31388 52332 31444 52334
rect 31836 52332 31892 52388
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 36428 53788 36484 53844
rect 34300 53676 34356 53732
rect 35868 53452 35924 53508
rect 34076 53004 34132 53060
rect 31724 51938 31780 51940
rect 31724 51886 31726 51938
rect 31726 51886 31778 51938
rect 31778 51886 31780 51938
rect 31724 51884 31780 51886
rect 30828 51490 30884 51492
rect 30828 51438 30830 51490
rect 30830 51438 30882 51490
rect 30882 51438 30884 51490
rect 30828 51436 30884 51438
rect 30716 51378 30772 51380
rect 30716 51326 30718 51378
rect 30718 51326 30770 51378
rect 30770 51326 30772 51378
rect 30716 51324 30772 51326
rect 30716 50428 30772 50484
rect 30828 51100 30884 51156
rect 30716 49810 30772 49812
rect 30716 49758 30718 49810
rect 30718 49758 30770 49810
rect 30770 49758 30772 49810
rect 30716 49756 30772 49758
rect 29932 49644 29988 49700
rect 30268 48972 30324 49028
rect 29820 48914 29876 48916
rect 29820 48862 29822 48914
rect 29822 48862 29874 48914
rect 29874 48862 29876 48914
rect 29820 48860 29876 48862
rect 29708 46620 29764 46676
rect 31276 50876 31332 50932
rect 31164 50540 31220 50596
rect 30940 50428 30996 50484
rect 32396 51436 32452 51492
rect 33292 51884 33348 51940
rect 31836 51378 31892 51380
rect 31836 51326 31838 51378
rect 31838 51326 31890 51378
rect 31890 51326 31892 51378
rect 31836 51324 31892 51326
rect 32284 50540 32340 50596
rect 35196 53058 35252 53060
rect 35196 53006 35198 53058
rect 35198 53006 35250 53058
rect 35250 53006 35252 53058
rect 35196 53004 35252 53006
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 36988 53730 37044 53732
rect 36988 53678 36990 53730
rect 36990 53678 37042 53730
rect 37042 53678 37044 53730
rect 36988 53676 37044 53678
rect 37100 53452 37156 53508
rect 38108 55186 38164 55188
rect 38108 55134 38110 55186
rect 38110 55134 38162 55186
rect 38162 55134 38164 55186
rect 38108 55132 38164 55134
rect 37548 53788 37604 53844
rect 37100 53004 37156 53060
rect 37884 53452 37940 53508
rect 34972 51996 35028 52052
rect 35756 52050 35812 52052
rect 35756 51998 35758 52050
rect 35758 51998 35810 52050
rect 35810 51998 35812 52050
rect 35756 51996 35812 51998
rect 32956 50540 33012 50596
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 31276 49644 31332 49700
rect 31948 49756 32004 49812
rect 31948 48748 32004 48804
rect 30380 47516 30436 47572
rect 32060 47628 32116 47684
rect 31500 46674 31556 46676
rect 31500 46622 31502 46674
rect 31502 46622 31554 46674
rect 31554 46622 31556 46674
rect 31500 46620 31556 46622
rect 29932 45052 29988 45108
rect 28476 41804 28532 41860
rect 28140 41020 28196 41076
rect 27916 39564 27972 39620
rect 30380 44716 30436 44772
rect 30268 44322 30324 44324
rect 30268 44270 30270 44322
rect 30270 44270 30322 44322
rect 30322 44270 30324 44322
rect 30268 44268 30324 44270
rect 29932 42700 29988 42756
rect 30716 43932 30772 43988
rect 30716 43484 30772 43540
rect 30828 43260 30884 43316
rect 29260 42642 29316 42644
rect 29260 42590 29262 42642
rect 29262 42590 29314 42642
rect 29314 42590 29316 42642
rect 29260 42588 29316 42590
rect 30492 42476 30548 42532
rect 29372 41916 29428 41972
rect 30492 41916 30548 41972
rect 29484 41074 29540 41076
rect 29484 41022 29486 41074
rect 29486 41022 29538 41074
rect 29538 41022 29540 41074
rect 29484 41020 29540 41022
rect 30156 41074 30212 41076
rect 30156 41022 30158 41074
rect 30158 41022 30210 41074
rect 30210 41022 30212 41074
rect 30156 41020 30212 41022
rect 30828 42754 30884 42756
rect 30828 42702 30830 42754
rect 30830 42702 30882 42754
rect 30882 42702 30884 42754
rect 30828 42700 30884 42702
rect 31164 43820 31220 43876
rect 32284 48076 32340 48132
rect 31388 45388 31444 45444
rect 32396 44994 32452 44996
rect 32396 44942 32398 44994
rect 32398 44942 32450 44994
rect 32450 44942 32452 44994
rect 32396 44940 32452 44942
rect 32284 44604 32340 44660
rect 31276 43484 31332 43540
rect 32060 43260 32116 43316
rect 31276 42754 31332 42756
rect 31276 42702 31278 42754
rect 31278 42702 31330 42754
rect 31330 42702 31332 42754
rect 31276 42700 31332 42702
rect 30940 42642 30996 42644
rect 30940 42590 30942 42642
rect 30942 42590 30994 42642
rect 30994 42590 30996 42642
rect 30940 42588 30996 42590
rect 31388 41804 31444 41860
rect 28700 40796 28756 40852
rect 29260 40796 29316 40852
rect 29036 40402 29092 40404
rect 29036 40350 29038 40402
rect 29038 40350 29090 40402
rect 29090 40350 29092 40402
rect 29036 40348 29092 40350
rect 29708 39788 29764 39844
rect 30268 39788 30324 39844
rect 29148 39394 29204 39396
rect 29148 39342 29150 39394
rect 29150 39342 29202 39394
rect 29202 39342 29204 39394
rect 29148 39340 29204 39342
rect 26572 36204 26628 36260
rect 26348 35698 26404 35700
rect 26348 35646 26350 35698
rect 26350 35646 26402 35698
rect 26402 35646 26404 35698
rect 26348 35644 26404 35646
rect 26684 35644 26740 35700
rect 26684 35420 26740 35476
rect 25788 34690 25844 34692
rect 25788 34638 25790 34690
rect 25790 34638 25842 34690
rect 25842 34638 25844 34690
rect 25788 34636 25844 34638
rect 26460 34690 26516 34692
rect 26460 34638 26462 34690
rect 26462 34638 26514 34690
rect 26514 34638 26516 34690
rect 26460 34636 26516 34638
rect 27020 35586 27076 35588
rect 27020 35534 27022 35586
rect 27022 35534 27074 35586
rect 27074 35534 27076 35586
rect 27020 35532 27076 35534
rect 26684 33964 26740 34020
rect 25116 30940 25172 30996
rect 25340 31948 25396 32004
rect 26348 32450 26404 32452
rect 26348 32398 26350 32450
rect 26350 32398 26402 32450
rect 26402 32398 26404 32450
rect 26348 32396 26404 32398
rect 26796 31724 26852 31780
rect 25452 30940 25508 30996
rect 25788 30994 25844 30996
rect 25788 30942 25790 30994
rect 25790 30942 25842 30994
rect 25842 30942 25844 30994
rect 25788 30940 25844 30942
rect 23548 28924 23604 28980
rect 22204 26796 22260 26852
rect 26236 30156 26292 30212
rect 24668 30098 24724 30100
rect 24668 30046 24670 30098
rect 24670 30046 24722 30098
rect 24722 30046 24724 30098
rect 24668 30044 24724 30046
rect 27244 34412 27300 34468
rect 28028 38162 28084 38164
rect 28028 38110 28030 38162
rect 28030 38110 28082 38162
rect 28082 38110 28084 38162
rect 28028 38108 28084 38110
rect 28700 37938 28756 37940
rect 28700 37886 28702 37938
rect 28702 37886 28754 37938
rect 28754 37886 28756 37938
rect 28700 37884 28756 37886
rect 27580 37436 27636 37492
rect 28700 37436 28756 37492
rect 27580 36258 27636 36260
rect 27580 36206 27582 36258
rect 27582 36206 27634 36258
rect 27634 36206 27636 36258
rect 27580 36204 27636 36206
rect 28700 37266 28756 37268
rect 28700 37214 28702 37266
rect 28702 37214 28754 37266
rect 28754 37214 28756 37266
rect 28700 37212 28756 37214
rect 27692 35810 27748 35812
rect 27692 35758 27694 35810
rect 27694 35758 27746 35810
rect 27746 35758 27748 35810
rect 27692 35756 27748 35758
rect 27692 33516 27748 33572
rect 28364 35138 28420 35140
rect 28364 35086 28366 35138
rect 28366 35086 28418 35138
rect 28418 35086 28420 35138
rect 28364 35084 28420 35086
rect 27916 33964 27972 34020
rect 27580 32562 27636 32564
rect 27580 32510 27582 32562
rect 27582 32510 27634 32562
rect 27634 32510 27636 32562
rect 27580 32508 27636 32510
rect 27468 31052 27524 31108
rect 27356 30716 27412 30772
rect 27468 30828 27524 30884
rect 26460 30044 26516 30100
rect 24444 29260 24500 29316
rect 25228 29314 25284 29316
rect 25228 29262 25230 29314
rect 25230 29262 25282 29314
rect 25282 29262 25284 29314
rect 25228 29260 25284 29262
rect 26572 28812 26628 28868
rect 26348 28700 26404 28756
rect 27356 29148 27412 29204
rect 27244 28866 27300 28868
rect 27244 28814 27246 28866
rect 27246 28814 27298 28866
rect 27298 28814 27300 28866
rect 27244 28812 27300 28814
rect 27356 28642 27412 28644
rect 27356 28590 27358 28642
rect 27358 28590 27410 28642
rect 27410 28590 27412 28642
rect 27356 28588 27412 28590
rect 23884 28476 23940 28532
rect 23100 28028 23156 28084
rect 22764 26796 22820 26852
rect 22204 25004 22260 25060
rect 22876 24444 22932 24500
rect 21980 23884 22036 23940
rect 22316 23996 22372 24052
rect 22204 23826 22260 23828
rect 22204 23774 22206 23826
rect 22206 23774 22258 23826
rect 22258 23774 22260 23826
rect 22204 23772 22260 23774
rect 22092 23660 22148 23716
rect 21980 23548 22036 23604
rect 21532 23100 21588 23156
rect 22764 23100 22820 23156
rect 23324 25394 23380 25396
rect 23324 25342 23326 25394
rect 23326 25342 23378 25394
rect 23378 25342 23380 25394
rect 23324 25340 23380 25342
rect 23100 24220 23156 24276
rect 23212 24892 23268 24948
rect 23212 23548 23268 23604
rect 25788 28364 25844 28420
rect 26460 28418 26516 28420
rect 26460 28366 26462 28418
rect 26462 28366 26514 28418
rect 26514 28366 26516 28418
rect 26460 28364 26516 28366
rect 28028 31500 28084 31556
rect 28252 32060 28308 32116
rect 27916 31052 27972 31108
rect 27916 30268 27972 30324
rect 27356 28140 27412 28196
rect 26012 27858 26068 27860
rect 26012 27806 26014 27858
rect 26014 27806 26066 27858
rect 26066 27806 26068 27858
rect 26012 27804 26068 27806
rect 26572 27804 26628 27860
rect 23996 27020 24052 27076
rect 25564 27746 25620 27748
rect 25564 27694 25566 27746
rect 25566 27694 25618 27746
rect 25618 27694 25620 27746
rect 25564 27692 25620 27694
rect 24444 27634 24500 27636
rect 24444 27582 24446 27634
rect 24446 27582 24498 27634
rect 24498 27582 24500 27634
rect 24444 27580 24500 27582
rect 25340 27634 25396 27636
rect 25340 27582 25342 27634
rect 25342 27582 25394 27634
rect 25394 27582 25396 27634
rect 25340 27580 25396 27582
rect 26124 27692 26180 27748
rect 25564 27132 25620 27188
rect 24220 26796 24276 26852
rect 25900 27074 25956 27076
rect 25900 27022 25902 27074
rect 25902 27022 25954 27074
rect 25954 27022 25956 27074
rect 25900 27020 25956 27022
rect 26124 27020 26180 27076
rect 25788 26348 25844 26404
rect 26012 26908 26068 26964
rect 24332 26290 24388 26292
rect 24332 26238 24334 26290
rect 24334 26238 24386 26290
rect 24386 26238 24388 26290
rect 24332 26236 24388 26238
rect 25452 26290 25508 26292
rect 25452 26238 25454 26290
rect 25454 26238 25506 26290
rect 25506 26238 25508 26290
rect 25452 26236 25508 26238
rect 26348 26514 26404 26516
rect 26348 26462 26350 26514
rect 26350 26462 26402 26514
rect 26402 26462 26404 26514
rect 26348 26460 26404 26462
rect 26796 27074 26852 27076
rect 26796 27022 26798 27074
rect 26798 27022 26850 27074
rect 26850 27022 26852 27074
rect 26796 27020 26852 27022
rect 27132 27804 27188 27860
rect 27356 27692 27412 27748
rect 27020 26962 27076 26964
rect 27020 26910 27022 26962
rect 27022 26910 27074 26962
rect 27074 26910 27076 26962
rect 27020 26908 27076 26910
rect 27244 26514 27300 26516
rect 27244 26462 27246 26514
rect 27246 26462 27298 26514
rect 27298 26462 27300 26514
rect 27244 26460 27300 26462
rect 26460 26178 26516 26180
rect 26460 26126 26462 26178
rect 26462 26126 26514 26178
rect 26514 26126 26516 26178
rect 26460 26124 26516 26126
rect 27356 26124 27412 26180
rect 23548 24892 23604 24948
rect 24220 25116 24276 25172
rect 23660 23996 23716 24052
rect 24108 24498 24164 24500
rect 24108 24446 24110 24498
rect 24110 24446 24162 24498
rect 24162 24446 24164 24498
rect 24108 24444 24164 24446
rect 23772 23772 23828 23828
rect 21644 22316 21700 22372
rect 22428 22428 22484 22484
rect 22652 22316 22708 22372
rect 23996 24108 24052 24164
rect 24108 23660 24164 23716
rect 23884 23154 23940 23156
rect 23884 23102 23886 23154
rect 23886 23102 23938 23154
rect 23938 23102 23940 23154
rect 23884 23100 23940 23102
rect 24556 23100 24612 23156
rect 22988 21532 23044 21588
rect 22652 21026 22708 21028
rect 22652 20974 22654 21026
rect 22654 20974 22706 21026
rect 22706 20974 22708 21026
rect 22652 20972 22708 20974
rect 23212 21474 23268 21476
rect 23212 21422 23214 21474
rect 23214 21422 23266 21474
rect 23266 21422 23268 21474
rect 23212 21420 23268 21422
rect 22428 20748 22484 20804
rect 23212 20748 23268 20804
rect 25340 23154 25396 23156
rect 25340 23102 25342 23154
rect 25342 23102 25394 23154
rect 25394 23102 25396 23154
rect 25340 23100 25396 23102
rect 24668 22428 24724 22484
rect 23436 21026 23492 21028
rect 23436 20974 23438 21026
rect 23438 20974 23490 21026
rect 23490 20974 23492 21026
rect 23436 20972 23492 20974
rect 21196 19964 21252 20020
rect 23548 21532 23604 21588
rect 24108 21586 24164 21588
rect 24108 21534 24110 21586
rect 24110 21534 24162 21586
rect 24162 21534 24164 21586
rect 24108 21532 24164 21534
rect 23772 21420 23828 21476
rect 22540 19516 22596 19572
rect 22988 19180 23044 19236
rect 20748 19068 20804 19124
rect 22540 19122 22596 19124
rect 22540 19070 22542 19122
rect 22542 19070 22594 19122
rect 22594 19070 22596 19122
rect 22540 19068 22596 19070
rect 21868 18956 21924 19012
rect 20188 18284 20244 18340
rect 19180 17500 19236 17556
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20412 17388 20468 17444
rect 21420 17442 21476 17444
rect 21420 17390 21422 17442
rect 21422 17390 21474 17442
rect 21474 17390 21476 17442
rect 21420 17388 21476 17390
rect 20188 15372 20244 15428
rect 17388 13916 17444 13972
rect 16828 13692 16884 13748
rect 17724 14418 17780 14420
rect 17724 14366 17726 14418
rect 17726 14366 17778 14418
rect 17778 14366 17780 14418
rect 17724 14364 17780 14366
rect 17612 13580 17668 13636
rect 18172 13746 18228 13748
rect 18172 13694 18174 13746
rect 18174 13694 18226 13746
rect 18226 13694 18228 13746
rect 18172 13692 18228 13694
rect 15932 12348 15988 12404
rect 17500 12402 17556 12404
rect 17500 12350 17502 12402
rect 17502 12350 17554 12402
rect 17554 12350 17556 12402
rect 17500 12348 17556 12350
rect 15484 11676 15540 11732
rect 16156 11506 16212 11508
rect 16156 11454 16158 11506
rect 16158 11454 16210 11506
rect 16210 11454 16212 11506
rect 16156 11452 16212 11454
rect 15372 9212 15428 9268
rect 16716 9884 16772 9940
rect 15596 9100 15652 9156
rect 15148 9042 15204 9044
rect 15148 8990 15150 9042
rect 15150 8990 15202 9042
rect 15202 8990 15204 9042
rect 15148 8988 15204 8990
rect 15708 8988 15764 9044
rect 17388 9714 17444 9716
rect 17388 9662 17390 9714
rect 17390 9662 17442 9714
rect 17442 9662 17444 9714
rect 17388 9660 17444 9662
rect 18172 9154 18228 9156
rect 18172 9102 18174 9154
rect 18174 9102 18226 9154
rect 18226 9102 18228 9154
rect 18172 9100 18228 9102
rect 14924 5852 14980 5908
rect 15708 5906 15764 5908
rect 15708 5854 15710 5906
rect 15710 5854 15762 5906
rect 15762 5854 15764 5906
rect 15708 5852 15764 5854
rect 16268 6524 16324 6580
rect 16380 6412 16436 6468
rect 20188 14418 20244 14420
rect 20188 14366 20190 14418
rect 20190 14366 20242 14418
rect 20242 14366 20244 14418
rect 20188 14364 20244 14366
rect 19740 14252 19796 14308
rect 19180 13634 19236 13636
rect 19180 13582 19182 13634
rect 19182 13582 19234 13634
rect 19234 13582 19236 13634
rect 19180 13580 19236 13582
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 20076 12684 20132 12740
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19180 11788 19236 11844
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 20300 10108 20356 10164
rect 19068 9884 19124 9940
rect 19404 9602 19460 9604
rect 19404 9550 19406 9602
rect 19406 9550 19458 9602
rect 19458 9550 19460 9602
rect 19404 9548 19460 9550
rect 20076 9602 20132 9604
rect 20076 9550 20078 9602
rect 20078 9550 20130 9602
rect 20130 9550 20132 9602
rect 20076 9548 20132 9550
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 18956 8428 19012 8484
rect 19404 8876 19460 8932
rect 19628 8764 19684 8820
rect 18508 7308 18564 7364
rect 19068 7362 19124 7364
rect 19068 7310 19070 7362
rect 19070 7310 19122 7362
rect 19122 7310 19124 7362
rect 19068 7308 19124 7310
rect 17388 6690 17444 6692
rect 17388 6638 17390 6690
rect 17390 6638 17442 6690
rect 17442 6638 17444 6690
rect 17388 6636 17444 6638
rect 16828 6300 16884 6356
rect 16940 6466 16996 6468
rect 16940 6414 16942 6466
rect 16942 6414 16994 6466
rect 16994 6414 16996 6466
rect 16940 6412 16996 6414
rect 16828 6130 16884 6132
rect 16828 6078 16830 6130
rect 16830 6078 16882 6130
rect 16882 6078 16884 6130
rect 16828 6076 16884 6078
rect 17948 6300 18004 6356
rect 16828 5852 16884 5908
rect 20076 8428 20132 8484
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 20076 7644 20132 7700
rect 19068 6076 19124 6132
rect 19516 6690 19572 6692
rect 19516 6638 19518 6690
rect 19518 6638 19570 6690
rect 19570 6638 19572 6690
rect 19516 6636 19572 6638
rect 19964 6690 20020 6692
rect 19964 6638 19966 6690
rect 19966 6638 20018 6690
rect 20018 6638 20020 6690
rect 19964 6636 20020 6638
rect 19292 6300 19348 6356
rect 19292 6076 19348 6132
rect 11228 4284 11284 4340
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 16044 5292 16100 5348
rect 14588 5180 14644 5236
rect 15932 5234 15988 5236
rect 15932 5182 15934 5234
rect 15934 5182 15986 5234
rect 15986 5182 15988 5234
rect 15932 5180 15988 5182
rect 16268 5740 16324 5796
rect 17724 5794 17780 5796
rect 17724 5742 17726 5794
rect 17726 5742 17778 5794
rect 17778 5742 17780 5794
rect 17724 5740 17780 5742
rect 17612 5180 17668 5236
rect 16716 5068 16772 5124
rect 13356 4284 13412 4340
rect 13020 4226 13076 4228
rect 13020 4174 13022 4226
rect 13022 4174 13074 4226
rect 13074 4174 13076 4226
rect 13020 4172 13076 4174
rect 17836 5068 17892 5124
rect 18172 5122 18228 5124
rect 18172 5070 18174 5122
rect 18174 5070 18226 5122
rect 18226 5070 18228 5122
rect 18172 5068 18228 5070
rect 18396 5122 18452 5124
rect 18396 5070 18398 5122
rect 18398 5070 18450 5122
rect 18450 5070 18452 5122
rect 18396 5068 18452 5070
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19404 5292 19460 5348
rect 17836 4844 17892 4900
rect 18620 4898 18676 4900
rect 18620 4846 18622 4898
rect 18622 4846 18674 4898
rect 18674 4846 18676 4898
rect 18620 4844 18676 4846
rect 19740 5068 19796 5124
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 12796 3500 12852 3556
rect 4732 3276 4788 3332
rect 5516 3330 5572 3332
rect 5516 3278 5518 3330
rect 5518 3278 5570 3330
rect 5570 3278 5572 3330
rect 5516 3276 5572 3278
rect 20524 14306 20580 14308
rect 20524 14254 20526 14306
rect 20526 14254 20578 14306
rect 20578 14254 20580 14306
rect 20524 14252 20580 14254
rect 20748 14530 20804 14532
rect 20748 14478 20750 14530
rect 20750 14478 20802 14530
rect 20802 14478 20804 14530
rect 20748 14476 20804 14478
rect 21420 13074 21476 13076
rect 21420 13022 21422 13074
rect 21422 13022 21474 13074
rect 21474 13022 21476 13074
rect 21420 13020 21476 13022
rect 21308 11676 21364 11732
rect 22316 18338 22372 18340
rect 22316 18286 22318 18338
rect 22318 18286 22370 18338
rect 22370 18286 22372 18338
rect 22316 18284 22372 18286
rect 23772 20636 23828 20692
rect 22764 18338 22820 18340
rect 22764 18286 22766 18338
rect 22766 18286 22818 18338
rect 22818 18286 22820 18338
rect 22764 18284 22820 18286
rect 23548 18396 23604 18452
rect 23324 17052 23380 17108
rect 22988 16604 23044 16660
rect 23884 17106 23940 17108
rect 23884 17054 23886 17106
rect 23886 17054 23938 17106
rect 23938 17054 23940 17106
rect 23884 17052 23940 17054
rect 23436 15820 23492 15876
rect 22764 15036 22820 15092
rect 22988 14642 23044 14644
rect 22988 14590 22990 14642
rect 22990 14590 23042 14642
rect 23042 14590 23044 14642
rect 22988 14588 23044 14590
rect 22764 14476 22820 14532
rect 21868 13692 21924 13748
rect 22540 13804 22596 13860
rect 22092 13020 22148 13076
rect 21980 12738 22036 12740
rect 21980 12686 21982 12738
rect 21982 12686 22034 12738
rect 22034 12686 22036 12738
rect 21980 12684 22036 12686
rect 22876 13020 22932 13076
rect 22988 14364 23044 14420
rect 23660 15090 23716 15092
rect 23660 15038 23662 15090
rect 23662 15038 23714 15090
rect 23714 15038 23716 15090
rect 23660 15036 23716 15038
rect 23884 15148 23940 15204
rect 24444 19180 24500 19236
rect 25676 22482 25732 22484
rect 25676 22430 25678 22482
rect 25678 22430 25730 22482
rect 25730 22430 25732 22482
rect 25676 22428 25732 22430
rect 25340 21420 25396 21476
rect 24108 18172 24164 18228
rect 26796 23042 26852 23044
rect 26796 22990 26798 23042
rect 26798 22990 26850 23042
rect 26850 22990 26852 23042
rect 26796 22988 26852 22990
rect 26012 21420 26068 21476
rect 25228 18450 25284 18452
rect 25228 18398 25230 18450
rect 25230 18398 25282 18450
rect 25282 18398 25284 18450
rect 25228 18396 25284 18398
rect 25340 18060 25396 18116
rect 24668 16994 24724 16996
rect 24668 16942 24670 16994
rect 24670 16942 24722 16994
rect 24722 16942 24724 16994
rect 24668 16940 24724 16942
rect 25340 16940 25396 16996
rect 24332 16604 24388 16660
rect 25900 20018 25956 20020
rect 25900 19966 25902 20018
rect 25902 19966 25954 20018
rect 25954 19966 25956 20018
rect 25900 19964 25956 19966
rect 25788 16492 25844 16548
rect 24332 16098 24388 16100
rect 24332 16046 24334 16098
rect 24334 16046 24386 16098
rect 24386 16046 24388 16098
rect 24332 16044 24388 16046
rect 25004 16098 25060 16100
rect 25004 16046 25006 16098
rect 25006 16046 25058 16098
rect 25058 16046 25060 16098
rect 25004 16044 25060 16046
rect 24332 15820 24388 15876
rect 23772 13916 23828 13972
rect 23660 13804 23716 13860
rect 23436 13746 23492 13748
rect 23436 13694 23438 13746
rect 23438 13694 23490 13746
rect 23490 13694 23492 13746
rect 23436 13692 23492 13694
rect 25676 15260 25732 15316
rect 27020 22428 27076 22484
rect 27356 22428 27412 22484
rect 26348 21420 26404 21476
rect 26796 21474 26852 21476
rect 26796 21422 26798 21474
rect 26798 21422 26850 21474
rect 26850 21422 26852 21474
rect 26796 21420 26852 21422
rect 27804 28140 27860 28196
rect 27580 26962 27636 26964
rect 27580 26910 27582 26962
rect 27582 26910 27634 26962
rect 27634 26910 27636 26962
rect 27580 26908 27636 26910
rect 28028 30716 28084 30772
rect 27916 25340 27972 25396
rect 27804 22988 27860 23044
rect 28140 29148 28196 29204
rect 28140 27692 28196 27748
rect 28476 31500 28532 31556
rect 28364 27858 28420 27860
rect 28364 27806 28366 27858
rect 28366 27806 28418 27858
rect 28418 27806 28420 27858
rect 28364 27804 28420 27806
rect 28700 30882 28756 30884
rect 28700 30830 28702 30882
rect 28702 30830 28754 30882
rect 28754 30830 28756 30882
rect 28700 30828 28756 30830
rect 28700 28364 28756 28420
rect 28700 27468 28756 27524
rect 28252 26348 28308 26404
rect 28140 26236 28196 26292
rect 28140 25228 28196 25284
rect 28364 26012 28420 26068
rect 30604 39340 30660 39396
rect 30380 38722 30436 38724
rect 30380 38670 30382 38722
rect 30382 38670 30434 38722
rect 30434 38670 30436 38722
rect 30380 38668 30436 38670
rect 32284 43260 32340 43316
rect 32284 42082 32340 42084
rect 32284 42030 32286 42082
rect 32286 42030 32338 42082
rect 32338 42030 32340 42082
rect 32284 42028 32340 42030
rect 32396 41970 32452 41972
rect 32396 41918 32398 41970
rect 32398 41918 32450 41970
rect 32450 41918 32452 41970
rect 32396 41916 32452 41918
rect 31836 41804 31892 41860
rect 32284 41858 32340 41860
rect 32284 41806 32286 41858
rect 32286 41806 32338 41858
rect 32338 41806 32340 41858
rect 32284 41804 32340 41806
rect 32508 38946 32564 38948
rect 32508 38894 32510 38946
rect 32510 38894 32562 38946
rect 32562 38894 32564 38946
rect 32508 38892 32564 38894
rect 31612 38668 31668 38724
rect 30156 38108 30212 38164
rect 29260 37938 29316 37940
rect 29260 37886 29262 37938
rect 29262 37886 29314 37938
rect 29314 37886 29316 37938
rect 29260 37884 29316 37886
rect 29036 37826 29092 37828
rect 29036 37774 29038 37826
rect 29038 37774 29090 37826
rect 29090 37774 29092 37826
rect 29036 37772 29092 37774
rect 29260 37548 29316 37604
rect 29148 37436 29204 37492
rect 29484 37266 29540 37268
rect 29484 37214 29486 37266
rect 29486 37214 29538 37266
rect 29538 37214 29540 37266
rect 29484 37212 29540 37214
rect 30156 37154 30212 37156
rect 30156 37102 30158 37154
rect 30158 37102 30210 37154
rect 30210 37102 30212 37154
rect 30156 37100 30212 37102
rect 29036 35922 29092 35924
rect 29036 35870 29038 35922
rect 29038 35870 29090 35922
rect 29090 35870 29092 35922
rect 29036 35868 29092 35870
rect 29596 35084 29652 35140
rect 31388 37436 31444 37492
rect 31276 36988 31332 37044
rect 30828 35756 30884 35812
rect 30492 35532 30548 35588
rect 29372 32732 29428 32788
rect 31164 33516 31220 33572
rect 29708 33346 29764 33348
rect 29708 33294 29710 33346
rect 29710 33294 29762 33346
rect 29762 33294 29764 33346
rect 29708 33292 29764 33294
rect 31164 32844 31220 32900
rect 29596 32508 29652 32564
rect 29260 32396 29316 32452
rect 29148 31890 29204 31892
rect 29148 31838 29150 31890
rect 29150 31838 29202 31890
rect 29202 31838 29204 31890
rect 29148 31836 29204 31838
rect 29484 31724 29540 31780
rect 29820 32732 29876 32788
rect 31612 33180 31668 33236
rect 30940 32674 30996 32676
rect 30940 32622 30942 32674
rect 30942 32622 30994 32674
rect 30994 32622 30996 32674
rect 30940 32620 30996 32622
rect 30156 30828 30212 30884
rect 29932 30210 29988 30212
rect 29932 30158 29934 30210
rect 29934 30158 29986 30210
rect 29986 30158 29988 30210
rect 29932 30156 29988 30158
rect 29932 29932 29988 29988
rect 29036 28642 29092 28644
rect 29036 28590 29038 28642
rect 29038 28590 29090 28642
rect 29090 28590 29092 28642
rect 29036 28588 29092 28590
rect 29372 28364 29428 28420
rect 30828 32284 30884 32340
rect 31052 32450 31108 32452
rect 31052 32398 31054 32450
rect 31054 32398 31106 32450
rect 31106 32398 31108 32450
rect 31052 32396 31108 32398
rect 31276 32284 31332 32340
rect 31500 31778 31556 31780
rect 31500 31726 31502 31778
rect 31502 31726 31554 31778
rect 31554 31726 31556 31778
rect 31500 31724 31556 31726
rect 32508 38556 32564 38612
rect 32060 37490 32116 37492
rect 32060 37438 32062 37490
rect 32062 37438 32114 37490
rect 32114 37438 32116 37490
rect 32060 37436 32116 37438
rect 31948 36988 32004 37044
rect 32396 37100 32452 37156
rect 32396 36652 32452 36708
rect 32620 36988 32676 37044
rect 31836 36092 31892 36148
rect 31948 35698 32004 35700
rect 31948 35646 31950 35698
rect 31950 35646 32002 35698
rect 32002 35646 32004 35698
rect 31948 35644 32004 35646
rect 32060 35586 32116 35588
rect 32060 35534 32062 35586
rect 32062 35534 32114 35586
rect 32114 35534 32116 35586
rect 32060 35532 32116 35534
rect 32172 33516 32228 33572
rect 32620 34636 32676 34692
rect 31948 33234 32004 33236
rect 31948 33182 31950 33234
rect 31950 33182 32002 33234
rect 32002 33182 32004 33234
rect 31948 33180 32004 33182
rect 31836 32844 31892 32900
rect 32732 34300 32788 34356
rect 31836 31612 31892 31668
rect 31724 31218 31780 31220
rect 31724 31166 31726 31218
rect 31726 31166 31778 31218
rect 31778 31166 31780 31218
rect 31724 31164 31780 31166
rect 31500 31052 31556 31108
rect 31052 30994 31108 30996
rect 31052 30942 31054 30994
rect 31054 30942 31106 30994
rect 31106 30942 31108 30994
rect 31052 30940 31108 30942
rect 31948 30994 32004 30996
rect 31948 30942 31950 30994
rect 31950 30942 32002 30994
rect 32002 30942 32004 30994
rect 31948 30940 32004 30942
rect 31836 30882 31892 30884
rect 31836 30830 31838 30882
rect 31838 30830 31890 30882
rect 31890 30830 31892 30882
rect 31836 30828 31892 30830
rect 30604 30210 30660 30212
rect 30604 30158 30606 30210
rect 30606 30158 30658 30210
rect 30658 30158 30660 30210
rect 30604 30156 30660 30158
rect 31052 28754 31108 28756
rect 31052 28702 31054 28754
rect 31054 28702 31106 28754
rect 31106 28702 31108 28754
rect 31052 28700 31108 28702
rect 32508 28700 32564 28756
rect 30268 28028 30324 28084
rect 30044 27692 30100 27748
rect 29820 27074 29876 27076
rect 29820 27022 29822 27074
rect 29822 27022 29874 27074
rect 29874 27022 29876 27074
rect 29820 27020 29876 27022
rect 29596 26236 29652 26292
rect 28812 25676 28868 25732
rect 28588 25228 28644 25284
rect 26460 20018 26516 20020
rect 26460 19966 26462 20018
rect 26462 19966 26514 20018
rect 26514 19966 26516 20018
rect 26460 19964 26516 19966
rect 26908 20018 26964 20020
rect 26908 19966 26910 20018
rect 26910 19966 26962 20018
rect 26962 19966 26964 20018
rect 26908 19964 26964 19966
rect 28812 23154 28868 23156
rect 28812 23102 28814 23154
rect 28814 23102 28866 23154
rect 28866 23102 28868 23154
rect 28812 23100 28868 23102
rect 29148 23042 29204 23044
rect 29148 22990 29150 23042
rect 29150 22990 29202 23042
rect 29202 22990 29204 23042
rect 29148 22988 29204 22990
rect 27916 20076 27972 20132
rect 26348 19852 26404 19908
rect 27692 20018 27748 20020
rect 27692 19966 27694 20018
rect 27694 19966 27746 20018
rect 27746 19966 27748 20018
rect 27692 19964 27748 19966
rect 28252 19906 28308 19908
rect 28252 19854 28254 19906
rect 28254 19854 28306 19906
rect 28306 19854 28308 19906
rect 28252 19852 28308 19854
rect 27356 19404 27412 19460
rect 27692 19516 27748 19572
rect 27356 19234 27412 19236
rect 27356 19182 27358 19234
rect 27358 19182 27410 19234
rect 27410 19182 27412 19234
rect 27356 19180 27412 19182
rect 27020 18172 27076 18228
rect 27580 17554 27636 17556
rect 27580 17502 27582 17554
rect 27582 17502 27634 17554
rect 27634 17502 27636 17554
rect 27580 17500 27636 17502
rect 26236 17052 26292 17108
rect 27916 17554 27972 17556
rect 27916 17502 27918 17554
rect 27918 17502 27970 17554
rect 27970 17502 27972 17554
rect 27916 17500 27972 17502
rect 27020 16492 27076 16548
rect 27804 16492 27860 16548
rect 28140 15372 28196 15428
rect 24668 14418 24724 14420
rect 24668 14366 24670 14418
rect 24670 14366 24722 14418
rect 24722 14366 24724 14418
rect 24668 14364 24724 14366
rect 24668 13970 24724 13972
rect 24668 13918 24670 13970
rect 24670 13918 24722 13970
rect 24722 13918 24724 13970
rect 24668 13916 24724 13918
rect 25228 13916 25284 13972
rect 25452 13858 25508 13860
rect 25452 13806 25454 13858
rect 25454 13806 25506 13858
rect 25506 13806 25508 13858
rect 25452 13804 25508 13806
rect 24780 13020 24836 13076
rect 22876 12796 22932 12852
rect 21532 11452 21588 11508
rect 21756 10332 21812 10388
rect 20748 9938 20804 9940
rect 20748 9886 20750 9938
rect 20750 9886 20802 9938
rect 20802 9886 20804 9938
rect 20748 9884 20804 9886
rect 25116 11506 25172 11508
rect 25116 11454 25118 11506
rect 25118 11454 25170 11506
rect 25170 11454 25172 11506
rect 25116 11452 25172 11454
rect 24780 11116 24836 11172
rect 24108 10722 24164 10724
rect 24108 10670 24110 10722
rect 24110 10670 24162 10722
rect 24162 10670 24164 10722
rect 24108 10668 24164 10670
rect 22204 10444 22260 10500
rect 22540 9996 22596 10052
rect 22876 10610 22932 10612
rect 22876 10558 22878 10610
rect 22878 10558 22930 10610
rect 22930 10558 22932 10610
rect 22876 10556 22932 10558
rect 22652 10332 22708 10388
rect 20972 9548 21028 9604
rect 21868 9548 21924 9604
rect 20748 8930 20804 8932
rect 20748 8878 20750 8930
rect 20750 8878 20802 8930
rect 20802 8878 20804 8930
rect 20748 8876 20804 8878
rect 20636 8818 20692 8820
rect 20636 8766 20638 8818
rect 20638 8766 20690 8818
rect 20690 8766 20692 8818
rect 20636 8764 20692 8766
rect 20412 7868 20468 7924
rect 20636 8428 20692 8484
rect 20412 5068 20468 5124
rect 21308 8428 21364 8484
rect 21980 6802 22036 6804
rect 21980 6750 21982 6802
rect 21982 6750 22034 6802
rect 22034 6750 22036 6802
rect 21980 6748 22036 6750
rect 22764 10108 22820 10164
rect 23884 10610 23940 10612
rect 23884 10558 23886 10610
rect 23886 10558 23938 10610
rect 23938 10558 23940 10610
rect 23884 10556 23940 10558
rect 23772 10498 23828 10500
rect 23772 10446 23774 10498
rect 23774 10446 23826 10498
rect 23826 10446 23828 10498
rect 23772 10444 23828 10446
rect 23436 9996 23492 10052
rect 23212 7980 23268 8036
rect 22876 6802 22932 6804
rect 22876 6750 22878 6802
rect 22878 6750 22930 6802
rect 22930 6750 22932 6802
rect 22876 6748 22932 6750
rect 22988 6690 23044 6692
rect 22988 6638 22990 6690
rect 22990 6638 23042 6690
rect 23042 6638 23044 6690
rect 22988 6636 23044 6638
rect 22764 6578 22820 6580
rect 22764 6526 22766 6578
rect 22766 6526 22818 6578
rect 22818 6526 22820 6578
rect 22764 6524 22820 6526
rect 23548 6524 23604 6580
rect 21756 6412 21812 6468
rect 21308 6130 21364 6132
rect 21308 6078 21310 6130
rect 21310 6078 21362 6130
rect 21362 6078 21364 6130
rect 21308 6076 21364 6078
rect 24556 8034 24612 8036
rect 24556 7982 24558 8034
rect 24558 7982 24610 8034
rect 24610 7982 24612 8034
rect 24556 7980 24612 7982
rect 24668 7308 24724 7364
rect 24780 7420 24836 7476
rect 24108 6636 24164 6692
rect 23884 6524 23940 6580
rect 20748 5122 20804 5124
rect 20748 5070 20750 5122
rect 20750 5070 20802 5122
rect 20802 5070 20804 5122
rect 20748 5068 20804 5070
rect 21644 5122 21700 5124
rect 21644 5070 21646 5122
rect 21646 5070 21698 5122
rect 21698 5070 21700 5122
rect 21644 5068 21700 5070
rect 22764 5292 22820 5348
rect 21420 4844 21476 4900
rect 21868 4898 21924 4900
rect 21868 4846 21870 4898
rect 21870 4846 21922 4898
rect 21922 4846 21924 4898
rect 21868 4844 21924 4846
rect 22876 5180 22932 5236
rect 20300 4060 20356 4116
rect 20860 3612 20916 3668
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 22092 3666 22148 3668
rect 22092 3614 22094 3666
rect 22094 3614 22146 3666
rect 22146 3614 22148 3666
rect 22092 3612 22148 3614
rect 21084 3554 21140 3556
rect 21084 3502 21086 3554
rect 21086 3502 21138 3554
rect 21138 3502 21140 3554
rect 21084 3500 21140 3502
rect 24108 5234 24164 5236
rect 24108 5182 24110 5234
rect 24110 5182 24162 5234
rect 24162 5182 24164 5234
rect 24108 5180 24164 5182
rect 23772 5068 23828 5124
rect 24892 8204 24948 8260
rect 24780 6412 24836 6468
rect 25340 11228 25396 11284
rect 25340 10668 25396 10724
rect 28140 15036 28196 15092
rect 26908 13746 26964 13748
rect 26908 13694 26910 13746
rect 26910 13694 26962 13746
rect 26962 13694 26964 13746
rect 26908 13692 26964 13694
rect 30828 27634 30884 27636
rect 30828 27582 30830 27634
rect 30830 27582 30882 27634
rect 30882 27582 30884 27634
rect 30828 27580 30884 27582
rect 31276 28082 31332 28084
rect 31276 28030 31278 28082
rect 31278 28030 31330 28082
rect 31330 28030 31332 28082
rect 31276 28028 31332 28030
rect 32172 28082 32228 28084
rect 32172 28030 32174 28082
rect 32174 28030 32226 28082
rect 32226 28030 32228 28082
rect 32172 28028 32228 28030
rect 31724 27916 31780 27972
rect 31164 27858 31220 27860
rect 31164 27806 31166 27858
rect 31166 27806 31218 27858
rect 31218 27806 31220 27858
rect 31164 27804 31220 27806
rect 31388 27746 31444 27748
rect 31388 27694 31390 27746
rect 31390 27694 31442 27746
rect 31442 27694 31444 27746
rect 31388 27692 31444 27694
rect 30156 25116 30212 25172
rect 30268 25340 30324 25396
rect 31612 26796 31668 26852
rect 31836 27804 31892 27860
rect 30716 26290 30772 26292
rect 30716 26238 30718 26290
rect 30718 26238 30770 26290
rect 30770 26238 30772 26290
rect 30716 26236 30772 26238
rect 31948 27074 32004 27076
rect 31948 27022 31950 27074
rect 31950 27022 32002 27074
rect 32002 27022 32004 27074
rect 31948 27020 32004 27022
rect 32172 26796 32228 26852
rect 30716 25564 30772 25620
rect 31388 25618 31444 25620
rect 31388 25566 31390 25618
rect 31390 25566 31442 25618
rect 31442 25566 31444 25618
rect 31388 25564 31444 25566
rect 31836 23772 31892 23828
rect 31948 23714 32004 23716
rect 31948 23662 31950 23714
rect 31950 23662 32002 23714
rect 32002 23662 32004 23714
rect 31948 23660 32004 23662
rect 29708 23436 29764 23492
rect 29260 19180 29316 19236
rect 29372 23100 29428 23156
rect 31500 23436 31556 23492
rect 29708 22988 29764 23044
rect 31276 23042 31332 23044
rect 31276 22990 31278 23042
rect 31278 22990 31330 23042
rect 31330 22990 31332 23042
rect 31276 22988 31332 22990
rect 32060 23324 32116 23380
rect 32508 23772 32564 23828
rect 31612 22764 31668 22820
rect 32508 22764 32564 22820
rect 32284 22652 32340 22708
rect 31500 22258 31556 22260
rect 31500 22206 31502 22258
rect 31502 22206 31554 22258
rect 31554 22206 31556 22258
rect 31500 22204 31556 22206
rect 32508 22204 32564 22260
rect 29820 20018 29876 20020
rect 29820 19966 29822 20018
rect 29822 19966 29874 20018
rect 29874 19966 29876 20018
rect 29820 19964 29876 19966
rect 29372 17500 29428 17556
rect 28364 14812 28420 14868
rect 26572 13356 26628 13412
rect 25788 13074 25844 13076
rect 25788 13022 25790 13074
rect 25790 13022 25842 13074
rect 25842 13022 25844 13074
rect 25788 13020 25844 13022
rect 26460 11282 26516 11284
rect 26460 11230 26462 11282
rect 26462 11230 26514 11282
rect 26514 11230 26516 11282
rect 26460 11228 26516 11230
rect 25676 11170 25732 11172
rect 25676 11118 25678 11170
rect 25678 11118 25730 11170
rect 25730 11118 25732 11170
rect 25676 11116 25732 11118
rect 26236 9996 26292 10052
rect 26684 10444 26740 10500
rect 27468 10498 27524 10500
rect 27468 10446 27470 10498
rect 27470 10446 27522 10498
rect 27522 10446 27524 10498
rect 27468 10444 27524 10446
rect 26796 10050 26852 10052
rect 26796 9998 26798 10050
rect 26798 9998 26850 10050
rect 26850 9998 26852 10050
rect 26796 9996 26852 9998
rect 27804 10050 27860 10052
rect 27804 9998 27806 10050
rect 27806 9998 27858 10050
rect 27858 9998 27860 10050
rect 27804 9996 27860 9998
rect 25564 8092 25620 8148
rect 26460 8370 26516 8372
rect 26460 8318 26462 8370
rect 26462 8318 26514 8370
rect 26514 8318 26516 8370
rect 26460 8316 26516 8318
rect 25788 8258 25844 8260
rect 25788 8206 25790 8258
rect 25790 8206 25842 8258
rect 25842 8206 25844 8258
rect 25788 8204 25844 8206
rect 25116 5964 25172 6020
rect 25228 6524 25284 6580
rect 24444 5906 24500 5908
rect 24444 5854 24446 5906
rect 24446 5854 24498 5906
rect 24498 5854 24500 5906
rect 24444 5852 24500 5854
rect 25452 5906 25508 5908
rect 25452 5854 25454 5906
rect 25454 5854 25506 5906
rect 25506 5854 25508 5906
rect 25452 5852 25508 5854
rect 24220 4956 24276 5012
rect 24332 4844 24388 4900
rect 23100 4172 23156 4228
rect 25228 4956 25284 5012
rect 25228 4060 25284 4116
rect 24892 3612 24948 3668
rect 26236 7474 26292 7476
rect 26236 7422 26238 7474
rect 26238 7422 26290 7474
rect 26290 7422 26292 7474
rect 26236 7420 26292 7422
rect 26236 7196 26292 7252
rect 28252 13356 28308 13412
rect 28028 13020 28084 13076
rect 28252 13132 28308 13188
rect 28588 15202 28644 15204
rect 28588 15150 28590 15202
rect 28590 15150 28642 15202
rect 28642 15150 28644 15202
rect 28588 15148 28644 15150
rect 30156 19906 30212 19908
rect 30156 19854 30158 19906
rect 30158 19854 30210 19906
rect 30210 19854 30212 19906
rect 30156 19852 30212 19854
rect 31500 20018 31556 20020
rect 31500 19966 31502 20018
rect 31502 19966 31554 20018
rect 31554 19966 31556 20018
rect 31500 19964 31556 19966
rect 32508 20300 32564 20356
rect 30828 19852 30884 19908
rect 31612 19122 31668 19124
rect 31612 19070 31614 19122
rect 31614 19070 31666 19122
rect 31666 19070 31668 19122
rect 31612 19068 31668 19070
rect 32284 19906 32340 19908
rect 32284 19854 32286 19906
rect 32286 19854 32338 19906
rect 32338 19854 32340 19906
rect 32284 19852 32340 19854
rect 30044 17052 30100 17108
rect 30716 17052 30772 17108
rect 32732 22370 32788 22372
rect 32732 22318 32734 22370
rect 32734 22318 32786 22370
rect 32786 22318 32788 22370
rect 32732 22316 32788 22318
rect 35868 50594 35924 50596
rect 35868 50542 35870 50594
rect 35870 50542 35922 50594
rect 35922 50542 35924 50594
rect 35868 50540 35924 50542
rect 35644 49980 35700 50036
rect 35532 49868 35588 49924
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 34636 48524 34692 48580
rect 34412 48242 34468 48244
rect 34412 48190 34414 48242
rect 34414 48190 34466 48242
rect 34466 48190 34468 48242
rect 34412 48188 34468 48190
rect 33292 48130 33348 48132
rect 33292 48078 33294 48130
rect 33294 48078 33346 48130
rect 33346 48078 33348 48130
rect 33292 48076 33348 48078
rect 33964 47570 34020 47572
rect 33964 47518 33966 47570
rect 33966 47518 34018 47570
rect 34018 47518 34020 47570
rect 33964 47516 34020 47518
rect 33068 46786 33124 46788
rect 33068 46734 33070 46786
rect 33070 46734 33122 46786
rect 33122 46734 33124 46786
rect 33068 46732 33124 46734
rect 33740 46786 33796 46788
rect 33740 46734 33742 46786
rect 33742 46734 33794 46786
rect 33794 46734 33796 46786
rect 33740 46732 33796 46734
rect 33404 46674 33460 46676
rect 33404 46622 33406 46674
rect 33406 46622 33458 46674
rect 33458 46622 33460 46674
rect 33404 46620 33460 46622
rect 33292 46060 33348 46116
rect 33740 44994 33796 44996
rect 33740 44942 33742 44994
rect 33742 44942 33794 44994
rect 33794 44942 33796 44994
rect 33740 44940 33796 44942
rect 33068 44604 33124 44660
rect 33628 43708 33684 43764
rect 33180 43260 33236 43316
rect 33068 41858 33124 41860
rect 33068 41806 33070 41858
rect 33070 41806 33122 41858
rect 33122 41806 33124 41858
rect 33068 41804 33124 41806
rect 33628 41858 33684 41860
rect 33628 41806 33630 41858
rect 33630 41806 33682 41858
rect 33682 41806 33684 41858
rect 33628 41804 33684 41806
rect 33404 38892 33460 38948
rect 33180 38556 33236 38612
rect 33180 36652 33236 36708
rect 33516 36988 33572 37044
rect 33292 36258 33348 36260
rect 33292 36206 33294 36258
rect 33294 36206 33346 36258
rect 33346 36206 33348 36258
rect 33292 36204 33348 36206
rect 33068 36092 33124 36148
rect 33068 35644 33124 35700
rect 34412 45164 34468 45220
rect 34748 48300 34804 48356
rect 34636 44492 34692 44548
rect 34636 43708 34692 43764
rect 34300 41916 34356 41972
rect 34300 40348 34356 40404
rect 35084 48242 35140 48244
rect 35084 48190 35086 48242
rect 35086 48190 35138 48242
rect 35138 48190 35140 48242
rect 35084 48188 35140 48190
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 37100 50594 37156 50596
rect 37100 50542 37102 50594
rect 37102 50542 37154 50594
rect 37154 50542 37156 50594
rect 37100 50540 37156 50542
rect 37996 53004 38052 53060
rect 37772 51490 37828 51492
rect 37772 51438 37774 51490
rect 37774 51438 37826 51490
rect 37826 51438 37828 51490
rect 37772 51436 37828 51438
rect 37548 51378 37604 51380
rect 37548 51326 37550 51378
rect 37550 51326 37602 51378
rect 37602 51326 37604 51378
rect 37548 51324 37604 51326
rect 38220 51378 38276 51380
rect 38220 51326 38222 51378
rect 38222 51326 38274 51378
rect 38274 51326 38276 51378
rect 38220 51324 38276 51326
rect 57596 56082 57652 56084
rect 57596 56030 57598 56082
rect 57598 56030 57650 56082
rect 57650 56030 57652 56082
rect 57596 56028 57652 56030
rect 58156 56082 58212 56084
rect 58156 56030 58158 56082
rect 58158 56030 58210 56082
rect 58210 56030 58212 56082
rect 58156 56028 58212 56030
rect 40236 55410 40292 55412
rect 40236 55358 40238 55410
rect 40238 55358 40290 55410
rect 40290 55358 40292 55410
rect 40236 55356 40292 55358
rect 41804 55356 41860 55412
rect 40684 55186 40740 55188
rect 40684 55134 40686 55186
rect 40686 55134 40738 55186
rect 40738 55134 40740 55186
rect 40684 55132 40740 55134
rect 40236 54738 40292 54740
rect 40236 54686 40238 54738
rect 40238 54686 40290 54738
rect 40290 54686 40292 54738
rect 40236 54684 40292 54686
rect 40124 54626 40180 54628
rect 40124 54574 40126 54626
rect 40126 54574 40178 54626
rect 40178 54574 40180 54626
rect 40124 54572 40180 54574
rect 39116 53842 39172 53844
rect 39116 53790 39118 53842
rect 39118 53790 39170 53842
rect 39170 53790 39172 53842
rect 39116 53788 39172 53790
rect 40012 53842 40068 53844
rect 40012 53790 40014 53842
rect 40014 53790 40066 53842
rect 40066 53790 40068 53842
rect 40012 53788 40068 53790
rect 39228 52892 39284 52948
rect 38780 52668 38836 52724
rect 41244 55298 41300 55300
rect 41244 55246 41246 55298
rect 41246 55246 41298 55298
rect 41298 55246 41300 55298
rect 41244 55244 41300 55246
rect 41020 54684 41076 54740
rect 42364 55298 42420 55300
rect 42364 55246 42366 55298
rect 42366 55246 42418 55298
rect 42418 55246 42420 55298
rect 42364 55244 42420 55246
rect 40908 54572 40964 54628
rect 42140 54626 42196 54628
rect 42140 54574 42142 54626
rect 42142 54574 42194 54626
rect 42194 54574 42196 54626
rect 42140 54572 42196 54574
rect 40796 53676 40852 53732
rect 41244 53900 41300 53956
rect 40012 53452 40068 53508
rect 40796 53506 40852 53508
rect 40796 53454 40798 53506
rect 40798 53454 40850 53506
rect 40850 53454 40852 53506
rect 40796 53452 40852 53454
rect 37100 50034 37156 50036
rect 37100 49982 37102 50034
rect 37102 49982 37154 50034
rect 37154 49982 37156 50034
rect 37100 49980 37156 49982
rect 36652 49586 36708 49588
rect 36652 49534 36654 49586
rect 36654 49534 36706 49586
rect 36706 49534 36708 49586
rect 36652 49532 36708 49534
rect 36204 48354 36260 48356
rect 36204 48302 36206 48354
rect 36206 48302 36258 48354
rect 36258 48302 36260 48354
rect 36204 48300 36260 48302
rect 36316 48412 36372 48468
rect 36092 47516 36148 47572
rect 36316 47346 36372 47348
rect 36316 47294 36318 47346
rect 36318 47294 36370 47346
rect 36370 47294 36372 47346
rect 36316 47292 36372 47294
rect 37212 48412 37268 48468
rect 37436 49532 37492 49588
rect 38444 51212 38500 51268
rect 37660 49922 37716 49924
rect 37660 49870 37662 49922
rect 37662 49870 37714 49922
rect 37714 49870 37716 49922
rect 37660 49868 37716 49870
rect 37548 49196 37604 49252
rect 37100 48076 37156 48132
rect 37212 48188 37268 48244
rect 37548 48076 37604 48132
rect 37884 47964 37940 48020
rect 37436 47068 37492 47124
rect 37100 46956 37156 47012
rect 37212 46844 37268 46900
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 37324 46284 37380 46340
rect 36204 45948 36260 46004
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 36316 43596 36372 43652
rect 35084 43372 35140 43428
rect 34076 39228 34132 39284
rect 34524 39228 34580 39284
rect 33964 38780 34020 38836
rect 34636 38108 34692 38164
rect 34860 38946 34916 38948
rect 34860 38894 34862 38946
rect 34862 38894 34914 38946
rect 34914 38894 34916 38946
rect 34860 38892 34916 38894
rect 34748 38780 34804 38836
rect 34188 37996 34244 38052
rect 33964 36258 34020 36260
rect 33964 36206 33966 36258
rect 33966 36206 34018 36258
rect 34018 36206 34020 36258
rect 33964 36204 34020 36206
rect 33852 36092 33908 36148
rect 33180 34860 33236 34916
rect 33292 34690 33348 34692
rect 33292 34638 33294 34690
rect 33294 34638 33346 34690
rect 33346 34638 33348 34690
rect 33292 34636 33348 34638
rect 33180 34300 33236 34356
rect 33292 33516 33348 33572
rect 33180 33068 33236 33124
rect 33852 33068 33908 33124
rect 33180 31218 33236 31220
rect 33180 31166 33182 31218
rect 33182 31166 33234 31218
rect 33234 31166 33236 31218
rect 33180 31164 33236 31166
rect 33180 30268 33236 30324
rect 33292 27858 33348 27860
rect 33292 27806 33294 27858
rect 33294 27806 33346 27858
rect 33346 27806 33348 27858
rect 33292 27804 33348 27806
rect 33068 27132 33124 27188
rect 33180 24220 33236 24276
rect 33180 23660 33236 23716
rect 33068 23324 33124 23380
rect 33180 23042 33236 23044
rect 33180 22990 33182 23042
rect 33182 22990 33234 23042
rect 33234 22990 33236 23042
rect 33180 22988 33236 22990
rect 33068 22652 33124 22708
rect 33180 22764 33236 22820
rect 34636 37772 34692 37828
rect 34300 36540 34356 36596
rect 34412 35196 34468 35252
rect 34412 34412 34468 34468
rect 34972 36316 35028 36372
rect 34300 33906 34356 33908
rect 34300 33854 34302 33906
rect 34302 33854 34354 33906
rect 34354 33854 34356 33906
rect 34300 33852 34356 33854
rect 34188 32956 34244 33012
rect 34972 35196 35028 35252
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 36428 42866 36484 42868
rect 36428 42814 36430 42866
rect 36430 42814 36482 42866
rect 36482 42814 36484 42866
rect 36428 42812 36484 42814
rect 35420 42140 35476 42196
rect 35308 41970 35364 41972
rect 35308 41918 35310 41970
rect 35310 41918 35362 41970
rect 35362 41918 35364 41970
rect 35308 41916 35364 41918
rect 35868 41804 35924 41860
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35756 40402 35812 40404
rect 35756 40350 35758 40402
rect 35758 40350 35810 40402
rect 35810 40350 35812 40402
rect 35756 40348 35812 40350
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 36428 41020 36484 41076
rect 37100 46002 37156 46004
rect 37100 45950 37102 46002
rect 37102 45950 37154 46002
rect 37154 45950 37156 46002
rect 37100 45948 37156 45950
rect 37212 41970 37268 41972
rect 37212 41918 37214 41970
rect 37214 41918 37266 41970
rect 37266 41918 37268 41970
rect 37212 41916 37268 41918
rect 38108 47068 38164 47124
rect 38332 48188 38388 48244
rect 38332 47852 38388 47908
rect 40348 50316 40404 50372
rect 38556 49756 38612 49812
rect 39676 49308 39732 49364
rect 39116 49250 39172 49252
rect 39116 49198 39118 49250
rect 39118 49198 39170 49250
rect 39170 49198 39172 49250
rect 39116 49196 39172 49198
rect 39564 49026 39620 49028
rect 39564 48974 39566 49026
rect 39566 48974 39618 49026
rect 39618 48974 39620 49026
rect 39564 48972 39620 48974
rect 40348 49026 40404 49028
rect 40348 48974 40350 49026
rect 40350 48974 40402 49026
rect 40402 48974 40404 49026
rect 40348 48972 40404 48974
rect 38556 48914 38612 48916
rect 38556 48862 38558 48914
rect 38558 48862 38610 48914
rect 38610 48862 38612 48914
rect 38556 48860 38612 48862
rect 39788 48802 39844 48804
rect 39788 48750 39790 48802
rect 39790 48750 39842 48802
rect 39842 48750 39844 48802
rect 39788 48748 39844 48750
rect 38444 46620 38500 46676
rect 38780 48636 38836 48692
rect 38668 47570 38724 47572
rect 38668 47518 38670 47570
rect 38670 47518 38722 47570
rect 38722 47518 38724 47570
rect 38668 47516 38724 47518
rect 38220 46284 38276 46340
rect 39676 48242 39732 48244
rect 39676 48190 39678 48242
rect 39678 48190 39730 48242
rect 39730 48190 39732 48242
rect 39676 48188 39732 48190
rect 39340 48130 39396 48132
rect 39340 48078 39342 48130
rect 39342 48078 39394 48130
rect 39394 48078 39396 48130
rect 39340 48076 39396 48078
rect 39228 46844 39284 46900
rect 40124 48524 40180 48580
rect 40348 48242 40404 48244
rect 40348 48190 40350 48242
rect 40350 48190 40402 48242
rect 40402 48190 40404 48242
rect 40348 48188 40404 48190
rect 40236 48018 40292 48020
rect 40236 47966 40238 48018
rect 40238 47966 40290 48018
rect 40290 47966 40292 48018
rect 40236 47964 40292 47966
rect 39900 46956 39956 47012
rect 41244 53676 41300 53732
rect 41132 52946 41188 52948
rect 41132 52894 41134 52946
rect 41134 52894 41186 52946
rect 41186 52894 41188 52946
rect 41132 52892 41188 52894
rect 41692 53788 41748 53844
rect 41356 52946 41412 52948
rect 41356 52894 41358 52946
rect 41358 52894 41410 52946
rect 41410 52894 41412 52946
rect 41356 52892 41412 52894
rect 41468 52722 41524 52724
rect 41468 52670 41470 52722
rect 41470 52670 41522 52722
rect 41522 52670 41524 52722
rect 41468 52668 41524 52670
rect 42140 53506 42196 53508
rect 42140 53454 42142 53506
rect 42142 53454 42194 53506
rect 42194 53454 42196 53506
rect 42140 53452 42196 53454
rect 42252 51884 42308 51940
rect 42252 51212 42308 51268
rect 41244 50316 41300 50372
rect 40908 49810 40964 49812
rect 40908 49758 40910 49810
rect 40910 49758 40962 49810
rect 40962 49758 40964 49810
rect 40908 49756 40964 49758
rect 41132 49810 41188 49812
rect 41132 49758 41134 49810
rect 41134 49758 41186 49810
rect 41186 49758 41188 49810
rect 41132 49756 41188 49758
rect 40572 48802 40628 48804
rect 40572 48750 40574 48802
rect 40574 48750 40626 48802
rect 40626 48750 40628 48802
rect 40572 48748 40628 48750
rect 40796 49026 40852 49028
rect 40796 48974 40798 49026
rect 40798 48974 40850 49026
rect 40850 48974 40852 49026
rect 40796 48972 40852 48974
rect 41804 49308 41860 49364
rect 41468 48802 41524 48804
rect 41468 48750 41470 48802
rect 41470 48750 41522 48802
rect 41522 48750 41524 48802
rect 41468 48748 41524 48750
rect 40684 48300 40740 48356
rect 42588 53900 42644 53956
rect 42476 52892 42532 52948
rect 45500 55244 45556 55300
rect 46060 55298 46116 55300
rect 46060 55246 46062 55298
rect 46062 55246 46114 55298
rect 46114 55246 46116 55298
rect 46060 55244 46116 55246
rect 46732 54684 46788 54740
rect 47404 54738 47460 54740
rect 47404 54686 47406 54738
rect 47406 54686 47458 54738
rect 47458 54686 47460 54738
rect 47404 54684 47460 54686
rect 43484 54348 43540 54404
rect 43036 53452 43092 53508
rect 44716 54402 44772 54404
rect 44716 54350 44718 54402
rect 44718 54350 44770 54402
rect 44770 54350 44772 54402
rect 44716 54348 44772 54350
rect 46508 53452 46564 53508
rect 43372 52892 43428 52948
rect 45052 53116 45108 53172
rect 43036 52332 43092 52388
rect 43708 52386 43764 52388
rect 43708 52334 43710 52386
rect 43710 52334 43762 52386
rect 43762 52334 43764 52386
rect 43708 52332 43764 52334
rect 47628 54514 47684 54516
rect 47628 54462 47630 54514
rect 47630 54462 47682 54514
rect 47682 54462 47684 54514
rect 47628 54460 47684 54462
rect 46732 53170 46788 53172
rect 46732 53118 46734 53170
rect 46734 53118 46786 53170
rect 46786 53118 46788 53170
rect 46732 53116 46788 53118
rect 45276 52892 45332 52948
rect 46284 52892 46340 52948
rect 45948 52386 46004 52388
rect 45948 52334 45950 52386
rect 45950 52334 46002 52386
rect 46002 52334 46004 52386
rect 45948 52332 46004 52334
rect 46956 52946 47012 52948
rect 46956 52894 46958 52946
rect 46958 52894 47010 52946
rect 47010 52894 47012 52946
rect 46956 52892 47012 52894
rect 42700 51884 42756 51940
rect 43260 51266 43316 51268
rect 43260 51214 43262 51266
rect 43262 51214 43314 51266
rect 43314 51214 43316 51266
rect 43260 51212 43316 51214
rect 42364 48972 42420 49028
rect 46844 51884 46900 51940
rect 48300 54402 48356 54404
rect 48300 54350 48302 54402
rect 48302 54350 48354 54402
rect 48354 54350 48356 54402
rect 48300 54348 48356 54350
rect 49308 55298 49364 55300
rect 49308 55246 49310 55298
rect 49310 55246 49362 55298
rect 49362 55246 49364 55298
rect 49308 55244 49364 55246
rect 51996 55244 52052 55300
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 48748 53506 48804 53508
rect 48748 53454 48750 53506
rect 48750 53454 48802 53506
rect 48802 53454 48804 53506
rect 48748 53452 48804 53454
rect 48076 53116 48132 53172
rect 48188 52220 48244 52276
rect 48412 52162 48468 52164
rect 48412 52110 48414 52162
rect 48414 52110 48466 52162
rect 48466 52110 48468 52162
rect 48412 52108 48468 52110
rect 49644 53452 49700 53508
rect 48860 52220 48916 52276
rect 45500 51212 45556 51268
rect 46172 51100 46228 51156
rect 46508 51100 46564 51156
rect 46060 49420 46116 49476
rect 46956 49420 47012 49476
rect 41244 48018 41300 48020
rect 41244 47966 41246 48018
rect 41246 47966 41298 48018
rect 41298 47966 41300 48018
rect 41244 47964 41300 47966
rect 42364 48802 42420 48804
rect 42364 48750 42366 48802
rect 42366 48750 42418 48802
rect 42418 48750 42420 48802
rect 42364 48748 42420 48750
rect 42700 48748 42756 48804
rect 42476 48300 42532 48356
rect 43596 48972 43652 49028
rect 43372 48914 43428 48916
rect 43372 48862 43374 48914
rect 43374 48862 43426 48914
rect 43426 48862 43428 48914
rect 43372 48860 43428 48862
rect 45388 49026 45444 49028
rect 45388 48974 45390 49026
rect 45390 48974 45442 49026
rect 45442 48974 45444 49026
rect 45388 48972 45444 48974
rect 44044 48860 44100 48916
rect 43260 48242 43316 48244
rect 43260 48190 43262 48242
rect 43262 48190 43314 48242
rect 43314 48190 43316 48242
rect 43260 48188 43316 48190
rect 43036 47852 43092 47908
rect 41132 46786 41188 46788
rect 41132 46734 41134 46786
rect 41134 46734 41186 46786
rect 41186 46734 41188 46786
rect 41132 46732 41188 46734
rect 41580 46674 41636 46676
rect 41580 46622 41582 46674
rect 41582 46622 41634 46674
rect 41634 46622 41636 46674
rect 41580 46620 41636 46622
rect 43820 48242 43876 48244
rect 43820 48190 43822 48242
rect 43822 48190 43874 48242
rect 43874 48190 43876 48242
rect 43820 48188 43876 48190
rect 44268 48636 44324 48692
rect 44268 48130 44324 48132
rect 44268 48078 44270 48130
rect 44270 48078 44322 48130
rect 44322 48078 44324 48130
rect 44268 48076 44324 48078
rect 43596 47346 43652 47348
rect 43596 47294 43598 47346
rect 43598 47294 43650 47346
rect 43650 47294 43652 47346
rect 43596 47292 43652 47294
rect 40460 45948 40516 46004
rect 37548 43484 37604 43540
rect 37772 44434 37828 44436
rect 37772 44382 37774 44434
rect 37774 44382 37826 44434
rect 37826 44382 37828 44434
rect 37772 44380 37828 44382
rect 40572 45276 40628 45332
rect 40124 45218 40180 45220
rect 40124 45166 40126 45218
rect 40126 45166 40178 45218
rect 40178 45166 40180 45218
rect 40124 45164 40180 45166
rect 39564 44380 39620 44436
rect 38220 43650 38276 43652
rect 38220 43598 38222 43650
rect 38222 43598 38274 43650
rect 38274 43598 38276 43650
rect 38220 43596 38276 43598
rect 38444 43596 38500 43652
rect 37660 42812 37716 42868
rect 38108 42924 38164 42980
rect 39340 43650 39396 43652
rect 39340 43598 39342 43650
rect 39342 43598 39394 43650
rect 39394 43598 39396 43650
rect 39340 43596 39396 43598
rect 40908 45164 40964 45220
rect 40572 44156 40628 44212
rect 37660 42364 37716 42420
rect 37884 42530 37940 42532
rect 37884 42478 37886 42530
rect 37886 42478 37938 42530
rect 37938 42478 37940 42530
rect 37884 42476 37940 42478
rect 37772 42140 37828 42196
rect 38556 43538 38612 43540
rect 38556 43486 38558 43538
rect 38558 43486 38610 43538
rect 38610 43486 38612 43538
rect 38556 43484 38612 43486
rect 38668 42530 38724 42532
rect 38668 42478 38670 42530
rect 38670 42478 38722 42530
rect 38722 42478 38724 42530
rect 38668 42476 38724 42478
rect 38332 42364 38388 42420
rect 37996 41970 38052 41972
rect 37996 41918 37998 41970
rect 37998 41918 38050 41970
rect 38050 41918 38052 41970
rect 37996 41916 38052 41918
rect 39004 42924 39060 42980
rect 39004 42140 39060 42196
rect 39564 42252 39620 42308
rect 37772 41692 37828 41748
rect 37324 41244 37380 41300
rect 37100 41074 37156 41076
rect 37100 41022 37102 41074
rect 37102 41022 37154 41074
rect 37154 41022 37156 41074
rect 37100 41020 37156 41022
rect 37324 40348 37380 40404
rect 36988 39900 37044 39956
rect 35308 39340 35364 39396
rect 36316 39394 36372 39396
rect 36316 39342 36318 39394
rect 36318 39342 36370 39394
rect 36370 39342 36372 39394
rect 36316 39340 36372 39342
rect 35756 39004 35812 39060
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35644 38050 35700 38052
rect 35644 37998 35646 38050
rect 35646 37998 35698 38050
rect 35698 37998 35700 38050
rect 35644 37996 35700 37998
rect 35532 37436 35588 37492
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35644 37212 35700 37268
rect 36652 39228 36708 39284
rect 36652 39004 36708 39060
rect 36316 38050 36372 38052
rect 36316 37998 36318 38050
rect 36318 37998 36370 38050
rect 36370 37998 36372 38050
rect 36316 37996 36372 37998
rect 35756 36540 35812 36596
rect 35980 37548 36036 37604
rect 36204 37266 36260 37268
rect 36204 37214 36206 37266
rect 36206 37214 36258 37266
rect 36258 37214 36260 37266
rect 36204 37212 36260 37214
rect 36428 37212 36484 37268
rect 35868 36988 35924 37044
rect 36316 37100 36372 37156
rect 36316 36540 36372 36596
rect 35196 36316 35252 36372
rect 35644 36370 35700 36372
rect 35644 36318 35646 36370
rect 35646 36318 35698 36370
rect 35698 36318 35700 36370
rect 35644 36316 35700 36318
rect 36316 36316 36372 36372
rect 36428 35698 36484 35700
rect 36428 35646 36430 35698
rect 36430 35646 36482 35698
rect 36482 35646 36484 35698
rect 36428 35644 36484 35646
rect 36204 35420 36260 35476
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 36316 34972 36372 35028
rect 34748 34914 34804 34916
rect 34748 34862 34750 34914
rect 34750 34862 34802 34914
rect 34802 34862 34804 34914
rect 34748 34860 34804 34862
rect 34636 34354 34692 34356
rect 34636 34302 34638 34354
rect 34638 34302 34690 34354
rect 34690 34302 34692 34354
rect 34636 34300 34692 34302
rect 34748 34636 34804 34692
rect 34524 32844 34580 32900
rect 34636 33852 34692 33908
rect 34188 32786 34244 32788
rect 34188 32734 34190 32786
rect 34190 32734 34242 32786
rect 34242 32734 34244 32786
rect 34188 32732 34244 32734
rect 34412 31890 34468 31892
rect 34412 31838 34414 31890
rect 34414 31838 34466 31890
rect 34466 31838 34468 31890
rect 34412 31836 34468 31838
rect 34636 31724 34692 31780
rect 34860 34076 34916 34132
rect 33852 31106 33908 31108
rect 33852 31054 33854 31106
rect 33854 31054 33906 31106
rect 33906 31054 33908 31106
rect 33852 31052 33908 31054
rect 33740 30994 33796 30996
rect 33740 30942 33742 30994
rect 33742 30942 33794 30994
rect 33794 30942 33796 30994
rect 33740 30940 33796 30942
rect 33516 30268 33572 30324
rect 34524 30994 34580 30996
rect 34524 30942 34526 30994
rect 34526 30942 34578 30994
rect 34578 30942 34580 30994
rect 34524 30940 34580 30942
rect 33852 28476 33908 28532
rect 34300 28476 34356 28532
rect 34412 28364 34468 28420
rect 33740 27970 33796 27972
rect 33740 27918 33742 27970
rect 33742 27918 33794 27970
rect 33794 27918 33796 27970
rect 33740 27916 33796 27918
rect 33516 27858 33572 27860
rect 33516 27806 33518 27858
rect 33518 27806 33570 27858
rect 33570 27806 33572 27858
rect 33516 27804 33572 27806
rect 33740 27580 33796 27636
rect 34860 31276 34916 31332
rect 34860 31106 34916 31108
rect 34860 31054 34862 31106
rect 34862 31054 34914 31106
rect 34914 31054 34916 31106
rect 34860 31052 34916 31054
rect 34860 30156 34916 30212
rect 34636 27580 34692 27636
rect 35084 34690 35140 34692
rect 35084 34638 35086 34690
rect 35086 34638 35138 34690
rect 35138 34638 35140 34690
rect 35084 34636 35140 34638
rect 35084 34300 35140 34356
rect 36092 34354 36148 34356
rect 36092 34302 36094 34354
rect 36094 34302 36146 34354
rect 36146 34302 36148 34354
rect 36092 34300 36148 34302
rect 35084 34130 35140 34132
rect 35084 34078 35086 34130
rect 35086 34078 35138 34130
rect 35138 34078 35140 34130
rect 35084 34076 35140 34078
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35532 33516 35588 33572
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 32002 35252 32004
rect 35196 31950 35198 32002
rect 35198 31950 35250 32002
rect 35250 31950 35252 32002
rect 35196 31948 35252 31950
rect 35084 31836 35140 31892
rect 35420 31724 35476 31780
rect 35868 34076 35924 34132
rect 35532 31218 35588 31220
rect 35532 31166 35534 31218
rect 35534 31166 35586 31218
rect 35586 31166 35588 31218
rect 35532 31164 35588 31166
rect 34748 27186 34804 27188
rect 34748 27134 34750 27186
rect 34750 27134 34802 27186
rect 34802 27134 34804 27186
rect 34748 27132 34804 27134
rect 34860 26962 34916 26964
rect 34860 26910 34862 26962
rect 34862 26910 34914 26962
rect 34914 26910 34916 26962
rect 34860 26908 34916 26910
rect 33740 23154 33796 23156
rect 33740 23102 33742 23154
rect 33742 23102 33794 23154
rect 33794 23102 33796 23154
rect 33740 23100 33796 23102
rect 33740 22316 33796 22372
rect 33404 22204 33460 22260
rect 33068 20076 33124 20132
rect 32956 19852 33012 19908
rect 34636 21420 34692 21476
rect 32956 19292 33012 19348
rect 34300 20076 34356 20132
rect 32172 18562 32228 18564
rect 32172 18510 32174 18562
rect 32174 18510 32226 18562
rect 32226 18510 32228 18562
rect 32172 18508 32228 18510
rect 32060 18284 32116 18340
rect 32172 17778 32228 17780
rect 32172 17726 32174 17778
rect 32174 17726 32226 17778
rect 32226 17726 32228 17778
rect 32172 17724 32228 17726
rect 32620 19068 32676 19124
rect 29596 16716 29652 16772
rect 30828 16770 30884 16772
rect 30828 16718 30830 16770
rect 30830 16718 30882 16770
rect 30882 16718 30884 16770
rect 30828 16716 30884 16718
rect 28924 15426 28980 15428
rect 28924 15374 28926 15426
rect 28926 15374 28978 15426
rect 28978 15374 28980 15426
rect 28924 15372 28980 15374
rect 28700 15036 28756 15092
rect 30828 15596 30884 15652
rect 29596 15036 29652 15092
rect 28476 13746 28532 13748
rect 28476 13694 28478 13746
rect 28478 13694 28530 13746
rect 28530 13694 28532 13746
rect 28476 13692 28532 13694
rect 28588 12962 28644 12964
rect 28588 12910 28590 12962
rect 28590 12910 28642 12962
rect 28642 12910 28644 12962
rect 28588 12908 28644 12910
rect 28140 10610 28196 10612
rect 28140 10558 28142 10610
rect 28142 10558 28194 10610
rect 28194 10558 28196 10610
rect 28140 10556 28196 10558
rect 32732 18284 32788 18340
rect 32620 16940 32676 16996
rect 29596 13468 29652 13524
rect 31164 15596 31220 15652
rect 29820 13074 29876 13076
rect 29820 13022 29822 13074
rect 29822 13022 29874 13074
rect 29874 13022 29876 13074
rect 29820 13020 29876 13022
rect 30156 12962 30212 12964
rect 30156 12910 30158 12962
rect 30158 12910 30210 12962
rect 30210 12910 30212 12962
rect 30156 12908 30212 12910
rect 30828 13186 30884 13188
rect 30828 13134 30830 13186
rect 30830 13134 30882 13186
rect 30882 13134 30884 13186
rect 30828 13132 30884 13134
rect 30716 12962 30772 12964
rect 30716 12910 30718 12962
rect 30718 12910 30770 12962
rect 30770 12910 30772 12962
rect 30716 12908 30772 12910
rect 31388 15260 31444 15316
rect 29708 12796 29764 12852
rect 30380 12850 30436 12852
rect 30380 12798 30382 12850
rect 30382 12798 30434 12850
rect 30434 12798 30436 12850
rect 30380 12796 30436 12798
rect 30828 12850 30884 12852
rect 30828 12798 30830 12850
rect 30830 12798 30882 12850
rect 30882 12798 30884 12850
rect 30828 12796 30884 12798
rect 31164 11394 31220 11396
rect 31164 11342 31166 11394
rect 31166 11342 31218 11394
rect 31218 11342 31220 11394
rect 31164 11340 31220 11342
rect 29372 10610 29428 10612
rect 29372 10558 29374 10610
rect 29374 10558 29426 10610
rect 29426 10558 29428 10610
rect 29372 10556 29428 10558
rect 30604 10444 30660 10500
rect 28140 9548 28196 9604
rect 27916 9436 27972 9492
rect 28588 9436 28644 9492
rect 26684 6972 26740 7028
rect 26460 6860 26516 6916
rect 25788 5964 25844 6020
rect 25788 5682 25844 5684
rect 25788 5630 25790 5682
rect 25790 5630 25842 5682
rect 25842 5630 25844 5682
rect 25788 5628 25844 5630
rect 26236 5964 26292 6020
rect 27132 7308 27188 7364
rect 27356 6972 27412 7028
rect 27580 6860 27636 6916
rect 26684 5628 26740 5684
rect 26572 5122 26628 5124
rect 26572 5070 26574 5122
rect 26574 5070 26626 5122
rect 26626 5070 26628 5122
rect 26572 5068 26628 5070
rect 26908 4172 26964 4228
rect 28140 4226 28196 4228
rect 28140 4174 28142 4226
rect 28142 4174 28194 4226
rect 28194 4174 28196 4226
rect 28140 4172 28196 4174
rect 25676 3724 25732 3780
rect 26124 3666 26180 3668
rect 26124 3614 26126 3666
rect 26126 3614 26178 3666
rect 26178 3614 26180 3666
rect 26124 3612 26180 3614
rect 29148 9548 29204 9604
rect 30044 9826 30100 9828
rect 30044 9774 30046 9826
rect 30046 9774 30098 9826
rect 30098 9774 30100 9826
rect 30044 9772 30100 9774
rect 29820 9660 29876 9716
rect 30380 9266 30436 9268
rect 30380 9214 30382 9266
rect 30382 9214 30434 9266
rect 30434 9214 30436 9266
rect 30380 9212 30436 9214
rect 28812 8316 28868 8372
rect 29484 7980 29540 8036
rect 30268 8034 30324 8036
rect 30268 7982 30270 8034
rect 30270 7982 30322 8034
rect 30322 7982 30324 8034
rect 30268 7980 30324 7982
rect 30044 7868 30100 7924
rect 29708 7362 29764 7364
rect 29708 7310 29710 7362
rect 29710 7310 29762 7362
rect 29762 7310 29764 7362
rect 29708 7308 29764 7310
rect 29820 7250 29876 7252
rect 29820 7198 29822 7250
rect 29822 7198 29874 7250
rect 29874 7198 29876 7250
rect 29820 7196 29876 7198
rect 30828 9772 30884 9828
rect 30716 9714 30772 9716
rect 30716 9662 30718 9714
rect 30718 9662 30770 9714
rect 30770 9662 30772 9714
rect 30716 9660 30772 9662
rect 31500 15148 31556 15204
rect 31948 15148 32004 15204
rect 32508 15202 32564 15204
rect 32508 15150 32510 15202
rect 32510 15150 32562 15202
rect 32562 15150 32564 15202
rect 32508 15148 32564 15150
rect 31836 13132 31892 13188
rect 31612 12962 31668 12964
rect 31612 12910 31614 12962
rect 31614 12910 31666 12962
rect 31666 12910 31668 12962
rect 31612 12908 31668 12910
rect 33628 18562 33684 18564
rect 33628 18510 33630 18562
rect 33630 18510 33682 18562
rect 33682 18510 33684 18562
rect 33628 18508 33684 18510
rect 33516 18450 33572 18452
rect 33516 18398 33518 18450
rect 33518 18398 33570 18450
rect 33570 18398 33572 18450
rect 33516 18396 33572 18398
rect 33180 17724 33236 17780
rect 34748 19122 34804 19124
rect 34748 19070 34750 19122
rect 34750 19070 34802 19122
rect 34802 19070 34804 19122
rect 34748 19068 34804 19070
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35084 28476 35140 28532
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35980 33516 36036 33572
rect 36540 33404 36596 33460
rect 36092 33292 36148 33348
rect 35980 31106 36036 31108
rect 35980 31054 35982 31106
rect 35982 31054 36034 31106
rect 36034 31054 36036 31106
rect 35980 31052 36036 31054
rect 37212 39058 37268 39060
rect 37212 39006 37214 39058
rect 37214 39006 37266 39058
rect 37266 39006 37268 39058
rect 37212 39004 37268 39006
rect 36988 38780 37044 38836
rect 38556 41692 38612 41748
rect 39116 40124 39172 40180
rect 38556 39900 38612 39956
rect 36876 37996 36932 38052
rect 37884 39058 37940 39060
rect 37884 39006 37886 39058
rect 37886 39006 37938 39058
rect 37938 39006 37940 39058
rect 37884 39004 37940 39006
rect 37884 38780 37940 38836
rect 37548 38220 37604 38276
rect 38668 39116 38724 39172
rect 37548 37548 37604 37604
rect 38108 37772 38164 37828
rect 38108 37548 38164 37604
rect 37100 37266 37156 37268
rect 37100 37214 37102 37266
rect 37102 37214 37154 37266
rect 37154 37214 37156 37266
rect 37100 37212 37156 37214
rect 36876 37100 36932 37156
rect 38220 37100 38276 37156
rect 37436 36204 37492 36260
rect 36764 34076 36820 34132
rect 36988 33852 37044 33908
rect 37100 33516 37156 33572
rect 36652 31164 36708 31220
rect 36316 30210 36372 30212
rect 36316 30158 36318 30210
rect 36318 30158 36370 30210
rect 36370 30158 36372 30210
rect 36316 30156 36372 30158
rect 36652 30940 36708 30996
rect 36988 29596 37044 29652
rect 36428 27916 36484 27972
rect 36652 28476 36708 28532
rect 36540 27804 36596 27860
rect 37212 33292 37268 33348
rect 37324 31836 37380 31892
rect 37660 35084 37716 35140
rect 37772 35026 37828 35028
rect 37772 34974 37774 35026
rect 37774 34974 37826 35026
rect 37826 34974 37828 35026
rect 37772 34972 37828 34974
rect 37660 33852 37716 33908
rect 37996 35420 38052 35476
rect 37884 33516 37940 33572
rect 38668 36876 38724 36932
rect 38444 35756 38500 35812
rect 39004 35698 39060 35700
rect 39004 35646 39006 35698
rect 39006 35646 39058 35698
rect 39058 35646 39060 35698
rect 39004 35644 39060 35646
rect 38892 35474 38948 35476
rect 38892 35422 38894 35474
rect 38894 35422 38946 35474
rect 38946 35422 38948 35474
rect 38892 35420 38948 35422
rect 38444 33516 38500 33572
rect 39228 38834 39284 38836
rect 39228 38782 39230 38834
rect 39230 38782 39282 38834
rect 39282 38782 39284 38834
rect 39228 38780 39284 38782
rect 40348 40796 40404 40852
rect 39900 40236 39956 40292
rect 40908 41298 40964 41300
rect 40908 41246 40910 41298
rect 40910 41246 40962 41298
rect 40962 41246 40964 41298
rect 40908 41244 40964 41246
rect 40908 40796 40964 40852
rect 40236 38780 40292 38836
rect 39788 37772 39844 37828
rect 40012 36876 40068 36932
rect 39452 35756 39508 35812
rect 39676 35698 39732 35700
rect 39676 35646 39678 35698
rect 39678 35646 39730 35698
rect 39730 35646 39732 35698
rect 39676 35644 39732 35646
rect 39228 33906 39284 33908
rect 39228 33854 39230 33906
rect 39230 33854 39282 33906
rect 39282 33854 39284 33906
rect 39228 33852 39284 33854
rect 38108 33404 38164 33460
rect 38444 33346 38500 33348
rect 38444 33294 38446 33346
rect 38446 33294 38498 33346
rect 38498 33294 38500 33346
rect 38444 33292 38500 33294
rect 38108 33122 38164 33124
rect 38108 33070 38110 33122
rect 38110 33070 38162 33122
rect 38162 33070 38164 33122
rect 38108 33068 38164 33070
rect 37548 31948 37604 32004
rect 38556 32732 38612 32788
rect 37324 30940 37380 30996
rect 37100 28364 37156 28420
rect 36540 27020 36596 27076
rect 35980 26684 36036 26740
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35980 24780 36036 24836
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35532 24108 35588 24164
rect 35308 23826 35364 23828
rect 35308 23774 35310 23826
rect 35310 23774 35362 23826
rect 35362 23774 35364 23826
rect 35308 23772 35364 23774
rect 35308 23324 35364 23380
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 36092 23884 36148 23940
rect 36204 24556 36260 24612
rect 35980 23324 36036 23380
rect 36652 26178 36708 26180
rect 36652 26126 36654 26178
rect 36654 26126 36706 26178
rect 36706 26126 36708 26178
rect 36652 26124 36708 26126
rect 36428 26012 36484 26068
rect 36428 23660 36484 23716
rect 37100 27074 37156 27076
rect 37100 27022 37102 27074
rect 37102 27022 37154 27074
rect 37154 27022 37156 27074
rect 37100 27020 37156 27022
rect 37436 30044 37492 30100
rect 37436 29650 37492 29652
rect 37436 29598 37438 29650
rect 37438 29598 37490 29650
rect 37490 29598 37492 29650
rect 37436 29596 37492 29598
rect 37324 27916 37380 27972
rect 38220 30156 38276 30212
rect 37772 29036 37828 29092
rect 37548 27634 37604 27636
rect 37548 27582 37550 27634
rect 37550 27582 37602 27634
rect 37602 27582 37604 27634
rect 37548 27580 37604 27582
rect 37996 29596 38052 29652
rect 40012 32732 40068 32788
rect 40460 39116 40516 39172
rect 40460 35026 40516 35028
rect 40460 34974 40462 35026
rect 40462 34974 40514 35026
rect 40514 34974 40516 35026
rect 40460 34972 40516 34974
rect 41916 45276 41972 45332
rect 43148 45948 43204 46004
rect 43036 44940 43092 44996
rect 42812 44322 42868 44324
rect 42812 44270 42814 44322
rect 42814 44270 42866 44322
rect 42866 44270 42868 44322
rect 42812 44268 42868 44270
rect 43484 45724 43540 45780
rect 43820 44994 43876 44996
rect 43820 44942 43822 44994
rect 43822 44942 43874 44994
rect 43874 44942 43876 44994
rect 43820 44940 43876 44942
rect 43148 44156 43204 44212
rect 42476 44098 42532 44100
rect 42476 44046 42478 44098
rect 42478 44046 42530 44098
rect 42530 44046 42532 44098
rect 42476 44044 42532 44046
rect 42588 43484 42644 43540
rect 42588 43260 42644 43316
rect 40908 40290 40964 40292
rect 40908 40238 40910 40290
rect 40910 40238 40962 40290
rect 40962 40238 40964 40290
rect 40908 40236 40964 40238
rect 41244 40178 41300 40180
rect 41244 40126 41246 40178
rect 41246 40126 41298 40178
rect 41298 40126 41300 40178
rect 41244 40124 41300 40126
rect 41692 40124 41748 40180
rect 43260 44044 43316 44100
rect 43820 44268 43876 44324
rect 43596 43820 43652 43876
rect 43260 43484 43316 43540
rect 43260 42700 43316 42756
rect 42364 40908 42420 40964
rect 41916 40236 41972 40292
rect 42588 40236 42644 40292
rect 41356 39564 41412 39620
rect 42140 39618 42196 39620
rect 42140 39566 42142 39618
rect 42142 39566 42194 39618
rect 42194 39566 42196 39618
rect 42140 39564 42196 39566
rect 43484 40236 43540 40292
rect 43596 42700 43652 42756
rect 44940 48242 44996 48244
rect 44940 48190 44942 48242
rect 44942 48190 44994 48242
rect 44994 48190 44996 48242
rect 44940 48188 44996 48190
rect 44492 47628 44548 47684
rect 45612 48636 45668 48692
rect 45276 48130 45332 48132
rect 45276 48078 45278 48130
rect 45278 48078 45330 48130
rect 45330 48078 45332 48130
rect 45276 48076 45332 48078
rect 46060 48466 46116 48468
rect 46060 48414 46062 48466
rect 46062 48414 46114 48466
rect 46114 48414 46116 48466
rect 46060 48412 46116 48414
rect 46172 48354 46228 48356
rect 46172 48302 46174 48354
rect 46174 48302 46226 48354
rect 46226 48302 46228 48354
rect 46172 48300 46228 48302
rect 46956 48242 47012 48244
rect 46956 48190 46958 48242
rect 46958 48190 47010 48242
rect 47010 48190 47012 48242
rect 46956 48188 47012 48190
rect 45948 48130 46004 48132
rect 45948 48078 45950 48130
rect 45950 48078 46002 48130
rect 46002 48078 46004 48130
rect 45948 48076 46004 48078
rect 45836 47516 45892 47572
rect 47180 48524 47236 48580
rect 47180 47740 47236 47796
rect 47292 48300 47348 48356
rect 46172 46674 46228 46676
rect 46172 46622 46174 46674
rect 46174 46622 46226 46674
rect 46226 46622 46228 46674
rect 46172 46620 46228 46622
rect 46620 46508 46676 46564
rect 44044 45778 44100 45780
rect 44044 45726 44046 45778
rect 44046 45726 44098 45778
rect 44098 45726 44100 45778
rect 44044 45724 44100 45726
rect 44268 45276 44324 45332
rect 45388 45276 45444 45332
rect 44044 44322 44100 44324
rect 44044 44270 44046 44322
rect 44046 44270 44098 44322
rect 44098 44270 44100 44322
rect 44044 44268 44100 44270
rect 44268 43708 44324 43764
rect 43708 41186 43764 41188
rect 43708 41134 43710 41186
rect 43710 41134 43762 41186
rect 43762 41134 43764 41186
rect 43708 41132 43764 41134
rect 43820 40962 43876 40964
rect 43820 40910 43822 40962
rect 43822 40910 43874 40962
rect 43874 40910 43876 40962
rect 43820 40908 43876 40910
rect 43820 39564 43876 39620
rect 43596 39452 43652 39508
rect 42364 39394 42420 39396
rect 42364 39342 42366 39394
rect 42366 39342 42418 39394
rect 42418 39342 42420 39394
rect 42364 39340 42420 39342
rect 43148 39394 43204 39396
rect 43148 39342 43150 39394
rect 43150 39342 43202 39394
rect 43202 39342 43204 39394
rect 43148 39340 43204 39342
rect 47068 45276 47124 45332
rect 47852 48300 47908 48356
rect 47516 48188 47572 48244
rect 49196 51996 49252 52052
rect 49532 52162 49588 52164
rect 49532 52110 49534 52162
rect 49534 52110 49586 52162
rect 49586 52110 49588 52162
rect 49532 52108 49588 52110
rect 49420 51884 49476 51940
rect 48972 49868 49028 49924
rect 49196 50652 49252 50708
rect 50876 53730 50932 53732
rect 50876 53678 50878 53730
rect 50878 53678 50930 53730
rect 50930 53678 50932 53730
rect 50876 53676 50932 53678
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 49980 53058 50036 53060
rect 49980 53006 49982 53058
rect 49982 53006 50034 53058
rect 50034 53006 50036 53058
rect 49980 53004 50036 53006
rect 50092 52946 50148 52948
rect 50092 52894 50094 52946
rect 50094 52894 50146 52946
rect 50146 52894 50148 52946
rect 50092 52892 50148 52894
rect 49308 49532 49364 49588
rect 48076 48354 48132 48356
rect 48076 48302 48078 48354
rect 48078 48302 48130 48354
rect 48130 48302 48132 48354
rect 48076 48300 48132 48302
rect 50316 52050 50372 52052
rect 50316 51998 50318 52050
rect 50318 51998 50370 52050
rect 50370 51998 50372 52050
rect 50316 51996 50372 51998
rect 50540 51884 50596 51940
rect 50092 50818 50148 50820
rect 50092 50766 50094 50818
rect 50094 50766 50146 50818
rect 50146 50766 50148 50818
rect 50092 50764 50148 50766
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 49980 50652 50036 50708
rect 50652 50652 50708 50708
rect 50764 51324 50820 51380
rect 50204 49922 50260 49924
rect 50204 49870 50206 49922
rect 50206 49870 50258 49922
rect 50258 49870 50260 49922
rect 50204 49868 50260 49870
rect 51660 53004 51716 53060
rect 50764 50428 50820 50484
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 51212 50764 51268 50820
rect 51548 50428 51604 50484
rect 50988 50204 51044 50260
rect 51548 49532 51604 49588
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 49532 48300 49588 48356
rect 49868 47292 49924 47348
rect 49644 46450 49700 46452
rect 49644 46398 49646 46450
rect 49646 46398 49698 46450
rect 49698 46398 49700 46450
rect 49644 46396 49700 46398
rect 49420 45612 49476 45668
rect 48188 44940 48244 44996
rect 44716 43426 44772 43428
rect 44716 43374 44718 43426
rect 44718 43374 44770 43426
rect 44770 43374 44772 43426
rect 44716 43372 44772 43374
rect 47068 44268 47124 44324
rect 45500 43372 45556 43428
rect 49084 44994 49140 44996
rect 49084 44942 49086 44994
rect 49086 44942 49138 44994
rect 49138 44942 49140 44994
rect 49084 44940 49140 44942
rect 50652 47516 50708 47572
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 50316 46674 50372 46676
rect 50316 46622 50318 46674
rect 50318 46622 50370 46674
rect 50370 46622 50372 46674
rect 50316 46620 50372 46622
rect 49868 45388 49924 45444
rect 50540 46620 50596 46676
rect 50540 45666 50596 45668
rect 50540 45614 50542 45666
rect 50542 45614 50594 45666
rect 50594 45614 50596 45666
rect 50540 45612 50596 45614
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 49756 44434 49812 44436
rect 49756 44382 49758 44434
rect 49758 44382 49810 44434
rect 49810 44382 49812 44434
rect 49756 44380 49812 44382
rect 49420 43484 49476 43540
rect 46732 42978 46788 42980
rect 46732 42926 46734 42978
rect 46734 42926 46786 42978
rect 46786 42926 46788 42978
rect 46732 42924 46788 42926
rect 49420 42924 49476 42980
rect 45500 42588 45556 42644
rect 44940 42476 44996 42532
rect 44828 42194 44884 42196
rect 44828 42142 44830 42194
rect 44830 42142 44882 42194
rect 44882 42142 44884 42194
rect 44828 42140 44884 42142
rect 44380 42028 44436 42084
rect 44492 41132 44548 41188
rect 45276 42194 45332 42196
rect 45276 42142 45278 42194
rect 45278 42142 45330 42194
rect 45330 42142 45332 42194
rect 45276 42140 45332 42142
rect 46172 42642 46228 42644
rect 46172 42590 46174 42642
rect 46174 42590 46226 42642
rect 46226 42590 46228 42642
rect 46172 42588 46228 42590
rect 45164 42082 45220 42084
rect 45164 42030 45166 42082
rect 45166 42030 45218 42082
rect 45218 42030 45220 42082
rect 45164 42028 45220 42030
rect 44156 40012 44212 40068
rect 43932 39004 43988 39060
rect 43596 38108 43652 38164
rect 43708 38444 43764 38500
rect 42028 37548 42084 37604
rect 43484 37324 43540 37380
rect 41580 36316 41636 36372
rect 41244 35138 41300 35140
rect 41244 35086 41246 35138
rect 41246 35086 41298 35138
rect 41298 35086 41300 35138
rect 41244 35084 41300 35086
rect 41580 35644 41636 35700
rect 41692 35084 41748 35140
rect 40348 31164 40404 31220
rect 40460 32060 40516 32116
rect 40348 30940 40404 30996
rect 39452 30268 39508 30324
rect 39340 30210 39396 30212
rect 39340 30158 39342 30210
rect 39342 30158 39394 30210
rect 39394 30158 39396 30210
rect 39340 30156 39396 30158
rect 39900 29932 39956 29988
rect 37100 26514 37156 26516
rect 37100 26462 37102 26514
rect 37102 26462 37154 26514
rect 37154 26462 37156 26514
rect 37100 26460 37156 26462
rect 37436 26124 37492 26180
rect 37324 26012 37380 26068
rect 36876 23826 36932 23828
rect 36876 23774 36878 23826
rect 36878 23774 36930 23826
rect 36930 23774 36932 23826
rect 36876 23772 36932 23774
rect 36876 23100 36932 23156
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 34524 18396 34580 18452
rect 35084 20748 35140 20804
rect 33852 18172 33908 18228
rect 33404 15148 33460 15204
rect 34076 15148 34132 15204
rect 33516 14364 33572 14420
rect 33068 13132 33124 13188
rect 34412 13692 34468 13748
rect 34300 13468 34356 13524
rect 33852 12962 33908 12964
rect 33852 12910 33854 12962
rect 33854 12910 33906 12962
rect 33906 12910 33908 12962
rect 33852 12908 33908 12910
rect 34636 12962 34692 12964
rect 34636 12910 34638 12962
rect 34638 12910 34690 12962
rect 34690 12910 34692 12962
rect 34636 12908 34692 12910
rect 33516 12796 33572 12852
rect 35980 20748 36036 20804
rect 35756 20636 35812 20692
rect 36540 21586 36596 21588
rect 36540 21534 36542 21586
rect 36542 21534 36594 21586
rect 36594 21534 36596 21586
rect 36540 21532 36596 21534
rect 36652 21474 36708 21476
rect 36652 21422 36654 21474
rect 36654 21422 36706 21474
rect 36706 21422 36708 21474
rect 36652 21420 36708 21422
rect 35980 20300 36036 20356
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35084 18338 35140 18340
rect 35084 18286 35086 18338
rect 35086 18286 35138 18338
rect 35138 18286 35140 18338
rect 35084 18284 35140 18286
rect 34972 18172 35028 18228
rect 35532 18172 35588 18228
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 36092 18284 36148 18340
rect 36204 17778 36260 17780
rect 36204 17726 36206 17778
rect 36206 17726 36258 17778
rect 36258 17726 36260 17778
rect 36204 17724 36260 17726
rect 35980 16044 36036 16100
rect 36428 15986 36484 15988
rect 36428 15934 36430 15986
rect 36430 15934 36482 15986
rect 36482 15934 36484 15986
rect 36428 15932 36484 15934
rect 36092 15820 36148 15876
rect 35308 15372 35364 15428
rect 35532 15260 35588 15316
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 34972 14306 35028 14308
rect 34972 14254 34974 14306
rect 34974 14254 35026 14306
rect 35026 14254 35028 14306
rect 34972 14252 35028 14254
rect 34860 13804 34916 13860
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 36316 15708 36372 15764
rect 35644 13804 35700 13860
rect 35532 12908 35588 12964
rect 35756 13468 35812 13524
rect 35980 13746 36036 13748
rect 35980 13694 35982 13746
rect 35982 13694 36034 13746
rect 36034 13694 36036 13746
rect 35980 13692 36036 13694
rect 34748 12684 34804 12740
rect 34636 11340 34692 11396
rect 35196 11900 35252 11956
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 36204 14306 36260 14308
rect 36204 14254 36206 14306
rect 36206 14254 36258 14306
rect 36258 14254 36260 14306
rect 36204 14252 36260 14254
rect 36204 13468 36260 13524
rect 36092 13020 36148 13076
rect 36652 15314 36708 15316
rect 36652 15262 36654 15314
rect 36654 15262 36706 15314
rect 36706 15262 36708 15314
rect 36652 15260 36708 15262
rect 37212 23714 37268 23716
rect 37212 23662 37214 23714
rect 37214 23662 37266 23714
rect 37266 23662 37268 23714
rect 37212 23660 37268 23662
rect 37212 23324 37268 23380
rect 37436 23938 37492 23940
rect 37436 23886 37438 23938
rect 37438 23886 37490 23938
rect 37490 23886 37492 23938
rect 37436 23884 37492 23886
rect 37100 21308 37156 21364
rect 37100 20524 37156 20580
rect 37436 21698 37492 21700
rect 37436 21646 37438 21698
rect 37438 21646 37490 21698
rect 37490 21646 37492 21698
rect 37436 21644 37492 21646
rect 37324 21532 37380 21588
rect 37884 26348 37940 26404
rect 37884 25618 37940 25620
rect 37884 25566 37886 25618
rect 37886 25566 37938 25618
rect 37938 25566 37940 25618
rect 37884 25564 37940 25566
rect 38556 27916 38612 27972
rect 38108 26514 38164 26516
rect 38108 26462 38110 26514
rect 38110 26462 38162 26514
rect 38162 26462 38164 26514
rect 38108 26460 38164 26462
rect 38108 25004 38164 25060
rect 39116 27634 39172 27636
rect 39116 27582 39118 27634
rect 39118 27582 39170 27634
rect 39170 27582 39172 27634
rect 39116 27580 39172 27582
rect 38556 26178 38612 26180
rect 38556 26126 38558 26178
rect 38558 26126 38610 26178
rect 38610 26126 38612 26178
rect 38556 26124 38612 26126
rect 39228 26796 39284 26852
rect 39004 26514 39060 26516
rect 39004 26462 39006 26514
rect 39006 26462 39058 26514
rect 39058 26462 39060 26514
rect 39004 26460 39060 26462
rect 38556 25228 38612 25284
rect 39564 25228 39620 25284
rect 38220 24892 38276 24948
rect 39116 25004 39172 25060
rect 37996 24834 38052 24836
rect 37996 24782 37998 24834
rect 37998 24782 38050 24834
rect 38050 24782 38052 24834
rect 37996 24780 38052 24782
rect 38332 24780 38388 24836
rect 37772 24668 37828 24724
rect 38668 24668 38724 24724
rect 38220 24556 38276 24612
rect 38108 23884 38164 23940
rect 38444 23436 38500 23492
rect 37996 21644 38052 21700
rect 37436 19740 37492 19796
rect 37324 19404 37380 19460
rect 37660 21362 37716 21364
rect 37660 21310 37662 21362
rect 37662 21310 37714 21362
rect 37714 21310 37716 21362
rect 37660 21308 37716 21310
rect 37884 20524 37940 20580
rect 37100 19068 37156 19124
rect 37212 18172 37268 18228
rect 37996 19404 38052 19460
rect 38668 23660 38724 23716
rect 38780 21810 38836 21812
rect 38780 21758 38782 21810
rect 38782 21758 38834 21810
rect 38834 21758 38836 21810
rect 38780 21756 38836 21758
rect 39340 24722 39396 24724
rect 39340 24670 39342 24722
rect 39342 24670 39394 24722
rect 39394 24670 39396 24722
rect 39340 24668 39396 24670
rect 39340 22428 39396 22484
rect 39116 21532 39172 21588
rect 38892 21420 38948 21476
rect 39228 20860 39284 20916
rect 39340 20578 39396 20580
rect 39340 20526 39342 20578
rect 39342 20526 39394 20578
rect 39394 20526 39396 20578
rect 39340 20524 39396 20526
rect 38444 19180 38500 19236
rect 38556 19404 38612 19460
rect 37996 19122 38052 19124
rect 37996 19070 37998 19122
rect 37998 19070 38050 19122
rect 38050 19070 38052 19122
rect 37996 19068 38052 19070
rect 38444 19010 38500 19012
rect 38444 18958 38446 19010
rect 38446 18958 38498 19010
rect 38498 18958 38500 19010
rect 38444 18956 38500 18958
rect 38332 18844 38388 18900
rect 37548 18172 37604 18228
rect 37660 16828 37716 16884
rect 35868 10780 35924 10836
rect 30604 7868 30660 7924
rect 30940 9714 30996 9716
rect 30940 9662 30942 9714
rect 30942 9662 30994 9714
rect 30994 9662 30996 9714
rect 30940 9660 30996 9662
rect 31388 9212 31444 9268
rect 31724 10444 31780 10500
rect 30380 7362 30436 7364
rect 30380 7310 30382 7362
rect 30382 7310 30434 7362
rect 30434 7310 30436 7362
rect 30380 7308 30436 7310
rect 32284 10498 32340 10500
rect 32284 10446 32286 10498
rect 32286 10446 32338 10498
rect 32338 10446 32340 10498
rect 32284 10444 32340 10446
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 33964 9714 34020 9716
rect 33964 9662 33966 9714
rect 33966 9662 34018 9714
rect 34018 9662 34020 9714
rect 33964 9660 34020 9662
rect 36988 14642 37044 14644
rect 36988 14590 36990 14642
rect 36990 14590 37042 14642
rect 37042 14590 37044 14642
rect 36988 14588 37044 14590
rect 37548 16044 37604 16100
rect 37100 13074 37156 13076
rect 37100 13022 37102 13074
rect 37102 13022 37154 13074
rect 37154 13022 37156 13074
rect 37100 13020 37156 13022
rect 36988 11900 37044 11956
rect 33292 8930 33348 8932
rect 33292 8878 33294 8930
rect 33294 8878 33346 8930
rect 33346 8878 33348 8930
rect 33292 8876 33348 8878
rect 33964 8258 34020 8260
rect 33964 8206 33966 8258
rect 33966 8206 34018 8258
rect 34018 8206 34020 8258
rect 33964 8204 34020 8206
rect 30828 7474 30884 7476
rect 30828 7422 30830 7474
rect 30830 7422 30882 7474
rect 30882 7422 30884 7474
rect 30828 7420 30884 7422
rect 31612 7474 31668 7476
rect 31612 7422 31614 7474
rect 31614 7422 31666 7474
rect 31666 7422 31668 7474
rect 31612 7420 31668 7422
rect 31164 7362 31220 7364
rect 31164 7310 31166 7362
rect 31166 7310 31218 7362
rect 31218 7310 31220 7362
rect 31164 7308 31220 7310
rect 30716 6972 30772 7028
rect 29708 5122 29764 5124
rect 29708 5070 29710 5122
rect 29710 5070 29762 5122
rect 29762 5070 29764 5122
rect 29708 5068 29764 5070
rect 30380 5068 30436 5124
rect 29260 4956 29316 5012
rect 34300 8876 34356 8932
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 34748 8258 34804 8260
rect 34748 8206 34750 8258
rect 34750 8206 34802 8258
rect 34802 8206 34804 8258
rect 34748 8204 34804 8206
rect 33852 7308 33908 7364
rect 34972 7868 35028 7924
rect 31836 6972 31892 7028
rect 33740 6972 33796 7028
rect 33516 6690 33572 6692
rect 33516 6638 33518 6690
rect 33518 6638 33570 6690
rect 33570 6638 33572 6690
rect 33516 6636 33572 6638
rect 34636 6748 34692 6804
rect 34636 6300 34692 6356
rect 33292 4562 33348 4564
rect 33292 4510 33294 4562
rect 33294 4510 33346 4562
rect 33346 4510 33348 4562
rect 33292 4508 33348 4510
rect 34972 6300 35028 6356
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35308 6860 35364 6916
rect 35980 6860 36036 6916
rect 35196 6300 35252 6356
rect 37660 15932 37716 15988
rect 37996 18284 38052 18340
rect 37884 17724 37940 17780
rect 38556 18562 38612 18564
rect 38556 18510 38558 18562
rect 38558 18510 38610 18562
rect 38610 18510 38612 18562
rect 38556 18508 38612 18510
rect 39116 18338 39172 18340
rect 39116 18286 39118 18338
rect 39118 18286 39170 18338
rect 39170 18286 39172 18338
rect 39116 18284 39172 18286
rect 38332 16098 38388 16100
rect 38332 16046 38334 16098
rect 38334 16046 38386 16098
rect 38386 16046 38388 16098
rect 38332 16044 38388 16046
rect 37772 15820 37828 15876
rect 38108 15874 38164 15876
rect 38108 15822 38110 15874
rect 38110 15822 38162 15874
rect 38162 15822 38164 15874
rect 38108 15820 38164 15822
rect 38444 15708 38500 15764
rect 37884 14588 37940 14644
rect 37996 14364 38052 14420
rect 37884 13186 37940 13188
rect 37884 13134 37886 13186
rect 37886 13134 37938 13186
rect 37938 13134 37940 13186
rect 37884 13132 37940 13134
rect 39116 13132 39172 13188
rect 37660 13074 37716 13076
rect 37660 13022 37662 13074
rect 37662 13022 37714 13074
rect 37714 13022 37716 13074
rect 37660 13020 37716 13022
rect 38668 13074 38724 13076
rect 38668 13022 38670 13074
rect 38670 13022 38722 13074
rect 38722 13022 38724 13074
rect 38668 13020 38724 13022
rect 37996 12124 38052 12180
rect 38220 11788 38276 11844
rect 38220 11116 38276 11172
rect 37436 10834 37492 10836
rect 37436 10782 37438 10834
rect 37438 10782 37490 10834
rect 37490 10782 37492 10834
rect 37436 10780 37492 10782
rect 39004 11116 39060 11172
rect 37324 10556 37380 10612
rect 37996 10556 38052 10612
rect 37660 9826 37716 9828
rect 37660 9774 37662 9826
rect 37662 9774 37714 9826
rect 37714 9774 37716 9826
rect 37660 9772 37716 9774
rect 39116 9884 39172 9940
rect 39228 11900 39284 11956
rect 39340 10610 39396 10612
rect 39340 10558 39342 10610
rect 39342 10558 39394 10610
rect 39394 10558 39396 10610
rect 39340 10556 39396 10558
rect 39228 9826 39284 9828
rect 39228 9774 39230 9826
rect 39230 9774 39282 9826
rect 39282 9774 39284 9826
rect 39228 9772 39284 9774
rect 39676 24892 39732 24948
rect 40348 25228 40404 25284
rect 40124 25004 40180 25060
rect 39900 24722 39956 24724
rect 39900 24670 39902 24722
rect 39902 24670 39954 24722
rect 39954 24670 39956 24722
rect 39900 24668 39956 24670
rect 39676 21756 39732 21812
rect 39788 21474 39844 21476
rect 39788 21422 39790 21474
rect 39790 21422 39842 21474
rect 39842 21422 39844 21474
rect 39788 21420 39844 21422
rect 39788 20914 39844 20916
rect 39788 20862 39790 20914
rect 39790 20862 39842 20914
rect 39842 20862 39844 20914
rect 39788 20860 39844 20862
rect 39900 14530 39956 14532
rect 39900 14478 39902 14530
rect 39902 14478 39954 14530
rect 39954 14478 39956 14530
rect 39900 14476 39956 14478
rect 40124 22764 40180 22820
rect 40124 22482 40180 22484
rect 40124 22430 40126 22482
rect 40126 22430 40178 22482
rect 40178 22430 40180 22482
rect 40124 22428 40180 22430
rect 40908 32060 40964 32116
rect 41804 34748 41860 34804
rect 41244 33068 41300 33124
rect 41356 33404 41412 33460
rect 41916 33458 41972 33460
rect 41916 33406 41918 33458
rect 41918 33406 41970 33458
rect 41970 33406 41972 33458
rect 41916 33404 41972 33406
rect 41468 32450 41524 32452
rect 41468 32398 41470 32450
rect 41470 32398 41522 32450
rect 41522 32398 41524 32450
rect 41468 32396 41524 32398
rect 41132 31724 41188 31780
rect 41580 31612 41636 31668
rect 40460 19852 40516 19908
rect 40348 18956 40404 19012
rect 40012 13356 40068 13412
rect 40124 18284 40180 18340
rect 40236 14476 40292 14532
rect 40460 18620 40516 18676
rect 40684 31164 40740 31220
rect 41356 31218 41412 31220
rect 41356 31166 41358 31218
rect 41358 31166 41410 31218
rect 41410 31166 41412 31218
rect 41356 31164 41412 31166
rect 42140 35698 42196 35700
rect 42140 35646 42142 35698
rect 42142 35646 42194 35698
rect 42194 35646 42196 35698
rect 42140 35644 42196 35646
rect 42364 35532 42420 35588
rect 42140 34972 42196 35028
rect 42364 34802 42420 34804
rect 42364 34750 42366 34802
rect 42366 34750 42418 34802
rect 42418 34750 42420 34802
rect 42364 34748 42420 34750
rect 42252 34690 42308 34692
rect 42252 34638 42254 34690
rect 42254 34638 42306 34690
rect 42306 34638 42308 34690
rect 42252 34636 42308 34638
rect 42028 33346 42084 33348
rect 42028 33294 42030 33346
rect 42030 33294 42082 33346
rect 42082 33294 42084 33346
rect 42028 33292 42084 33294
rect 42140 34524 42196 34580
rect 43372 36594 43428 36596
rect 43372 36542 43374 36594
rect 43374 36542 43426 36594
rect 43426 36542 43428 36594
rect 43372 36540 43428 36542
rect 42700 36316 42756 36372
rect 42588 35586 42644 35588
rect 42588 35534 42590 35586
rect 42590 35534 42642 35586
rect 42642 35534 42644 35586
rect 42588 35532 42644 35534
rect 42588 34802 42644 34804
rect 42588 34750 42590 34802
rect 42590 34750 42642 34802
rect 42642 34750 42644 34802
rect 42588 34748 42644 34750
rect 43036 36258 43092 36260
rect 43036 36206 43038 36258
rect 43038 36206 43090 36258
rect 43090 36206 43092 36258
rect 43036 36204 43092 36206
rect 43372 35532 43428 35588
rect 42588 34524 42644 34580
rect 41804 31890 41860 31892
rect 41804 31838 41806 31890
rect 41806 31838 41858 31890
rect 41858 31838 41860 31890
rect 41804 31836 41860 31838
rect 41132 30994 41188 30996
rect 41132 30942 41134 30994
rect 41134 30942 41186 30994
rect 41186 30942 41188 30994
rect 41132 30940 41188 30942
rect 40908 30828 40964 30884
rect 41468 30268 41524 30324
rect 40796 29986 40852 29988
rect 40796 29934 40798 29986
rect 40798 29934 40850 29986
rect 40850 29934 40852 29986
rect 40796 29932 40852 29934
rect 42028 28754 42084 28756
rect 42028 28702 42030 28754
rect 42030 28702 42082 28754
rect 42082 28702 42084 28754
rect 42028 28700 42084 28702
rect 41692 27746 41748 27748
rect 41692 27694 41694 27746
rect 41694 27694 41746 27746
rect 41746 27694 41748 27746
rect 41692 27692 41748 27694
rect 41020 26796 41076 26852
rect 40908 25004 40964 25060
rect 40796 24892 40852 24948
rect 41468 25228 41524 25284
rect 41132 23826 41188 23828
rect 41132 23774 41134 23826
rect 41134 23774 41186 23826
rect 41186 23774 41188 23826
rect 41132 23772 41188 23774
rect 40908 21756 40964 21812
rect 40684 20860 40740 20916
rect 41468 24444 41524 24500
rect 41692 23772 41748 23828
rect 41580 22428 41636 22484
rect 42476 33234 42532 33236
rect 42476 33182 42478 33234
rect 42478 33182 42530 33234
rect 42530 33182 42532 33234
rect 42476 33180 42532 33182
rect 42700 33292 42756 33348
rect 42588 32450 42644 32452
rect 42588 32398 42590 32450
rect 42590 32398 42642 32450
rect 42642 32398 42644 32450
rect 42588 32396 42644 32398
rect 42364 31724 42420 31780
rect 42588 31218 42644 31220
rect 42588 31166 42590 31218
rect 42590 31166 42642 31218
rect 42642 31166 42644 31218
rect 42588 31164 42644 31166
rect 42700 31612 42756 31668
rect 42476 30882 42532 30884
rect 42476 30830 42478 30882
rect 42478 30830 42530 30882
rect 42530 30830 42532 30882
rect 42476 30828 42532 30830
rect 42812 28700 42868 28756
rect 43260 34914 43316 34916
rect 43260 34862 43262 34914
rect 43262 34862 43314 34914
rect 43314 34862 43316 34914
rect 43260 34860 43316 34862
rect 43148 34636 43204 34692
rect 42588 27580 42644 27636
rect 42476 21644 42532 21700
rect 41356 21586 41412 21588
rect 41356 21534 41358 21586
rect 41358 21534 41410 21586
rect 41410 21534 41412 21586
rect 41356 21532 41412 21534
rect 41020 18956 41076 19012
rect 40684 18396 40740 18452
rect 41020 17724 41076 17780
rect 41692 18450 41748 18452
rect 41692 18398 41694 18450
rect 41694 18398 41746 18450
rect 41746 18398 41748 18450
rect 41692 18396 41748 18398
rect 41916 20130 41972 20132
rect 41916 20078 41918 20130
rect 41918 20078 41970 20130
rect 41970 20078 41972 20130
rect 41916 20076 41972 20078
rect 42364 20130 42420 20132
rect 42364 20078 42366 20130
rect 42366 20078 42418 20130
rect 42418 20078 42420 20130
rect 42364 20076 42420 20078
rect 42588 19740 42644 19796
rect 42140 19346 42196 19348
rect 42140 19294 42142 19346
rect 42142 19294 42194 19346
rect 42194 19294 42196 19346
rect 42140 19292 42196 19294
rect 41916 18620 41972 18676
rect 42252 18620 42308 18676
rect 42924 25394 42980 25396
rect 42924 25342 42926 25394
rect 42926 25342 42978 25394
rect 42978 25342 42980 25394
rect 42924 25340 42980 25342
rect 42924 21474 42980 21476
rect 42924 21422 42926 21474
rect 42926 21422 42978 21474
rect 42978 21422 42980 21474
rect 42924 21420 42980 21422
rect 43484 28754 43540 28756
rect 43484 28702 43486 28754
rect 43486 28702 43538 28754
rect 43538 28702 43540 28754
rect 43484 28700 43540 28702
rect 43932 38780 43988 38836
rect 43820 38332 43876 38388
rect 44268 38162 44324 38164
rect 44268 38110 44270 38162
rect 44270 38110 44322 38162
rect 44322 38110 44324 38162
rect 44268 38108 44324 38110
rect 43820 37324 43876 37380
rect 45724 40908 45780 40964
rect 46060 40402 46116 40404
rect 46060 40350 46062 40402
rect 46062 40350 46114 40402
rect 46114 40350 46116 40402
rect 46060 40348 46116 40350
rect 46284 40290 46340 40292
rect 46284 40238 46286 40290
rect 46286 40238 46338 40290
rect 46338 40238 46340 40290
rect 46284 40236 46340 40238
rect 46620 40236 46676 40292
rect 45388 39788 45444 39844
rect 45724 38834 45780 38836
rect 45724 38782 45726 38834
rect 45726 38782 45778 38834
rect 45778 38782 45780 38834
rect 45724 38780 45780 38782
rect 49756 42700 49812 42756
rect 47964 42082 48020 42084
rect 47964 42030 47966 42082
rect 47966 42030 48018 42082
rect 48018 42030 48020 42082
rect 47964 42028 48020 42030
rect 46956 40236 47012 40292
rect 47516 41804 47572 41860
rect 46620 38892 46676 38948
rect 46844 39004 46900 39060
rect 45052 38332 45108 38388
rect 46284 38834 46340 38836
rect 46284 38782 46286 38834
rect 46286 38782 46338 38834
rect 46338 38782 46340 38834
rect 46284 38780 46340 38782
rect 45948 37772 46004 37828
rect 44716 36540 44772 36596
rect 44828 36652 44884 36708
rect 44940 36428 44996 36484
rect 43820 36204 43876 36260
rect 43932 34860 43988 34916
rect 44716 33180 44772 33236
rect 44716 32450 44772 32452
rect 44716 32398 44718 32450
rect 44718 32398 44770 32450
rect 44770 32398 44772 32450
rect 44716 32396 44772 32398
rect 45276 35532 45332 35588
rect 48972 41970 49028 41972
rect 48972 41918 48974 41970
rect 48974 41918 49026 41970
rect 49026 41918 49028 41970
rect 48972 41916 49028 41918
rect 48076 41746 48132 41748
rect 48076 41694 48078 41746
rect 48078 41694 48130 41746
rect 48130 41694 48132 41746
rect 48076 41692 48132 41694
rect 49084 41692 49140 41748
rect 48748 40962 48804 40964
rect 48748 40910 48750 40962
rect 48750 40910 48802 40962
rect 48802 40910 48804 40962
rect 48748 40908 48804 40910
rect 49308 40908 49364 40964
rect 47516 40348 47572 40404
rect 48748 39788 48804 39844
rect 47852 39228 47908 39284
rect 47516 38892 47572 38948
rect 47740 38722 47796 38724
rect 47740 38670 47742 38722
rect 47742 38670 47794 38722
rect 47794 38670 47796 38722
rect 47740 38668 47796 38670
rect 47404 38444 47460 38500
rect 47180 37772 47236 37828
rect 48748 39228 48804 39284
rect 49756 40236 49812 40292
rect 50204 44268 50260 44324
rect 50316 45276 50372 45332
rect 50092 43596 50148 43652
rect 50876 45276 50932 45332
rect 50988 45164 51044 45220
rect 51100 47570 51156 47572
rect 51100 47518 51102 47570
rect 51102 47518 51154 47570
rect 51154 47518 51156 47570
rect 51100 47516 51156 47518
rect 50428 44380 50484 44436
rect 49980 39788 50036 39844
rect 50092 40460 50148 40516
rect 49420 39394 49476 39396
rect 49420 39342 49422 39394
rect 49422 39342 49474 39394
rect 49474 39342 49476 39394
rect 49420 39340 49476 39342
rect 47964 38444 48020 38500
rect 48860 38834 48916 38836
rect 48860 38782 48862 38834
rect 48862 38782 48914 38834
rect 48914 38782 48916 38834
rect 48860 38780 48916 38782
rect 49084 39004 49140 39060
rect 48188 37436 48244 37492
rect 48748 38050 48804 38052
rect 48748 37998 48750 38050
rect 48750 37998 48802 38050
rect 48802 37998 48804 38050
rect 48748 37996 48804 37998
rect 48300 37100 48356 37156
rect 46284 36316 46340 36372
rect 46844 36370 46900 36372
rect 46844 36318 46846 36370
rect 46846 36318 46898 36370
rect 46898 36318 46900 36370
rect 46844 36316 46900 36318
rect 47180 36204 47236 36260
rect 47516 35698 47572 35700
rect 47516 35646 47518 35698
rect 47518 35646 47570 35698
rect 47570 35646 47572 35698
rect 47516 35644 47572 35646
rect 47852 35308 47908 35364
rect 46844 35084 46900 35140
rect 44940 33180 44996 33236
rect 44380 31778 44436 31780
rect 44380 31726 44382 31778
rect 44382 31726 44434 31778
rect 44434 31726 44436 31778
rect 44380 31724 44436 31726
rect 45836 31836 45892 31892
rect 46060 34748 46116 34804
rect 47068 33740 47124 33796
rect 46620 33180 46676 33236
rect 46508 32060 46564 32116
rect 45612 30882 45668 30884
rect 45612 30830 45614 30882
rect 45614 30830 45666 30882
rect 45666 30830 45668 30882
rect 45612 30828 45668 30830
rect 46060 30828 46116 30884
rect 45612 30268 45668 30324
rect 43708 28028 43764 28084
rect 44044 28812 44100 28868
rect 44604 29202 44660 29204
rect 44604 29150 44606 29202
rect 44606 29150 44658 29202
rect 44658 29150 44660 29202
rect 44604 29148 44660 29150
rect 44492 28700 44548 28756
rect 44940 28700 44996 28756
rect 43708 27804 43764 27860
rect 44268 28642 44324 28644
rect 44268 28590 44270 28642
rect 44270 28590 44322 28642
rect 44322 28590 44324 28642
rect 44268 28588 44324 28590
rect 44380 27858 44436 27860
rect 44380 27806 44382 27858
rect 44382 27806 44434 27858
rect 44434 27806 44436 27858
rect 44380 27804 44436 27806
rect 45052 28252 45108 28308
rect 46060 29148 46116 29204
rect 46956 31052 47012 31108
rect 46956 30268 47012 30324
rect 46172 29036 46228 29092
rect 46396 29372 46452 29428
rect 46396 28700 46452 28756
rect 46620 29314 46676 29316
rect 46620 29262 46622 29314
rect 46622 29262 46674 29314
rect 46674 29262 46676 29314
rect 46620 29260 46676 29262
rect 46172 28418 46228 28420
rect 46172 28366 46174 28418
rect 46174 28366 46226 28418
rect 46226 28366 46228 28418
rect 46172 28364 46228 28366
rect 43372 25340 43428 25396
rect 43372 21698 43428 21700
rect 43372 21646 43374 21698
rect 43374 21646 43426 21698
rect 43426 21646 43428 21698
rect 43372 21644 43428 21646
rect 43148 20076 43204 20132
rect 42812 19852 42868 19908
rect 43148 19852 43204 19908
rect 42588 19180 42644 19236
rect 42476 18172 42532 18228
rect 41468 16882 41524 16884
rect 41468 16830 41470 16882
rect 41470 16830 41522 16882
rect 41522 16830 41524 16882
rect 41468 16828 41524 16830
rect 41804 16828 41860 16884
rect 41916 16940 41972 16996
rect 41804 16044 41860 16100
rect 40908 14530 40964 14532
rect 40908 14478 40910 14530
rect 40910 14478 40962 14530
rect 40962 14478 40964 14530
rect 40908 14476 40964 14478
rect 41692 13970 41748 13972
rect 41692 13918 41694 13970
rect 41694 13918 41746 13970
rect 41746 13918 41748 13970
rect 41692 13916 41748 13918
rect 40348 13692 40404 13748
rect 40908 13468 40964 13524
rect 40460 12460 40516 12516
rect 40012 12066 40068 12068
rect 40012 12014 40014 12066
rect 40014 12014 40066 12066
rect 40066 12014 40068 12066
rect 40012 12012 40068 12014
rect 40012 10610 40068 10612
rect 40012 10558 40014 10610
rect 40014 10558 40066 10610
rect 40066 10558 40068 10610
rect 40012 10556 40068 10558
rect 39452 9660 39508 9716
rect 38108 9548 38164 9604
rect 39340 9602 39396 9604
rect 39340 9550 39342 9602
rect 39342 9550 39394 9602
rect 39394 9550 39396 9602
rect 39340 9548 39396 9550
rect 39116 9436 39172 9492
rect 39564 9100 39620 9156
rect 40236 9660 40292 9716
rect 40124 9154 40180 9156
rect 40124 9102 40126 9154
rect 40126 9102 40178 9154
rect 40178 9102 40180 9154
rect 40124 9100 40180 9102
rect 40236 8818 40292 8820
rect 40236 8766 40238 8818
rect 40238 8766 40290 8818
rect 40290 8766 40292 8818
rect 40236 8764 40292 8766
rect 37324 7756 37380 7812
rect 39228 7644 39284 7700
rect 38220 7196 38276 7252
rect 36316 6188 36372 6244
rect 34412 4562 34468 4564
rect 34412 4510 34414 4562
rect 34414 4510 34466 4562
rect 34466 4510 34468 4562
rect 34412 4508 34468 4510
rect 34524 4956 34580 5012
rect 32172 4396 32228 4452
rect 33180 4450 33236 4452
rect 33180 4398 33182 4450
rect 33182 4398 33234 4450
rect 33234 4398 33236 4450
rect 33180 4396 33236 4398
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 37212 6188 37268 6244
rect 39116 7250 39172 7252
rect 39116 7198 39118 7250
rect 39118 7198 39170 7250
rect 39170 7198 39172 7250
rect 39116 7196 39172 7198
rect 37548 5906 37604 5908
rect 37548 5854 37550 5906
rect 37550 5854 37602 5906
rect 37602 5854 37604 5906
rect 37548 5852 37604 5854
rect 38556 5852 38612 5908
rect 39228 5010 39284 5012
rect 39228 4958 39230 5010
rect 39230 4958 39282 5010
rect 39282 4958 39284 5010
rect 39228 4956 39284 4958
rect 40348 8540 40404 8596
rect 39900 7698 39956 7700
rect 39900 7646 39902 7698
rect 39902 7646 39954 7698
rect 39954 7646 39956 7698
rect 39900 7644 39956 7646
rect 40908 12460 40964 12516
rect 41356 13244 41412 13300
rect 41468 13746 41524 13748
rect 41468 13694 41470 13746
rect 41470 13694 41522 13746
rect 41522 13694 41524 13746
rect 41468 13692 41524 13694
rect 41356 12572 41412 12628
rect 41356 12402 41412 12404
rect 41356 12350 41358 12402
rect 41358 12350 41410 12402
rect 41410 12350 41412 12402
rect 41356 12348 41412 12350
rect 40572 11900 40628 11956
rect 41580 12178 41636 12180
rect 41580 12126 41582 12178
rect 41582 12126 41634 12178
rect 41634 12126 41636 12178
rect 41580 12124 41636 12126
rect 41244 12066 41300 12068
rect 41244 12014 41246 12066
rect 41246 12014 41298 12066
rect 41298 12014 41300 12066
rect 41244 12012 41300 12014
rect 41132 11900 41188 11956
rect 40908 10668 40964 10724
rect 41916 13858 41972 13860
rect 41916 13806 41918 13858
rect 41918 13806 41970 13858
rect 41970 13806 41972 13858
rect 41916 13804 41972 13806
rect 42028 13244 42084 13300
rect 42140 13916 42196 13972
rect 41916 12572 41972 12628
rect 42812 15372 42868 15428
rect 42700 13916 42756 13972
rect 42140 12402 42196 12404
rect 42140 12350 42142 12402
rect 42142 12350 42194 12402
rect 42194 12350 42196 12402
rect 42140 12348 42196 12350
rect 41916 11900 41972 11956
rect 42700 13522 42756 13524
rect 42700 13470 42702 13522
rect 42702 13470 42754 13522
rect 42754 13470 42756 13522
rect 42700 13468 42756 13470
rect 42476 13244 42532 13300
rect 42364 12402 42420 12404
rect 42364 12350 42366 12402
rect 42366 12350 42418 12402
rect 42418 12350 42420 12402
rect 42364 12348 42420 12350
rect 43036 19234 43092 19236
rect 43036 19182 43038 19234
rect 43038 19182 43090 19234
rect 43090 19182 43092 19234
rect 43036 19180 43092 19182
rect 43036 18620 43092 18676
rect 43260 18396 43316 18452
rect 43260 18060 43316 18116
rect 43260 16940 43316 16996
rect 42924 12348 42980 12404
rect 42476 11900 42532 11956
rect 41580 10722 41636 10724
rect 41580 10670 41582 10722
rect 41582 10670 41634 10722
rect 41634 10670 41636 10722
rect 41580 10668 41636 10670
rect 41468 9714 41524 9716
rect 41468 9662 41470 9714
rect 41470 9662 41522 9714
rect 41522 9662 41524 9714
rect 41468 9660 41524 9662
rect 39676 7474 39732 7476
rect 39676 7422 39678 7474
rect 39678 7422 39730 7474
rect 39730 7422 39732 7474
rect 39676 7420 39732 7422
rect 40908 9436 40964 9492
rect 41244 9602 41300 9604
rect 41244 9550 41246 9602
rect 41246 9550 41298 9602
rect 41298 9550 41300 9602
rect 41244 9548 41300 9550
rect 41244 8540 41300 8596
rect 41356 8316 41412 8372
rect 42476 10780 42532 10836
rect 42924 10668 42980 10724
rect 42588 9996 42644 10052
rect 42252 9884 42308 9940
rect 43036 9100 43092 9156
rect 43484 19010 43540 19012
rect 43484 18958 43486 19010
rect 43486 18958 43538 19010
rect 43538 18958 43540 19010
rect 43484 18956 43540 18958
rect 43484 15874 43540 15876
rect 43484 15822 43486 15874
rect 43486 15822 43538 15874
rect 43538 15822 43540 15874
rect 43484 15820 43540 15822
rect 43484 13468 43540 13524
rect 43932 24444 43988 24500
rect 44268 22482 44324 22484
rect 44268 22430 44270 22482
rect 44270 22430 44322 22482
rect 44322 22430 44324 22482
rect 44268 22428 44324 22430
rect 44604 21532 44660 21588
rect 44156 20524 44212 20580
rect 43932 19010 43988 19012
rect 43932 18958 43934 19010
rect 43934 18958 43986 19010
rect 43986 18958 43988 19010
rect 43932 18956 43988 18958
rect 44940 24610 44996 24612
rect 44940 24558 44942 24610
rect 44942 24558 44994 24610
rect 44994 24558 44996 24610
rect 44940 24556 44996 24558
rect 45276 23938 45332 23940
rect 45276 23886 45278 23938
rect 45278 23886 45330 23938
rect 45330 23886 45332 23938
rect 45276 23884 45332 23886
rect 45612 27746 45668 27748
rect 45612 27694 45614 27746
rect 45614 27694 45666 27746
rect 45666 27694 45668 27746
rect 45612 27692 45668 27694
rect 46620 26290 46676 26292
rect 46620 26238 46622 26290
rect 46622 26238 46674 26290
rect 46674 26238 46676 26290
rect 46620 26236 46676 26238
rect 45948 23938 46004 23940
rect 45948 23886 45950 23938
rect 45950 23886 46002 23938
rect 46002 23886 46004 23938
rect 45948 23884 46004 23886
rect 46396 23938 46452 23940
rect 46396 23886 46398 23938
rect 46398 23886 46450 23938
rect 46450 23886 46452 23938
rect 46396 23884 46452 23886
rect 45724 23826 45780 23828
rect 45724 23774 45726 23826
rect 45726 23774 45778 23826
rect 45778 23774 45780 23826
rect 45724 23772 45780 23774
rect 46060 22988 46116 23044
rect 45388 21586 45444 21588
rect 45388 21534 45390 21586
rect 45390 21534 45442 21586
rect 45442 21534 45444 21586
rect 45388 21532 45444 21534
rect 44716 19292 44772 19348
rect 44492 19180 44548 19236
rect 44268 19010 44324 19012
rect 44268 18958 44270 19010
rect 44270 18958 44322 19010
rect 44322 18958 44324 19010
rect 44268 18956 44324 18958
rect 43820 18060 43876 18116
rect 44156 17500 44212 17556
rect 45276 18956 45332 19012
rect 47740 32562 47796 32564
rect 47740 32510 47742 32562
rect 47742 32510 47794 32562
rect 47794 32510 47796 32562
rect 47740 32508 47796 32510
rect 47740 32060 47796 32116
rect 47292 31948 47348 32004
rect 47516 31218 47572 31220
rect 47516 31166 47518 31218
rect 47518 31166 47570 31218
rect 47570 31166 47572 31218
rect 47516 31164 47572 31166
rect 47404 31106 47460 31108
rect 47404 31054 47406 31106
rect 47406 31054 47458 31106
rect 47458 31054 47460 31106
rect 47404 31052 47460 31054
rect 47180 29426 47236 29428
rect 47180 29374 47182 29426
rect 47182 29374 47234 29426
rect 47234 29374 47236 29426
rect 47180 29372 47236 29374
rect 47180 28642 47236 28644
rect 47180 28590 47182 28642
rect 47182 28590 47234 28642
rect 47234 28590 47236 28642
rect 47180 28588 47236 28590
rect 47516 29260 47572 29316
rect 47964 31500 48020 31556
rect 48188 31164 48244 31220
rect 48188 30716 48244 30772
rect 47180 27804 47236 27860
rect 47628 28252 47684 28308
rect 47740 27858 47796 27860
rect 47740 27806 47742 27858
rect 47742 27806 47794 27858
rect 47794 27806 47796 27858
rect 47740 27804 47796 27806
rect 47628 27746 47684 27748
rect 47628 27694 47630 27746
rect 47630 27694 47682 27746
rect 47682 27694 47684 27746
rect 47628 27692 47684 27694
rect 48748 37548 48804 37604
rect 48860 37490 48916 37492
rect 48860 37438 48862 37490
rect 48862 37438 48914 37490
rect 48914 37438 48916 37490
rect 48860 37436 48916 37438
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 51772 51212 51828 51268
rect 51324 44492 51380 44548
rect 51996 47180 52052 47236
rect 51548 45276 51604 45332
rect 50764 43538 50820 43540
rect 50764 43486 50766 43538
rect 50766 43486 50818 43538
rect 50818 43486 50820 43538
rect 50764 43484 50820 43486
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 51884 45164 51940 45220
rect 51772 44322 51828 44324
rect 51772 44270 51774 44322
rect 51774 44270 51826 44322
rect 51826 44270 51828 44322
rect 51772 44268 51828 44270
rect 51324 42700 51380 42756
rect 51772 42588 51828 42644
rect 50764 41804 50820 41860
rect 51548 42028 51604 42084
rect 51212 41186 51268 41188
rect 51212 41134 51214 41186
rect 51214 41134 51266 41186
rect 51266 41134 51268 41186
rect 51212 41132 51268 41134
rect 52108 46786 52164 46788
rect 52108 46734 52110 46786
rect 52110 46734 52162 46786
rect 52162 46734 52164 46786
rect 52108 46732 52164 46734
rect 52108 44492 52164 44548
rect 52668 55298 52724 55300
rect 52668 55246 52670 55298
rect 52670 55246 52722 55298
rect 52722 55246 52724 55298
rect 52668 55244 52724 55246
rect 53452 55186 53508 55188
rect 53452 55134 53454 55186
rect 53454 55134 53506 55186
rect 53506 55134 53508 55186
rect 53452 55132 53508 55134
rect 54460 55132 54516 55188
rect 54572 54460 54628 54516
rect 52892 54348 52948 54404
rect 52780 53842 52836 53844
rect 52780 53790 52782 53842
rect 52782 53790 52834 53842
rect 52834 53790 52836 53842
rect 52780 53788 52836 53790
rect 54236 53900 54292 53956
rect 53676 53788 53732 53844
rect 54348 53788 54404 53844
rect 54908 53900 54964 53956
rect 53228 53564 53284 53620
rect 54012 53618 54068 53620
rect 54012 53566 54014 53618
rect 54014 53566 54066 53618
rect 54066 53566 54068 53618
rect 54012 53564 54068 53566
rect 53004 52108 53060 52164
rect 52444 47740 52500 47796
rect 53788 51266 53844 51268
rect 53788 51214 53790 51266
rect 53790 51214 53842 51266
rect 53842 51214 53844 51266
rect 53788 51212 53844 51214
rect 55356 53900 55412 53956
rect 55020 53730 55076 53732
rect 55020 53678 55022 53730
rect 55022 53678 55074 53730
rect 55074 53678 55076 53730
rect 55020 53676 55076 53678
rect 56252 54572 56308 54628
rect 55244 53506 55300 53508
rect 55244 53454 55246 53506
rect 55246 53454 55298 53506
rect 55298 53454 55300 53506
rect 55244 53452 55300 53454
rect 54796 52946 54852 52948
rect 54796 52894 54798 52946
rect 54798 52894 54850 52946
rect 54850 52894 54852 52946
rect 54796 52892 54852 52894
rect 55244 52892 55300 52948
rect 55468 52946 55524 52948
rect 55468 52894 55470 52946
rect 55470 52894 55522 52946
rect 55522 52894 55524 52946
rect 55468 52892 55524 52894
rect 55244 52274 55300 52276
rect 55244 52222 55246 52274
rect 55246 52222 55298 52274
rect 55298 52222 55300 52274
rect 55244 52220 55300 52222
rect 55916 51884 55972 51940
rect 56140 52220 56196 52276
rect 55356 51378 55412 51380
rect 55356 51326 55358 51378
rect 55358 51326 55410 51378
rect 55410 51326 55412 51378
rect 55356 51324 55412 51326
rect 54572 50428 54628 50484
rect 55244 50428 55300 50484
rect 52556 47516 52612 47572
rect 52780 47234 52836 47236
rect 52780 47182 52782 47234
rect 52782 47182 52834 47234
rect 52834 47182 52836 47234
rect 52780 47180 52836 47182
rect 52780 46620 52836 46676
rect 52892 45500 52948 45556
rect 53004 46732 53060 46788
rect 52780 45218 52836 45220
rect 52780 45166 52782 45218
rect 52782 45166 52834 45218
rect 52834 45166 52836 45218
rect 52780 45164 52836 45166
rect 53116 46396 53172 46452
rect 52444 43596 52500 43652
rect 55804 49868 55860 49924
rect 53900 47346 53956 47348
rect 53900 47294 53902 47346
rect 53902 47294 53954 47346
rect 53954 47294 53956 47346
rect 53900 47292 53956 47294
rect 53452 45890 53508 45892
rect 53452 45838 53454 45890
rect 53454 45838 53506 45890
rect 53506 45838 53508 45890
rect 53452 45836 53508 45838
rect 53340 45724 53396 45780
rect 55580 47292 55636 47348
rect 54236 46956 54292 47012
rect 53900 45778 53956 45780
rect 53900 45726 53902 45778
rect 53902 45726 53954 45778
rect 53954 45726 53956 45778
rect 53900 45724 53956 45726
rect 55468 46786 55524 46788
rect 55468 46734 55470 46786
rect 55470 46734 55522 46786
rect 55522 46734 55524 46786
rect 55468 46732 55524 46734
rect 55692 46956 55748 47012
rect 53564 45388 53620 45444
rect 53676 45612 53732 45668
rect 54012 45500 54068 45556
rect 52892 42754 52948 42756
rect 52892 42702 52894 42754
rect 52894 42702 52946 42754
rect 52946 42702 52948 42754
rect 52892 42700 52948 42702
rect 52780 42642 52836 42644
rect 52780 42590 52782 42642
rect 52782 42590 52834 42642
rect 52834 42590 52836 42642
rect 52780 42588 52836 42590
rect 51884 41916 51940 41972
rect 51772 41858 51828 41860
rect 51772 41806 51774 41858
rect 51774 41806 51826 41858
rect 51826 41806 51828 41858
rect 51772 41804 51828 41806
rect 51660 41132 51716 41188
rect 51884 40962 51940 40964
rect 51884 40910 51886 40962
rect 51886 40910 51938 40962
rect 51938 40910 51940 40962
rect 51884 40908 51940 40910
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 50428 40348 50484 40404
rect 51884 40402 51940 40404
rect 51884 40350 51886 40402
rect 51886 40350 51938 40402
rect 51938 40350 51940 40402
rect 51884 40348 51940 40350
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 50540 38050 50596 38052
rect 50540 37998 50542 38050
rect 50542 37998 50594 38050
rect 50594 37998 50596 38050
rect 50540 37996 50596 37998
rect 52332 41132 52388 41188
rect 52332 40626 52388 40628
rect 52332 40574 52334 40626
rect 52334 40574 52386 40626
rect 52386 40574 52388 40626
rect 52332 40572 52388 40574
rect 52220 40124 52276 40180
rect 52108 39900 52164 39956
rect 52556 40908 52612 40964
rect 52668 40348 52724 40404
rect 52780 40572 52836 40628
rect 53340 41804 53396 41860
rect 53900 45052 53956 45108
rect 54348 45836 54404 45892
rect 54796 45724 54852 45780
rect 54572 45666 54628 45668
rect 54572 45614 54574 45666
rect 54574 45614 54626 45666
rect 54626 45614 54628 45666
rect 54572 45612 54628 45614
rect 54572 45388 54628 45444
rect 55244 46674 55300 46676
rect 55244 46622 55246 46674
rect 55246 46622 55298 46674
rect 55298 46622 55300 46674
rect 55244 46620 55300 46622
rect 55356 46562 55412 46564
rect 55356 46510 55358 46562
rect 55358 46510 55410 46562
rect 55410 46510 55412 46562
rect 55356 46508 55412 46510
rect 54236 45052 54292 45108
rect 55244 45164 55300 45220
rect 54908 45052 54964 45108
rect 54460 43820 54516 43876
rect 54572 43708 54628 43764
rect 55468 43820 55524 43876
rect 55132 43708 55188 43764
rect 54236 40626 54292 40628
rect 54236 40574 54238 40626
rect 54238 40574 54290 40626
rect 54290 40574 54292 40626
rect 54236 40572 54292 40574
rect 53676 40460 53732 40516
rect 52668 39676 52724 39732
rect 52668 39004 52724 39060
rect 52108 38722 52164 38724
rect 52108 38670 52110 38722
rect 52110 38670 52162 38722
rect 52162 38670 52164 38722
rect 52108 38668 52164 38670
rect 51884 37996 51940 38052
rect 49756 37548 49812 37604
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 48972 37100 49028 37156
rect 48748 36482 48804 36484
rect 48748 36430 48750 36482
rect 48750 36430 48802 36482
rect 48802 36430 48804 36482
rect 48748 36428 48804 36430
rect 48972 35810 49028 35812
rect 48972 35758 48974 35810
rect 48974 35758 49026 35810
rect 49026 35758 49028 35810
rect 48972 35756 49028 35758
rect 49644 36204 49700 36260
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 51212 35756 51268 35812
rect 49980 35308 50036 35364
rect 50204 34914 50260 34916
rect 50204 34862 50206 34914
rect 50206 34862 50258 34914
rect 50258 34862 50260 34914
rect 50204 34860 50260 34862
rect 50764 34860 50820 34916
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 49196 34076 49252 34132
rect 48412 31724 48468 31780
rect 48636 32508 48692 32564
rect 48748 32396 48804 32452
rect 48412 30940 48468 30996
rect 52108 36594 52164 36596
rect 52108 36542 52110 36594
rect 52110 36542 52162 36594
rect 52162 36542 52164 36594
rect 52108 36540 52164 36542
rect 51548 34860 51604 34916
rect 50316 33234 50372 33236
rect 50316 33182 50318 33234
rect 50318 33182 50370 33234
rect 50370 33182 50372 33234
rect 50316 33180 50372 33182
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 50764 32786 50820 32788
rect 50764 32734 50766 32786
rect 50766 32734 50818 32786
rect 50818 32734 50820 32786
rect 50764 32732 50820 32734
rect 53228 40402 53284 40404
rect 53228 40350 53230 40402
rect 53230 40350 53282 40402
rect 53282 40350 53284 40402
rect 53228 40348 53284 40350
rect 55132 41916 55188 41972
rect 55692 43708 55748 43764
rect 56812 53452 56868 53508
rect 56588 52946 56644 52948
rect 56588 52894 56590 52946
rect 56590 52894 56642 52946
rect 56642 52894 56644 52946
rect 56588 52892 56644 52894
rect 57036 51884 57092 51940
rect 57372 50204 57428 50260
rect 57484 49980 57540 50036
rect 57932 50482 57988 50484
rect 57932 50430 57934 50482
rect 57934 50430 57986 50482
rect 57986 50430 57988 50482
rect 57932 50428 57988 50430
rect 56588 49922 56644 49924
rect 56588 49870 56590 49922
rect 56590 49870 56642 49922
rect 56642 49870 56644 49922
rect 56588 49868 56644 49870
rect 56700 49196 56756 49252
rect 56364 47292 56420 47348
rect 57596 49810 57652 49812
rect 57596 49758 57598 49810
rect 57598 49758 57650 49810
rect 57650 49758 57652 49810
rect 57596 49756 57652 49758
rect 58156 50204 58212 50260
rect 58156 49196 58212 49252
rect 57036 46786 57092 46788
rect 57036 46734 57038 46786
rect 57038 46734 57090 46786
rect 57090 46734 57092 46786
rect 57036 46732 57092 46734
rect 56700 46620 56756 46676
rect 57260 46620 57316 46676
rect 56140 45052 56196 45108
rect 56588 45666 56644 45668
rect 56588 45614 56590 45666
rect 56590 45614 56642 45666
rect 56642 45614 56644 45666
rect 56588 45612 56644 45614
rect 56364 43932 56420 43988
rect 57484 46060 57540 46116
rect 56140 43260 56196 43316
rect 55580 41916 55636 41972
rect 54460 40348 54516 40404
rect 53452 40290 53508 40292
rect 53452 40238 53454 40290
rect 53454 40238 53506 40290
rect 53506 40238 53508 40290
rect 53452 40236 53508 40238
rect 52892 40124 52948 40180
rect 54348 40012 54404 40068
rect 52892 39564 52948 39620
rect 53676 39730 53732 39732
rect 53676 39678 53678 39730
rect 53678 39678 53730 39730
rect 53730 39678 53732 39730
rect 53676 39676 53732 39678
rect 53116 39004 53172 39060
rect 52780 36594 52836 36596
rect 52780 36542 52782 36594
rect 52782 36542 52834 36594
rect 52834 36542 52836 36594
rect 52780 36540 52836 36542
rect 52892 36316 52948 36372
rect 52668 36204 52724 36260
rect 52220 34972 52276 35028
rect 52220 33964 52276 34020
rect 51884 33346 51940 33348
rect 51884 33294 51886 33346
rect 51886 33294 51938 33346
rect 51938 33294 51940 33346
rect 51884 33292 51940 33294
rect 52108 33122 52164 33124
rect 52108 33070 52110 33122
rect 52110 33070 52162 33122
rect 52162 33070 52164 33122
rect 52108 33068 52164 33070
rect 51884 32732 51940 32788
rect 51996 32674 52052 32676
rect 51996 32622 51998 32674
rect 51998 32622 52050 32674
rect 52050 32622 52052 32674
rect 51996 32620 52052 32622
rect 49084 32562 49140 32564
rect 49084 32510 49086 32562
rect 49086 32510 49138 32562
rect 49138 32510 49140 32562
rect 49084 32508 49140 32510
rect 49756 32562 49812 32564
rect 49756 32510 49758 32562
rect 49758 32510 49810 32562
rect 49810 32510 49812 32562
rect 49756 32508 49812 32510
rect 50540 32562 50596 32564
rect 50540 32510 50542 32562
rect 50542 32510 50594 32562
rect 50594 32510 50596 32562
rect 50540 32508 50596 32510
rect 51660 32562 51716 32564
rect 51660 32510 51662 32562
rect 51662 32510 51714 32562
rect 51714 32510 51716 32562
rect 51660 32508 51716 32510
rect 49644 32450 49700 32452
rect 49644 32398 49646 32450
rect 49646 32398 49698 32450
rect 49698 32398 49700 32450
rect 49644 32396 49700 32398
rect 49532 31836 49588 31892
rect 49196 31554 49252 31556
rect 49196 31502 49198 31554
rect 49198 31502 49250 31554
rect 49250 31502 49252 31554
rect 49196 31500 49252 31502
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 48748 31164 48804 31220
rect 48972 30994 49028 30996
rect 48972 30942 48974 30994
rect 48974 30942 49026 30994
rect 49026 30942 49028 30994
rect 48972 30940 49028 30942
rect 48524 30156 48580 30212
rect 48524 29372 48580 29428
rect 48412 28418 48468 28420
rect 48412 28366 48414 28418
rect 48414 28366 48466 28418
rect 48466 28366 48468 28418
rect 48412 28364 48468 28366
rect 48636 28252 48692 28308
rect 48636 26908 48692 26964
rect 49308 30770 49364 30772
rect 49308 30718 49310 30770
rect 49310 30718 49362 30770
rect 49362 30718 49364 30770
rect 49308 30716 49364 30718
rect 49532 30156 49588 30212
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 49644 29650 49700 29652
rect 49644 29598 49646 29650
rect 49646 29598 49698 29650
rect 49698 29598 49700 29650
rect 49644 29596 49700 29598
rect 49532 29484 49588 29540
rect 49308 29426 49364 29428
rect 49308 29374 49310 29426
rect 49310 29374 49362 29426
rect 49362 29374 49364 29426
rect 49308 29372 49364 29374
rect 50764 29538 50820 29540
rect 50764 29486 50766 29538
rect 50766 29486 50818 29538
rect 50818 29486 50820 29538
rect 50764 29484 50820 29486
rect 52892 34972 52948 35028
rect 53116 36988 53172 37044
rect 53900 36988 53956 37044
rect 53116 36092 53172 36148
rect 53116 35308 53172 35364
rect 53340 33964 53396 34020
rect 53004 33516 53060 33572
rect 52556 33068 52612 33124
rect 52780 33234 52836 33236
rect 52780 33182 52782 33234
rect 52782 33182 52834 33234
rect 52834 33182 52836 33234
rect 52780 33180 52836 33182
rect 52556 32562 52612 32564
rect 52556 32510 52558 32562
rect 52558 32510 52610 32562
rect 52610 32510 52612 32562
rect 52556 32508 52612 32510
rect 52332 32396 52388 32452
rect 52668 31890 52724 31892
rect 52668 31838 52670 31890
rect 52670 31838 52722 31890
rect 52722 31838 52724 31890
rect 52668 31836 52724 31838
rect 52892 32508 52948 32564
rect 52892 32284 52948 32340
rect 53004 32732 53060 32788
rect 53116 32620 53172 32676
rect 53340 32338 53396 32340
rect 53340 32286 53342 32338
rect 53342 32286 53394 32338
rect 53394 32286 53396 32338
rect 53340 32284 53396 32286
rect 53228 31778 53284 31780
rect 53228 31726 53230 31778
rect 53230 31726 53282 31778
rect 53282 31726 53284 31778
rect 53228 31724 53284 31726
rect 54012 36092 54068 36148
rect 55244 40290 55300 40292
rect 55244 40238 55246 40290
rect 55246 40238 55298 40290
rect 55298 40238 55300 40290
rect 55244 40236 55300 40238
rect 54796 40124 54852 40180
rect 54908 39676 54964 39732
rect 54572 39340 54628 39396
rect 54572 39116 54628 39172
rect 54908 39452 54964 39508
rect 54460 38220 54516 38276
rect 54348 36988 54404 37044
rect 54348 36258 54404 36260
rect 54348 36206 54350 36258
rect 54350 36206 54402 36258
rect 54402 36206 54404 36258
rect 54348 36204 54404 36206
rect 55692 40572 55748 40628
rect 57484 44380 57540 44436
rect 56924 43820 56980 43876
rect 56924 43314 56980 43316
rect 56924 43262 56926 43314
rect 56926 43262 56978 43314
rect 56978 43262 56980 43314
rect 56924 43260 56980 43262
rect 56812 41916 56868 41972
rect 58268 44492 58324 44548
rect 58156 44434 58212 44436
rect 58156 44382 58158 44434
rect 58158 44382 58210 44434
rect 58210 44382 58212 44434
rect 58156 44380 58212 44382
rect 56140 40348 56196 40404
rect 58156 41916 58212 41972
rect 57596 40236 57652 40292
rect 55244 39618 55300 39620
rect 55244 39566 55246 39618
rect 55246 39566 55298 39618
rect 55298 39566 55300 39618
rect 55244 39564 55300 39566
rect 55804 39116 55860 39172
rect 55468 39058 55524 39060
rect 55468 39006 55470 39058
rect 55470 39006 55522 39058
rect 55522 39006 55524 39058
rect 55468 39004 55524 39006
rect 55916 39058 55972 39060
rect 55916 39006 55918 39058
rect 55918 39006 55970 39058
rect 55970 39006 55972 39058
rect 55916 39004 55972 39006
rect 57484 40124 57540 40180
rect 57820 39004 57876 39060
rect 58044 40236 58100 40292
rect 57148 38108 57204 38164
rect 58268 40124 58324 40180
rect 58156 38668 58212 38724
rect 54908 37212 54964 37268
rect 55244 37154 55300 37156
rect 55244 37102 55246 37154
rect 55246 37102 55298 37154
rect 55298 37102 55300 37154
rect 55244 37100 55300 37102
rect 55356 36540 55412 36596
rect 57820 37212 57876 37268
rect 56588 37154 56644 37156
rect 56588 37102 56590 37154
rect 56590 37102 56642 37154
rect 56642 37102 56644 37154
rect 56588 37100 56644 37102
rect 56700 36988 56756 37044
rect 56028 36540 56084 36596
rect 54908 36370 54964 36372
rect 54908 36318 54910 36370
rect 54910 36318 54962 36370
rect 54962 36318 54964 36370
rect 54908 36316 54964 36318
rect 54796 36092 54852 36148
rect 54684 35698 54740 35700
rect 54684 35646 54686 35698
rect 54686 35646 54738 35698
rect 54738 35646 54740 35698
rect 54684 35644 54740 35646
rect 54236 35308 54292 35364
rect 54124 34018 54180 34020
rect 54124 33966 54126 34018
rect 54126 33966 54178 34018
rect 54178 33966 54180 34018
rect 54124 33964 54180 33966
rect 54572 33740 54628 33796
rect 53564 33068 53620 33124
rect 53900 32338 53956 32340
rect 53900 32286 53902 32338
rect 53902 32286 53954 32338
rect 53954 32286 53956 32338
rect 53900 32284 53956 32286
rect 54236 32786 54292 32788
rect 54236 32734 54238 32786
rect 54238 32734 54290 32786
rect 54290 32734 54292 32786
rect 54236 32732 54292 32734
rect 54460 32562 54516 32564
rect 54460 32510 54462 32562
rect 54462 32510 54514 32562
rect 54514 32510 54516 32562
rect 54460 32508 54516 32510
rect 55132 35810 55188 35812
rect 55132 35758 55134 35810
rect 55134 35758 55186 35810
rect 55186 35758 55188 35810
rect 55132 35756 55188 35758
rect 54796 35586 54852 35588
rect 54796 35534 54798 35586
rect 54798 35534 54850 35586
rect 54850 35534 54852 35586
rect 54796 35532 54852 35534
rect 54796 33740 54852 33796
rect 54796 33458 54852 33460
rect 54796 33406 54798 33458
rect 54798 33406 54850 33458
rect 54850 33406 54852 33458
rect 54796 33404 54852 33406
rect 53676 31836 53732 31892
rect 53676 31666 53732 31668
rect 53676 31614 53678 31666
rect 53678 31614 53730 31666
rect 53730 31614 53732 31666
rect 53676 31612 53732 31614
rect 52220 30268 52276 30324
rect 49196 25900 49252 25956
rect 49868 26962 49924 26964
rect 49868 26910 49870 26962
rect 49870 26910 49922 26962
rect 49922 26910 49924 26962
rect 49868 26908 49924 26910
rect 50652 29426 50708 29428
rect 50652 29374 50654 29426
rect 50654 29374 50706 29426
rect 50706 29374 50708 29426
rect 50652 29372 50708 29374
rect 51548 29650 51604 29652
rect 51548 29598 51550 29650
rect 51550 29598 51602 29650
rect 51602 29598 51604 29650
rect 51548 29596 51604 29598
rect 53676 30322 53732 30324
rect 53676 30270 53678 30322
rect 53678 30270 53730 30322
rect 53730 30270 53732 30322
rect 53676 30268 53732 30270
rect 53788 29986 53844 29988
rect 53788 29934 53790 29986
rect 53790 29934 53842 29986
rect 53842 29934 53844 29986
rect 53788 29932 53844 29934
rect 54012 30210 54068 30212
rect 54012 30158 54014 30210
rect 54014 30158 54066 30210
rect 54066 30158 54068 30210
rect 54012 30156 54068 30158
rect 51996 28700 52052 28756
rect 51324 28642 51380 28644
rect 51324 28590 51326 28642
rect 51326 28590 51378 28642
rect 51378 28590 51380 28642
rect 51324 28588 51380 28590
rect 51548 28642 51604 28644
rect 51548 28590 51550 28642
rect 51550 28590 51602 28642
rect 51602 28590 51604 28642
rect 51548 28588 51604 28590
rect 52780 29372 52836 29428
rect 52668 28642 52724 28644
rect 52668 28590 52670 28642
rect 52670 28590 52722 28642
rect 52722 28590 52724 28642
rect 52668 28588 52724 28590
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 50092 26962 50148 26964
rect 50092 26910 50094 26962
rect 50094 26910 50146 26962
rect 50146 26910 50148 26962
rect 50092 26908 50148 26910
rect 50652 26850 50708 26852
rect 50652 26798 50654 26850
rect 50654 26798 50706 26850
rect 50706 26798 50708 26850
rect 50652 26796 50708 26798
rect 50316 26460 50372 26516
rect 49868 25900 49924 25956
rect 48300 25564 48356 25620
rect 49084 24892 49140 24948
rect 49308 24834 49364 24836
rect 49308 24782 49310 24834
rect 49310 24782 49362 24834
rect 49362 24782 49364 24834
rect 49308 24780 49364 24782
rect 48748 24444 48804 24500
rect 49756 25116 49812 25172
rect 50092 25676 50148 25732
rect 49084 23938 49140 23940
rect 49084 23886 49086 23938
rect 49086 23886 49138 23938
rect 49138 23886 49140 23938
rect 49084 23884 49140 23886
rect 49980 23884 50036 23940
rect 48076 23042 48132 23044
rect 48076 22990 48078 23042
rect 48078 22990 48130 23042
rect 48130 22990 48132 23042
rect 48076 22988 48132 22990
rect 47964 22652 48020 22708
rect 48300 22540 48356 22596
rect 48748 23100 48804 23156
rect 48860 22764 48916 22820
rect 49196 23154 49252 23156
rect 49196 23102 49198 23154
rect 49198 23102 49250 23154
rect 49250 23102 49252 23154
rect 49196 23100 49252 23102
rect 48972 22652 49028 22708
rect 48748 22428 48804 22484
rect 49420 23154 49476 23156
rect 49420 23102 49422 23154
rect 49422 23102 49474 23154
rect 49474 23102 49476 23154
rect 49420 23100 49476 23102
rect 48972 22316 49028 22372
rect 48188 21474 48244 21476
rect 48188 21422 48190 21474
rect 48190 21422 48242 21474
rect 48242 21422 48244 21474
rect 48188 21420 48244 21422
rect 49756 22764 49812 22820
rect 49308 22316 49364 22372
rect 49532 22652 49588 22708
rect 49980 22652 50036 22708
rect 49420 21474 49476 21476
rect 49420 21422 49422 21474
rect 49422 21422 49474 21474
rect 49474 21422 49476 21474
rect 49420 21420 49476 21422
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 50652 26402 50708 26404
rect 50652 26350 50654 26402
rect 50654 26350 50706 26402
rect 50706 26350 50708 26402
rect 50652 26348 50708 26350
rect 51212 27692 51268 27748
rect 52108 27074 52164 27076
rect 52108 27022 52110 27074
rect 52110 27022 52162 27074
rect 52162 27022 52164 27074
rect 52108 27020 52164 27022
rect 51324 26908 51380 26964
rect 52892 27074 52948 27076
rect 52892 27022 52894 27074
rect 52894 27022 52946 27074
rect 52946 27022 52948 27074
rect 52892 27020 52948 27022
rect 52108 26460 52164 26516
rect 53900 28754 53956 28756
rect 53900 28702 53902 28754
rect 53902 28702 53954 28754
rect 53954 28702 53956 28754
rect 53900 28700 53956 28702
rect 54460 31890 54516 31892
rect 54460 31838 54462 31890
rect 54462 31838 54514 31890
rect 54514 31838 54516 31890
rect 54460 31836 54516 31838
rect 54236 31612 54292 31668
rect 54796 31666 54852 31668
rect 54796 31614 54798 31666
rect 54798 31614 54850 31666
rect 54850 31614 54852 31666
rect 54796 31612 54852 31614
rect 54684 30828 54740 30884
rect 55132 35308 55188 35364
rect 54348 30210 54404 30212
rect 54348 30158 54350 30210
rect 54350 30158 54402 30210
rect 54402 30158 54404 30210
rect 54348 30156 54404 30158
rect 54236 29484 54292 29540
rect 54908 29932 54964 29988
rect 54908 28700 54964 28756
rect 54124 27746 54180 27748
rect 54124 27694 54126 27746
rect 54126 27694 54178 27746
rect 54178 27694 54180 27746
rect 54124 27692 54180 27694
rect 51100 26348 51156 26404
rect 50540 25676 50596 25732
rect 52108 26124 52164 26180
rect 50764 25506 50820 25508
rect 50764 25454 50766 25506
rect 50766 25454 50818 25506
rect 50818 25454 50820 25506
rect 50764 25452 50820 25454
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 51772 25394 51828 25396
rect 51772 25342 51774 25394
rect 51774 25342 51826 25394
rect 51826 25342 51828 25394
rect 51772 25340 51828 25342
rect 51212 24892 51268 24948
rect 51548 25282 51604 25284
rect 51548 25230 51550 25282
rect 51550 25230 51602 25282
rect 51602 25230 51604 25282
rect 51548 25228 51604 25230
rect 51324 24668 51380 24724
rect 51324 24108 51380 24164
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 52892 26012 52948 26068
rect 52668 25394 52724 25396
rect 52668 25342 52670 25394
rect 52670 25342 52722 25394
rect 52722 25342 52724 25394
rect 52668 25340 52724 25342
rect 52220 25228 52276 25284
rect 52780 24668 52836 24724
rect 51772 23154 51828 23156
rect 51772 23102 51774 23154
rect 51774 23102 51826 23154
rect 51826 23102 51828 23154
rect 51772 23100 51828 23102
rect 51212 22316 51268 22372
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 52108 22316 52164 22372
rect 53340 26290 53396 26292
rect 53340 26238 53342 26290
rect 53342 26238 53394 26290
rect 53394 26238 53396 26290
rect 53340 26236 53396 26238
rect 53004 24668 53060 24724
rect 53788 24162 53844 24164
rect 53788 24110 53790 24162
rect 53790 24110 53842 24162
rect 53842 24110 53844 24162
rect 53788 24108 53844 24110
rect 53004 23772 53060 23828
rect 53900 23100 53956 23156
rect 52892 22764 52948 22820
rect 52780 22594 52836 22596
rect 52780 22542 52782 22594
rect 52782 22542 52834 22594
rect 52834 22542 52836 22594
rect 52780 22540 52836 22542
rect 52780 22316 52836 22372
rect 50876 20524 50932 20580
rect 52220 20524 52276 20580
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 49196 19964 49252 20020
rect 45500 19234 45556 19236
rect 45500 19182 45502 19234
rect 45502 19182 45554 19234
rect 45554 19182 45556 19234
rect 45500 19180 45556 19182
rect 45388 18284 45444 18340
rect 45276 17500 45332 17556
rect 44044 15986 44100 15988
rect 44044 15934 44046 15986
rect 44046 15934 44098 15986
rect 44098 15934 44100 15986
rect 44044 15932 44100 15934
rect 43820 13804 43876 13860
rect 44268 14588 44324 14644
rect 43596 9996 43652 10052
rect 43372 9212 43428 9268
rect 44268 9660 44324 9716
rect 43708 9154 43764 9156
rect 43708 9102 43710 9154
rect 43710 9102 43762 9154
rect 43762 9102 43764 9154
rect 43708 9100 43764 9102
rect 42140 8370 42196 8372
rect 42140 8318 42142 8370
rect 42142 8318 42194 8370
rect 42194 8318 42196 8370
rect 42140 8316 42196 8318
rect 40908 7474 40964 7476
rect 40908 7422 40910 7474
rect 40910 7422 40962 7474
rect 40962 7422 40964 7474
rect 40908 7420 40964 7422
rect 42252 7756 42308 7812
rect 41580 7474 41636 7476
rect 41580 7422 41582 7474
rect 41582 7422 41634 7474
rect 41634 7422 41636 7474
rect 41580 7420 41636 7422
rect 42252 6972 42308 7028
rect 41132 6636 41188 6692
rect 42252 6748 42308 6804
rect 42700 6690 42756 6692
rect 42700 6638 42702 6690
rect 42702 6638 42754 6690
rect 42754 6638 42756 6690
rect 42700 6636 42756 6638
rect 43148 6748 43204 6804
rect 44268 8988 44324 9044
rect 44156 7420 44212 7476
rect 43484 6972 43540 7028
rect 43708 6860 43764 6916
rect 40236 6524 40292 6580
rect 41132 5852 41188 5908
rect 39564 4396 39620 4452
rect 41020 5180 41076 5236
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 28588 3612 28644 3668
rect 38892 3612 38948 3668
rect 28140 3500 28196 3556
rect 36652 3554 36708 3556
rect 36652 3502 36654 3554
rect 36654 3502 36706 3554
rect 36706 3502 36708 3554
rect 36652 3500 36708 3502
rect 40796 3666 40852 3668
rect 40796 3614 40798 3666
rect 40798 3614 40850 3666
rect 40850 3614 40852 3666
rect 40796 3612 40852 3614
rect 41132 5068 41188 5124
rect 42700 5234 42756 5236
rect 42700 5182 42702 5234
rect 42702 5182 42754 5234
rect 42754 5182 42756 5234
rect 42700 5180 42756 5182
rect 43036 4060 43092 4116
rect 43148 3724 43204 3780
rect 44044 6412 44100 6468
rect 43596 5068 43652 5124
rect 43484 3612 43540 3668
rect 46620 19234 46676 19236
rect 46620 19182 46622 19234
rect 46622 19182 46674 19234
rect 46674 19182 46676 19234
rect 46620 19180 46676 19182
rect 45724 18338 45780 18340
rect 45724 18286 45726 18338
rect 45726 18286 45778 18338
rect 45778 18286 45780 18338
rect 45724 18284 45780 18286
rect 46956 17778 47012 17780
rect 46956 17726 46958 17778
rect 46958 17726 47010 17778
rect 47010 17726 47012 17778
rect 46956 17724 47012 17726
rect 48636 19346 48692 19348
rect 48636 19294 48638 19346
rect 48638 19294 48690 19346
rect 48690 19294 48692 19346
rect 48636 19292 48692 19294
rect 48300 19122 48356 19124
rect 48300 19070 48302 19122
rect 48302 19070 48354 19122
rect 48354 19070 48356 19122
rect 48300 19068 48356 19070
rect 49196 18956 49252 19012
rect 47964 18620 48020 18676
rect 49420 19292 49476 19348
rect 49868 20018 49924 20020
rect 49868 19966 49870 20018
rect 49870 19966 49922 20018
rect 49922 19966 49924 20018
rect 49868 19964 49924 19966
rect 49532 19068 49588 19124
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 49420 18508 49476 18564
rect 50428 18508 50484 18564
rect 48188 18172 48244 18228
rect 48748 18172 48804 18228
rect 45724 16940 45780 16996
rect 46172 16882 46228 16884
rect 46172 16830 46174 16882
rect 46174 16830 46226 16882
rect 46226 16830 46228 16882
rect 46172 16828 46228 16830
rect 47852 17724 47908 17780
rect 46732 16828 46788 16884
rect 47516 16882 47572 16884
rect 47516 16830 47518 16882
rect 47518 16830 47570 16882
rect 47570 16830 47572 16882
rect 47516 16828 47572 16830
rect 47292 16770 47348 16772
rect 47292 16718 47294 16770
rect 47294 16718 47346 16770
rect 47346 16718 47348 16770
rect 47292 16716 47348 16718
rect 48748 16940 48804 16996
rect 48188 16716 48244 16772
rect 46844 15932 46900 15988
rect 46732 15820 46788 15876
rect 45052 14642 45108 14644
rect 45052 14590 45054 14642
rect 45054 14590 45106 14642
rect 45106 14590 45108 14642
rect 45052 14588 45108 14590
rect 44828 13804 44884 13860
rect 45724 13692 45780 13748
rect 45388 13132 45444 13188
rect 45052 12738 45108 12740
rect 45052 12686 45054 12738
rect 45054 12686 45106 12738
rect 45106 12686 45108 12738
rect 45052 12684 45108 12686
rect 45164 12290 45220 12292
rect 45164 12238 45166 12290
rect 45166 12238 45218 12290
rect 45218 12238 45220 12290
rect 45164 12236 45220 12238
rect 46956 14476 47012 14532
rect 46284 13746 46340 13748
rect 46284 13694 46286 13746
rect 46286 13694 46338 13746
rect 46338 13694 46340 13746
rect 46284 13692 46340 13694
rect 45948 13356 46004 13412
rect 46396 12796 46452 12852
rect 45948 12684 46004 12740
rect 45724 12236 45780 12292
rect 45836 12012 45892 12068
rect 48300 16658 48356 16660
rect 48300 16606 48302 16658
rect 48302 16606 48354 16658
rect 48354 16606 48356 16658
rect 48300 16604 48356 16606
rect 48188 16210 48244 16212
rect 48188 16158 48190 16210
rect 48190 16158 48242 16210
rect 48242 16158 48244 16210
rect 48188 16156 48244 16158
rect 47180 13132 47236 13188
rect 46732 12290 46788 12292
rect 46732 12238 46734 12290
rect 46734 12238 46786 12290
rect 46786 12238 46788 12290
rect 46732 12236 46788 12238
rect 46844 12684 46900 12740
rect 46620 12178 46676 12180
rect 46620 12126 46622 12178
rect 46622 12126 46674 12178
rect 46674 12126 46676 12178
rect 46620 12124 46676 12126
rect 46508 10892 46564 10948
rect 45836 10780 45892 10836
rect 45612 10444 45668 10500
rect 47292 12348 47348 12404
rect 47068 12236 47124 12292
rect 46956 11618 47012 11620
rect 46956 11566 46958 11618
rect 46958 11566 47010 11618
rect 47010 11566 47012 11618
rect 46956 11564 47012 11566
rect 48860 16210 48916 16212
rect 48860 16158 48862 16210
rect 48862 16158 48914 16210
rect 48914 16158 48916 16210
rect 48860 16156 48916 16158
rect 49644 16156 49700 16212
rect 48748 15314 48804 15316
rect 48748 15262 48750 15314
rect 48750 15262 48802 15314
rect 48802 15262 48804 15314
rect 48748 15260 48804 15262
rect 48188 15202 48244 15204
rect 48188 15150 48190 15202
rect 48190 15150 48242 15202
rect 48242 15150 48244 15202
rect 48188 15148 48244 15150
rect 48972 15202 49028 15204
rect 48972 15150 48974 15202
rect 48974 15150 49026 15202
rect 49026 15150 49028 15202
rect 48972 15148 49028 15150
rect 49756 15202 49812 15204
rect 49756 15150 49758 15202
rect 49758 15150 49810 15202
rect 49810 15150 49812 15202
rect 49756 15148 49812 15150
rect 49308 14700 49364 14756
rect 48636 14530 48692 14532
rect 48636 14478 48638 14530
rect 48638 14478 48690 14530
rect 48690 14478 48692 14530
rect 48636 14476 48692 14478
rect 48076 13746 48132 13748
rect 48076 13694 48078 13746
rect 48078 13694 48130 13746
rect 48130 13694 48132 13746
rect 48076 13692 48132 13694
rect 47740 12348 47796 12404
rect 47964 12124 48020 12180
rect 52108 19234 52164 19236
rect 52108 19182 52110 19234
rect 52110 19182 52162 19234
rect 52162 19182 52164 19234
rect 52108 19180 52164 19182
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 51436 17836 51492 17892
rect 52108 17612 52164 17668
rect 51884 17388 51940 17444
rect 51212 16828 51268 16884
rect 51660 16828 51716 16884
rect 50988 16210 51044 16212
rect 50988 16158 50990 16210
rect 50990 16158 51042 16210
rect 51042 16158 51044 16210
rect 50988 16156 51044 16158
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 50540 14530 50596 14532
rect 50540 14478 50542 14530
rect 50542 14478 50594 14530
rect 50594 14478 50596 14530
rect 50540 14476 50596 14478
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 49308 13746 49364 13748
rect 49308 13694 49310 13746
rect 49310 13694 49362 13746
rect 49362 13694 49364 13746
rect 49308 13692 49364 13694
rect 49532 13746 49588 13748
rect 49532 13694 49534 13746
rect 49534 13694 49586 13746
rect 49586 13694 49588 13746
rect 49532 13692 49588 13694
rect 49196 13468 49252 13524
rect 49084 12908 49140 12964
rect 48972 12402 49028 12404
rect 48972 12350 48974 12402
rect 48974 12350 49026 12402
rect 49026 12350 49028 12402
rect 48972 12348 49028 12350
rect 48188 12236 48244 12292
rect 48076 11676 48132 11732
rect 48188 12012 48244 12068
rect 49196 12572 49252 12628
rect 49308 12236 49364 12292
rect 49756 13580 49812 13636
rect 50092 13522 50148 13524
rect 50092 13470 50094 13522
rect 50094 13470 50146 13522
rect 50146 13470 50148 13522
rect 50092 13468 50148 13470
rect 49756 12796 49812 12852
rect 49980 12684 50036 12740
rect 50204 12572 50260 12628
rect 51212 13916 51268 13972
rect 50540 13746 50596 13748
rect 50540 13694 50542 13746
rect 50542 13694 50594 13746
rect 50594 13694 50596 13746
rect 50540 13692 50596 13694
rect 50988 12962 51044 12964
rect 50988 12910 50990 12962
rect 50990 12910 51042 12962
rect 51042 12910 51044 12962
rect 50988 12908 51044 12910
rect 50876 12738 50932 12740
rect 50876 12686 50878 12738
rect 50878 12686 50930 12738
rect 50930 12686 50932 12738
rect 50876 12684 50932 12686
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 49420 12124 49476 12180
rect 50204 12124 50260 12180
rect 49084 12012 49140 12068
rect 48748 11564 48804 11620
rect 46956 10780 47012 10836
rect 47180 10892 47236 10948
rect 46732 10444 46788 10500
rect 47404 10386 47460 10388
rect 47404 10334 47406 10386
rect 47406 10334 47458 10386
rect 47458 10334 47460 10386
rect 47404 10332 47460 10334
rect 48748 10386 48804 10388
rect 48748 10334 48750 10386
rect 48750 10334 48802 10386
rect 48802 10334 48804 10386
rect 48748 10332 48804 10334
rect 47740 10050 47796 10052
rect 47740 9998 47742 10050
rect 47742 9998 47794 10050
rect 47794 9998 47796 10050
rect 47740 9996 47796 9998
rect 46172 9042 46228 9044
rect 46172 8990 46174 9042
rect 46174 8990 46226 9042
rect 46226 8990 46228 9042
rect 46172 8988 46228 8990
rect 45612 6748 45668 6804
rect 45724 7980 45780 8036
rect 47964 9826 48020 9828
rect 47964 9774 47966 9826
rect 47966 9774 48018 9826
rect 48018 9774 48020 9826
rect 47964 9772 48020 9774
rect 48860 9996 48916 10052
rect 48076 9154 48132 9156
rect 48076 9102 48078 9154
rect 48078 9102 48130 9154
rect 48130 9102 48132 9154
rect 48076 9100 48132 9102
rect 48188 9042 48244 9044
rect 48188 8990 48190 9042
rect 48190 8990 48242 9042
rect 48242 8990 48244 9042
rect 48188 8988 48244 8990
rect 49084 9772 49140 9828
rect 50876 11676 50932 11732
rect 50204 11394 50260 11396
rect 50204 11342 50206 11394
rect 50206 11342 50258 11394
rect 50258 11342 50260 11394
rect 50204 11340 50260 11342
rect 51884 14812 51940 14868
rect 52892 20524 52948 20580
rect 53900 21586 53956 21588
rect 53900 21534 53902 21586
rect 53902 21534 53954 21586
rect 53954 21534 53956 21586
rect 53900 21532 53956 21534
rect 53004 19292 53060 19348
rect 52556 19180 52612 19236
rect 53788 19346 53844 19348
rect 53788 19294 53790 19346
rect 53790 19294 53842 19346
rect 53842 19294 53844 19346
rect 53788 19292 53844 19294
rect 53116 19122 53172 19124
rect 53116 19070 53118 19122
rect 53118 19070 53170 19122
rect 53170 19070 53172 19122
rect 53116 19068 53172 19070
rect 52668 18956 52724 19012
rect 52892 17666 52948 17668
rect 52892 17614 52894 17666
rect 52894 17614 52946 17666
rect 52946 17614 52948 17666
rect 52892 17612 52948 17614
rect 52780 17500 52836 17556
rect 54236 26796 54292 26852
rect 54908 26796 54964 26852
rect 55020 29484 55076 29540
rect 54348 26402 54404 26404
rect 54348 26350 54350 26402
rect 54350 26350 54402 26402
rect 54402 26350 54404 26402
rect 54348 26348 54404 26350
rect 55020 26348 55076 26404
rect 54124 26290 54180 26292
rect 54124 26238 54126 26290
rect 54126 26238 54178 26290
rect 54178 26238 54180 26290
rect 54124 26236 54180 26238
rect 54908 25676 54964 25732
rect 54572 24722 54628 24724
rect 54572 24670 54574 24722
rect 54574 24670 54626 24722
rect 54626 24670 54628 24722
rect 54572 24668 54628 24670
rect 54460 24556 54516 24612
rect 56028 35698 56084 35700
rect 56028 35646 56030 35698
rect 56030 35646 56082 35698
rect 56082 35646 56084 35698
rect 56028 35644 56084 35646
rect 55468 35586 55524 35588
rect 55468 35534 55470 35586
rect 55470 35534 55522 35586
rect 55522 35534 55524 35586
rect 55468 35532 55524 35534
rect 56700 35308 56756 35364
rect 55244 33740 55300 33796
rect 56028 33458 56084 33460
rect 56028 33406 56030 33458
rect 56030 33406 56082 33458
rect 56082 33406 56084 33458
rect 56028 33404 56084 33406
rect 57372 32786 57428 32788
rect 57372 32734 57374 32786
rect 57374 32734 57426 32786
rect 57426 32734 57428 32786
rect 57372 32732 57428 32734
rect 56028 31666 56084 31668
rect 56028 31614 56030 31666
rect 56030 31614 56082 31666
rect 56082 31614 56084 31666
rect 56028 31612 56084 31614
rect 55244 25676 55300 25732
rect 54796 25282 54852 25284
rect 54796 25230 54798 25282
rect 54798 25230 54850 25282
rect 54850 25230 54852 25282
rect 54796 25228 54852 25230
rect 58156 35756 58212 35812
rect 58156 33292 58212 33348
rect 58156 32786 58212 32788
rect 58156 32734 58158 32786
rect 58158 32734 58210 32786
rect 58210 32734 58212 32786
rect 58156 32732 58212 32734
rect 58156 31724 58212 31780
rect 58156 28754 58212 28756
rect 58156 28702 58158 28754
rect 58158 28702 58210 28754
rect 58210 28702 58212 28754
rect 58156 28700 58212 28702
rect 55468 26796 55524 26852
rect 57596 26796 57652 26852
rect 58156 26796 58212 26852
rect 55692 26290 55748 26292
rect 55692 26238 55694 26290
rect 55694 26238 55746 26290
rect 55746 26238 55748 26290
rect 55692 26236 55748 26238
rect 55692 25564 55748 25620
rect 58156 25618 58212 25620
rect 58156 25566 58158 25618
rect 58158 25566 58210 25618
rect 58210 25566 58212 25618
rect 58156 25564 58212 25566
rect 54796 24332 54852 24388
rect 54684 22764 54740 22820
rect 55132 24498 55188 24500
rect 55132 24446 55134 24498
rect 55134 24446 55186 24498
rect 55186 24446 55188 24498
rect 55132 24444 55188 24446
rect 56028 25228 56084 25284
rect 55580 24610 55636 24612
rect 55580 24558 55582 24610
rect 55582 24558 55634 24610
rect 55634 24558 55636 24610
rect 55580 24556 55636 24558
rect 55804 24498 55860 24500
rect 55804 24446 55806 24498
rect 55806 24446 55858 24498
rect 55858 24446 55860 24498
rect 55804 24444 55860 24446
rect 56924 24722 56980 24724
rect 56924 24670 56926 24722
rect 56926 24670 56978 24722
rect 56978 24670 56980 24722
rect 56924 24668 56980 24670
rect 56028 24444 56084 24500
rect 55244 23154 55300 23156
rect 55244 23102 55246 23154
rect 55246 23102 55298 23154
rect 55298 23102 55300 23154
rect 55244 23100 55300 23102
rect 55244 22764 55300 22820
rect 55244 21532 55300 21588
rect 55692 22428 55748 22484
rect 56588 24332 56644 24388
rect 56924 23996 56980 24052
rect 58156 24050 58212 24052
rect 58156 23998 58158 24050
rect 58158 23998 58210 24050
rect 58210 23998 58212 24050
rect 58156 23996 58212 23998
rect 58156 22482 58212 22484
rect 58156 22430 58158 22482
rect 58158 22430 58210 22482
rect 58210 22430 58212 22482
rect 58156 22428 58212 22430
rect 57820 21698 57876 21700
rect 57820 21646 57822 21698
rect 57822 21646 57874 21698
rect 57874 21646 57876 21698
rect 57820 21644 57876 21646
rect 58156 21084 58212 21140
rect 54908 20076 54964 20132
rect 54012 19180 54068 19236
rect 54460 19292 54516 19348
rect 53228 17388 53284 17444
rect 54012 17388 54068 17444
rect 52444 16940 52500 16996
rect 52668 16604 52724 16660
rect 54684 19906 54740 19908
rect 54684 19854 54686 19906
rect 54686 19854 54738 19906
rect 54738 19854 54740 19906
rect 54684 19852 54740 19854
rect 54684 19234 54740 19236
rect 54684 19182 54686 19234
rect 54686 19182 54738 19234
rect 54738 19182 54740 19234
rect 54684 19180 54740 19182
rect 54460 19122 54516 19124
rect 54460 19070 54462 19122
rect 54462 19070 54514 19122
rect 54514 19070 54516 19122
rect 54460 19068 54516 19070
rect 54796 19010 54852 19012
rect 54796 18958 54798 19010
rect 54798 18958 54850 19010
rect 54850 18958 54852 19010
rect 54796 18956 54852 18958
rect 56140 20130 56196 20132
rect 56140 20078 56142 20130
rect 56142 20078 56194 20130
rect 56194 20078 56196 20130
rect 56140 20076 56196 20078
rect 55468 19906 55524 19908
rect 55468 19854 55470 19906
rect 55470 19854 55522 19906
rect 55522 19854 55524 19906
rect 55468 19852 55524 19854
rect 58156 19346 58212 19348
rect 58156 19294 58158 19346
rect 58158 19294 58210 19346
rect 58210 19294 58212 19346
rect 58156 19292 58212 19294
rect 55132 18956 55188 19012
rect 55468 18396 55524 18452
rect 55916 19180 55972 19236
rect 55244 18284 55300 18340
rect 53788 15986 53844 15988
rect 53788 15934 53790 15986
rect 53790 15934 53842 15986
rect 53842 15934 53844 15986
rect 53788 15932 53844 15934
rect 52444 15036 52500 15092
rect 52780 15036 52836 15092
rect 51884 14588 51940 14644
rect 51996 14476 52052 14532
rect 51996 13970 52052 13972
rect 51996 13918 51998 13970
rect 51998 13918 52050 13970
rect 52050 13918 52052 13970
rect 51996 13916 52052 13918
rect 52444 13746 52500 13748
rect 52444 13694 52446 13746
rect 52446 13694 52498 13746
rect 52498 13694 52500 13746
rect 52444 13692 52500 13694
rect 51884 13634 51940 13636
rect 51884 13582 51886 13634
rect 51886 13582 51938 13634
rect 51938 13582 51940 13634
rect 51884 13580 51940 13582
rect 52892 13580 52948 13636
rect 53452 15036 53508 15092
rect 54012 16156 54068 16212
rect 54572 15986 54628 15988
rect 54572 15934 54574 15986
rect 54574 15934 54626 15986
rect 54626 15934 54628 15986
rect 54572 15932 54628 15934
rect 54348 15148 54404 15204
rect 53340 14530 53396 14532
rect 53340 14478 53342 14530
rect 53342 14478 53394 14530
rect 53394 14478 53396 14530
rect 53340 14476 53396 14478
rect 53228 13692 53284 13748
rect 52892 13356 52948 13412
rect 52108 12290 52164 12292
rect 52108 12238 52110 12290
rect 52110 12238 52162 12290
rect 52162 12238 52164 12290
rect 52108 12236 52164 12238
rect 52892 12850 52948 12852
rect 52892 12798 52894 12850
rect 52894 12798 52946 12850
rect 52946 12798 52948 12850
rect 52892 12796 52948 12798
rect 52780 12684 52836 12740
rect 52780 12236 52836 12292
rect 53340 13356 53396 13412
rect 53340 12796 53396 12852
rect 53340 11954 53396 11956
rect 53340 11902 53342 11954
rect 53342 11902 53394 11954
rect 53394 11902 53396 11954
rect 53340 11900 53396 11902
rect 53116 11452 53172 11508
rect 50316 11116 50372 11172
rect 50092 10722 50148 10724
rect 50092 10670 50094 10722
rect 50094 10670 50146 10722
rect 50146 10670 50148 10722
rect 50092 10668 50148 10670
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 53900 12738 53956 12740
rect 53900 12686 53902 12738
rect 53902 12686 53954 12738
rect 53954 12686 53956 12738
rect 53900 12684 53956 12686
rect 51436 11282 51492 11284
rect 51436 11230 51438 11282
rect 51438 11230 51490 11282
rect 51490 11230 51492 11282
rect 51436 11228 51492 11230
rect 53004 11228 53060 11284
rect 51324 11170 51380 11172
rect 51324 11118 51326 11170
rect 51326 11118 51378 11170
rect 51378 11118 51380 11170
rect 51324 11116 51380 11118
rect 50988 10668 51044 10724
rect 50540 9826 50596 9828
rect 50540 9774 50542 9826
rect 50542 9774 50594 9826
rect 50594 9774 50596 9826
rect 50540 9772 50596 9774
rect 51324 9772 51380 9828
rect 49644 9436 49700 9492
rect 48972 9042 49028 9044
rect 48972 8990 48974 9042
rect 48974 8990 49026 9042
rect 49026 8990 49028 9042
rect 48972 8988 49028 8990
rect 47628 8482 47684 8484
rect 47628 8430 47630 8482
rect 47630 8430 47682 8482
rect 47682 8430 47684 8482
rect 47628 8428 47684 8430
rect 49644 9100 49700 9156
rect 48748 8428 48804 8484
rect 49980 9436 50036 9492
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 51660 9548 51716 9604
rect 50092 9100 50148 9156
rect 49980 8764 50036 8820
rect 51212 9042 51268 9044
rect 51212 8990 51214 9042
rect 51214 8990 51266 9042
rect 51266 8990 51268 9042
rect 51212 8988 51268 8990
rect 46284 7868 46340 7924
rect 45948 7474 46004 7476
rect 45948 7422 45950 7474
rect 45950 7422 46002 7474
rect 46002 7422 46004 7474
rect 45948 7420 46004 7422
rect 44380 6636 44436 6692
rect 45052 6690 45108 6692
rect 45052 6638 45054 6690
rect 45054 6638 45106 6690
rect 45106 6638 45108 6690
rect 45052 6636 45108 6638
rect 45388 6524 45444 6580
rect 44828 6412 44884 6468
rect 45388 6300 45444 6356
rect 45500 6636 45556 6692
rect 46172 6636 46228 6692
rect 46060 6578 46116 6580
rect 46060 6526 46062 6578
rect 46062 6526 46114 6578
rect 46114 6526 46116 6578
rect 46060 6524 46116 6526
rect 45612 6466 45668 6468
rect 45612 6414 45614 6466
rect 45614 6414 45666 6466
rect 45666 6414 45668 6466
rect 45612 6412 45668 6414
rect 45500 6076 45556 6132
rect 46396 6300 46452 6356
rect 47068 8034 47124 8036
rect 47068 7982 47070 8034
rect 47070 7982 47122 8034
rect 47122 7982 47124 8034
rect 47068 7980 47124 7982
rect 47628 8034 47684 8036
rect 47628 7982 47630 8034
rect 47630 7982 47682 8034
rect 47682 7982 47684 8034
rect 47628 7980 47684 7982
rect 47292 7868 47348 7924
rect 49644 7868 49700 7924
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 51436 8204 51492 8260
rect 47180 6690 47236 6692
rect 47180 6638 47182 6690
rect 47182 6638 47234 6690
rect 47234 6638 47236 6690
rect 47180 6636 47236 6638
rect 46956 6524 47012 6580
rect 46620 6466 46676 6468
rect 46620 6414 46622 6466
rect 46622 6414 46674 6466
rect 46674 6414 46676 6466
rect 46620 6412 46676 6414
rect 48972 6914 49028 6916
rect 48972 6862 48974 6914
rect 48974 6862 49026 6914
rect 49026 6862 49028 6914
rect 48972 6860 49028 6862
rect 49644 6860 49700 6916
rect 49308 6748 49364 6804
rect 47404 6524 47460 6580
rect 46956 5964 47012 6020
rect 47852 6018 47908 6020
rect 47852 5966 47854 6018
rect 47854 5966 47906 6018
rect 47906 5966 47908 6018
rect 47852 5964 47908 5966
rect 47404 5906 47460 5908
rect 47404 5854 47406 5906
rect 47406 5854 47458 5906
rect 47458 5854 47460 5906
rect 47404 5852 47460 5854
rect 46620 5740 46676 5796
rect 47964 5794 48020 5796
rect 47964 5742 47966 5794
rect 47966 5742 48018 5794
rect 48018 5742 48020 5794
rect 47964 5740 48020 5742
rect 49644 6130 49700 6132
rect 49644 6078 49646 6130
rect 49646 6078 49698 6130
rect 49698 6078 49700 6130
rect 49644 6076 49700 6078
rect 50092 6914 50148 6916
rect 50092 6862 50094 6914
rect 50094 6862 50146 6914
rect 50146 6862 50148 6914
rect 50092 6860 50148 6862
rect 50988 7644 51044 7700
rect 50204 6748 50260 6804
rect 50764 6748 50820 6804
rect 52780 9548 52836 9604
rect 52892 9154 52948 9156
rect 52892 9102 52894 9154
rect 52894 9102 52946 9154
rect 52946 9102 52948 9154
rect 52892 9100 52948 9102
rect 52332 8764 52388 8820
rect 52220 7084 52276 7140
rect 52892 8258 52948 8260
rect 52892 8206 52894 8258
rect 52894 8206 52946 8258
rect 52946 8206 52948 8258
rect 52892 8204 52948 8206
rect 52332 6972 52388 7028
rect 52668 6860 52724 6916
rect 52780 6972 52836 7028
rect 52108 6636 52164 6692
rect 51100 6578 51156 6580
rect 51100 6526 51102 6578
rect 51102 6526 51154 6578
rect 51154 6526 51156 6578
rect 51100 6524 51156 6526
rect 50092 6076 50148 6132
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 49980 5852 50036 5908
rect 50316 5906 50372 5908
rect 50316 5854 50318 5906
rect 50318 5854 50370 5906
rect 50370 5854 50372 5906
rect 50316 5852 50372 5854
rect 49084 5740 49140 5796
rect 49308 5122 49364 5124
rect 49308 5070 49310 5122
rect 49310 5070 49362 5122
rect 49362 5070 49364 5122
rect 49308 5068 49364 5070
rect 44940 5010 44996 5012
rect 44940 4958 44942 5010
rect 44942 4958 44994 5010
rect 44994 4958 44996 5010
rect 44940 4956 44996 4958
rect 46508 4956 46564 5012
rect 46060 4898 46116 4900
rect 46060 4846 46062 4898
rect 46062 4846 46114 4898
rect 46114 4846 46116 4898
rect 46060 4844 46116 4846
rect 45388 4114 45444 4116
rect 45388 4062 45390 4114
rect 45390 4062 45442 4114
rect 45442 4062 45444 4114
rect 45388 4060 45444 4062
rect 44492 3724 44548 3780
rect 44380 3666 44436 3668
rect 44380 3614 44382 3666
rect 44382 3614 44434 3666
rect 44434 3614 44436 3666
rect 44380 3612 44436 3614
rect 47404 4844 47460 4900
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 47404 3554 47460 3556
rect 47404 3502 47406 3554
rect 47406 3502 47458 3554
rect 47458 3502 47460 3554
rect 47404 3500 47460 3502
rect 45052 3388 45108 3444
rect 53564 9100 53620 9156
rect 54012 11954 54068 11956
rect 54012 11902 54014 11954
rect 54014 11902 54066 11954
rect 54066 11902 54068 11954
rect 54012 11900 54068 11902
rect 54012 11452 54068 11508
rect 54236 12684 54292 12740
rect 54236 11788 54292 11844
rect 54012 10220 54068 10276
rect 54012 8370 54068 8372
rect 54012 8318 54014 8370
rect 54014 8318 54066 8370
rect 54066 8318 54068 8370
rect 54012 8316 54068 8318
rect 53116 8204 53172 8260
rect 53900 8258 53956 8260
rect 53900 8206 53902 8258
rect 53902 8206 53954 8258
rect 53954 8206 53956 8258
rect 53900 8204 53956 8206
rect 53116 7586 53172 7588
rect 53116 7534 53118 7586
rect 53118 7534 53170 7586
rect 53170 7534 53172 7586
rect 53116 7532 53172 7534
rect 53340 7644 53396 7700
rect 54460 12738 54516 12740
rect 54460 12686 54462 12738
rect 54462 12686 54514 12738
rect 54514 12686 54516 12738
rect 54460 12684 54516 12686
rect 55356 16828 55412 16884
rect 54908 14588 54964 14644
rect 58156 16210 58212 16212
rect 58156 16158 58158 16210
rect 58158 16158 58210 16210
rect 58210 16158 58212 16210
rect 58156 16156 58212 16158
rect 57820 15426 57876 15428
rect 57820 15374 57822 15426
rect 57822 15374 57874 15426
rect 57874 15374 57876 15426
rect 57820 15372 57876 15374
rect 57596 15314 57652 15316
rect 57596 15262 57598 15314
rect 57598 15262 57650 15314
rect 57650 15262 57652 15314
rect 57596 15260 57652 15262
rect 58156 15314 58212 15316
rect 58156 15262 58158 15314
rect 58158 15262 58210 15314
rect 58210 15262 58212 15314
rect 58156 15260 58212 15262
rect 58156 14812 58212 14868
rect 56028 14642 56084 14644
rect 56028 14590 56030 14642
rect 56030 14590 56082 14642
rect 56082 14590 56084 14642
rect 56028 14588 56084 14590
rect 54908 14306 54964 14308
rect 54908 14254 54910 14306
rect 54910 14254 54962 14306
rect 54962 14254 54964 14306
rect 54908 14252 54964 14254
rect 55692 14252 55748 14308
rect 54684 12572 54740 12628
rect 55132 12572 55188 12628
rect 54460 12460 54516 12516
rect 55020 12460 55076 12516
rect 54572 12178 54628 12180
rect 54572 12126 54574 12178
rect 54574 12126 54626 12178
rect 54626 12126 54628 12178
rect 54572 12124 54628 12126
rect 58156 12796 58212 12852
rect 55356 12178 55412 12180
rect 55356 12126 55358 12178
rect 55358 12126 55410 12178
rect 55410 12126 55412 12178
rect 55356 12124 55412 12126
rect 55244 11506 55300 11508
rect 55244 11454 55246 11506
rect 55246 11454 55298 11506
rect 55298 11454 55300 11506
rect 55244 11452 55300 11454
rect 55692 11452 55748 11508
rect 57372 11506 57428 11508
rect 57372 11454 57374 11506
rect 57374 11454 57426 11506
rect 57426 11454 57428 11506
rect 57372 11452 57428 11454
rect 55468 11340 55524 11396
rect 55132 9548 55188 9604
rect 55244 10220 55300 10276
rect 54572 9042 54628 9044
rect 54572 8990 54574 9042
rect 54574 8990 54626 9042
rect 54626 8990 54628 9042
rect 54572 8988 54628 8990
rect 58044 11394 58100 11396
rect 58044 11342 58046 11394
rect 58046 11342 58098 11394
rect 58098 11342 58100 11394
rect 58044 11340 58100 11342
rect 57596 9436 57652 9492
rect 57820 9266 57876 9268
rect 57820 9214 57822 9266
rect 57822 9214 57874 9266
rect 57874 9214 57876 9266
rect 57820 9212 57876 9214
rect 55468 9100 55524 9156
rect 54460 8818 54516 8820
rect 54460 8766 54462 8818
rect 54462 8766 54514 8818
rect 54514 8766 54516 8818
rect 54460 8764 54516 8766
rect 54348 8540 54404 8596
rect 54236 8092 54292 8148
rect 52892 6748 52948 6804
rect 53116 6860 53172 6916
rect 53340 6914 53396 6916
rect 53340 6862 53342 6914
rect 53342 6862 53394 6914
rect 53394 6862 53396 6914
rect 53340 6860 53396 6862
rect 54348 8316 54404 8372
rect 54908 8316 54964 8372
rect 56588 9042 56644 9044
rect 56588 8990 56590 9042
rect 56590 8990 56642 9042
rect 56642 8990 56644 9042
rect 56588 8988 56644 8990
rect 58156 9436 58212 9492
rect 54908 8146 54964 8148
rect 54908 8094 54910 8146
rect 54910 8094 54962 8146
rect 54962 8094 54964 8146
rect 54908 8092 54964 8094
rect 54348 7586 54404 7588
rect 54348 7534 54350 7586
rect 54350 7534 54402 7586
rect 54402 7534 54404 7586
rect 54348 7532 54404 7534
rect 55356 7474 55412 7476
rect 55356 7422 55358 7474
rect 55358 7422 55410 7474
rect 55410 7422 55412 7474
rect 55356 7420 55412 7422
rect 56588 7474 56644 7476
rect 56588 7422 56590 7474
rect 56590 7422 56642 7474
rect 56642 7422 56644 7474
rect 56588 7420 56644 7422
rect 54124 7084 54180 7140
rect 53564 6972 53620 7028
rect 54236 6860 54292 6916
rect 54796 7196 54852 7252
rect 55244 6802 55300 6804
rect 55244 6750 55246 6802
rect 55246 6750 55298 6802
rect 55298 6750 55300 6802
rect 55244 6748 55300 6750
rect 56028 6636 56084 6692
rect 53452 5180 53508 5236
rect 51324 4898 51380 4900
rect 51324 4846 51326 4898
rect 51326 4846 51378 4898
rect 51378 4846 51380 4898
rect 51324 4844 51380 4846
rect 52668 4844 52724 4900
rect 58044 6690 58100 6692
rect 58044 6638 58046 6690
rect 58046 6638 58098 6690
rect 58098 6638 58100 6690
rect 58044 6636 58100 6638
rect 54684 5234 54740 5236
rect 54684 5182 54686 5234
rect 54686 5182 54738 5234
rect 54738 5182 54740 5234
rect 54684 5180 54740 5182
rect 57820 4450 57876 4452
rect 57820 4398 57822 4450
rect 57822 4398 57874 4450
rect 57874 4398 57876 4450
rect 57820 4396 57876 4398
rect 58156 3612 58212 3668
rect 48860 3500 48916 3556
rect 48972 3442 49028 3444
rect 48972 3390 48974 3442
rect 48974 3390 49026 3442
rect 49026 3390 49028 3442
rect 48972 3388 49028 3390
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
<< metal3 >>
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 59200 56084 60000 56112
rect 57586 56028 57596 56084
rect 57652 56028 58156 56084
rect 58212 56028 60000 56084
rect 59200 56000 60000 56028
rect 23062 55916 23100 55972
rect 23156 55916 23166 55972
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 25778 55356 25788 55412
rect 25844 55356 27132 55412
rect 27188 55356 27524 55412
rect 40226 55356 40236 55412
rect 40292 55356 41804 55412
rect 41860 55356 41870 55412
rect 22978 55244 22988 55300
rect 23044 55244 25452 55300
rect 25508 55244 25518 55300
rect 27468 55188 27524 55356
rect 32050 55244 32060 55300
rect 32116 55244 33516 55300
rect 33572 55244 34076 55300
rect 34132 55244 34142 55300
rect 41234 55244 41244 55300
rect 41300 55244 42364 55300
rect 42420 55244 42430 55300
rect 45490 55244 45500 55300
rect 45556 55244 46060 55300
rect 46116 55244 49308 55300
rect 49364 55244 51996 55300
rect 52052 55244 52668 55300
rect 52724 55244 52734 55300
rect 18274 55132 18284 55188
rect 18340 55132 22764 55188
rect 22820 55132 22830 55188
rect 26114 55132 26124 55188
rect 26180 55132 26684 55188
rect 26740 55132 26908 55188
rect 27458 55132 27468 55188
rect 27524 55132 27534 55188
rect 29810 55132 29820 55188
rect 29876 55132 31276 55188
rect 31332 55132 31342 55188
rect 38098 55132 38108 55188
rect 38164 55132 40684 55188
rect 40740 55132 40750 55188
rect 53442 55132 53452 55188
rect 53508 55132 54460 55188
rect 54516 55132 54526 55188
rect 26852 55076 26908 55132
rect 26852 55020 27356 55076
rect 27412 55020 31388 55076
rect 31444 55020 31454 55076
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 27458 54684 27468 54740
rect 27524 54684 28252 54740
rect 28308 54684 28318 54740
rect 40226 54684 40236 54740
rect 40292 54684 41020 54740
rect 41076 54684 41086 54740
rect 46722 54684 46732 54740
rect 46788 54684 47404 54740
rect 47460 54684 47470 54740
rect 40114 54572 40124 54628
rect 40180 54572 40908 54628
rect 40964 54572 42140 54628
rect 42196 54572 42206 54628
rect 54572 54572 56252 54628
rect 56308 54572 56318 54628
rect 54572 54516 54628 54572
rect 23090 54460 23100 54516
rect 23156 54460 23548 54516
rect 23604 54460 23614 54516
rect 26852 54460 29036 54516
rect 29092 54460 29102 54516
rect 47618 54460 47628 54516
rect 47684 54460 54572 54516
rect 54628 54460 54638 54516
rect 26852 54404 26908 54460
rect 20290 54348 20300 54404
rect 20356 54348 21308 54404
rect 21364 54348 21374 54404
rect 24770 54348 24780 54404
rect 24836 54348 26908 54404
rect 43474 54348 43484 54404
rect 43540 54348 44716 54404
rect 44772 54348 44782 54404
rect 48290 54348 48300 54404
rect 48356 54348 52892 54404
rect 52948 54348 52958 54404
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 20962 54012 20972 54068
rect 21028 54012 21868 54068
rect 21924 54012 22540 54068
rect 22596 54012 22606 54068
rect 26898 54012 26908 54068
rect 26964 54012 29764 54068
rect 27580 53900 29484 53956
rect 29540 53900 29550 53956
rect 27580 53844 27636 53900
rect 29708 53844 29764 54012
rect 41234 53900 41244 53956
rect 41300 53900 42588 53956
rect 42644 53900 42654 53956
rect 54226 53900 54236 53956
rect 54292 53900 54908 53956
rect 54964 53900 55356 53956
rect 55412 53900 55422 53956
rect 21634 53788 21644 53844
rect 21700 53788 21980 53844
rect 22036 53788 27636 53844
rect 28130 53788 28140 53844
rect 28196 53788 29372 53844
rect 29428 53788 29438 53844
rect 29698 53788 29708 53844
rect 29764 53788 31836 53844
rect 31892 53788 31902 53844
rect 36418 53788 36428 53844
rect 36484 53788 37548 53844
rect 37604 53788 39116 53844
rect 39172 53788 40012 53844
rect 40068 53788 41692 53844
rect 41748 53788 41758 53844
rect 50876 53788 52780 53844
rect 52836 53788 52846 53844
rect 53666 53788 53676 53844
rect 53732 53788 54348 53844
rect 54404 53788 54414 53844
rect 27580 53732 27636 53788
rect 50876 53732 50932 53788
rect 52780 53732 52836 53788
rect 18162 53676 18172 53732
rect 18228 53676 20188 53732
rect 20244 53676 20254 53732
rect 20402 53676 20412 53732
rect 20468 53676 21868 53732
rect 21924 53676 21934 53732
rect 22082 53676 22092 53732
rect 22148 53676 22876 53732
rect 22932 53676 22942 53732
rect 23874 53676 23884 53732
rect 23940 53676 25228 53732
rect 25284 53676 25294 53732
rect 27570 53676 27580 53732
rect 27636 53676 27646 53732
rect 28242 53676 28252 53732
rect 28308 53676 28318 53732
rect 34290 53676 34300 53732
rect 34356 53676 36988 53732
rect 37044 53676 37054 53732
rect 40786 53676 40796 53732
rect 40852 53676 41244 53732
rect 41300 53676 41310 53732
rect 50866 53676 50876 53732
rect 50932 53676 50942 53732
rect 52780 53676 55020 53732
rect 55076 53676 55086 53732
rect 22092 53620 22148 53676
rect 28252 53620 28308 53676
rect 21410 53564 21420 53620
rect 21476 53564 22148 53620
rect 26338 53564 26348 53620
rect 26404 53564 28308 53620
rect 53218 53564 53228 53620
rect 53284 53564 54012 53620
rect 54068 53564 54078 53620
rect 22978 53452 22988 53508
rect 23044 53452 25452 53508
rect 25508 53452 25518 53508
rect 26450 53452 26460 53508
rect 26516 53452 27244 53508
rect 27300 53452 27310 53508
rect 27906 53452 27916 53508
rect 27972 53452 30604 53508
rect 30660 53452 30670 53508
rect 35858 53452 35868 53508
rect 35924 53452 37100 53508
rect 37156 53452 37884 53508
rect 37940 53452 37950 53508
rect 40002 53452 40012 53508
rect 40068 53452 40796 53508
rect 40852 53452 40862 53508
rect 42130 53452 42140 53508
rect 42196 53452 43036 53508
rect 43092 53452 43102 53508
rect 46498 53452 46508 53508
rect 46564 53452 48748 53508
rect 48804 53452 49644 53508
rect 49700 53452 49710 53508
rect 55234 53452 55244 53508
rect 55300 53452 56812 53508
rect 56868 53452 56878 53508
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 45042 53116 45052 53172
rect 45108 53116 46732 53172
rect 46788 53116 48076 53172
rect 48132 53116 48142 53172
rect 34066 53004 34076 53060
rect 34132 53004 35196 53060
rect 35252 53004 37100 53060
rect 37156 53004 37996 53060
rect 38052 53004 38062 53060
rect 49970 53004 49980 53060
rect 50036 53004 51660 53060
rect 51716 53004 51726 53060
rect 19058 52892 19068 52948
rect 19124 52892 24668 52948
rect 24724 52892 24734 52948
rect 28354 52892 28364 52948
rect 28420 52892 29260 52948
rect 29316 52892 29326 52948
rect 39218 52892 39228 52948
rect 39284 52892 41132 52948
rect 41188 52892 41198 52948
rect 41346 52892 41356 52948
rect 41412 52892 42476 52948
rect 42532 52892 43372 52948
rect 43428 52892 45276 52948
rect 45332 52892 45342 52948
rect 46274 52892 46284 52948
rect 46340 52892 46956 52948
rect 47012 52892 50092 52948
rect 50148 52892 50158 52948
rect 54786 52892 54796 52948
rect 54852 52892 55244 52948
rect 55300 52892 55310 52948
rect 55458 52892 55468 52948
rect 55524 52892 56588 52948
rect 56644 52892 56654 52948
rect 17490 52780 17500 52836
rect 17556 52780 22652 52836
rect 22708 52780 22718 52836
rect 38770 52668 38780 52724
rect 38836 52668 41468 52724
rect 41524 52668 41534 52724
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 31378 52332 31388 52388
rect 31444 52332 31836 52388
rect 31892 52332 31902 52388
rect 43026 52332 43036 52388
rect 43092 52332 43708 52388
rect 43764 52332 45948 52388
rect 46004 52332 46014 52388
rect 18050 52220 18060 52276
rect 18116 52220 19404 52276
rect 19460 52220 19964 52276
rect 20020 52220 20030 52276
rect 48178 52220 48188 52276
rect 48244 52220 48860 52276
rect 48916 52220 48926 52276
rect 55234 52220 55244 52276
rect 55300 52220 56140 52276
rect 56196 52220 56206 52276
rect 22978 52108 22988 52164
rect 23044 52108 23996 52164
rect 24052 52108 24556 52164
rect 24612 52108 25788 52164
rect 25844 52108 25854 52164
rect 48402 52108 48412 52164
rect 48468 52108 49532 52164
rect 49588 52108 49598 52164
rect 49756 52108 53004 52164
rect 53060 52108 53070 52164
rect 49756 52052 49812 52108
rect 50316 52052 50372 52108
rect 15922 51996 15932 52052
rect 15988 51996 20300 52052
rect 20356 51996 20366 52052
rect 34962 51996 34972 52052
rect 35028 51996 35756 52052
rect 35812 51996 35822 52052
rect 49186 51996 49196 52052
rect 49252 51996 49812 52052
rect 50306 51996 50316 52052
rect 50372 51996 50382 52052
rect 31714 51884 31724 51940
rect 31780 51884 33292 51940
rect 33348 51884 33358 51940
rect 42242 51884 42252 51940
rect 42308 51884 42700 51940
rect 42756 51884 42766 51940
rect 46834 51884 46844 51940
rect 46900 51884 49420 51940
rect 49476 51884 50540 51940
rect 50596 51884 55916 51940
rect 55972 51884 57036 51940
rect 57092 51884 57102 51940
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 30370 51436 30380 51492
rect 30436 51436 30828 51492
rect 30884 51436 32396 51492
rect 32452 51436 32462 51492
rect 37762 51436 37772 51492
rect 37828 51436 38668 51492
rect 38612 51380 38668 51436
rect 20402 51324 20412 51380
rect 20468 51324 21084 51380
rect 21140 51324 22988 51380
rect 23044 51324 23772 51380
rect 23828 51324 23838 51380
rect 30706 51324 30716 51380
rect 30772 51324 31836 51380
rect 31892 51324 31902 51380
rect 37538 51324 37548 51380
rect 37604 51324 38220 51380
rect 38276 51324 38286 51380
rect 38612 51324 50764 51380
rect 50820 51324 55356 51380
rect 55412 51324 55422 51380
rect 38220 51268 38276 51324
rect 19618 51212 19628 51268
rect 19684 51212 20636 51268
rect 20692 51212 20702 51268
rect 23314 51212 23324 51268
rect 23380 51212 23996 51268
rect 24052 51212 24062 51268
rect 38220 51212 38444 51268
rect 38500 51212 42252 51268
rect 42308 51212 42318 51268
rect 43250 51212 43260 51268
rect 43316 51212 45500 51268
rect 45556 51212 45566 51268
rect 51762 51212 51772 51268
rect 51828 51212 53788 51268
rect 53844 51212 53854 51268
rect 42252 51156 42308 51212
rect 16146 51100 16156 51156
rect 16212 51100 21196 51156
rect 21252 51100 21262 51156
rect 28354 51100 28364 51156
rect 28420 51100 30828 51156
rect 30884 51100 30894 51156
rect 42252 51100 46172 51156
rect 46228 51100 46508 51156
rect 46564 51100 46574 51156
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 27122 50876 27132 50932
rect 27188 50876 30492 50932
rect 30548 50876 31276 50932
rect 31332 50876 31342 50932
rect 28690 50764 28700 50820
rect 28756 50764 30156 50820
rect 30212 50764 30222 50820
rect 50082 50764 50092 50820
rect 50148 50764 51212 50820
rect 51268 50764 51278 50820
rect 19058 50652 19068 50708
rect 19124 50652 21308 50708
rect 21364 50652 21374 50708
rect 22754 50652 22764 50708
rect 22820 50652 29484 50708
rect 29540 50652 29550 50708
rect 49186 50652 49196 50708
rect 49252 50652 49980 50708
rect 50036 50652 50652 50708
rect 50708 50652 50718 50708
rect 26338 50540 26348 50596
rect 26404 50540 26908 50596
rect 26964 50540 31164 50596
rect 31220 50540 31230 50596
rect 32274 50540 32284 50596
rect 32340 50540 32956 50596
rect 33012 50540 35868 50596
rect 35924 50540 37100 50596
rect 37156 50540 37166 50596
rect 20178 50428 20188 50484
rect 20244 50428 21980 50484
rect 22036 50428 22046 50484
rect 25890 50428 25900 50484
rect 25956 50428 28252 50484
rect 28308 50428 28318 50484
rect 28578 50428 28588 50484
rect 28644 50428 29932 50484
rect 29988 50428 30716 50484
rect 30772 50428 30940 50484
rect 30996 50428 31006 50484
rect 50754 50428 50764 50484
rect 50820 50428 51548 50484
rect 51604 50428 51614 50484
rect 54562 50428 54572 50484
rect 54628 50428 55244 50484
rect 55300 50428 57932 50484
rect 57988 50428 57998 50484
rect 18386 50316 18396 50372
rect 18452 50316 21532 50372
rect 21588 50316 23324 50372
rect 23380 50316 23390 50372
rect 40338 50316 40348 50372
rect 40404 50316 41244 50372
rect 41300 50316 41310 50372
rect 50988 50260 51044 50428
rect 59200 50260 60000 50288
rect 50978 50204 50988 50260
rect 51044 50204 51054 50260
rect 57362 50204 57372 50260
rect 57428 50204 58156 50260
rect 58212 50204 60000 50260
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 59200 50176 60000 50204
rect 26226 50092 26236 50148
rect 26292 50092 26908 50148
rect 26964 50092 26974 50148
rect 35634 49980 35644 50036
rect 35700 49980 37100 50036
rect 37156 49980 57484 50036
rect 57540 49980 57550 50036
rect 35522 49868 35532 49924
rect 35588 49868 37660 49924
rect 37716 49868 43708 49924
rect 48962 49868 48972 49924
rect 49028 49868 50204 49924
rect 50260 49868 50270 49924
rect 55794 49868 55804 49924
rect 55860 49868 56588 49924
rect 56644 49868 56654 49924
rect 43652 49812 43708 49868
rect 14354 49756 14364 49812
rect 14420 49756 15372 49812
rect 15428 49756 15438 49812
rect 24546 49756 24556 49812
rect 24612 49756 25676 49812
rect 25732 49756 25742 49812
rect 30706 49756 30716 49812
rect 30772 49756 31948 49812
rect 32004 49756 32014 49812
rect 38546 49756 38556 49812
rect 38612 49756 40908 49812
rect 40964 49756 40974 49812
rect 41122 49756 41132 49812
rect 41188 49756 41198 49812
rect 43652 49756 57596 49812
rect 57652 49756 57662 49812
rect 25330 49644 25340 49700
rect 25396 49644 26124 49700
rect 26180 49644 26572 49700
rect 26628 49644 26638 49700
rect 29922 49644 29932 49700
rect 29988 49644 31276 49700
rect 31332 49644 31342 49700
rect 26310 49532 26348 49588
rect 26404 49532 26414 49588
rect 36642 49532 36652 49588
rect 36708 49532 37436 49588
rect 37492 49532 37502 49588
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 41132 49364 41188 49756
rect 49298 49532 49308 49588
rect 49364 49532 51548 49588
rect 51604 49532 51614 49588
rect 46050 49420 46060 49476
rect 46116 49420 46956 49476
rect 47012 49420 47022 49476
rect 25890 49308 25900 49364
rect 25956 49308 26348 49364
rect 26404 49308 26414 49364
rect 39666 49308 39676 49364
rect 39732 49308 41804 49364
rect 41860 49308 41870 49364
rect 37538 49196 37548 49252
rect 37604 49196 39116 49252
rect 39172 49196 39182 49252
rect 56690 49196 56700 49252
rect 56756 49196 58156 49252
rect 58212 49196 58222 49252
rect 18946 49084 18956 49140
rect 19012 49084 19964 49140
rect 20020 49084 20030 49140
rect 28018 48972 28028 49028
rect 28084 48972 30268 49028
rect 30324 48972 30334 49028
rect 20738 48860 20748 48916
rect 20804 48860 21644 48916
rect 21700 48860 22092 48916
rect 22148 48860 22158 48916
rect 27794 48860 27804 48916
rect 27860 48860 29820 48916
rect 29876 48860 29886 48916
rect 38536 48860 38556 48916
rect 38612 48804 38668 49196
rect 39554 48972 39564 49028
rect 39620 48972 40348 49028
rect 40404 48972 40414 49028
rect 40786 48972 40796 49028
rect 40852 48972 42364 49028
rect 42420 48972 42430 49028
rect 43586 48972 43596 49028
rect 43652 48972 45388 49028
rect 45444 48972 45454 49028
rect 43362 48860 43372 48916
rect 43428 48860 44044 48916
rect 44100 48860 44110 48916
rect 43372 48804 43428 48860
rect 8082 48748 8092 48804
rect 8148 48748 10444 48804
rect 10500 48748 10510 48804
rect 19628 48748 19740 48804
rect 19796 48748 19806 48804
rect 20066 48748 20076 48804
rect 20132 48748 21420 48804
rect 21476 48748 22876 48804
rect 22932 48748 22942 48804
rect 31938 48748 31948 48804
rect 32004 48748 34692 48804
rect 38612 48748 38836 48804
rect 39778 48748 39788 48804
rect 39844 48748 40572 48804
rect 40628 48748 40638 48804
rect 41458 48748 41468 48804
rect 41524 48748 42364 48804
rect 42420 48748 42430 48804
rect 42690 48748 42700 48804
rect 42756 48748 43428 48804
rect 19628 48468 19684 48748
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 34636 48580 34692 48748
rect 38780 48692 38836 48748
rect 38770 48636 38780 48692
rect 38836 48636 38846 48692
rect 44258 48636 44268 48692
rect 44324 48636 45612 48692
rect 45668 48636 45678 48692
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 34626 48524 34636 48580
rect 34692 48524 34702 48580
rect 40114 48524 40124 48580
rect 40180 48524 47180 48580
rect 47236 48524 47246 48580
rect 19628 48412 21644 48468
rect 21700 48412 22540 48468
rect 22596 48412 22606 48468
rect 36306 48412 36316 48468
rect 36372 48412 37212 48468
rect 37268 48412 37278 48468
rect 46050 48412 46060 48468
rect 46116 48412 48132 48468
rect 48076 48356 48132 48412
rect 8306 48300 8316 48356
rect 8372 48300 9548 48356
rect 9604 48300 9614 48356
rect 34738 48300 34748 48356
rect 34804 48300 36204 48356
rect 36260 48300 36270 48356
rect 40674 48300 40684 48356
rect 40740 48300 42476 48356
rect 42532 48300 42542 48356
rect 46162 48300 46172 48356
rect 46228 48300 47292 48356
rect 47348 48300 47852 48356
rect 47908 48300 47918 48356
rect 48066 48300 48076 48356
rect 48132 48300 49532 48356
rect 49588 48300 49598 48356
rect 26786 48188 26796 48244
rect 26852 48188 29036 48244
rect 29092 48188 29102 48244
rect 34402 48188 34412 48244
rect 34468 48188 35084 48244
rect 35140 48188 35150 48244
rect 37202 48188 37212 48244
rect 37268 48188 38332 48244
rect 38388 48188 39676 48244
rect 39732 48188 39742 48244
rect 40338 48188 40348 48244
rect 40404 48188 40414 48244
rect 43250 48188 43260 48244
rect 43316 48188 43820 48244
rect 43876 48188 43886 48244
rect 44930 48188 44940 48244
rect 44996 48188 46956 48244
rect 47012 48188 47516 48244
rect 47572 48188 47582 48244
rect 40348 48132 40404 48188
rect 6850 48076 6860 48132
rect 6916 48076 9660 48132
rect 9716 48076 9726 48132
rect 14690 48076 14700 48132
rect 14756 48076 15932 48132
rect 15988 48076 15998 48132
rect 32274 48076 32284 48132
rect 32340 48076 33292 48132
rect 33348 48076 37100 48132
rect 37156 48076 37166 48132
rect 37538 48076 37548 48132
rect 37604 48076 39340 48132
rect 39396 48076 39406 48132
rect 40348 48076 44268 48132
rect 44324 48076 44334 48132
rect 45266 48076 45276 48132
rect 45332 48076 45948 48132
rect 46004 48076 46014 48132
rect 37100 48020 37156 48076
rect 37100 47964 37884 48020
rect 37940 47964 37950 48020
rect 40226 47964 40236 48020
rect 40292 47964 41244 48020
rect 41300 47964 41310 48020
rect 38322 47852 38332 47908
rect 38388 47852 43036 47908
rect 43092 47852 43102 47908
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 47170 47740 47180 47796
rect 47236 47740 52444 47796
rect 52500 47740 52510 47796
rect 16034 47628 16044 47684
rect 16100 47628 17612 47684
rect 17668 47628 32060 47684
rect 32116 47628 32126 47684
rect 38668 47628 44492 47684
rect 44548 47628 44558 47684
rect 38668 47572 38724 47628
rect 6178 47516 6188 47572
rect 6244 47516 6972 47572
rect 7028 47516 7038 47572
rect 28578 47516 28588 47572
rect 28644 47516 30380 47572
rect 30436 47516 30446 47572
rect 33954 47516 33964 47572
rect 34020 47516 36092 47572
rect 36148 47516 36158 47572
rect 38658 47516 38668 47572
rect 38724 47516 38734 47572
rect 43652 47516 45836 47572
rect 45892 47516 45902 47572
rect 50642 47516 50652 47572
rect 50708 47516 51100 47572
rect 51156 47516 52556 47572
rect 52612 47516 52622 47572
rect 11330 47404 11340 47460
rect 11396 47404 14588 47460
rect 14644 47404 14654 47460
rect 17042 47404 17052 47460
rect 17108 47404 17500 47460
rect 17556 47404 17948 47460
rect 18004 47404 18620 47460
rect 18676 47404 18686 47460
rect 19954 47404 19964 47460
rect 20020 47404 21532 47460
rect 21588 47404 21598 47460
rect 13458 47292 13468 47348
rect 13524 47292 15260 47348
rect 15316 47292 15820 47348
rect 15876 47292 15886 47348
rect 23062 47292 23100 47348
rect 23156 47292 23166 47348
rect 36306 47292 36316 47348
rect 36372 47292 36382 47348
rect 43586 47292 43596 47348
rect 43652 47292 43708 47516
rect 49858 47292 49868 47348
rect 49924 47292 53900 47348
rect 53956 47292 53966 47348
rect 55570 47292 55580 47348
rect 55636 47292 56364 47348
rect 56420 47292 56430 47348
rect 10434 47180 10444 47236
rect 10500 47180 11004 47236
rect 11060 47180 11070 47236
rect 16258 47180 16268 47236
rect 16324 47180 16940 47236
rect 16996 47180 17006 47236
rect 17378 47180 17388 47236
rect 17444 47180 17948 47236
rect 18004 47180 20188 47236
rect 20244 47180 21196 47236
rect 21252 47180 21262 47236
rect 21746 47180 21756 47236
rect 21812 47180 22876 47236
rect 22932 47180 24108 47236
rect 24164 47180 24174 47236
rect 36316 47124 36372 47292
rect 51986 47180 51996 47236
rect 52052 47180 52780 47236
rect 52836 47180 52846 47236
rect 21522 47068 21532 47124
rect 21588 47068 23212 47124
rect 23268 47068 23278 47124
rect 36316 47068 37436 47124
rect 37492 47068 38108 47124
rect 38164 47068 38174 47124
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 37090 46956 37100 47012
rect 37156 46956 39900 47012
rect 39956 46956 39966 47012
rect 54226 46956 54236 47012
rect 54292 46956 55692 47012
rect 55748 46956 55758 47012
rect 22642 46844 22652 46900
rect 22708 46844 26460 46900
rect 26516 46844 28588 46900
rect 28644 46844 28654 46900
rect 37202 46844 37212 46900
rect 37268 46844 39228 46900
rect 39284 46844 39294 46900
rect 18610 46732 18620 46788
rect 18676 46732 33068 46788
rect 33124 46732 33740 46788
rect 33796 46732 41132 46788
rect 41188 46732 41198 46788
rect 52098 46732 52108 46788
rect 52164 46732 53004 46788
rect 53060 46732 53070 46788
rect 55458 46732 55468 46788
rect 55524 46732 57036 46788
rect 57092 46732 57102 46788
rect 18722 46620 18732 46676
rect 18788 46620 19628 46676
rect 19684 46620 24332 46676
rect 24388 46620 25228 46676
rect 25284 46620 25294 46676
rect 25778 46620 25788 46676
rect 25844 46620 25854 46676
rect 26898 46620 26908 46676
rect 26964 46620 28364 46676
rect 28420 46620 28430 46676
rect 29698 46620 29708 46676
rect 29764 46620 31500 46676
rect 31556 46620 31566 46676
rect 33394 46620 33404 46676
rect 33460 46620 38444 46676
rect 38500 46620 38510 46676
rect 41570 46620 41580 46676
rect 41636 46620 46172 46676
rect 46228 46620 46238 46676
rect 50306 46620 50316 46676
rect 50372 46620 50540 46676
rect 50596 46620 50606 46676
rect 52770 46620 52780 46676
rect 52836 46620 55244 46676
rect 55300 46620 56420 46676
rect 56690 46620 56700 46676
rect 56756 46620 57260 46676
rect 57316 46620 57326 46676
rect 6290 46508 6300 46564
rect 6356 46508 7644 46564
rect 7700 46508 7710 46564
rect 25788 46452 25844 46620
rect 56364 46564 56420 46620
rect 26114 46508 26124 46564
rect 26180 46508 26796 46564
rect 26852 46508 26862 46564
rect 46610 46508 46620 46564
rect 46676 46508 55356 46564
rect 55412 46508 55422 46564
rect 56364 46508 57540 46564
rect 15026 46396 15036 46452
rect 15092 46396 16156 46452
rect 16212 46396 16222 46452
rect 25788 46396 26908 46452
rect 26964 46396 26974 46452
rect 49634 46396 49644 46452
rect 49700 46396 53116 46452
rect 53172 46396 53182 46452
rect 37314 46284 37324 46340
rect 37380 46284 38220 46340
rect 38276 46284 38286 46340
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 57484 46116 57540 46508
rect 18610 46060 18620 46116
rect 18676 46060 21420 46116
rect 21476 46060 33292 46116
rect 33348 46060 33358 46116
rect 57474 46060 57484 46116
rect 57540 46060 57550 46116
rect 7186 45948 7196 46004
rect 7252 45948 7980 46004
rect 8036 45948 8046 46004
rect 36194 45948 36204 46004
rect 36260 45948 37100 46004
rect 37156 45948 40460 46004
rect 40516 45948 43148 46004
rect 43204 45948 43214 46004
rect 4162 45836 4172 45892
rect 4228 45836 6748 45892
rect 6804 45836 9548 45892
rect 9604 45836 9614 45892
rect 21746 45836 21756 45892
rect 21812 45836 24108 45892
rect 24164 45836 24174 45892
rect 53442 45836 53452 45892
rect 53508 45836 54348 45892
rect 54404 45836 55468 45892
rect 11666 45724 11676 45780
rect 11732 45724 12572 45780
rect 12628 45724 12638 45780
rect 14242 45724 14252 45780
rect 14308 45724 15260 45780
rect 15316 45724 19516 45780
rect 19572 45724 19582 45780
rect 23426 45724 23436 45780
rect 23492 45724 25564 45780
rect 25620 45724 25630 45780
rect 43474 45724 43484 45780
rect 43540 45724 44044 45780
rect 44100 45724 44110 45780
rect 53330 45724 53340 45780
rect 53396 45724 53900 45780
rect 53956 45724 54796 45780
rect 54852 45724 54862 45780
rect 55412 45668 55468 45836
rect 12674 45612 12684 45668
rect 12740 45612 13244 45668
rect 13300 45612 14700 45668
rect 14756 45612 14766 45668
rect 49410 45612 49420 45668
rect 49476 45612 50540 45668
rect 50596 45612 50606 45668
rect 53666 45612 53676 45668
rect 53732 45612 54572 45668
rect 54628 45612 54638 45668
rect 55412 45612 56588 45668
rect 56644 45612 56654 45668
rect 7410 45500 7420 45556
rect 7476 45500 7756 45556
rect 7812 45500 11340 45556
rect 11396 45500 13916 45556
rect 13972 45500 13982 45556
rect 23426 45500 23436 45556
rect 23492 45500 25340 45556
rect 25396 45500 25406 45556
rect 52882 45500 52892 45556
rect 52948 45500 54012 45556
rect 54068 45500 54078 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 28354 45388 28364 45444
rect 28420 45388 31388 45444
rect 31444 45388 31454 45444
rect 49858 45388 49868 45444
rect 49924 45388 49934 45444
rect 53554 45388 53564 45444
rect 53620 45388 54572 45444
rect 54628 45388 54638 45444
rect 49868 45332 49924 45388
rect 12450 45276 12460 45332
rect 12516 45276 13020 45332
rect 13076 45276 14364 45332
rect 14420 45276 14430 45332
rect 14690 45276 14700 45332
rect 14756 45276 15484 45332
rect 15540 45276 15550 45332
rect 26898 45276 26908 45332
rect 26964 45276 27692 45332
rect 27748 45276 27758 45332
rect 40562 45276 40572 45332
rect 40628 45276 41916 45332
rect 41972 45276 41982 45332
rect 44258 45276 44268 45332
rect 44324 45276 45388 45332
rect 45444 45276 47068 45332
rect 47124 45276 47134 45332
rect 49868 45276 50316 45332
rect 50372 45276 50382 45332
rect 50866 45276 50876 45332
rect 50932 45276 51548 45332
rect 51604 45276 51614 45332
rect 8530 45164 8540 45220
rect 8596 45164 9660 45220
rect 9716 45164 9726 45220
rect 14578 45164 14588 45220
rect 14644 45164 16660 45220
rect 23650 45164 23660 45220
rect 23716 45164 26348 45220
rect 26404 45164 27020 45220
rect 27076 45164 27086 45220
rect 34402 45164 34412 45220
rect 34468 45164 40124 45220
rect 40180 45164 40908 45220
rect 40964 45164 40974 45220
rect 50978 45164 50988 45220
rect 51044 45164 51884 45220
rect 51940 45164 52780 45220
rect 52836 45164 55244 45220
rect 55300 45164 55310 45220
rect 16604 45108 16660 45164
rect 8194 45052 8204 45108
rect 8260 45052 9884 45108
rect 9940 45052 9950 45108
rect 11218 45052 11228 45108
rect 11284 45052 12236 45108
rect 12292 45052 13020 45108
rect 13076 45052 13086 45108
rect 13346 45052 13356 45108
rect 13412 45052 14700 45108
rect 14756 45052 14766 45108
rect 15092 45052 15372 45108
rect 15428 45052 15438 45108
rect 16594 45052 16604 45108
rect 16660 45052 16670 45108
rect 22642 45052 22652 45108
rect 22708 45052 23772 45108
rect 23828 45052 23838 45108
rect 26450 45052 26460 45108
rect 26516 45052 28588 45108
rect 28644 45052 28654 45108
rect 29922 45052 29932 45108
rect 29988 45052 29998 45108
rect 53890 45052 53900 45108
rect 53956 45052 54236 45108
rect 54292 45052 54302 45108
rect 54898 45052 54908 45108
rect 54964 45052 56140 45108
rect 56196 45052 56206 45108
rect 15092 44996 15148 45052
rect 10546 44940 10556 44996
rect 10612 44940 12012 44996
rect 12068 44940 15148 44996
rect 19842 44828 19852 44884
rect 19908 44828 20412 44884
rect 20468 44828 20478 44884
rect 29932 44772 29988 45052
rect 32386 44940 32396 44996
rect 32452 44940 33740 44996
rect 33796 44940 33806 44996
rect 43026 44940 43036 44996
rect 43092 44940 43820 44996
rect 43876 44940 43886 44996
rect 48178 44940 48188 44996
rect 48244 44940 49084 44996
rect 49140 44940 49150 44996
rect 29932 44716 30380 44772
rect 30436 44716 30446 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 32274 44604 32284 44660
rect 32340 44604 33068 44660
rect 33124 44604 33134 44660
rect 34598 44492 34636 44548
rect 34692 44492 34702 44548
rect 51314 44492 51324 44548
rect 51380 44492 52108 44548
rect 52164 44492 52174 44548
rect 58258 44492 58268 44548
rect 58324 44492 58548 44548
rect 58492 44436 58548 44492
rect 59200 44436 60000 44464
rect 7634 44380 7644 44436
rect 7700 44380 8540 44436
rect 8596 44380 8606 44436
rect 10658 44380 10668 44436
rect 10724 44380 14252 44436
rect 14308 44380 18284 44436
rect 18340 44380 18350 44436
rect 37762 44380 37772 44436
rect 37828 44380 39564 44436
rect 39620 44380 39630 44436
rect 49746 44380 49756 44436
rect 49812 44380 50428 44436
rect 50484 44380 50494 44436
rect 57474 44380 57484 44436
rect 57540 44380 58156 44436
rect 58212 44380 58222 44436
rect 58492 44380 60000 44436
rect 7858 44268 7868 44324
rect 7924 44268 8316 44324
rect 8372 44212 8428 44324
rect 14130 44268 14140 44324
rect 14196 44268 16268 44324
rect 16324 44268 16334 44324
rect 22866 44268 22876 44324
rect 22932 44268 25788 44324
rect 25844 44268 25854 44324
rect 27682 44268 27692 44324
rect 27748 44268 30268 44324
rect 30324 44268 30334 44324
rect 42802 44268 42812 44324
rect 42868 44268 43820 44324
rect 43876 44268 43886 44324
rect 44034 44268 44044 44324
rect 44100 44268 47068 44324
rect 47124 44268 47134 44324
rect 49756 44212 49812 44380
rect 59200 44352 60000 44380
rect 50194 44268 50204 44324
rect 50260 44268 51772 44324
rect 51828 44268 51838 44324
rect 8372 44156 9548 44212
rect 9604 44156 9614 44212
rect 26450 44156 26460 44212
rect 26516 44156 27804 44212
rect 27860 44156 40572 44212
rect 40628 44156 40638 44212
rect 43138 44156 43148 44212
rect 43204 44156 49812 44212
rect 9090 44044 9100 44100
rect 9156 44044 9996 44100
rect 10052 44044 11116 44100
rect 11172 44044 11182 44100
rect 14802 44044 14812 44100
rect 14868 44044 16044 44100
rect 16100 44044 16110 44100
rect 42466 44044 42476 44100
rect 42532 44044 43260 44100
rect 43316 44044 43326 44100
rect 8418 43932 8428 43988
rect 8484 43932 9436 43988
rect 9492 43932 10220 43988
rect 10276 43932 10668 43988
rect 10724 43932 10734 43988
rect 30706 43932 30716 43988
rect 30772 43932 30782 43988
rect 54460 43932 56364 43988
rect 56420 43932 56430 43988
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 30716 43876 30772 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 54460 43876 54516 43932
rect 4722 43820 4732 43876
rect 4788 43820 8204 43876
rect 8260 43820 10108 43876
rect 10164 43820 10174 43876
rect 30716 43820 31164 43876
rect 31220 43820 43596 43876
rect 43652 43764 43708 43876
rect 54450 43820 54460 43876
rect 54516 43820 54526 43876
rect 55458 43820 55468 43876
rect 55524 43820 56924 43876
rect 56980 43820 56990 43876
rect 16594 43708 16604 43764
rect 16660 43708 17948 43764
rect 18004 43708 18014 43764
rect 33618 43708 33628 43764
rect 33684 43708 34636 43764
rect 34692 43708 34702 43764
rect 43652 43708 44268 43764
rect 44324 43708 44334 43764
rect 54562 43708 54572 43764
rect 54628 43708 55132 43764
rect 55188 43708 55692 43764
rect 55748 43708 55758 43764
rect 14690 43596 14700 43652
rect 14756 43596 15372 43652
rect 15428 43596 15438 43652
rect 16370 43596 16380 43652
rect 16436 43596 17388 43652
rect 17444 43596 18732 43652
rect 18788 43596 18798 43652
rect 23762 43596 23772 43652
rect 23828 43596 25452 43652
rect 25508 43596 25518 43652
rect 36306 43596 36316 43652
rect 36372 43596 38220 43652
rect 38276 43596 38286 43652
rect 38434 43596 38444 43652
rect 38500 43596 39340 43652
rect 39396 43596 39406 43652
rect 50082 43596 50092 43652
rect 50148 43596 52444 43652
rect 52500 43596 52510 43652
rect 7634 43484 7644 43540
rect 7700 43484 10332 43540
rect 10388 43484 10398 43540
rect 16380 43428 16436 43596
rect 30706 43484 30716 43540
rect 30772 43484 31276 43540
rect 31332 43484 31342 43540
rect 37538 43484 37548 43540
rect 37604 43484 38556 43540
rect 38612 43484 38622 43540
rect 42578 43484 42588 43540
rect 42644 43484 43260 43540
rect 43316 43484 43326 43540
rect 49410 43484 49420 43540
rect 49476 43484 50764 43540
rect 50820 43484 50830 43540
rect 10434 43372 10444 43428
rect 10500 43372 13580 43428
rect 13636 43372 16436 43428
rect 21410 43372 21420 43428
rect 21476 43372 35084 43428
rect 35140 43372 44716 43428
rect 44772 43372 45500 43428
rect 45556 43372 45566 43428
rect 25106 43260 25116 43316
rect 25172 43260 25564 43316
rect 25620 43260 25630 43316
rect 30818 43260 30828 43316
rect 30884 43260 32060 43316
rect 32116 43260 32126 43316
rect 32274 43260 32284 43316
rect 32340 43260 33180 43316
rect 33236 43260 42588 43316
rect 42644 43260 42654 43316
rect 56130 43260 56140 43316
rect 56196 43260 56924 43316
rect 56980 43260 56990 43316
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 38098 42924 38108 42980
rect 38164 42924 39004 42980
rect 39060 42924 39070 42980
rect 46722 42924 46732 42980
rect 46788 42924 49420 42980
rect 49476 42924 49486 42980
rect 26450 42812 26460 42868
rect 26516 42812 27244 42868
rect 27300 42812 27310 42868
rect 36418 42812 36428 42868
rect 36484 42812 37660 42868
rect 37716 42812 37726 42868
rect 14354 42700 14364 42756
rect 14420 42700 15820 42756
rect 15876 42700 15886 42756
rect 20738 42700 20748 42756
rect 20804 42700 21420 42756
rect 21476 42700 21486 42756
rect 29922 42700 29932 42756
rect 29988 42700 30828 42756
rect 30884 42700 30894 42756
rect 31266 42700 31276 42756
rect 31332 42700 31342 42756
rect 43250 42700 43260 42756
rect 43316 42700 43596 42756
rect 43652 42700 43662 42756
rect 49746 42700 49756 42756
rect 49812 42700 51324 42756
rect 51380 42700 52892 42756
rect 52948 42700 52958 42756
rect 31276 42644 31332 42700
rect 29250 42588 29260 42644
rect 29316 42588 30940 42644
rect 30996 42588 31006 42644
rect 31164 42588 31332 42644
rect 45490 42588 45500 42644
rect 45556 42588 46172 42644
rect 46228 42588 46238 42644
rect 51762 42588 51772 42644
rect 51828 42588 52780 42644
rect 52836 42588 52846 42644
rect 31164 42532 31220 42588
rect 12674 42476 12684 42532
rect 12740 42476 13916 42532
rect 13972 42476 13982 42532
rect 21186 42476 21196 42532
rect 21252 42476 21980 42532
rect 22036 42476 22046 42532
rect 30482 42476 30492 42532
rect 30548 42476 31220 42532
rect 37874 42476 37884 42532
rect 37940 42476 38668 42532
rect 38724 42476 44940 42532
rect 44996 42476 45006 42532
rect 37650 42364 37660 42420
rect 37716 42364 38332 42420
rect 38388 42364 38668 42420
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 38612 42308 38668 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 38612 42252 39564 42308
rect 39620 42252 39630 42308
rect 25330 42140 25340 42196
rect 25396 42140 25676 42196
rect 25732 42140 25742 42196
rect 35410 42140 35420 42196
rect 35476 42140 37772 42196
rect 37828 42140 37838 42196
rect 38994 42140 39004 42196
rect 39060 42140 43484 42196
rect 43540 42140 44828 42196
rect 44884 42140 45276 42196
rect 45332 42140 45342 42196
rect 14466 42028 14476 42084
rect 14532 42028 15820 42084
rect 15876 42028 15886 42084
rect 26002 42028 26012 42084
rect 26068 42028 27692 42084
rect 27748 42028 27758 42084
rect 32274 42028 32284 42084
rect 32340 42028 33684 42084
rect 44370 42028 44380 42084
rect 44436 42028 45164 42084
rect 45220 42028 47964 42084
rect 48020 42028 51548 42084
rect 51604 42028 51614 42084
rect 10322 41916 10332 41972
rect 10388 41916 11340 41972
rect 11396 41916 12012 41972
rect 12068 41916 12078 41972
rect 15092 41916 15372 41972
rect 15428 41916 15438 41972
rect 22082 41916 22092 41972
rect 22148 41916 23996 41972
rect 24052 41916 24062 41972
rect 24210 41916 24220 41972
rect 24276 41916 24668 41972
rect 24724 41916 25788 41972
rect 25844 41916 25854 41972
rect 26226 41916 26236 41972
rect 26292 41916 26908 41972
rect 26964 41916 26974 41972
rect 27234 41916 27244 41972
rect 27300 41916 29372 41972
rect 29428 41916 29438 41972
rect 30482 41916 30492 41972
rect 30548 41916 32396 41972
rect 32452 41916 32462 41972
rect 15092 41748 15148 41916
rect 33628 41860 33684 42028
rect 34290 41916 34300 41972
rect 34356 41916 35308 41972
rect 35364 41916 35374 41972
rect 37202 41916 37212 41972
rect 37268 41916 37996 41972
rect 38052 41916 38062 41972
rect 48962 41916 48972 41972
rect 49028 41916 51884 41972
rect 51940 41916 51950 41972
rect 55122 41916 55132 41972
rect 55188 41916 55580 41972
rect 55636 41916 55646 41972
rect 56802 41916 56812 41972
rect 56868 41916 58156 41972
rect 58212 41916 58222 41972
rect 23314 41804 23324 41860
rect 23380 41804 23772 41860
rect 23828 41804 23838 41860
rect 28466 41804 28476 41860
rect 28532 41804 31388 41860
rect 31444 41804 31836 41860
rect 31892 41804 31902 41860
rect 32274 41804 32284 41860
rect 32340 41804 33068 41860
rect 33124 41804 33134 41860
rect 33618 41804 33628 41860
rect 33684 41804 35868 41860
rect 35924 41804 35934 41860
rect 47506 41804 47516 41860
rect 47572 41804 50764 41860
rect 50820 41804 50830 41860
rect 51762 41804 51772 41860
rect 51828 41804 53340 41860
rect 53396 41804 53406 41860
rect 10098 41692 10108 41748
rect 10164 41692 11340 41748
rect 11396 41692 15148 41748
rect 23874 41692 23884 41748
rect 23940 41692 24444 41748
rect 24500 41692 26124 41748
rect 26180 41692 26190 41748
rect 37762 41692 37772 41748
rect 37828 41692 38556 41748
rect 38612 41692 38622 41748
rect 48066 41692 48076 41748
rect 48132 41692 49084 41748
rect 49140 41692 49150 41748
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 19842 41356 19852 41412
rect 19908 41356 24108 41412
rect 24164 41356 25340 41412
rect 25396 41356 25406 41412
rect 17602 41244 17612 41300
rect 17668 41244 26012 41300
rect 26068 41244 26078 41300
rect 37314 41244 37324 41300
rect 37380 41244 40908 41300
rect 40964 41244 40974 41300
rect 16370 41132 16380 41188
rect 16436 41132 17500 41188
rect 17556 41132 18508 41188
rect 18564 41132 18574 41188
rect 25778 41132 25788 41188
rect 25844 41132 27468 41188
rect 27524 41132 27534 41188
rect 43698 41132 43708 41188
rect 43764 41132 44492 41188
rect 44548 41132 51212 41188
rect 51268 41132 51660 41188
rect 51716 41132 52332 41188
rect 52388 41132 52398 41188
rect 26338 41020 26348 41076
rect 26404 41020 26684 41076
rect 26740 41020 28140 41076
rect 28196 41020 28206 41076
rect 29026 41020 29036 41076
rect 29092 41020 29484 41076
rect 29540 41020 30156 41076
rect 30212 41020 30222 41076
rect 36418 41020 36428 41076
rect 36484 41020 37100 41076
rect 37156 41020 37166 41076
rect 29036 40964 29092 41020
rect 25890 40908 25900 40964
rect 25956 40908 26908 40964
rect 26964 40908 26974 40964
rect 27794 40908 27804 40964
rect 27860 40908 29092 40964
rect 42354 40908 42364 40964
rect 42420 40908 43820 40964
rect 43876 40908 43886 40964
rect 45714 40908 45724 40964
rect 45780 40908 48748 40964
rect 48804 40908 49308 40964
rect 49364 40908 49374 40964
rect 51874 40908 51884 40964
rect 51940 40908 52556 40964
rect 52612 40908 52622 40964
rect 28690 40796 28700 40852
rect 28756 40796 29260 40852
rect 29316 40796 40348 40852
rect 40404 40796 40908 40852
rect 40964 40796 40974 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 4946 40572 4956 40628
rect 5012 40572 9660 40628
rect 9716 40572 10444 40628
rect 10500 40572 10510 40628
rect 15250 40572 15260 40628
rect 15316 40572 16604 40628
rect 16660 40572 16670 40628
rect 18946 40572 18956 40628
rect 19012 40572 19628 40628
rect 19684 40572 19694 40628
rect 52322 40572 52332 40628
rect 52388 40572 52780 40628
rect 52836 40572 54236 40628
rect 54292 40572 55692 40628
rect 55748 40572 55758 40628
rect 1810 40460 1820 40516
rect 1876 40460 8316 40516
rect 8372 40460 8428 40516
rect 8484 40460 8494 40516
rect 24770 40460 24780 40516
rect 24836 40460 26012 40516
rect 26068 40460 26078 40516
rect 50082 40460 50092 40516
rect 50148 40460 53676 40516
rect 53732 40460 53742 40516
rect 14242 40348 14252 40404
rect 14308 40348 16156 40404
rect 16212 40348 16222 40404
rect 16594 40348 16604 40404
rect 16660 40348 17500 40404
rect 17556 40348 17566 40404
rect 25330 40348 25340 40404
rect 25396 40348 29036 40404
rect 29092 40348 29102 40404
rect 34290 40348 34300 40404
rect 34356 40348 35756 40404
rect 35812 40348 37324 40404
rect 37380 40348 37390 40404
rect 46050 40348 46060 40404
rect 46116 40348 47516 40404
rect 47572 40348 47582 40404
rect 50418 40348 50428 40404
rect 50484 40348 51884 40404
rect 51940 40348 52668 40404
rect 52724 40348 52734 40404
rect 53218 40348 53228 40404
rect 53284 40348 54460 40404
rect 54516 40348 54526 40404
rect 56130 40348 56140 40404
rect 56196 40348 56206 40404
rect 56140 40292 56196 40348
rect 12786 40236 12796 40292
rect 12852 40236 16492 40292
rect 16548 40236 16558 40292
rect 17266 40236 17276 40292
rect 17332 40236 18172 40292
rect 18228 40236 18620 40292
rect 18676 40236 19068 40292
rect 19124 40236 19134 40292
rect 24434 40236 24444 40292
rect 24500 40236 25004 40292
rect 25060 40236 25070 40292
rect 39890 40236 39900 40292
rect 39956 40236 40908 40292
rect 40964 40236 40974 40292
rect 41906 40236 41916 40292
rect 41972 40236 42588 40292
rect 42644 40236 43484 40292
rect 43540 40236 43550 40292
rect 46274 40236 46284 40292
rect 46340 40236 46620 40292
rect 46676 40236 46956 40292
rect 47012 40236 47022 40292
rect 49746 40236 49756 40292
rect 49812 40236 53452 40292
rect 53508 40236 55244 40292
rect 55300 40236 56196 40292
rect 57586 40236 57596 40292
rect 57652 40236 58044 40292
rect 58100 40236 58110 40292
rect 20402 40124 20412 40180
rect 20468 40124 20860 40180
rect 20916 40124 24556 40180
rect 24612 40124 24622 40180
rect 39106 40124 39116 40180
rect 39172 40124 41244 40180
rect 41300 40124 41692 40180
rect 41748 40124 41758 40180
rect 52210 40124 52220 40180
rect 52276 40124 52892 40180
rect 52948 40124 52958 40180
rect 54786 40124 54796 40180
rect 54852 40124 57484 40180
rect 57540 40124 58268 40180
rect 58324 40124 58334 40180
rect 44146 40012 44156 40068
rect 44212 40012 54348 40068
rect 54404 40012 54414 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 36978 39900 36988 39956
rect 37044 39900 38556 39956
rect 38612 39900 52108 39956
rect 52164 39900 52174 39956
rect 21522 39788 21532 39844
rect 21588 39788 22316 39844
rect 22372 39788 22382 39844
rect 29698 39788 29708 39844
rect 29764 39788 30268 39844
rect 30324 39788 45388 39844
rect 45444 39788 45454 39844
rect 48738 39788 48748 39844
rect 48804 39788 49980 39844
rect 50036 39788 50046 39844
rect 22418 39676 22428 39732
rect 22484 39676 24332 39732
rect 24388 39676 24398 39732
rect 52658 39676 52668 39732
rect 52724 39676 53676 39732
rect 53732 39676 54908 39732
rect 54964 39676 54974 39732
rect 17154 39564 17164 39620
rect 17220 39564 17836 39620
rect 17892 39564 23884 39620
rect 23940 39564 23950 39620
rect 24210 39564 24220 39620
rect 24276 39564 24556 39620
rect 24612 39564 25340 39620
rect 25396 39564 26908 39620
rect 26964 39564 27916 39620
rect 27972 39564 27982 39620
rect 41346 39564 41356 39620
rect 41412 39564 42140 39620
rect 42196 39564 43820 39620
rect 43876 39564 43886 39620
rect 52882 39564 52892 39620
rect 52948 39564 55244 39620
rect 55300 39564 55310 39620
rect 23884 39508 23940 39564
rect 16930 39452 16940 39508
rect 16996 39452 18844 39508
rect 18900 39452 18910 39508
rect 23884 39452 24444 39508
rect 24500 39452 24510 39508
rect 24882 39452 24892 39508
rect 24948 39452 26012 39508
rect 26068 39452 26078 39508
rect 43586 39452 43596 39508
rect 43652 39452 54908 39508
rect 54964 39452 54974 39508
rect 7298 39340 7308 39396
rect 7364 39340 9324 39396
rect 9380 39340 9390 39396
rect 14802 39340 14812 39396
rect 14868 39340 17052 39396
rect 17108 39340 17118 39396
rect 21970 39340 21980 39396
rect 22036 39340 29148 39396
rect 29204 39340 30604 39396
rect 30660 39340 30670 39396
rect 35298 39340 35308 39396
rect 35364 39340 36316 39396
rect 36372 39340 42364 39396
rect 42420 39340 43148 39396
rect 43204 39340 43214 39396
rect 49410 39340 49420 39396
rect 49476 39340 54572 39396
rect 54628 39340 54638 39396
rect 34066 39228 34076 39284
rect 34132 39228 34524 39284
rect 34580 39228 36652 39284
rect 36708 39228 36718 39284
rect 47842 39228 47852 39284
rect 47908 39228 48748 39284
rect 48804 39228 48814 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 8372 39116 8540 39172
rect 8596 39116 11004 39172
rect 11060 39116 11070 39172
rect 24434 39116 24444 39172
rect 24500 39116 38668 39172
rect 38724 39116 40460 39172
rect 40516 39116 40526 39172
rect 43652 39116 50484 39172
rect 54562 39116 54572 39172
rect 54628 39116 55804 39172
rect 55860 39116 55870 39172
rect 5282 39004 5292 39060
rect 5348 39004 6580 39060
rect 2482 38892 2492 38948
rect 2548 38892 6356 38948
rect 6300 38836 6356 38892
rect 5730 38780 5740 38836
rect 5796 38780 5806 38836
rect 6290 38780 6300 38836
rect 6356 38780 6366 38836
rect 5740 38612 5796 38780
rect 6524 38724 6580 39004
rect 8372 38836 8428 39116
rect 43652 39060 43708 39116
rect 50428 39060 50484 39116
rect 8866 39004 8876 39060
rect 8932 39004 8942 39060
rect 32508 39004 35756 39060
rect 35812 39004 35822 39060
rect 36642 39004 36652 39060
rect 36708 39004 37212 39060
rect 37268 39004 37884 39060
rect 37940 39004 37950 39060
rect 38612 39004 43708 39060
rect 43922 39004 43932 39060
rect 43988 39004 46844 39060
rect 46900 39004 49084 39060
rect 49140 39004 49150 39060
rect 50428 39004 52668 39060
rect 52724 39004 53116 39060
rect 53172 39004 53182 39060
rect 55458 39004 55468 39060
rect 55524 39004 55916 39060
rect 55972 39004 57820 39060
rect 57876 39004 57886 39060
rect 8876 38836 8932 39004
rect 32508 38948 32564 39004
rect 38612 38948 38668 39004
rect 23090 38892 23100 38948
rect 23156 38892 26796 38948
rect 26852 38892 32508 38948
rect 32564 38892 32574 38948
rect 33394 38892 33404 38948
rect 33460 38892 34860 38948
rect 34916 38892 34926 38948
rect 37212 38892 38668 38948
rect 45724 38892 46620 38948
rect 46676 38892 47516 38948
rect 47572 38892 47582 38948
rect 6738 38780 6748 38836
rect 6804 38780 7196 38836
rect 7252 38780 8428 38836
rect 8652 38780 8932 38836
rect 12562 38780 12572 38836
rect 12628 38780 13468 38836
rect 13524 38780 13534 38836
rect 18498 38780 18508 38836
rect 18564 38780 19180 38836
rect 19236 38780 19246 38836
rect 33954 38780 33964 38836
rect 34020 38780 34748 38836
rect 34804 38780 36988 38836
rect 37044 38780 37054 38836
rect 8652 38724 8708 38780
rect 37212 38724 37268 38892
rect 45724 38836 45780 38892
rect 37874 38780 37884 38836
rect 37940 38780 39228 38836
rect 39284 38780 39294 38836
rect 40226 38780 40236 38836
rect 40292 38780 43932 38836
rect 43988 38780 43998 38836
rect 45714 38780 45724 38836
rect 45780 38780 45790 38836
rect 46274 38780 46284 38836
rect 46340 38780 48860 38836
rect 48916 38780 48926 38836
rect 6524 38668 7532 38724
rect 7588 38668 8204 38724
rect 8260 38668 8708 38724
rect 8866 38668 8876 38724
rect 8932 38668 11676 38724
rect 11732 38668 11742 38724
rect 18050 38668 18060 38724
rect 18116 38668 18844 38724
rect 18900 38668 18910 38724
rect 19058 38668 19068 38724
rect 19124 38668 20076 38724
rect 20132 38668 23436 38724
rect 23492 38668 26964 38724
rect 27570 38668 27580 38724
rect 27636 38668 30380 38724
rect 30436 38668 30446 38724
rect 31602 38668 31612 38724
rect 31668 38668 37268 38724
rect 47730 38668 47740 38724
rect 47796 38668 52108 38724
rect 52164 38668 52174 38724
rect 58146 38668 58156 38724
rect 58212 38668 58222 38724
rect 26908 38612 26964 38668
rect 58156 38612 58212 38668
rect 59200 38612 60000 38640
rect 5740 38556 7756 38612
rect 7812 38556 7822 38612
rect 17042 38556 17052 38612
rect 17108 38556 17948 38612
rect 18004 38556 18014 38612
rect 26908 38556 27020 38612
rect 27076 38556 27086 38612
rect 32498 38556 32508 38612
rect 32564 38556 33180 38612
rect 33236 38556 33246 38612
rect 58156 38556 60000 38612
rect 59200 38528 60000 38556
rect 5170 38444 5180 38500
rect 5236 38444 6188 38500
rect 6244 38444 6254 38500
rect 43698 38444 43708 38500
rect 43764 38444 47404 38500
rect 47460 38444 47964 38500
rect 48020 38444 48030 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 43810 38332 43820 38388
rect 43876 38332 45052 38388
rect 45108 38332 45118 38388
rect 37538 38220 37548 38276
rect 37604 38220 54460 38276
rect 54516 38220 54526 38276
rect 2482 38108 2492 38164
rect 2548 38108 5852 38164
rect 5908 38108 5918 38164
rect 21186 38108 21196 38164
rect 21252 38108 23660 38164
rect 23716 38108 23726 38164
rect 28018 38108 28028 38164
rect 28084 38108 30156 38164
rect 30212 38108 30222 38164
rect 34188 38108 34636 38164
rect 34692 38108 34702 38164
rect 43586 38108 43596 38164
rect 43652 38108 44268 38164
rect 44324 38108 57148 38164
rect 57204 38108 57214 38164
rect 34188 38052 34244 38108
rect 5618 37996 5628 38052
rect 5684 37996 6860 38052
rect 6916 37996 8876 38052
rect 8932 37996 9660 38052
rect 9716 37996 9726 38052
rect 34178 37996 34188 38052
rect 34244 37996 34254 38052
rect 35634 37996 35644 38052
rect 35700 37996 36316 38052
rect 36372 37996 36876 38052
rect 36932 37996 36942 38052
rect 48738 37996 48748 38052
rect 48804 37996 50540 38052
rect 50596 37996 51884 38052
rect 51940 37996 51950 38052
rect 28690 37884 28700 37940
rect 28756 37884 29260 37940
rect 29316 37884 29326 37940
rect 5170 37772 5180 37828
rect 5236 37772 6748 37828
rect 6804 37772 6814 37828
rect 23986 37772 23996 37828
rect 24052 37772 29036 37828
rect 29092 37772 29102 37828
rect 34598 37772 34636 37828
rect 34692 37772 34702 37828
rect 38098 37772 38108 37828
rect 38164 37772 39788 37828
rect 39844 37772 45948 37828
rect 46004 37772 47180 37828
rect 47236 37772 47246 37828
rect 27010 37660 27020 37716
rect 27076 37660 38668 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 38612 37604 38668 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 29250 37548 29260 37604
rect 29316 37548 35980 37604
rect 36036 37548 37548 37604
rect 37604 37548 38108 37604
rect 38164 37548 38174 37604
rect 38612 37548 42028 37604
rect 42084 37548 42094 37604
rect 48738 37548 48748 37604
rect 48804 37548 49756 37604
rect 49812 37548 49822 37604
rect 11666 37436 11676 37492
rect 11732 37436 12348 37492
rect 12404 37436 27580 37492
rect 27636 37436 27646 37492
rect 28690 37436 28700 37492
rect 28756 37436 29148 37492
rect 29204 37436 29214 37492
rect 31378 37436 31388 37492
rect 31444 37436 32060 37492
rect 32116 37436 32126 37492
rect 35522 37436 35532 37492
rect 35588 37436 36484 37492
rect 48178 37436 48188 37492
rect 48244 37436 48860 37492
rect 48916 37436 48926 37492
rect 36428 37268 36484 37436
rect 43474 37324 43484 37380
rect 43540 37324 43820 37380
rect 43876 37324 43886 37380
rect 12562 37212 12572 37268
rect 12628 37212 16492 37268
rect 16548 37212 16558 37268
rect 19506 37212 19516 37268
rect 19572 37212 20524 37268
rect 20580 37212 20590 37268
rect 22530 37212 22540 37268
rect 22596 37212 22988 37268
rect 23044 37212 23054 37268
rect 24098 37212 24108 37268
rect 24164 37212 28700 37268
rect 28756 37212 28766 37268
rect 29474 37212 29484 37268
rect 29540 37212 35476 37268
rect 35634 37212 35644 37268
rect 35700 37212 36204 37268
rect 36260 37212 36270 37268
rect 36418 37212 36428 37268
rect 36484 37212 37100 37268
rect 37156 37212 37166 37268
rect 54898 37212 54908 37268
rect 54964 37212 57820 37268
rect 57876 37212 57886 37268
rect 35420 37156 35476 37212
rect 19730 37100 19740 37156
rect 19796 37100 20188 37156
rect 20244 37100 20254 37156
rect 20626 37100 20636 37156
rect 20692 37100 23548 37156
rect 23604 37100 23614 37156
rect 30146 37100 30156 37156
rect 30212 37100 32396 37156
rect 32452 37100 32462 37156
rect 35420 37100 36316 37156
rect 36372 37100 36382 37156
rect 36866 37100 36876 37156
rect 36932 37100 38220 37156
rect 38276 37100 38286 37156
rect 48290 37100 48300 37156
rect 48356 37100 48972 37156
rect 49028 37100 49038 37156
rect 55234 37100 55244 37156
rect 55300 37100 56588 37156
rect 56644 37100 56654 37156
rect 7634 36988 7644 37044
rect 7700 36988 8652 37044
rect 8708 36988 8718 37044
rect 12114 36988 12124 37044
rect 12180 36988 31276 37044
rect 31332 36988 31342 37044
rect 31938 36988 31948 37044
rect 32004 36988 32620 37044
rect 32676 36988 33516 37044
rect 33572 36988 35868 37044
rect 35924 36988 35934 37044
rect 53106 36988 53116 37044
rect 53172 36988 53900 37044
rect 53956 36988 53966 37044
rect 54338 36988 54348 37044
rect 54404 36988 56700 37044
rect 56756 36988 56766 37044
rect 12124 36932 12180 36988
rect 10546 36876 10556 36932
rect 10612 36876 12180 36932
rect 38658 36876 38668 36932
rect 38724 36876 40012 36932
rect 40068 36876 40078 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 32386 36652 32396 36708
rect 32452 36652 33180 36708
rect 33236 36652 43484 36708
rect 43540 36652 44828 36708
rect 44884 36652 44894 36708
rect 34290 36540 34300 36596
rect 34356 36540 35756 36596
rect 35812 36540 35822 36596
rect 36306 36540 36316 36596
rect 36372 36540 43372 36596
rect 43428 36540 44716 36596
rect 44772 36540 44782 36596
rect 52098 36540 52108 36596
rect 52164 36540 52780 36596
rect 52836 36540 52846 36596
rect 55346 36540 55356 36596
rect 55412 36540 56028 36596
rect 56084 36540 56094 36596
rect 16034 36428 16044 36484
rect 16100 36428 16604 36484
rect 16660 36428 16670 36484
rect 25442 36428 25452 36484
rect 25508 36428 38668 36484
rect 44930 36428 44940 36484
rect 44996 36428 48748 36484
rect 48804 36428 48814 36484
rect 2482 36316 2492 36372
rect 2548 36316 4508 36372
rect 4564 36316 4574 36372
rect 14130 36316 14140 36372
rect 14196 36316 15148 36372
rect 15204 36316 15214 36372
rect 24994 36316 25004 36372
rect 25060 36316 26124 36372
rect 26180 36316 26190 36372
rect 26786 36316 26796 36372
rect 26852 36316 26908 36428
rect 38612 36372 38668 36428
rect 34962 36316 34972 36372
rect 35028 36316 35196 36372
rect 35252 36316 35262 36372
rect 35634 36316 35644 36372
rect 35700 36316 36316 36372
rect 36372 36316 36382 36372
rect 38612 36316 41580 36372
rect 41636 36316 41646 36372
rect 42690 36316 42700 36372
rect 42756 36316 46284 36372
rect 46340 36316 46844 36372
rect 46900 36316 46910 36372
rect 52882 36316 52892 36372
rect 52948 36316 54908 36372
rect 54964 36316 54974 36372
rect 4722 36204 4732 36260
rect 4788 36204 5516 36260
rect 5572 36204 5582 36260
rect 13234 36204 13244 36260
rect 13300 36204 13804 36260
rect 13860 36204 13870 36260
rect 20066 36204 20076 36260
rect 20132 36204 21196 36260
rect 21252 36204 21262 36260
rect 26562 36204 26572 36260
rect 26628 36204 27580 36260
rect 27636 36204 27646 36260
rect 33282 36204 33292 36260
rect 33348 36204 33964 36260
rect 34020 36204 37436 36260
rect 37492 36204 37502 36260
rect 43026 36204 43036 36260
rect 43092 36204 43820 36260
rect 43876 36204 43886 36260
rect 47170 36204 47180 36260
rect 47236 36204 49644 36260
rect 49700 36204 52668 36260
rect 52724 36204 54348 36260
rect 54404 36204 54414 36260
rect 26852 36092 31836 36148
rect 31892 36092 33068 36148
rect 33124 36092 33134 36148
rect 33842 36092 33852 36148
rect 33908 36092 33918 36148
rect 53106 36092 53116 36148
rect 53172 36092 54012 36148
rect 54068 36092 54796 36148
rect 54852 36092 54862 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 26852 35924 26908 36092
rect 33852 36036 33908 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 8082 35868 8092 35924
rect 8148 35868 8428 35924
rect 13346 35868 13356 35924
rect 13412 35868 14252 35924
rect 14308 35868 14924 35924
rect 14980 35868 26908 35924
rect 27244 35980 33908 36036
rect 8372 35812 8428 35868
rect 27244 35812 27300 35980
rect 28998 35868 29036 35924
rect 29092 35868 29102 35924
rect 4162 35756 4172 35812
rect 4228 35756 5068 35812
rect 5124 35756 5134 35812
rect 6066 35756 6076 35812
rect 6132 35756 7756 35812
rect 7812 35756 7822 35812
rect 8372 35756 8876 35812
rect 8932 35756 8942 35812
rect 15138 35756 15148 35812
rect 15204 35756 16268 35812
rect 16324 35756 16334 35812
rect 17490 35756 17500 35812
rect 17556 35756 27300 35812
rect 27682 35756 27692 35812
rect 27748 35756 30828 35812
rect 30884 35756 30894 35812
rect 38434 35756 38444 35812
rect 38500 35756 39452 35812
rect 39508 35756 39518 35812
rect 48962 35756 48972 35812
rect 49028 35756 51212 35812
rect 51268 35756 51278 35812
rect 55122 35756 55132 35812
rect 55188 35756 58156 35812
rect 58212 35756 58222 35812
rect 27692 35700 27748 35756
rect 4834 35644 4844 35700
rect 4900 35644 5516 35700
rect 5572 35644 5582 35700
rect 7522 35644 7532 35700
rect 7588 35644 8764 35700
rect 8820 35644 8830 35700
rect 9314 35644 9324 35700
rect 9380 35644 9884 35700
rect 9940 35644 9950 35700
rect 12674 35644 12684 35700
rect 12740 35644 13580 35700
rect 13636 35644 13646 35700
rect 14578 35644 14588 35700
rect 14644 35644 16156 35700
rect 16212 35644 16716 35700
rect 16772 35644 16782 35700
rect 26338 35644 26348 35700
rect 26404 35644 26414 35700
rect 26674 35644 26684 35700
rect 26740 35644 27748 35700
rect 31938 35644 31948 35700
rect 32004 35644 33068 35700
rect 33124 35644 36428 35700
rect 36484 35644 36494 35700
rect 38994 35644 39004 35700
rect 39060 35644 39676 35700
rect 39732 35644 39742 35700
rect 41570 35644 41580 35700
rect 41636 35644 42140 35700
rect 42196 35644 47516 35700
rect 47572 35644 47582 35700
rect 54674 35644 54684 35700
rect 54740 35644 56028 35700
rect 56084 35644 56094 35700
rect 13580 35588 13636 35644
rect 26348 35588 26404 35644
rect 13580 35532 15372 35588
rect 15428 35532 15438 35588
rect 26348 35532 27020 35588
rect 27076 35532 27086 35588
rect 30482 35532 30492 35588
rect 30548 35532 32060 35588
rect 32116 35532 32126 35588
rect 42354 35532 42364 35588
rect 42420 35532 42588 35588
rect 42644 35532 43372 35588
rect 43428 35532 45276 35588
rect 45332 35532 45342 35588
rect 54786 35532 54796 35588
rect 54852 35532 55468 35588
rect 55524 35532 55534 35588
rect 23650 35420 23660 35476
rect 23716 35420 26012 35476
rect 26068 35420 26684 35476
rect 26740 35420 26750 35476
rect 36194 35420 36204 35476
rect 36260 35420 37996 35476
rect 38052 35420 38892 35476
rect 38948 35420 38958 35476
rect 5058 35308 5068 35364
rect 5124 35308 5134 35364
rect 14914 35308 14924 35364
rect 14980 35308 15484 35364
rect 15540 35308 15550 35364
rect 47842 35308 47852 35364
rect 47908 35308 49980 35364
rect 50036 35308 53116 35364
rect 53172 35308 53182 35364
rect 54226 35308 54236 35364
rect 54292 35308 55132 35364
rect 55188 35308 56700 35364
rect 56756 35308 56766 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 5068 35252 5124 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 5068 35196 6076 35252
rect 6132 35196 6142 35252
rect 11330 35196 11340 35252
rect 11396 35196 11788 35252
rect 11844 35196 12572 35252
rect 12628 35196 13916 35252
rect 13972 35196 13982 35252
rect 15698 35196 15708 35252
rect 15764 35196 16380 35252
rect 16436 35196 16446 35252
rect 34402 35196 34412 35252
rect 34468 35196 34972 35252
rect 35028 35196 35038 35252
rect 4834 35084 4844 35140
rect 4900 35084 5964 35140
rect 6020 35084 6030 35140
rect 28354 35084 28364 35140
rect 28420 35084 29596 35140
rect 29652 35084 37660 35140
rect 37716 35084 37726 35140
rect 41234 35084 41244 35140
rect 41300 35084 41692 35140
rect 41748 35084 46844 35140
rect 46900 35084 46910 35140
rect 9650 34972 9660 35028
rect 9716 34972 10556 35028
rect 10612 34972 10622 35028
rect 36306 34972 36316 35028
rect 36372 34972 37772 35028
rect 37828 34972 37838 35028
rect 40450 34972 40460 35028
rect 40516 34972 42140 35028
rect 42196 34972 42206 35028
rect 52210 34972 52220 35028
rect 52276 34972 52892 35028
rect 52948 34972 52958 35028
rect 17378 34860 17388 34916
rect 17444 34860 19180 34916
rect 19236 34860 20860 34916
rect 20916 34860 20926 34916
rect 33170 34860 33180 34916
rect 33236 34860 34748 34916
rect 34804 34860 34814 34916
rect 43250 34860 43260 34916
rect 43316 34860 43932 34916
rect 43988 34860 43998 34916
rect 50194 34860 50204 34916
rect 50260 34860 50764 34916
rect 50820 34860 51548 34916
rect 51604 34860 51614 34916
rect 4610 34748 4620 34804
rect 4676 34748 5628 34804
rect 5684 34748 5694 34804
rect 41794 34748 41804 34804
rect 41860 34748 42364 34804
rect 42420 34748 42430 34804
rect 42578 34748 42588 34804
rect 42644 34748 46060 34804
rect 46116 34748 46126 34804
rect 2482 34636 2492 34692
rect 2548 34636 5740 34692
rect 5796 34636 5806 34692
rect 25778 34636 25788 34692
rect 25844 34636 26460 34692
rect 26516 34636 26526 34692
rect 32610 34636 32620 34692
rect 32676 34636 33292 34692
rect 33348 34636 33358 34692
rect 34738 34636 34748 34692
rect 34804 34636 35084 34692
rect 35140 34636 35150 34692
rect 42242 34636 42252 34692
rect 42308 34636 43148 34692
rect 43204 34636 43214 34692
rect 42130 34524 42140 34580
rect 42196 34524 42588 34580
rect 42644 34524 42654 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 27234 34412 27244 34468
rect 27300 34412 34412 34468
rect 34468 34412 34478 34468
rect 32722 34300 32732 34356
rect 32788 34300 33180 34356
rect 33236 34300 33246 34356
rect 34626 34300 34636 34356
rect 34692 34300 35084 34356
rect 35140 34300 35150 34356
rect 36082 34300 36092 34356
rect 36148 34300 36158 34356
rect 36092 34244 36148 34300
rect 20514 34188 20524 34244
rect 20580 34188 36148 34244
rect 8194 34076 8204 34132
rect 8260 34076 9660 34132
rect 9716 34076 9726 34132
rect 16370 34076 16380 34132
rect 16436 34076 19516 34132
rect 19572 34076 19582 34132
rect 20290 34076 20300 34132
rect 20356 34076 21868 34132
rect 21924 34076 21934 34132
rect 34850 34076 34860 34132
rect 34916 34076 35084 34132
rect 35140 34076 35150 34132
rect 35858 34076 35868 34132
rect 35924 34076 36764 34132
rect 36820 34076 49196 34132
rect 49252 34076 49262 34132
rect 16482 33964 16492 34020
rect 16548 33964 17388 34020
rect 17444 33964 17454 34020
rect 26674 33964 26684 34020
rect 26740 33964 27916 34020
rect 27972 33964 27982 34020
rect 52210 33964 52220 34020
rect 52276 33964 53340 34020
rect 53396 33964 54124 34020
rect 54180 33964 54190 34020
rect 16034 33852 16044 33908
rect 16100 33852 19516 33908
rect 19572 33852 19582 33908
rect 34290 33852 34300 33908
rect 34356 33852 34636 33908
rect 34692 33852 34702 33908
rect 36978 33852 36988 33908
rect 37044 33852 37660 33908
rect 37716 33852 39228 33908
rect 39284 33852 39294 33908
rect 47058 33740 47068 33796
rect 47124 33740 54572 33796
rect 54628 33740 54796 33796
rect 54852 33740 55244 33796
rect 55300 33740 55310 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 6402 33516 6412 33572
rect 6468 33516 6860 33572
rect 6916 33516 7532 33572
rect 7588 33516 7598 33572
rect 11330 33516 11340 33572
rect 11396 33516 12348 33572
rect 12404 33516 12414 33572
rect 27682 33516 27692 33572
rect 27748 33516 31164 33572
rect 31220 33516 31230 33572
rect 32162 33516 32172 33572
rect 32228 33516 33292 33572
rect 33348 33516 35532 33572
rect 35588 33516 35980 33572
rect 36036 33516 36046 33572
rect 37090 33516 37100 33572
rect 37156 33516 37884 33572
rect 37940 33516 38444 33572
rect 38500 33516 38510 33572
rect 52098 33516 52108 33572
rect 52164 33516 53004 33572
rect 53060 33516 53070 33572
rect 20850 33404 20860 33460
rect 20916 33404 25228 33460
rect 25284 33404 26908 33460
rect 36530 33404 36540 33460
rect 36596 33404 38108 33460
rect 38164 33404 38174 33460
rect 41346 33404 41356 33460
rect 41412 33404 41916 33460
rect 41972 33404 41982 33460
rect 54786 33404 54796 33460
rect 54852 33404 56028 33460
rect 56084 33404 56094 33460
rect 26852 33348 26908 33404
rect 1810 33292 1820 33348
rect 1876 33292 4956 33348
rect 5012 33292 6972 33348
rect 7028 33292 7038 33348
rect 26852 33292 29708 33348
rect 29764 33292 29774 33348
rect 36082 33292 36092 33348
rect 36148 33292 37212 33348
rect 37268 33292 38444 33348
rect 38500 33292 38510 33348
rect 42018 33292 42028 33348
rect 42084 33292 42700 33348
rect 42756 33292 42766 33348
rect 51874 33292 51884 33348
rect 51940 33292 58156 33348
rect 58212 33292 58222 33348
rect 20290 33180 20300 33236
rect 20356 33180 22428 33236
rect 22484 33180 22494 33236
rect 31602 33180 31612 33236
rect 31668 33180 31948 33236
rect 32004 33180 32014 33236
rect 42466 33180 42476 33236
rect 42532 33180 44716 33236
rect 44772 33180 44782 33236
rect 44930 33180 44940 33236
rect 44996 33180 46620 33236
rect 46676 33180 46686 33236
rect 50306 33180 50316 33236
rect 50372 33180 52780 33236
rect 52836 33180 52846 33236
rect 14690 33068 14700 33124
rect 14756 33068 16492 33124
rect 16548 33068 16558 33124
rect 33170 33068 33180 33124
rect 33236 33068 33852 33124
rect 33908 33068 33918 33124
rect 38098 33068 38108 33124
rect 38164 33068 41244 33124
rect 41300 33068 41310 33124
rect 52098 33068 52108 33124
rect 52164 33068 52556 33124
rect 52612 33068 53564 33124
rect 53620 33068 53630 33124
rect 34150 32956 34188 33012
rect 34244 32956 34254 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 22754 32844 22764 32900
rect 22820 32844 24108 32900
rect 24164 32844 24174 32900
rect 31154 32844 31164 32900
rect 31220 32844 31836 32900
rect 31892 32844 31902 32900
rect 34486 32844 34524 32900
rect 34580 32844 34590 32900
rect 59200 32788 60000 32816
rect 4610 32732 4620 32788
rect 4676 32732 5180 32788
rect 5236 32732 5964 32788
rect 6020 32732 6030 32788
rect 16370 32732 16380 32788
rect 16436 32732 17388 32788
rect 17444 32732 17454 32788
rect 22530 32732 22540 32788
rect 22596 32732 23548 32788
rect 23604 32732 23614 32788
rect 29362 32732 29372 32788
rect 29428 32732 29820 32788
rect 29876 32732 34188 32788
rect 34244 32732 38556 32788
rect 38612 32732 40012 32788
rect 40068 32732 40078 32788
rect 50754 32732 50764 32788
rect 50820 32732 51884 32788
rect 51940 32732 51950 32788
rect 52994 32732 53004 32788
rect 53060 32732 54236 32788
rect 54292 32732 54302 32788
rect 57362 32732 57372 32788
rect 57428 32732 58156 32788
rect 58212 32732 60000 32788
rect 59200 32704 60000 32732
rect 22306 32620 22316 32676
rect 22372 32620 24444 32676
rect 24500 32620 30940 32676
rect 30996 32620 31006 32676
rect 51986 32620 51996 32676
rect 52052 32620 53116 32676
rect 53172 32620 53182 32676
rect 4162 32508 4172 32564
rect 4228 32508 4956 32564
rect 5012 32508 6076 32564
rect 6132 32508 6142 32564
rect 22418 32508 22428 32564
rect 22484 32508 24108 32564
rect 24164 32508 26908 32564
rect 27570 32508 27580 32564
rect 27636 32508 29596 32564
rect 29652 32508 29662 32564
rect 47730 32508 47740 32564
rect 47796 32508 48636 32564
rect 48692 32508 49084 32564
rect 49140 32508 49150 32564
rect 49746 32508 49756 32564
rect 49812 32508 50540 32564
rect 50596 32508 50606 32564
rect 51650 32508 51660 32564
rect 51716 32508 52556 32564
rect 52612 32508 52622 32564
rect 52882 32508 52892 32564
rect 52948 32508 54460 32564
rect 54516 32508 54526 32564
rect 2482 32396 2492 32452
rect 2548 32396 5068 32452
rect 5124 32396 5134 32452
rect 21746 32396 21756 32452
rect 21812 32396 22092 32452
rect 22148 32396 22158 32452
rect 24210 32396 24220 32452
rect 24276 32396 26348 32452
rect 26404 32396 26414 32452
rect 26852 32340 26908 32508
rect 29250 32396 29260 32452
rect 29316 32396 31052 32452
rect 31108 32396 31118 32452
rect 41458 32396 41468 32452
rect 41524 32396 42588 32452
rect 42644 32396 42654 32452
rect 44706 32396 44716 32452
rect 44772 32396 48748 32452
rect 48804 32396 49644 32452
rect 49700 32396 49710 32452
rect 52294 32396 52332 32452
rect 52388 32396 52398 32452
rect 26852 32284 30828 32340
rect 30884 32284 31276 32340
rect 31332 32284 31342 32340
rect 49532 32284 52892 32340
rect 52948 32284 52958 32340
rect 53330 32284 53340 32340
rect 53396 32284 53900 32340
rect 53956 32284 53966 32340
rect 18946 32172 18956 32228
rect 19012 32172 21308 32228
rect 21364 32172 21868 32228
rect 21924 32172 23324 32228
rect 23380 32172 23390 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 28242 32060 28252 32116
rect 28308 32060 28318 32116
rect 40450 32060 40460 32116
rect 40516 32060 40908 32116
rect 40964 32060 40974 32116
rect 46498 32060 46508 32116
rect 46564 32060 47740 32116
rect 47796 32060 47806 32116
rect 24098 31948 24108 32004
rect 24164 31948 25340 32004
rect 25396 31948 25406 32004
rect 28252 31892 28308 32060
rect 35186 31948 35196 32004
rect 35252 31948 37548 32004
rect 37604 31948 37614 32004
rect 47282 31948 47292 32004
rect 47348 31948 47358 32004
rect 47292 31892 47348 31948
rect 49532 31892 49588 32284
rect 16482 31836 16492 31892
rect 16548 31836 16828 31892
rect 16884 31836 16894 31892
rect 28252 31836 29148 31892
rect 29204 31836 29214 31892
rect 34402 31836 34412 31892
rect 34468 31836 35084 31892
rect 35140 31836 35150 31892
rect 37314 31836 37324 31892
rect 37380 31836 41804 31892
rect 41860 31836 41870 31892
rect 45826 31836 45836 31892
rect 45892 31836 49532 31892
rect 49588 31836 49598 31892
rect 52658 31836 52668 31892
rect 52724 31836 53508 31892
rect 53666 31836 53676 31892
rect 53732 31836 54460 31892
rect 54516 31836 54526 31892
rect 53452 31780 53508 31836
rect 7298 31724 7308 31780
rect 7364 31724 8204 31780
rect 8260 31724 8270 31780
rect 22418 31724 22428 31780
rect 22484 31724 22988 31780
rect 23044 31724 26796 31780
rect 26852 31724 26862 31780
rect 29474 31724 29484 31780
rect 29540 31724 31500 31780
rect 31556 31724 31566 31780
rect 34626 31724 34636 31780
rect 34692 31724 35420 31780
rect 35476 31724 35486 31780
rect 41122 31724 41132 31780
rect 41188 31724 42364 31780
rect 42420 31724 42430 31780
rect 44370 31724 44380 31780
rect 44436 31724 48412 31780
rect 48468 31724 48478 31780
rect 50372 31724 53228 31780
rect 53284 31724 53294 31780
rect 53452 31724 58156 31780
rect 58212 31724 58222 31780
rect 7858 31612 7868 31668
rect 7924 31612 8652 31668
rect 8708 31612 8718 31668
rect 11218 31612 11228 31668
rect 11284 31612 12124 31668
rect 12180 31612 12190 31668
rect 20402 31612 20412 31668
rect 20468 31612 22316 31668
rect 22372 31612 22382 31668
rect 31826 31612 31836 31668
rect 31892 31612 41580 31668
rect 41636 31612 42700 31668
rect 42756 31612 42766 31668
rect 50372 31556 50428 31724
rect 53666 31612 53676 31668
rect 53732 31612 54236 31668
rect 54292 31612 54302 31668
rect 54786 31612 54796 31668
rect 54852 31612 56028 31668
rect 56084 31612 56094 31668
rect 4050 31500 4060 31556
rect 4116 31500 4732 31556
rect 4788 31500 5628 31556
rect 5684 31500 5694 31556
rect 28018 31500 28028 31556
rect 28084 31500 28476 31556
rect 28532 31500 28542 31556
rect 47954 31500 47964 31556
rect 48020 31500 49196 31556
rect 49252 31500 50428 31556
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 34850 31276 34860 31332
rect 34916 31276 35588 31332
rect 35532 31220 35588 31276
rect 5954 31164 5964 31220
rect 6020 31164 7532 31220
rect 7588 31164 8204 31220
rect 8260 31164 8270 31220
rect 17154 31164 17164 31220
rect 17220 31164 17836 31220
rect 17892 31164 17902 31220
rect 31714 31164 31724 31220
rect 31780 31164 33180 31220
rect 33236 31164 33246 31220
rect 35522 31164 35532 31220
rect 35588 31164 36652 31220
rect 36708 31164 36718 31220
rect 40338 31164 40348 31220
rect 40404 31164 40684 31220
rect 40740 31164 40750 31220
rect 41346 31164 41356 31220
rect 41412 31164 42588 31220
rect 42644 31164 42654 31220
rect 47506 31164 47516 31220
rect 47572 31164 48188 31220
rect 48244 31164 48748 31220
rect 48804 31164 48814 31220
rect 8204 31108 8260 31164
rect 4498 31052 4508 31108
rect 4564 31052 6188 31108
rect 6244 31052 6254 31108
rect 8204 31052 9548 31108
rect 9604 31052 9614 31108
rect 27458 31052 27468 31108
rect 27524 31052 27916 31108
rect 27972 31052 27982 31108
rect 31490 31052 31500 31108
rect 31556 31052 33852 31108
rect 33908 31052 34860 31108
rect 34916 31052 35980 31108
rect 36036 31052 36046 31108
rect 46946 31052 46956 31108
rect 47012 31052 47404 31108
rect 47460 31052 47470 31108
rect 25106 30940 25116 30996
rect 25172 30940 25452 30996
rect 25508 30940 25788 30996
rect 25844 30940 25854 30996
rect 31042 30940 31052 30996
rect 31108 30940 31948 30996
rect 32004 30940 33740 30996
rect 33796 30940 34524 30996
rect 34580 30940 34590 30996
rect 36642 30940 36652 30996
rect 36708 30940 37324 30996
rect 37380 30940 37390 30996
rect 40338 30940 40348 30996
rect 40404 30940 41132 30996
rect 41188 30940 48412 30996
rect 48468 30940 48972 30996
rect 49028 30940 49038 30996
rect 2482 30828 2492 30884
rect 2548 30828 4956 30884
rect 5012 30828 5022 30884
rect 16482 30828 16492 30884
rect 16548 30828 17500 30884
rect 17556 30828 17566 30884
rect 27458 30828 27468 30884
rect 27524 30828 28700 30884
rect 28756 30828 28766 30884
rect 30146 30828 30156 30884
rect 30212 30828 31836 30884
rect 31892 30828 31902 30884
rect 40898 30828 40908 30884
rect 40964 30828 42476 30884
rect 42532 30828 42542 30884
rect 45602 30828 45612 30884
rect 45668 30828 46060 30884
rect 46116 30828 54684 30884
rect 54740 30828 54750 30884
rect 27346 30716 27356 30772
rect 27412 30716 28028 30772
rect 28084 30716 28094 30772
rect 48178 30716 48188 30772
rect 48244 30716 49308 30772
rect 49364 30716 49374 30772
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 8418 30268 8428 30324
rect 8484 30268 10556 30324
rect 10612 30268 11564 30324
rect 11620 30268 11630 30324
rect 27906 30268 27916 30324
rect 27972 30268 33180 30324
rect 33236 30268 33516 30324
rect 33572 30268 33582 30324
rect 39442 30268 39452 30324
rect 39508 30268 41468 30324
rect 41524 30268 41534 30324
rect 45602 30268 45612 30324
rect 45668 30268 46956 30324
rect 47012 30268 47022 30324
rect 52210 30268 52220 30324
rect 52276 30268 53676 30324
rect 53732 30268 53742 30324
rect 8530 30156 8540 30212
rect 8596 30156 9548 30212
rect 9604 30156 9614 30212
rect 15922 30156 15932 30212
rect 15988 30156 16380 30212
rect 16436 30156 16716 30212
rect 16772 30156 17612 30212
rect 17668 30156 17678 30212
rect 26226 30156 26236 30212
rect 26292 30156 26908 30212
rect 29922 30156 29932 30212
rect 29988 30156 30604 30212
rect 30660 30156 30670 30212
rect 34850 30156 34860 30212
rect 34916 30156 36316 30212
rect 36372 30156 36382 30212
rect 38210 30156 38220 30212
rect 38276 30156 39340 30212
rect 39396 30156 39406 30212
rect 48514 30156 48524 30212
rect 48580 30156 49532 30212
rect 49588 30156 49598 30212
rect 54002 30156 54012 30212
rect 54068 30156 54348 30212
rect 54404 30156 54414 30212
rect 26852 30100 26908 30156
rect 8978 30044 8988 30100
rect 9044 30044 10668 30100
rect 10724 30044 11676 30100
rect 11732 30044 11742 30100
rect 16930 30044 16940 30100
rect 16996 30044 17948 30100
rect 18004 30044 19292 30100
rect 19348 30044 19358 30100
rect 24658 30044 24668 30100
rect 24724 30044 26460 30100
rect 26516 30044 26526 30100
rect 26852 30044 37436 30100
rect 37492 30044 37502 30100
rect 4946 29932 4956 29988
rect 5012 29932 5740 29988
rect 5796 29932 5806 29988
rect 7410 29932 7420 29988
rect 7476 29932 29932 29988
rect 29988 29932 29998 29988
rect 39890 29932 39900 29988
rect 39956 29932 40796 29988
rect 40852 29932 40862 29988
rect 53778 29932 53788 29988
rect 53844 29932 54908 29988
rect 54964 29932 54974 29988
rect 6514 29820 6524 29876
rect 6580 29820 7084 29876
rect 7140 29820 7756 29876
rect 7812 29820 18508 29876
rect 18564 29820 19068 29876
rect 19124 29820 19134 29876
rect 20402 29820 20412 29876
rect 20468 29820 34188 29876
rect 34244 29820 34254 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 5842 29596 5852 29652
rect 5908 29596 8540 29652
rect 8596 29596 8606 29652
rect 13794 29596 13804 29652
rect 13860 29596 16268 29652
rect 16324 29596 16334 29652
rect 19394 29596 19404 29652
rect 19460 29596 19852 29652
rect 19908 29596 20524 29652
rect 20580 29596 36988 29652
rect 37044 29596 37436 29652
rect 37492 29596 37996 29652
rect 38052 29596 38062 29652
rect 49634 29596 49644 29652
rect 49700 29596 51548 29652
rect 51604 29596 51614 29652
rect 49522 29484 49532 29540
rect 49588 29484 50764 29540
rect 50820 29484 50830 29540
rect 54226 29484 54236 29540
rect 54292 29484 55020 29540
rect 55076 29484 55086 29540
rect 8614 29372 8652 29428
rect 8708 29372 8718 29428
rect 46386 29372 46396 29428
rect 46452 29372 47180 29428
rect 47236 29372 47246 29428
rect 48514 29372 48524 29428
rect 48580 29372 49308 29428
rect 49364 29372 49374 29428
rect 50642 29372 50652 29428
rect 50708 29372 52780 29428
rect 52836 29372 52846 29428
rect 24434 29260 24444 29316
rect 24500 29260 25228 29316
rect 25284 29260 25294 29316
rect 34514 29260 34524 29316
rect 34580 29260 46620 29316
rect 46676 29260 47516 29316
rect 47572 29260 47582 29316
rect 27346 29148 27356 29204
rect 27412 29148 28140 29204
rect 28196 29148 37828 29204
rect 44594 29148 44604 29204
rect 44660 29148 46060 29204
rect 46116 29148 46126 29204
rect 37772 29092 37828 29148
rect 37762 29036 37772 29092
rect 37828 29036 46172 29092
rect 46228 29036 46238 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 15138 28924 15148 28980
rect 15204 28924 22316 28980
rect 22372 28924 23548 28980
rect 23604 28924 23614 28980
rect 22082 28812 22092 28868
rect 22148 28812 26572 28868
rect 26628 28812 26638 28868
rect 26852 28812 27244 28868
rect 27300 28812 27310 28868
rect 44034 28812 44044 28868
rect 44100 28812 44996 28868
rect 26852 28756 26908 28812
rect 44940 28756 44996 28812
rect 7858 28700 7868 28756
rect 7924 28700 9772 28756
rect 9828 28700 9838 28756
rect 12114 28700 12124 28756
rect 12180 28700 18396 28756
rect 18452 28700 18462 28756
rect 26338 28700 26348 28756
rect 26404 28700 26908 28756
rect 31042 28700 31052 28756
rect 31108 28700 32508 28756
rect 32564 28700 32574 28756
rect 42018 28700 42028 28756
rect 42084 28700 42812 28756
rect 42868 28700 43484 28756
rect 43540 28700 44492 28756
rect 44548 28700 44558 28756
rect 44930 28700 44940 28756
rect 44996 28700 46396 28756
rect 46452 28700 46462 28756
rect 51324 28700 51996 28756
rect 52052 28700 53900 28756
rect 53956 28700 53966 28756
rect 54898 28700 54908 28756
rect 54964 28700 58156 28756
rect 58212 28700 58222 28756
rect 51324 28644 51380 28700
rect 6850 28588 6860 28644
rect 6916 28588 7532 28644
rect 7588 28588 7598 28644
rect 8978 28588 8988 28644
rect 9044 28588 9660 28644
rect 9716 28588 10668 28644
rect 10724 28588 10734 28644
rect 10882 28588 10892 28644
rect 10948 28588 12012 28644
rect 12068 28588 12078 28644
rect 27346 28588 27356 28644
rect 27412 28588 29036 28644
rect 29092 28588 29102 28644
rect 44258 28588 44268 28644
rect 44324 28588 47180 28644
rect 47236 28588 47246 28644
rect 51314 28588 51324 28644
rect 51380 28588 51390 28644
rect 51538 28588 51548 28644
rect 51604 28588 52668 28644
rect 52724 28588 52734 28644
rect 7970 28476 7980 28532
rect 8036 28476 8652 28532
rect 8708 28476 8718 28532
rect 16370 28476 16380 28532
rect 16436 28476 16716 28532
rect 16772 28476 18732 28532
rect 18788 28476 18798 28532
rect 23874 28476 23884 28532
rect 23940 28476 33852 28532
rect 33908 28476 33918 28532
rect 34290 28476 34300 28532
rect 34356 28476 35084 28532
rect 35140 28476 36652 28532
rect 36708 28476 36718 28532
rect 11330 28364 11340 28420
rect 11396 28364 13020 28420
rect 13076 28364 13086 28420
rect 25778 28364 25788 28420
rect 25844 28364 26460 28420
rect 26516 28364 26908 28420
rect 28690 28364 28700 28420
rect 28756 28364 29372 28420
rect 29428 28364 34412 28420
rect 34468 28364 37100 28420
rect 37156 28364 37166 28420
rect 46162 28364 46172 28420
rect 46228 28364 48412 28420
rect 48468 28364 48478 28420
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 26852 28196 26908 28364
rect 45042 28252 45052 28308
rect 45108 28252 45118 28308
rect 47618 28252 47628 28308
rect 47684 28252 48636 28308
rect 48692 28252 48702 28308
rect 8082 28140 8092 28196
rect 8148 28140 8764 28196
rect 8820 28140 8830 28196
rect 26852 28140 27356 28196
rect 27412 28140 27804 28196
rect 27860 28140 31332 28196
rect 31276 28084 31332 28140
rect 20962 28028 20972 28084
rect 21028 28028 23100 28084
rect 23156 28028 30268 28084
rect 30324 28028 30334 28084
rect 31266 28028 31276 28084
rect 31332 28028 32172 28084
rect 32228 28028 43708 28084
rect 43764 28028 43774 28084
rect 31714 27916 31724 27972
rect 31780 27916 33740 27972
rect 33796 27916 33806 27972
rect 36418 27916 36428 27972
rect 36484 27916 37324 27972
rect 37380 27916 38556 27972
rect 38612 27916 38622 27972
rect 45052 27860 45108 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 3826 27804 3836 27860
rect 3892 27804 4844 27860
rect 4900 27804 4910 27860
rect 8642 27804 8652 27860
rect 8708 27804 10892 27860
rect 10948 27804 11228 27860
rect 11284 27804 11900 27860
rect 11956 27804 11966 27860
rect 26002 27804 26012 27860
rect 26068 27804 26572 27860
rect 26628 27804 27132 27860
rect 27188 27804 28364 27860
rect 28420 27804 28430 27860
rect 31154 27804 31164 27860
rect 31220 27804 31836 27860
rect 31892 27804 33292 27860
rect 33348 27804 33358 27860
rect 33506 27804 33516 27860
rect 33572 27804 36540 27860
rect 36596 27804 36606 27860
rect 43698 27804 43708 27860
rect 43764 27804 44380 27860
rect 44436 27804 47180 27860
rect 47236 27804 47740 27860
rect 47796 27804 47806 27860
rect 2482 27692 2492 27748
rect 2548 27692 3948 27748
rect 4004 27692 4014 27748
rect 14690 27692 14700 27748
rect 14756 27692 16268 27748
rect 16324 27692 16334 27748
rect 17714 27692 17724 27748
rect 17780 27692 19292 27748
rect 19348 27692 19358 27748
rect 25554 27692 25564 27748
rect 25620 27692 26124 27748
rect 26180 27692 26190 27748
rect 27346 27692 27356 27748
rect 27412 27692 28140 27748
rect 28196 27692 28206 27748
rect 30034 27692 30044 27748
rect 30100 27692 31388 27748
rect 31444 27692 31454 27748
rect 41682 27692 41692 27748
rect 41748 27692 45612 27748
rect 45668 27692 45678 27748
rect 47618 27692 47628 27748
rect 47684 27692 51212 27748
rect 51268 27692 51278 27748
rect 54086 27692 54124 27748
rect 54180 27692 54190 27748
rect 4498 27580 4508 27636
rect 4564 27580 4956 27636
rect 5012 27580 5022 27636
rect 8530 27580 8540 27636
rect 8596 27580 9660 27636
rect 9716 27580 10220 27636
rect 10276 27580 10668 27636
rect 10724 27580 21308 27636
rect 21364 27580 21374 27636
rect 24434 27580 24444 27636
rect 24500 27580 25340 27636
rect 25396 27580 25406 27636
rect 30818 27580 30828 27636
rect 30884 27580 33740 27636
rect 33796 27580 33806 27636
rect 33964 27580 34636 27636
rect 34692 27580 37548 27636
rect 37604 27580 37614 27636
rect 39106 27580 39116 27636
rect 39172 27580 42588 27636
rect 42644 27580 42654 27636
rect 33964 27524 34020 27580
rect 28690 27468 28700 27524
rect 28756 27468 34020 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 21634 27132 21644 27188
rect 21700 27132 25564 27188
rect 25620 27132 25630 27188
rect 33058 27132 33068 27188
rect 33124 27132 34748 27188
rect 34804 27132 34814 27188
rect 4946 27020 4956 27076
rect 5012 27020 5628 27076
rect 5684 27020 6524 27076
rect 6580 27020 7308 27076
rect 7364 27020 7374 27076
rect 9090 27020 9100 27076
rect 9156 27020 10556 27076
rect 10612 27020 11116 27076
rect 11172 27020 11182 27076
rect 23986 27020 23996 27076
rect 24052 27020 25900 27076
rect 25956 27020 25966 27076
rect 26114 27020 26124 27076
rect 26180 27020 26796 27076
rect 26852 27020 26862 27076
rect 29810 27020 29820 27076
rect 29876 27020 31948 27076
rect 32004 27020 32014 27076
rect 36530 27020 36540 27076
rect 36596 27020 37100 27076
rect 37156 27020 37166 27076
rect 52098 27020 52108 27076
rect 52164 27020 52892 27076
rect 52948 27020 52958 27076
rect 59200 26964 60000 26992
rect 4386 26908 4396 26964
rect 4452 26908 7196 26964
rect 7252 26908 7980 26964
rect 8036 26908 8046 26964
rect 26002 26908 26012 26964
rect 26068 26908 27020 26964
rect 27076 26908 27580 26964
rect 27636 26908 29652 26964
rect 34850 26908 34860 26964
rect 34916 26908 34926 26964
rect 48626 26908 48636 26964
rect 48692 26908 49868 26964
rect 49924 26908 49934 26964
rect 50082 26908 50092 26964
rect 50148 26908 51324 26964
rect 51380 26908 51390 26964
rect 58156 26908 60000 26964
rect 5852 26852 5908 26908
rect 29596 26852 29652 26908
rect 5618 26796 5628 26852
rect 5684 26796 5908 26852
rect 22194 26796 22204 26852
rect 22260 26796 22764 26852
rect 22820 26796 24220 26852
rect 24276 26796 24286 26852
rect 29596 26796 31612 26852
rect 31668 26796 32172 26852
rect 32228 26796 32238 26852
rect 34860 26740 34916 26908
rect 58156 26852 58212 26908
rect 59200 26880 60000 26908
rect 39218 26796 39228 26852
rect 39284 26796 41020 26852
rect 41076 26796 41086 26852
rect 50642 26796 50652 26852
rect 50708 26796 50988 26852
rect 51044 26796 51054 26852
rect 54226 26796 54236 26852
rect 54292 26796 54908 26852
rect 54964 26796 55468 26852
rect 55524 26796 55534 26852
rect 57586 26796 57596 26852
rect 57652 26796 58156 26852
rect 58212 26796 58222 26852
rect 34860 26684 35980 26740
rect 36036 26684 36046 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 3266 26460 3276 26516
rect 3332 26460 4732 26516
rect 4788 26460 5740 26516
rect 5796 26460 5806 26516
rect 26338 26460 26348 26516
rect 26404 26460 27244 26516
rect 27300 26460 27310 26516
rect 37090 26460 37100 26516
rect 37156 26460 38108 26516
rect 38164 26460 39004 26516
rect 39060 26460 39070 26516
rect 47012 26460 50316 26516
rect 50372 26460 52108 26516
rect 52164 26460 52174 26516
rect 3154 26348 3164 26404
rect 3220 26348 5180 26404
rect 5236 26348 5246 26404
rect 20066 26348 20076 26404
rect 20132 26348 25788 26404
rect 25844 26348 25854 26404
rect 28242 26348 28252 26404
rect 28308 26348 37884 26404
rect 37940 26348 37950 26404
rect 47012 26292 47068 26460
rect 50642 26348 50652 26404
rect 50708 26348 51100 26404
rect 51156 26348 51166 26404
rect 54338 26348 54348 26404
rect 54404 26348 55020 26404
rect 55076 26348 55086 26404
rect 4946 26236 4956 26292
rect 5012 26236 8876 26292
rect 8932 26236 9772 26292
rect 9828 26236 9838 26292
rect 24322 26236 24332 26292
rect 24388 26236 25452 26292
rect 25508 26236 25518 26292
rect 28130 26236 28140 26292
rect 28196 26236 29596 26292
rect 29652 26236 30716 26292
rect 30772 26236 30782 26292
rect 46610 26236 46620 26292
rect 46676 26236 47068 26292
rect 53330 26236 53340 26292
rect 53396 26236 54124 26292
rect 54180 26236 55692 26292
rect 55748 26236 55758 26292
rect 26450 26124 26460 26180
rect 26516 26124 27356 26180
rect 27412 26124 27422 26180
rect 36642 26124 36652 26180
rect 36708 26124 37436 26180
rect 37492 26124 38556 26180
rect 38612 26124 38622 26180
rect 52070 26124 52108 26180
rect 52164 26124 52174 26180
rect 28354 26012 28364 26068
rect 28420 26012 36428 26068
rect 36484 26012 37324 26068
rect 37380 26012 37390 26068
rect 52322 26012 52332 26068
rect 52388 26012 52892 26068
rect 52948 26012 52958 26068
rect 8978 25900 8988 25956
rect 9044 25900 10892 25956
rect 10948 25900 10958 25956
rect 49186 25900 49196 25956
rect 49252 25900 49868 25956
rect 49924 25900 49934 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 28802 25676 28812 25732
rect 28868 25676 28878 25732
rect 50082 25676 50092 25732
rect 50148 25676 50540 25732
rect 50596 25676 50606 25732
rect 54898 25676 54908 25732
rect 54964 25676 55244 25732
rect 55300 25676 55310 25732
rect 5170 25564 5180 25620
rect 5236 25564 6580 25620
rect 8418 25564 8428 25620
rect 8484 25564 8764 25620
rect 8820 25564 8830 25620
rect 6524 25508 6580 25564
rect 28812 25508 28868 25676
rect 30706 25564 30716 25620
rect 30772 25564 31388 25620
rect 31444 25564 31454 25620
rect 37874 25564 37884 25620
rect 37940 25564 48300 25620
rect 48356 25564 48366 25620
rect 55682 25564 55692 25620
rect 55748 25564 58156 25620
rect 58212 25564 58222 25620
rect 4274 25452 4284 25508
rect 4340 25452 5628 25508
rect 5684 25452 5694 25508
rect 6514 25452 6524 25508
rect 6580 25452 6590 25508
rect 28812 25452 38668 25508
rect 50754 25452 50764 25508
rect 50820 25452 50988 25508
rect 51044 25452 51054 25508
rect 38612 25396 38668 25452
rect 6626 25340 6636 25396
rect 6692 25340 7420 25396
rect 7476 25340 7868 25396
rect 7924 25340 8316 25396
rect 8372 25340 8382 25396
rect 23314 25340 23324 25396
rect 23380 25340 27916 25396
rect 27972 25340 30268 25396
rect 30324 25340 30334 25396
rect 38612 25340 42924 25396
rect 42980 25340 43372 25396
rect 43428 25340 43438 25396
rect 51762 25340 51772 25396
rect 51828 25340 52668 25396
rect 52724 25340 52734 25396
rect 2482 25228 2492 25284
rect 2548 25228 3836 25284
rect 3892 25228 3902 25284
rect 18050 25228 18060 25284
rect 18116 25228 19180 25284
rect 19236 25228 20244 25284
rect 28130 25228 28140 25284
rect 28196 25228 28588 25284
rect 28644 25228 28654 25284
rect 38546 25228 38556 25284
rect 38612 25228 39564 25284
rect 39620 25228 39630 25284
rect 40338 25228 40348 25284
rect 40404 25228 41468 25284
rect 41524 25228 51548 25284
rect 51604 25228 52220 25284
rect 52276 25228 52286 25284
rect 54786 25228 54796 25284
rect 54852 25228 56028 25284
rect 56084 25228 56094 25284
rect 5058 25116 5068 25172
rect 5124 25116 7980 25172
rect 8036 25116 8046 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 20188 25060 20244 25228
rect 24210 25116 24220 25172
rect 24276 25116 30156 25172
rect 30212 25116 30222 25172
rect 49746 25116 49756 25172
rect 49812 25116 49822 25172
rect 49756 25060 49812 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 20188 25004 22204 25060
rect 22260 25004 22270 25060
rect 38098 25004 38108 25060
rect 38164 25004 39116 25060
rect 39172 25004 40124 25060
rect 40180 25004 40908 25060
rect 40964 25004 40974 25060
rect 44156 25004 49812 25060
rect 23202 24892 23212 24948
rect 23268 24892 23548 24948
rect 23604 24892 23614 24948
rect 38210 24892 38220 24948
rect 38276 24892 39676 24948
rect 39732 24892 40796 24948
rect 40852 24892 40862 24948
rect 44156 24836 44212 25004
rect 49074 24892 49084 24948
rect 49140 24892 51212 24948
rect 51268 24892 51278 24948
rect 35970 24780 35980 24836
rect 36036 24780 37996 24836
rect 38052 24780 38062 24836
rect 38322 24780 38332 24836
rect 38388 24780 44212 24836
rect 49298 24780 49308 24836
rect 49364 24780 49374 24836
rect 49308 24724 49364 24780
rect 1810 24668 1820 24724
rect 1876 24668 5068 24724
rect 5124 24668 5134 24724
rect 10098 24668 10108 24724
rect 10164 24668 10780 24724
rect 10836 24668 13916 24724
rect 13972 24668 15036 24724
rect 15092 24668 15102 24724
rect 37762 24668 37772 24724
rect 37828 24668 38668 24724
rect 38724 24668 39340 24724
rect 39396 24668 39900 24724
rect 39956 24668 39966 24724
rect 49308 24668 51324 24724
rect 51380 24668 51390 24724
rect 52770 24668 52780 24724
rect 52836 24668 53004 24724
rect 53060 24668 54572 24724
rect 54628 24668 56924 24724
rect 56980 24668 56990 24724
rect 11442 24556 11452 24612
rect 11508 24556 12348 24612
rect 12404 24556 12414 24612
rect 14690 24556 14700 24612
rect 14756 24556 15932 24612
rect 15988 24556 15998 24612
rect 17826 24556 17836 24612
rect 17892 24556 18620 24612
rect 18676 24556 19292 24612
rect 19348 24556 19358 24612
rect 36194 24556 36204 24612
rect 36260 24556 38220 24612
rect 38276 24556 38286 24612
rect 44930 24556 44940 24612
rect 44996 24556 54460 24612
rect 54516 24556 55580 24612
rect 55636 24556 56084 24612
rect 56028 24500 56084 24556
rect 22866 24444 22876 24500
rect 22932 24444 24108 24500
rect 24164 24444 24174 24500
rect 41458 24444 41468 24500
rect 41524 24444 43932 24500
rect 43988 24444 48748 24500
rect 48804 24444 48814 24500
rect 55122 24444 55132 24500
rect 55188 24444 55804 24500
rect 55860 24444 55870 24500
rect 56018 24444 56028 24500
rect 56084 24444 56094 24500
rect 54786 24332 54796 24388
rect 54852 24332 56588 24388
rect 56644 24332 56654 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 23090 24220 23100 24276
rect 23156 24220 33180 24276
rect 33236 24220 33246 24276
rect 33180 24164 33236 24220
rect 8614 24108 8652 24164
rect 8708 24108 8718 24164
rect 19618 24108 19628 24164
rect 19684 24108 23996 24164
rect 24052 24108 24062 24164
rect 33180 24108 35532 24164
rect 35588 24108 35598 24164
rect 51314 24108 51324 24164
rect 51380 24108 53788 24164
rect 53844 24108 53854 24164
rect 20738 23996 20748 24052
rect 20804 23996 22316 24052
rect 22372 23996 23660 24052
rect 23716 23996 23726 24052
rect 56914 23996 56924 24052
rect 56980 23996 58156 24052
rect 58212 23996 58222 24052
rect 14578 23884 14588 23940
rect 14644 23884 15036 23940
rect 15092 23884 21980 23940
rect 22036 23884 22046 23940
rect 36082 23884 36092 23940
rect 36148 23884 37436 23940
rect 37492 23884 37502 23940
rect 38098 23884 38108 23940
rect 38164 23884 45276 23940
rect 45332 23884 45948 23940
rect 46004 23884 46396 23940
rect 46452 23884 46462 23940
rect 49074 23884 49084 23940
rect 49140 23884 49980 23940
rect 50036 23884 50046 23940
rect 12674 23772 12684 23828
rect 12740 23772 14140 23828
rect 14196 23772 14206 23828
rect 22194 23772 22204 23828
rect 22260 23772 23772 23828
rect 23828 23772 23838 23828
rect 31826 23772 31836 23828
rect 31892 23772 32508 23828
rect 32564 23772 32574 23828
rect 35298 23772 35308 23828
rect 35364 23772 36876 23828
rect 36932 23772 36942 23828
rect 41122 23772 41132 23828
rect 41188 23772 41692 23828
rect 41748 23772 41758 23828
rect 45714 23772 45724 23828
rect 45780 23772 53004 23828
rect 53060 23772 53070 23828
rect 9650 23660 9660 23716
rect 9716 23660 9884 23716
rect 9940 23660 10220 23716
rect 10276 23660 10286 23716
rect 22082 23660 22092 23716
rect 22148 23660 24108 23716
rect 24164 23660 24174 23716
rect 31938 23660 31948 23716
rect 32004 23660 33180 23716
rect 33236 23660 33246 23716
rect 36418 23660 36428 23716
rect 36484 23660 37212 23716
rect 37268 23660 37278 23716
rect 38612 23604 38668 23716
rect 38724 23660 38734 23716
rect 21970 23548 21980 23604
rect 22036 23548 23212 23604
rect 23268 23548 23278 23604
rect 38444 23548 38668 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 38444 23492 38500 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 29698 23436 29708 23492
rect 29764 23436 31500 23492
rect 31556 23436 31566 23492
rect 38434 23436 38444 23492
rect 38500 23436 38510 23492
rect 32050 23324 32060 23380
rect 32116 23324 33068 23380
rect 33124 23324 35308 23380
rect 35364 23324 35980 23380
rect 36036 23324 37212 23380
rect 37268 23324 37278 23380
rect 16706 23100 16716 23156
rect 16772 23100 17164 23156
rect 17220 23100 17948 23156
rect 18004 23100 18014 23156
rect 19506 23100 19516 23156
rect 19572 23100 19582 23156
rect 19842 23100 19852 23156
rect 19908 23100 21532 23156
rect 21588 23100 21598 23156
rect 22754 23100 22764 23156
rect 22820 23100 23884 23156
rect 23940 23100 24556 23156
rect 24612 23100 25340 23156
rect 25396 23100 25406 23156
rect 28802 23100 28812 23156
rect 28868 23100 29372 23156
rect 29428 23100 33740 23156
rect 33796 23100 36876 23156
rect 36932 23100 36942 23156
rect 48738 23100 48748 23156
rect 48804 23100 49196 23156
rect 49252 23100 49262 23156
rect 49410 23100 49420 23156
rect 49476 23100 51772 23156
rect 51828 23100 51838 23156
rect 53890 23100 53900 23156
rect 53956 23100 55244 23156
rect 55300 23100 55310 23156
rect 19516 23044 19572 23100
rect 19516 22988 20188 23044
rect 26786 22988 26796 23044
rect 26852 22988 27804 23044
rect 27860 22988 27870 23044
rect 29138 22988 29148 23044
rect 29204 22988 29708 23044
rect 29764 22988 29774 23044
rect 31266 22988 31276 23044
rect 31332 22988 33180 23044
rect 33236 22988 33246 23044
rect 46050 22988 46060 23044
rect 46116 22988 48076 23044
rect 48132 22988 48142 23044
rect 20132 22932 20188 22988
rect 4610 22876 4620 22932
rect 4676 22876 5628 22932
rect 5684 22876 5694 22932
rect 12338 22876 12348 22932
rect 12404 22876 13468 22932
rect 13524 22876 13534 22932
rect 13794 22876 13804 22932
rect 13860 22876 14140 22932
rect 14196 22876 19628 22932
rect 19684 22876 19694 22932
rect 20132 22876 20300 22932
rect 20356 22876 20366 22932
rect 31602 22764 31612 22820
rect 31668 22764 32508 22820
rect 32564 22764 33180 22820
rect 33236 22764 33246 22820
rect 40114 22764 40124 22820
rect 40180 22764 48860 22820
rect 48916 22764 49756 22820
rect 49812 22764 49822 22820
rect 52882 22764 52892 22820
rect 52948 22764 54684 22820
rect 54740 22764 55244 22820
rect 55300 22764 55310 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 32274 22652 32284 22708
rect 32340 22652 33068 22708
rect 33124 22652 33134 22708
rect 47954 22652 47964 22708
rect 48020 22652 48972 22708
rect 49028 22652 49532 22708
rect 49588 22652 49980 22708
rect 50036 22652 50046 22708
rect 2482 22540 2492 22596
rect 2548 22540 4732 22596
rect 4788 22540 4798 22596
rect 17602 22540 17612 22596
rect 17668 22540 17948 22596
rect 18004 22540 18014 22596
rect 48290 22540 48300 22596
rect 48356 22540 52780 22596
rect 52836 22540 52846 22596
rect 3378 22428 3388 22484
rect 3444 22428 3948 22484
rect 4004 22428 4956 22484
rect 5012 22428 22428 22484
rect 22484 22428 22494 22484
rect 24658 22428 24668 22484
rect 24724 22428 25676 22484
rect 25732 22428 27020 22484
rect 27076 22428 27356 22484
rect 27412 22428 27422 22484
rect 39330 22428 39340 22484
rect 39396 22428 40124 22484
rect 40180 22428 40190 22484
rect 41570 22428 41580 22484
rect 41636 22428 44268 22484
rect 44324 22428 48748 22484
rect 48804 22428 48814 22484
rect 55682 22428 55692 22484
rect 55748 22428 58156 22484
rect 58212 22428 58222 22484
rect 5954 22316 5964 22372
rect 6020 22316 12348 22372
rect 12404 22316 12414 22372
rect 17714 22316 17724 22372
rect 17780 22316 21644 22372
rect 21700 22316 22652 22372
rect 22708 22316 22718 22372
rect 32722 22316 32732 22372
rect 32788 22316 33740 22372
rect 33796 22316 33806 22372
rect 48962 22316 48972 22372
rect 49028 22316 49308 22372
rect 49364 22316 49374 22372
rect 51202 22316 51212 22372
rect 51268 22316 52108 22372
rect 52164 22316 52780 22372
rect 52836 22316 52846 22372
rect 31490 22204 31500 22260
rect 31556 22204 32508 22260
rect 32564 22204 33404 22260
rect 33460 22204 33470 22260
rect 4834 22092 4844 22148
rect 4900 22092 6188 22148
rect 6244 22092 6860 22148
rect 6916 22092 6926 22148
rect 16146 21980 16156 22036
rect 16212 21980 16716 22036
rect 16772 21980 16782 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 10770 21756 10780 21812
rect 10836 21756 12796 21812
rect 12852 21756 12862 21812
rect 13458 21756 13468 21812
rect 13524 21756 14700 21812
rect 14756 21756 14766 21812
rect 38770 21756 38780 21812
rect 38836 21756 39676 21812
rect 39732 21756 40908 21812
rect 40964 21756 40974 21812
rect 1810 21644 1820 21700
rect 1876 21644 6412 21700
rect 6468 21644 6478 21700
rect 37426 21644 37436 21700
rect 37492 21644 37996 21700
rect 38052 21644 38062 21700
rect 42466 21644 42476 21700
rect 42532 21644 43372 21700
rect 43428 21644 57820 21700
rect 57876 21644 57886 21700
rect 13234 21532 13244 21588
rect 13300 21532 14476 21588
rect 14532 21532 16604 21588
rect 16660 21532 17388 21588
rect 17444 21532 17454 21588
rect 22978 21532 22988 21588
rect 23044 21532 23548 21588
rect 23604 21532 24108 21588
rect 24164 21532 24174 21588
rect 36530 21532 36540 21588
rect 36596 21532 37324 21588
rect 37380 21532 37390 21588
rect 39106 21532 39116 21588
rect 39172 21532 41356 21588
rect 41412 21532 41422 21588
rect 44594 21532 44604 21588
rect 44660 21532 45388 21588
rect 45444 21532 45454 21588
rect 53890 21532 53900 21588
rect 53956 21532 55244 21588
rect 55300 21532 55310 21588
rect 23202 21420 23212 21476
rect 23268 21420 23772 21476
rect 23828 21420 23838 21476
rect 25330 21420 25340 21476
rect 25396 21420 26012 21476
rect 26068 21420 26348 21476
rect 26404 21420 26796 21476
rect 26852 21420 26862 21476
rect 34626 21420 34636 21476
rect 34692 21420 36652 21476
rect 36708 21420 36718 21476
rect 38882 21420 38892 21476
rect 38948 21420 39788 21476
rect 39844 21420 42924 21476
rect 42980 21420 42990 21476
rect 48178 21420 48188 21476
rect 48244 21420 49420 21476
rect 49476 21420 49486 21476
rect 37090 21308 37100 21364
rect 37156 21308 37660 21364
rect 37716 21308 37726 21364
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 59200 21140 60000 21168
rect 58146 21084 58156 21140
rect 58212 21084 60000 21140
rect 59200 21056 60000 21084
rect 17938 20972 17948 21028
rect 18004 20972 18284 21028
rect 18340 20972 19180 21028
rect 19236 20972 19246 21028
rect 22642 20972 22652 21028
rect 22708 20972 23436 21028
rect 23492 20972 23502 21028
rect 39218 20860 39228 20916
rect 39284 20860 39788 20916
rect 39844 20860 40684 20916
rect 40740 20860 40750 20916
rect 12674 20748 12684 20804
rect 12740 20748 13132 20804
rect 13188 20748 13468 20804
rect 13524 20748 14140 20804
rect 14196 20748 14206 20804
rect 22418 20748 22428 20804
rect 22484 20748 23212 20804
rect 23268 20748 23828 20804
rect 35074 20748 35084 20804
rect 35140 20748 35980 20804
rect 36036 20748 36046 20804
rect 23772 20692 23828 20748
rect 5058 20636 5068 20692
rect 5124 20636 7308 20692
rect 7364 20636 7374 20692
rect 23762 20636 23772 20692
rect 23828 20636 23838 20692
rect 35746 20636 35756 20692
rect 35812 20636 38668 20692
rect 38612 20580 38668 20636
rect 12898 20524 12908 20580
rect 12964 20524 13692 20580
rect 13748 20524 13758 20580
rect 37090 20524 37100 20580
rect 37156 20524 37884 20580
rect 37940 20524 37950 20580
rect 38612 20524 39340 20580
rect 39396 20524 44156 20580
rect 44212 20524 44222 20580
rect 50866 20524 50876 20580
rect 50932 20524 52220 20580
rect 52276 20524 52892 20580
rect 52948 20524 52958 20580
rect 6626 20412 6636 20468
rect 6692 20412 6972 20468
rect 7028 20412 15148 20468
rect 15204 20412 15820 20468
rect 15876 20412 15886 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 8642 20300 8652 20356
rect 8708 20300 13580 20356
rect 13636 20300 13646 20356
rect 32498 20300 32508 20356
rect 32564 20300 35980 20356
rect 36036 20300 36046 20356
rect 13570 20076 13580 20132
rect 13636 20076 14028 20132
rect 14084 20076 14094 20132
rect 17602 20076 17612 20132
rect 17668 20076 18844 20132
rect 18900 20076 19404 20132
rect 19460 20076 19470 20132
rect 20132 20076 20524 20132
rect 20580 20076 27916 20132
rect 27972 20076 27982 20132
rect 33058 20076 33068 20132
rect 33124 20076 34300 20132
rect 34356 20076 34366 20132
rect 41906 20076 41916 20132
rect 41972 20076 42364 20132
rect 42420 20076 43148 20132
rect 43204 20076 43214 20132
rect 54898 20076 54908 20132
rect 54964 20076 56140 20132
rect 56196 20076 56206 20132
rect 4498 19964 4508 20020
rect 4564 19964 6300 20020
rect 6356 19964 6366 20020
rect 20066 19964 20076 20020
rect 20132 19964 20188 20076
rect 21186 19964 21196 20020
rect 21252 19964 25900 20020
rect 25956 19964 25966 20020
rect 26450 19964 26460 20020
rect 26516 19964 26908 20020
rect 26964 19964 27692 20020
rect 27748 19964 27758 20020
rect 29810 19964 29820 20020
rect 29876 19964 31500 20020
rect 31556 19964 31566 20020
rect 49186 19964 49196 20020
rect 49252 19964 49868 20020
rect 49924 19964 49934 20020
rect 25900 19908 25956 19964
rect 10322 19852 10332 19908
rect 10388 19852 13916 19908
rect 13972 19852 13982 19908
rect 25900 19852 26348 19908
rect 26404 19852 26414 19908
rect 28242 19852 28252 19908
rect 28308 19852 28318 19908
rect 30146 19852 30156 19908
rect 30212 19852 30828 19908
rect 30884 19852 30894 19908
rect 32274 19852 32284 19908
rect 32340 19852 32956 19908
rect 33012 19852 33022 19908
rect 35308 19852 40460 19908
rect 40516 19852 40526 19908
rect 42802 19852 42812 19908
rect 42868 19852 43148 19908
rect 43204 19852 43214 19908
rect 54674 19852 54684 19908
rect 54740 19852 55468 19908
rect 55524 19852 55534 19908
rect 28252 19796 28308 19852
rect 35308 19796 35364 19852
rect 8754 19740 8764 19796
rect 8820 19740 9996 19796
rect 10052 19740 10062 19796
rect 16594 19740 16604 19796
rect 16660 19740 17388 19796
rect 17444 19740 17454 19796
rect 28252 19740 35364 19796
rect 37426 19740 37436 19796
rect 37492 19740 42588 19796
rect 42644 19740 42654 19796
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 22530 19516 22540 19572
rect 22596 19516 27692 19572
rect 27748 19516 27758 19572
rect 27346 19404 27356 19460
rect 27412 19404 37324 19460
rect 37380 19404 37390 19460
rect 37986 19404 37996 19460
rect 38052 19404 38556 19460
rect 38612 19404 38622 19460
rect 14914 19292 14924 19348
rect 14980 19292 16492 19348
rect 16548 19292 16558 19348
rect 32946 19292 32956 19348
rect 33012 19292 42140 19348
rect 42196 19292 44716 19348
rect 44772 19292 44782 19348
rect 48626 19292 48636 19348
rect 48692 19292 49420 19348
rect 49476 19292 49486 19348
rect 52994 19292 53004 19348
rect 53060 19292 53788 19348
rect 53844 19292 53854 19348
rect 54450 19292 54460 19348
rect 54516 19292 58156 19348
rect 58212 19292 58222 19348
rect 22978 19180 22988 19236
rect 23044 19180 24444 19236
rect 24500 19180 24510 19236
rect 27346 19180 27356 19236
rect 27412 19180 29260 19236
rect 29316 19180 29326 19236
rect 38406 19180 38444 19236
rect 38500 19180 38510 19236
rect 42578 19180 42588 19236
rect 42644 19180 43036 19236
rect 43092 19180 43102 19236
rect 44482 19180 44492 19236
rect 44548 19180 45500 19236
rect 45556 19180 46620 19236
rect 46676 19180 46686 19236
rect 52098 19180 52108 19236
rect 52164 19180 52556 19236
rect 52612 19180 52622 19236
rect 54002 19180 54012 19236
rect 54068 19180 54684 19236
rect 54740 19180 55916 19236
rect 55972 19180 55982 19236
rect 20738 19068 20748 19124
rect 20804 19068 22540 19124
rect 22596 19068 22606 19124
rect 31602 19068 31612 19124
rect 31668 19068 32620 19124
rect 32676 19068 32686 19124
rect 34738 19068 34748 19124
rect 34804 19068 37100 19124
rect 37156 19068 37996 19124
rect 38052 19068 38062 19124
rect 48290 19068 48300 19124
rect 48356 19068 49532 19124
rect 49588 19068 53116 19124
rect 53172 19068 54460 19124
rect 54516 19068 54526 19124
rect 13570 18956 13580 19012
rect 13636 18956 14252 19012
rect 14308 18956 14318 19012
rect 18162 18956 18172 19012
rect 18228 18956 21868 19012
rect 21924 18956 21934 19012
rect 38434 18956 38444 19012
rect 38500 18956 40348 19012
rect 40404 18956 41020 19012
rect 41076 18956 41086 19012
rect 43474 18956 43484 19012
rect 43540 18956 43932 19012
rect 43988 18956 43998 19012
rect 44258 18956 44268 19012
rect 44324 18956 45276 19012
rect 45332 18956 45342 19012
rect 49186 18956 49196 19012
rect 49252 18956 52668 19012
rect 52724 18956 54796 19012
rect 54852 18956 55132 19012
rect 55188 18956 55198 19012
rect 38322 18844 38332 18900
rect 38388 18844 38398 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 16482 18620 16492 18676
rect 16548 18620 17388 18676
rect 17444 18620 17454 18676
rect 18274 18620 18284 18676
rect 18340 18620 19068 18676
rect 19124 18620 19134 18676
rect 38332 18564 38388 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 40450 18620 40460 18676
rect 40516 18620 41916 18676
rect 41972 18620 41982 18676
rect 42242 18620 42252 18676
rect 42308 18620 43036 18676
rect 43092 18620 47964 18676
rect 48020 18620 48030 18676
rect 17938 18508 17948 18564
rect 18004 18508 18396 18564
rect 18452 18508 18956 18564
rect 19012 18508 19022 18564
rect 32162 18508 32172 18564
rect 32228 18508 33628 18564
rect 33684 18508 33694 18564
rect 38332 18508 38556 18564
rect 38612 18508 38622 18564
rect 49410 18508 49420 18564
rect 49476 18508 50428 18564
rect 50484 18508 50494 18564
rect 7410 18396 7420 18452
rect 7476 18396 9660 18452
rect 9716 18396 10220 18452
rect 10276 18396 10286 18452
rect 13458 18396 13468 18452
rect 13524 18396 13692 18452
rect 13748 18396 13758 18452
rect 14018 18396 14028 18452
rect 14084 18396 14700 18452
rect 14756 18396 16716 18452
rect 16772 18396 17612 18452
rect 17668 18396 17678 18452
rect 23538 18396 23548 18452
rect 23604 18396 25228 18452
rect 25284 18396 25294 18452
rect 33506 18396 33516 18452
rect 33572 18396 34524 18452
rect 34580 18396 34590 18452
rect 34748 18396 40684 18452
rect 40740 18396 40750 18452
rect 41682 18396 41692 18452
rect 41748 18396 43260 18452
rect 43316 18396 43326 18452
rect 55458 18396 55468 18452
rect 55524 18396 55534 18452
rect 34748 18340 34804 18396
rect 55468 18340 55524 18396
rect 3154 18284 3164 18340
rect 3220 18284 3612 18340
rect 3668 18284 3678 18340
rect 4498 18284 4508 18340
rect 4564 18284 6636 18340
rect 6692 18284 7756 18340
rect 7812 18284 7822 18340
rect 10994 18284 11004 18340
rect 11060 18284 14476 18340
rect 14532 18284 14542 18340
rect 20178 18284 20188 18340
rect 20244 18284 22316 18340
rect 22372 18284 22764 18340
rect 22820 18284 22830 18340
rect 32050 18284 32060 18340
rect 32116 18284 32732 18340
rect 32788 18284 34804 18340
rect 35074 18284 35084 18340
rect 35140 18284 36092 18340
rect 36148 18284 36158 18340
rect 37986 18284 37996 18340
rect 38052 18284 38444 18340
rect 38500 18284 39116 18340
rect 39172 18284 40124 18340
rect 40180 18284 40190 18340
rect 45378 18284 45388 18340
rect 45444 18284 45724 18340
rect 45780 18284 45790 18340
rect 55234 18284 55244 18340
rect 55300 18284 55524 18340
rect 22764 18228 22820 18284
rect 6850 18172 6860 18228
rect 6916 18172 7980 18228
rect 8036 18172 8046 18228
rect 14130 18172 14140 18228
rect 14196 18172 16044 18228
rect 16100 18172 16110 18228
rect 22764 18172 24108 18228
rect 24164 18172 24174 18228
rect 25340 18172 27020 18228
rect 27076 18172 27086 18228
rect 33842 18172 33852 18228
rect 33908 18172 34972 18228
rect 35028 18172 35038 18228
rect 35522 18172 35532 18228
rect 35588 18172 37212 18228
rect 37268 18172 37548 18228
rect 37604 18172 37614 18228
rect 42466 18172 42476 18228
rect 42532 18172 48188 18228
rect 48244 18172 48748 18228
rect 48804 18172 48814 18228
rect 25340 18116 25396 18172
rect 25330 18060 25340 18116
rect 25396 18060 25406 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 26852 17892 26908 18172
rect 43250 18060 43260 18116
rect 43316 18060 43820 18116
rect 43876 18060 43886 18116
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 26852 17836 31836 17892
rect 31892 17836 51436 17892
rect 51492 17836 51502 17892
rect 32162 17724 32172 17780
rect 32228 17724 33180 17780
rect 33236 17724 33246 17780
rect 36194 17724 36204 17780
rect 36260 17724 37884 17780
rect 37940 17724 37950 17780
rect 41010 17724 41020 17780
rect 41076 17724 46956 17780
rect 47012 17724 47852 17780
rect 47908 17724 47918 17780
rect 17826 17612 17836 17668
rect 17892 17612 18620 17668
rect 18676 17612 18686 17668
rect 52098 17612 52108 17668
rect 52164 17612 52892 17668
rect 52948 17612 52958 17668
rect 6402 17500 6412 17556
rect 6468 17500 6748 17556
rect 6804 17500 7420 17556
rect 7476 17500 7486 17556
rect 18050 17500 18060 17556
rect 18116 17500 19180 17556
rect 19236 17500 19246 17556
rect 27570 17500 27580 17556
rect 27636 17500 27916 17556
rect 27972 17500 29372 17556
rect 29428 17500 29438 17556
rect 44146 17500 44156 17556
rect 44212 17500 45276 17556
rect 45332 17500 52780 17556
rect 52836 17500 52846 17556
rect 15922 17388 15932 17444
rect 15988 17388 20412 17444
rect 20468 17388 21420 17444
rect 21476 17388 21486 17444
rect 51874 17388 51884 17444
rect 51940 17388 53228 17444
rect 53284 17388 54012 17444
rect 54068 17388 54078 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 15138 17052 15148 17108
rect 15204 17052 15708 17108
rect 15764 17052 15774 17108
rect 23314 17052 23324 17108
rect 23380 17052 23884 17108
rect 23940 17052 26236 17108
rect 26292 17052 26302 17108
rect 30034 17052 30044 17108
rect 30100 17052 30716 17108
rect 30772 17052 30782 17108
rect 24658 16940 24668 16996
rect 24724 16940 25340 16996
rect 25396 16940 25406 16996
rect 32610 16940 32620 16996
rect 32676 16940 41916 16996
rect 41972 16940 43260 16996
rect 43316 16940 43326 16996
rect 45714 16940 45724 16996
rect 45780 16940 48748 16996
rect 48804 16940 48814 16996
rect 52434 16940 52444 16996
rect 52500 16940 54460 16996
rect 54516 16940 54526 16996
rect 13794 16828 13804 16884
rect 13860 16828 15260 16884
rect 15316 16828 16828 16884
rect 16884 16828 16894 16884
rect 37650 16828 37660 16884
rect 37716 16828 41468 16884
rect 41524 16828 41804 16884
rect 41860 16828 46172 16884
rect 46228 16828 46238 16884
rect 46722 16828 46732 16884
rect 46788 16828 47516 16884
rect 47572 16828 47582 16884
rect 51202 16828 51212 16884
rect 51268 16828 51660 16884
rect 51716 16828 55356 16884
rect 55412 16828 55422 16884
rect 16034 16716 16044 16772
rect 16100 16716 18284 16772
rect 18340 16716 18350 16772
rect 29586 16716 29596 16772
rect 29652 16716 30828 16772
rect 30884 16716 30894 16772
rect 47282 16716 47292 16772
rect 47348 16716 48188 16772
rect 48244 16716 48254 16772
rect 14802 16604 14812 16660
rect 14868 16604 15372 16660
rect 15428 16604 22988 16660
rect 23044 16604 24332 16660
rect 24388 16604 24398 16660
rect 48290 16604 48300 16660
rect 48356 16604 52668 16660
rect 52724 16604 52734 16660
rect 9202 16492 9212 16548
rect 9268 16492 25788 16548
rect 25844 16492 27020 16548
rect 27076 16492 27804 16548
rect 27860 16492 27870 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 14690 16156 14700 16212
rect 14756 16156 17052 16212
rect 17108 16156 17118 16212
rect 48178 16156 48188 16212
rect 48244 16156 48860 16212
rect 48916 16156 48926 16212
rect 49634 16156 49644 16212
rect 49700 16156 50988 16212
rect 51044 16156 51054 16212
rect 54002 16156 54012 16212
rect 54068 16156 58156 16212
rect 58212 16156 58222 16212
rect 7970 16044 7980 16100
rect 8036 16044 8540 16100
rect 8596 16044 8876 16100
rect 8932 16044 8942 16100
rect 10322 16044 10332 16100
rect 10388 16044 11676 16100
rect 11732 16044 11742 16100
rect 14466 16044 14476 16100
rect 14532 16044 15036 16100
rect 15092 16044 15102 16100
rect 24322 16044 24332 16100
rect 24388 16044 25004 16100
rect 25060 16044 25070 16100
rect 35970 16044 35980 16100
rect 36036 16044 37548 16100
rect 37604 16044 37614 16100
rect 38322 16044 38332 16100
rect 38388 16044 41804 16100
rect 41860 16044 41870 16100
rect 36418 15932 36428 15988
rect 36484 15932 37660 15988
rect 37716 15932 37726 15988
rect 44034 15932 44044 15988
rect 44100 15932 46844 15988
rect 46900 15932 46910 15988
rect 53778 15932 53788 15988
rect 53844 15932 54572 15988
rect 54628 15932 54638 15988
rect 5506 15820 5516 15876
rect 5572 15820 6972 15876
rect 7028 15820 7038 15876
rect 23426 15820 23436 15876
rect 23492 15820 24332 15876
rect 24388 15820 24398 15876
rect 36082 15820 36092 15876
rect 36148 15820 37772 15876
rect 37828 15820 38108 15876
rect 38164 15820 38174 15876
rect 43474 15820 43484 15876
rect 43540 15820 46732 15876
rect 46788 15820 46798 15876
rect 8530 15708 8540 15764
rect 8596 15708 9548 15764
rect 9604 15708 9614 15764
rect 36306 15708 36316 15764
rect 36372 15708 38444 15764
rect 38500 15708 38510 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 30818 15596 30828 15652
rect 30884 15596 31164 15652
rect 31220 15596 31230 15652
rect 10098 15484 10108 15540
rect 10164 15484 11004 15540
rect 11060 15484 11070 15540
rect 6738 15372 6748 15428
rect 6804 15372 7420 15428
rect 7476 15372 7980 15428
rect 8036 15372 8046 15428
rect 9986 15372 9996 15428
rect 10052 15372 10556 15428
rect 10612 15372 20188 15428
rect 20244 15372 20254 15428
rect 28130 15372 28140 15428
rect 28196 15372 28924 15428
rect 28980 15372 35308 15428
rect 35364 15372 35374 15428
rect 42802 15372 42812 15428
rect 42868 15372 57820 15428
rect 57876 15372 57886 15428
rect 59200 15316 60000 15344
rect 25666 15260 25676 15316
rect 25732 15260 31388 15316
rect 31444 15260 31454 15316
rect 35522 15260 35532 15316
rect 35588 15260 36652 15316
rect 36708 15260 36718 15316
rect 48738 15260 48748 15316
rect 48804 15260 49812 15316
rect 57586 15260 57596 15316
rect 57652 15260 58156 15316
rect 58212 15260 60000 15316
rect 49756 15204 49812 15260
rect 59200 15232 60000 15260
rect 8194 15148 8204 15204
rect 8260 15148 9772 15204
rect 9828 15148 9838 15204
rect 11106 15148 11116 15204
rect 11172 15148 13356 15204
rect 13412 15148 13422 15204
rect 23874 15148 23884 15204
rect 23940 15148 28588 15204
rect 28644 15148 28654 15204
rect 31490 15148 31500 15204
rect 31556 15148 31948 15204
rect 32004 15148 32508 15204
rect 32564 15148 33404 15204
rect 33460 15148 34076 15204
rect 34132 15148 34142 15204
rect 48178 15148 48188 15204
rect 48244 15148 48972 15204
rect 49028 15148 49038 15204
rect 49746 15148 49756 15204
rect 49812 15148 54348 15204
rect 54404 15148 54414 15204
rect 22754 15036 22764 15092
rect 22820 15036 23660 15092
rect 23716 15036 23726 15092
rect 28130 15036 28140 15092
rect 28196 15036 28420 15092
rect 28690 15036 28700 15092
rect 28756 15036 29596 15092
rect 29652 15036 29662 15092
rect 52434 15036 52444 15092
rect 52500 15036 52780 15092
rect 52836 15036 53452 15092
rect 53508 15036 53518 15092
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 28364 14868 28420 15036
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 28354 14812 28364 14868
rect 28420 14812 28430 14868
rect 50372 14812 51884 14868
rect 51940 14812 58156 14868
rect 58212 14812 58222 14868
rect 50372 14756 50428 14812
rect 49298 14700 49308 14756
rect 49364 14700 50428 14756
rect 16706 14588 16716 14644
rect 16772 14588 22988 14644
rect 23044 14588 23054 14644
rect 36978 14588 36988 14644
rect 37044 14588 37884 14644
rect 37940 14588 37950 14644
rect 44258 14588 44268 14644
rect 44324 14588 45052 14644
rect 45108 14588 45118 14644
rect 50540 14588 51884 14644
rect 51940 14588 51950 14644
rect 54898 14588 54908 14644
rect 54964 14588 56028 14644
rect 56084 14588 56094 14644
rect 50540 14532 50596 14588
rect 13234 14476 13244 14532
rect 13300 14476 14028 14532
rect 14084 14476 15484 14532
rect 15540 14476 15550 14532
rect 20738 14476 20748 14532
rect 20804 14476 22764 14532
rect 22820 14476 22830 14532
rect 39890 14476 39900 14532
rect 39956 14476 40236 14532
rect 40292 14476 40908 14532
rect 40964 14476 40974 14532
rect 46946 14476 46956 14532
rect 47012 14476 48636 14532
rect 48692 14476 50540 14532
rect 50596 14476 50606 14532
rect 51986 14476 51996 14532
rect 52052 14476 53340 14532
rect 53396 14476 53406 14532
rect 17714 14364 17724 14420
rect 17780 14364 20188 14420
rect 20244 14364 20254 14420
rect 22978 14364 22988 14420
rect 23044 14364 24668 14420
rect 24724 14364 24734 14420
rect 33506 14364 33516 14420
rect 33572 14364 37996 14420
rect 38052 14364 38062 14420
rect 15250 14252 15260 14308
rect 15316 14252 16492 14308
rect 16548 14252 16558 14308
rect 19730 14252 19740 14308
rect 19796 14252 20524 14308
rect 20580 14252 20590 14308
rect 34962 14252 34972 14308
rect 35028 14252 36204 14308
rect 36260 14252 36270 14308
rect 54898 14252 54908 14308
rect 54964 14252 55692 14308
rect 55748 14252 55758 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 4162 13916 4172 13972
rect 4228 13916 4620 13972
rect 4676 13916 5068 13972
rect 5124 13916 6636 13972
rect 6692 13916 6702 13972
rect 15474 13916 15484 13972
rect 15540 13916 16380 13972
rect 16436 13916 17388 13972
rect 17444 13916 17454 13972
rect 23762 13916 23772 13972
rect 23828 13916 24668 13972
rect 24724 13916 25228 13972
rect 25284 13916 25294 13972
rect 41682 13916 41692 13972
rect 41748 13916 42140 13972
rect 42196 13916 42700 13972
rect 42756 13916 42766 13972
rect 51202 13916 51212 13972
rect 51268 13916 51996 13972
rect 52052 13916 52062 13972
rect 16258 13804 16268 13860
rect 16324 13804 22540 13860
rect 22596 13804 22606 13860
rect 23650 13804 23660 13860
rect 23716 13804 25452 13860
rect 25508 13804 25518 13860
rect 34850 13804 34860 13860
rect 34916 13804 35644 13860
rect 35700 13804 35710 13860
rect 41906 13804 41916 13860
rect 41972 13804 43820 13860
rect 43876 13804 44828 13860
rect 44884 13804 44894 13860
rect 13682 13692 13692 13748
rect 13748 13692 15708 13748
rect 15764 13692 15774 13748
rect 16818 13692 16828 13748
rect 16884 13692 18172 13748
rect 18228 13692 21868 13748
rect 21924 13692 23436 13748
rect 23492 13692 26908 13748
rect 26964 13692 28476 13748
rect 28532 13692 28542 13748
rect 34402 13692 34412 13748
rect 34468 13692 35980 13748
rect 36036 13692 36046 13748
rect 40338 13692 40348 13748
rect 40404 13692 41468 13748
rect 41524 13692 41534 13748
rect 45714 13692 45724 13748
rect 45780 13692 46284 13748
rect 46340 13692 46350 13748
rect 48066 13692 48076 13748
rect 48132 13692 49308 13748
rect 49364 13692 49374 13748
rect 49522 13692 49532 13748
rect 49588 13692 50540 13748
rect 50596 13692 50606 13748
rect 52434 13692 52444 13748
rect 52500 13692 53228 13748
rect 53284 13692 53294 13748
rect 3266 13580 3276 13636
rect 3332 13580 3724 13636
rect 3780 13580 3790 13636
rect 13234 13580 13244 13636
rect 13300 13580 13580 13636
rect 13636 13580 13646 13636
rect 17602 13580 17612 13636
rect 17668 13580 19180 13636
rect 19236 13580 19246 13636
rect 49746 13580 49756 13636
rect 49812 13580 51884 13636
rect 51940 13580 52892 13636
rect 52948 13580 52958 13636
rect 3042 13468 3052 13524
rect 3108 13468 3948 13524
rect 4004 13468 4014 13524
rect 28588 13468 29596 13524
rect 29652 13468 29662 13524
rect 34290 13468 34300 13524
rect 34356 13468 35756 13524
rect 35812 13468 35822 13524
rect 36194 13468 36204 13524
rect 36260 13468 40908 13524
rect 40964 13468 40974 13524
rect 42690 13468 42700 13524
rect 42756 13468 43484 13524
rect 43540 13468 43550 13524
rect 49186 13468 49196 13524
rect 49252 13468 50092 13524
rect 50148 13468 50158 13524
rect 28588 13412 28644 13468
rect 26562 13356 26572 13412
rect 26628 13356 28252 13412
rect 28308 13356 28644 13412
rect 40002 13356 40012 13412
rect 40068 13356 45948 13412
rect 46004 13356 46014 13412
rect 52882 13356 52892 13412
rect 52948 13356 53340 13412
rect 53396 13356 53406 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 41346 13244 41356 13300
rect 41412 13244 42028 13300
rect 42084 13244 42476 13300
rect 42532 13244 42542 13300
rect 28242 13132 28252 13188
rect 28308 13132 30828 13188
rect 30884 13132 31836 13188
rect 31892 13132 31902 13188
rect 33058 13132 33068 13188
rect 33124 13132 37884 13188
rect 37940 13132 39116 13188
rect 39172 13132 39182 13188
rect 45378 13132 45388 13188
rect 45444 13132 47180 13188
rect 47236 13132 47246 13188
rect 21410 13020 21420 13076
rect 21476 13020 22092 13076
rect 22148 13020 22876 13076
rect 22932 13020 22942 13076
rect 24770 13020 24780 13076
rect 24836 13020 25788 13076
rect 25844 13020 25854 13076
rect 28018 13020 28028 13076
rect 28084 13020 29820 13076
rect 29876 13020 29886 13076
rect 36082 13020 36092 13076
rect 36148 13020 37100 13076
rect 37156 13020 37166 13076
rect 37650 13020 37660 13076
rect 37716 13020 38668 13076
rect 38724 13020 38734 13076
rect 26852 12908 28588 12964
rect 28644 12908 28654 12964
rect 30146 12908 30156 12964
rect 30212 12908 30716 12964
rect 30772 12908 30782 12964
rect 31602 12908 31612 12964
rect 31668 12908 33852 12964
rect 33908 12908 34636 12964
rect 34692 12908 35532 12964
rect 35588 12908 35598 12964
rect 49074 12908 49084 12964
rect 49140 12908 50988 12964
rect 51044 12908 51054 12964
rect 26852 12852 26908 12908
rect 22866 12796 22876 12852
rect 22932 12796 26908 12852
rect 29698 12796 29708 12852
rect 29764 12796 30380 12852
rect 30436 12796 30828 12852
rect 30884 12796 33516 12852
rect 33572 12796 33582 12852
rect 46386 12796 46396 12852
rect 46452 12796 49756 12852
rect 49812 12796 49822 12852
rect 52882 12796 52892 12852
rect 52948 12796 53340 12852
rect 53396 12796 58156 12852
rect 58212 12796 58222 12852
rect 2482 12684 2492 12740
rect 2548 12684 4396 12740
rect 4452 12684 4462 12740
rect 20066 12684 20076 12740
rect 20132 12684 21980 12740
rect 22036 12684 34748 12740
rect 34804 12684 45052 12740
rect 45108 12684 45118 12740
rect 45938 12684 45948 12740
rect 46004 12684 46844 12740
rect 46900 12684 46910 12740
rect 49970 12684 49980 12740
rect 50036 12684 50876 12740
rect 50932 12684 50942 12740
rect 52770 12684 52780 12740
rect 52836 12684 53900 12740
rect 53956 12684 53966 12740
rect 54226 12684 54236 12740
rect 54292 12684 54460 12740
rect 54516 12684 54526 12740
rect 8194 12572 8204 12628
rect 8260 12572 10220 12628
rect 10276 12572 13468 12628
rect 13524 12572 13916 12628
rect 13972 12572 13982 12628
rect 41346 12572 41356 12628
rect 41412 12572 41916 12628
rect 41972 12572 49196 12628
rect 49252 12572 50204 12628
rect 50260 12572 50270 12628
rect 54674 12572 54684 12628
rect 54740 12572 55132 12628
rect 55188 12572 55198 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 40450 12460 40460 12516
rect 40516 12460 40908 12516
rect 40964 12460 42420 12516
rect 54422 12460 54460 12516
rect 54516 12460 55020 12516
rect 55076 12460 55086 12516
rect 42364 12404 42420 12460
rect 8306 12348 8316 12404
rect 8372 12348 9436 12404
rect 9492 12348 9502 12404
rect 15922 12348 15932 12404
rect 15988 12348 17500 12404
rect 17556 12348 17566 12404
rect 41346 12348 41356 12404
rect 41412 12348 42140 12404
rect 42196 12348 42206 12404
rect 42354 12348 42364 12404
rect 42420 12348 42924 12404
rect 42980 12348 42990 12404
rect 47282 12348 47292 12404
rect 47348 12348 47740 12404
rect 47796 12348 48972 12404
rect 49028 12348 49038 12404
rect 3332 12236 4844 12292
rect 4900 12236 6300 12292
rect 6356 12236 6366 12292
rect 14252 12236 14924 12292
rect 14980 12236 14990 12292
rect 45154 12236 45164 12292
rect 45220 12236 45724 12292
rect 45780 12236 45790 12292
rect 46722 12236 46732 12292
rect 46788 12236 47068 12292
rect 47124 12236 47134 12292
rect 48178 12236 48188 12292
rect 48244 12236 49308 12292
rect 49364 12236 49374 12292
rect 52098 12236 52108 12292
rect 52164 12236 52780 12292
rect 52836 12236 52846 12292
rect 3332 12068 3388 12236
rect 14252 12180 14308 12236
rect 45724 12180 45780 12236
rect 8642 12124 8652 12180
rect 8708 12124 9212 12180
rect 9268 12124 9772 12180
rect 9828 12124 9996 12180
rect 10052 12124 10062 12180
rect 12226 12124 12236 12180
rect 12292 12124 13468 12180
rect 13524 12124 14252 12180
rect 14308 12124 14318 12180
rect 14578 12124 14588 12180
rect 14644 12124 15596 12180
rect 15652 12124 15662 12180
rect 37986 12124 37996 12180
rect 38052 12124 41580 12180
rect 41636 12124 41646 12180
rect 45724 12124 46620 12180
rect 46676 12124 46686 12180
rect 47954 12124 47964 12180
rect 48020 12124 49420 12180
rect 49476 12124 50204 12180
rect 50260 12124 50270 12180
rect 54562 12124 54572 12180
rect 54628 12124 55356 12180
rect 55412 12124 55422 12180
rect 41580 12068 41636 12124
rect 1810 12012 1820 12068
rect 1876 12012 3388 12068
rect 10770 12012 10780 12068
rect 10836 12012 12348 12068
rect 12404 12012 12414 12068
rect 40002 12012 40012 12068
rect 40068 12012 41244 12068
rect 41300 12012 41310 12068
rect 41580 12012 45836 12068
rect 45892 12012 45902 12068
rect 48178 12012 48188 12068
rect 48244 12012 49084 12068
rect 49140 12012 49150 12068
rect 35186 11900 35196 11956
rect 35252 11900 36988 11956
rect 37044 11900 37054 11956
rect 39218 11900 39228 11956
rect 39284 11900 40572 11956
rect 40628 11900 41132 11956
rect 41188 11900 41198 11956
rect 41906 11900 41916 11956
rect 41972 11900 42476 11956
rect 42532 11900 42542 11956
rect 53330 11900 53340 11956
rect 53396 11900 54012 11956
rect 54068 11900 54078 11956
rect 10322 11788 10332 11844
rect 10388 11788 14028 11844
rect 14084 11788 14700 11844
rect 14756 11788 14766 11844
rect 19170 11788 19180 11844
rect 19236 11788 19246 11844
rect 38210 11788 38220 11844
rect 38276 11788 54236 11844
rect 54292 11788 54302 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 19180 11732 19236 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 15474 11676 15484 11732
rect 15540 11676 21308 11732
rect 21364 11676 21374 11732
rect 48066 11676 48076 11732
rect 48132 11676 50876 11732
rect 50932 11676 50942 11732
rect 46946 11564 46956 11620
rect 47012 11564 48748 11620
rect 48804 11564 48814 11620
rect 4834 11452 4844 11508
rect 4900 11452 5740 11508
rect 5796 11452 5806 11508
rect 7074 11452 7084 11508
rect 7140 11452 8428 11508
rect 8484 11452 8494 11508
rect 12786 11452 12796 11508
rect 12852 11452 13580 11508
rect 13636 11452 13646 11508
rect 14914 11452 14924 11508
rect 14980 11452 16156 11508
rect 16212 11452 16222 11508
rect 21522 11452 21532 11508
rect 21588 11452 25116 11508
rect 25172 11452 25182 11508
rect 53106 11452 53116 11508
rect 53172 11452 54012 11508
rect 54068 11452 55244 11508
rect 55300 11452 55310 11508
rect 55682 11452 55692 11508
rect 55748 11452 57372 11508
rect 57428 11452 57438 11508
rect 4610 11340 4620 11396
rect 4676 11340 5852 11396
rect 5908 11340 5918 11396
rect 12898 11340 12908 11396
rect 12964 11340 13692 11396
rect 13748 11340 14476 11396
rect 14532 11340 14542 11396
rect 31154 11340 31164 11396
rect 31220 11340 34636 11396
rect 34692 11340 34702 11396
rect 50194 11340 50204 11396
rect 50260 11340 50428 11396
rect 55458 11340 55468 11396
rect 55524 11340 58044 11396
rect 58100 11340 58110 11396
rect 50372 11284 50428 11340
rect 3938 11228 3948 11284
rect 4004 11228 5628 11284
rect 5684 11228 5694 11284
rect 25330 11228 25340 11284
rect 25396 11228 26460 11284
rect 26516 11228 26526 11284
rect 50372 11228 51436 11284
rect 51492 11228 53004 11284
rect 53060 11228 53070 11284
rect 8754 11116 8764 11172
rect 8820 11116 9324 11172
rect 9380 11116 14924 11172
rect 14980 11116 14990 11172
rect 24770 11116 24780 11172
rect 24836 11116 25676 11172
rect 25732 11116 31836 11172
rect 31892 11116 38220 11172
rect 38276 11116 39004 11172
rect 39060 11116 39070 11172
rect 50306 11116 50316 11172
rect 50372 11116 51324 11172
rect 51380 11116 51390 11172
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 46498 10892 46508 10948
rect 46564 10892 47180 10948
rect 47236 10892 47246 10948
rect 4162 10780 4172 10836
rect 4228 10780 5516 10836
rect 5572 10780 5582 10836
rect 35858 10780 35868 10836
rect 35924 10780 37436 10836
rect 37492 10780 37502 10836
rect 42466 10780 42476 10836
rect 42532 10780 45836 10836
rect 45892 10780 46956 10836
rect 47012 10780 47022 10836
rect 24098 10668 24108 10724
rect 24164 10668 25340 10724
rect 25396 10668 25406 10724
rect 40898 10668 40908 10724
rect 40964 10668 41580 10724
rect 41636 10668 42924 10724
rect 42980 10668 42990 10724
rect 50082 10668 50092 10724
rect 50148 10668 50988 10724
rect 51044 10668 51054 10724
rect 5618 10556 5628 10612
rect 5684 10556 5964 10612
rect 6020 10556 6030 10612
rect 22866 10556 22876 10612
rect 22932 10556 23884 10612
rect 23940 10556 23950 10612
rect 28130 10556 28140 10612
rect 28196 10556 29372 10612
rect 29428 10556 29438 10612
rect 37314 10556 37324 10612
rect 37380 10556 37996 10612
rect 38052 10556 39340 10612
rect 39396 10556 40012 10612
rect 40068 10556 40078 10612
rect 5628 10444 5740 10500
rect 5796 10444 5806 10500
rect 22194 10444 22204 10500
rect 22260 10444 23772 10500
rect 23828 10444 23838 10500
rect 26674 10444 26684 10500
rect 26740 10444 27468 10500
rect 27524 10444 27534 10500
rect 30594 10444 30604 10500
rect 30660 10444 31724 10500
rect 31780 10444 32284 10500
rect 32340 10444 32350 10500
rect 45602 10444 45612 10500
rect 45668 10444 46732 10500
rect 46788 10444 46798 10500
rect 5628 10276 5684 10444
rect 21746 10332 21756 10388
rect 21812 10332 22652 10388
rect 22708 10332 22718 10388
rect 47394 10332 47404 10388
rect 47460 10332 48748 10388
rect 48804 10332 48814 10388
rect 5618 10220 5628 10276
rect 5684 10220 5694 10276
rect 54002 10220 54012 10276
rect 54068 10220 55244 10276
rect 55300 10220 55310 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 20290 10108 20300 10164
rect 20356 10108 22764 10164
rect 22820 10108 22830 10164
rect 22530 9996 22540 10052
rect 22596 9996 23436 10052
rect 23492 9996 26236 10052
rect 26292 9996 26302 10052
rect 26786 9996 26796 10052
rect 26852 9996 27804 10052
rect 27860 9996 27870 10052
rect 42578 9996 42588 10052
rect 42644 9996 43596 10052
rect 43652 9996 47740 10052
rect 47796 9996 47806 10052
rect 48850 9996 48860 10052
rect 48916 9996 50428 10052
rect 16706 9884 16716 9940
rect 16772 9884 19068 9940
rect 19124 9884 20748 9940
rect 20804 9884 20814 9940
rect 39106 9884 39116 9940
rect 39172 9884 42252 9940
rect 42308 9884 42318 9940
rect 50372 9828 50428 9996
rect 30034 9772 30044 9828
rect 30100 9772 30828 9828
rect 30884 9772 30894 9828
rect 37650 9772 37660 9828
rect 37716 9772 39228 9828
rect 39284 9772 39294 9828
rect 47954 9772 47964 9828
rect 48020 9772 49084 9828
rect 49140 9772 49150 9828
rect 50372 9772 50540 9828
rect 50596 9772 51324 9828
rect 51380 9772 51390 9828
rect 6178 9660 6188 9716
rect 6244 9660 6860 9716
rect 6916 9660 6926 9716
rect 10098 9660 10108 9716
rect 10164 9660 13580 9716
rect 13636 9660 17388 9716
rect 17444 9660 17454 9716
rect 29810 9660 29820 9716
rect 29876 9660 30716 9716
rect 30772 9660 30782 9716
rect 30930 9660 30940 9716
rect 30996 9660 33964 9716
rect 34020 9660 34030 9716
rect 39442 9660 39452 9716
rect 39508 9660 40236 9716
rect 40292 9660 41300 9716
rect 41458 9660 41468 9716
rect 41524 9660 44268 9716
rect 44324 9660 44334 9716
rect 30940 9604 30996 9660
rect 41244 9604 41300 9660
rect 19394 9548 19404 9604
rect 19460 9548 20076 9604
rect 20132 9548 20972 9604
rect 21028 9548 21868 9604
rect 21924 9548 21934 9604
rect 28130 9548 28140 9604
rect 28196 9548 29148 9604
rect 29204 9548 30996 9604
rect 38098 9548 38108 9604
rect 38164 9548 39340 9604
rect 39396 9548 39406 9604
rect 41234 9548 41244 9604
rect 41300 9548 41310 9604
rect 51650 9548 51660 9604
rect 51716 9548 52780 9604
rect 52836 9548 55132 9604
rect 55188 9548 55198 9604
rect 59200 9492 60000 9520
rect 27906 9436 27916 9492
rect 27972 9436 28588 9492
rect 28644 9436 28654 9492
rect 39106 9436 39116 9492
rect 39172 9436 40908 9492
rect 40964 9436 40974 9492
rect 49634 9436 49644 9492
rect 49700 9436 49980 9492
rect 50036 9436 50046 9492
rect 57586 9436 57596 9492
rect 57652 9436 58156 9492
rect 58212 9436 60000 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 59200 9408 60000 9436
rect 2930 9212 2940 9268
rect 2996 9212 6076 9268
rect 6132 9212 6142 9268
rect 10210 9212 10220 9268
rect 10276 9212 10668 9268
rect 10724 9212 15372 9268
rect 15428 9212 15438 9268
rect 30370 9212 30380 9268
rect 30436 9212 31388 9268
rect 31444 9212 31454 9268
rect 43362 9212 43372 9268
rect 43428 9212 57820 9268
rect 57876 9212 57886 9268
rect 7298 9100 7308 9156
rect 7364 9100 8764 9156
rect 8820 9100 9772 9156
rect 9828 9100 9838 9156
rect 15586 9100 15596 9156
rect 15652 9100 18172 9156
rect 18228 9100 18238 9156
rect 39554 9100 39564 9156
rect 39620 9100 40124 9156
rect 40180 9100 40190 9156
rect 43026 9100 43036 9156
rect 43092 9100 43708 9156
rect 43764 9100 43774 9156
rect 48066 9100 48076 9156
rect 48132 9100 49644 9156
rect 49700 9100 49710 9156
rect 50082 9100 50092 9156
rect 50148 9100 52892 9156
rect 52948 9100 52958 9156
rect 53554 9100 53564 9156
rect 53620 9100 55468 9156
rect 55524 9100 55534 9156
rect 6290 8988 6300 9044
rect 6356 8988 6636 9044
rect 6692 8988 8428 9044
rect 8484 8988 9212 9044
rect 9268 8988 9278 9044
rect 15138 8988 15148 9044
rect 15204 8988 15708 9044
rect 15764 8988 26908 9044
rect 44258 8988 44268 9044
rect 44324 8988 46172 9044
rect 46228 8988 46238 9044
rect 48178 8988 48188 9044
rect 48244 8988 48972 9044
rect 49028 8988 49038 9044
rect 50372 8988 51212 9044
rect 51268 8988 51278 9044
rect 54562 8988 54572 9044
rect 54628 8988 56588 9044
rect 56644 8988 56654 9044
rect 19394 8876 19404 8932
rect 19460 8876 20748 8932
rect 20804 8876 20814 8932
rect 19618 8764 19628 8820
rect 19684 8764 20636 8820
rect 20692 8764 20702 8820
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 18946 8428 18956 8484
rect 19012 8428 20076 8484
rect 20132 8428 20636 8484
rect 20692 8428 21308 8484
rect 21364 8428 21374 8484
rect 26852 8372 26908 8988
rect 33282 8876 33292 8932
rect 33348 8876 34300 8932
rect 34356 8876 34366 8932
rect 50372 8820 50428 8988
rect 40226 8764 40236 8820
rect 40292 8764 49980 8820
rect 50036 8764 50428 8820
rect 52322 8764 52332 8820
rect 52388 8764 54460 8820
rect 54516 8764 54526 8820
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 40338 8540 40348 8596
rect 40404 8540 41244 8596
rect 41300 8540 41310 8596
rect 54310 8540 54348 8596
rect 54404 8540 54414 8596
rect 47618 8428 47628 8484
rect 47684 8428 48748 8484
rect 48804 8428 48814 8484
rect 8642 8316 8652 8372
rect 8708 8316 10332 8372
rect 10388 8316 10398 8372
rect 26450 8316 26460 8372
rect 26516 8316 28812 8372
rect 28868 8316 28878 8372
rect 41346 8316 41356 8372
rect 41412 8316 42140 8372
rect 42196 8316 42206 8372
rect 54002 8316 54012 8372
rect 54068 8316 54348 8372
rect 54404 8316 54908 8372
rect 54964 8316 54974 8372
rect 24882 8204 24892 8260
rect 24948 8204 25788 8260
rect 25844 8204 25854 8260
rect 33954 8204 33964 8260
rect 34020 8204 34748 8260
rect 34804 8204 34814 8260
rect 51426 8204 51436 8260
rect 51492 8204 52892 8260
rect 52948 8204 52958 8260
rect 53106 8204 53116 8260
rect 53172 8204 53900 8260
rect 53956 8204 53966 8260
rect 7746 8092 7756 8148
rect 7812 8092 8988 8148
rect 9044 8092 9054 8148
rect 12674 8092 12684 8148
rect 12740 8092 25564 8148
rect 25620 8092 25630 8148
rect 54226 8092 54236 8148
rect 54292 8092 54908 8148
rect 54964 8092 54974 8148
rect 23202 7980 23212 8036
rect 23268 7980 24556 8036
rect 24612 7980 24622 8036
rect 29474 7980 29484 8036
rect 29540 7980 30268 8036
rect 30324 7980 30334 8036
rect 45714 7980 45724 8036
rect 45780 7980 47068 8036
rect 47124 7980 47628 8036
rect 47684 7980 47694 8036
rect 20188 7868 20412 7924
rect 20468 7868 20478 7924
rect 30034 7868 30044 7924
rect 30100 7868 30604 7924
rect 30660 7868 34972 7924
rect 35028 7868 35038 7924
rect 46274 7868 46284 7924
rect 46340 7868 47292 7924
rect 47348 7868 49644 7924
rect 49700 7868 49710 7924
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 20188 7700 20244 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 37314 7756 37324 7812
rect 37380 7756 42252 7812
rect 42308 7756 42318 7812
rect 20066 7644 20076 7700
rect 20132 7644 20244 7700
rect 39218 7644 39228 7700
rect 39284 7644 39900 7700
rect 39956 7644 39966 7700
rect 50978 7644 50988 7700
rect 51044 7644 53340 7700
rect 53396 7644 53406 7700
rect 53106 7532 53116 7588
rect 53172 7532 54348 7588
rect 54404 7532 54414 7588
rect 5954 7420 5964 7476
rect 6020 7420 7756 7476
rect 7812 7420 7822 7476
rect 24770 7420 24780 7476
rect 24836 7420 26236 7476
rect 26292 7420 26302 7476
rect 30818 7420 30828 7476
rect 30884 7420 31612 7476
rect 31668 7420 31678 7476
rect 39666 7420 39676 7476
rect 39732 7420 40908 7476
rect 40964 7420 40974 7476
rect 41570 7420 41580 7476
rect 41636 7420 44156 7476
rect 44212 7420 45948 7476
rect 46004 7420 46014 7476
rect 55346 7420 55356 7476
rect 55412 7420 56588 7476
rect 56644 7420 56654 7476
rect 18498 7308 18508 7364
rect 18564 7308 19068 7364
rect 19124 7308 24668 7364
rect 24724 7308 27132 7364
rect 27188 7308 27198 7364
rect 29698 7308 29708 7364
rect 29764 7308 30380 7364
rect 30436 7308 30446 7364
rect 31154 7308 31164 7364
rect 31220 7308 33852 7364
rect 33908 7308 33918 7364
rect 31164 7252 31220 7308
rect 26226 7196 26236 7252
rect 26292 7196 26908 7252
rect 29810 7196 29820 7252
rect 29876 7196 31220 7252
rect 38210 7196 38220 7252
rect 38276 7196 39116 7252
rect 39172 7196 39182 7252
rect 54338 7196 54348 7252
rect 54404 7196 54796 7252
rect 54852 7196 54862 7252
rect 26852 7140 26908 7196
rect 26852 7084 33796 7140
rect 52210 7084 52220 7140
rect 52276 7084 54124 7140
rect 54180 7084 54190 7140
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 33740 7028 33796 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 26674 6972 26684 7028
rect 26740 6972 27356 7028
rect 27412 6972 30716 7028
rect 30772 6972 31836 7028
rect 31892 6972 31902 7028
rect 33730 6972 33740 7028
rect 33796 6972 33806 7028
rect 42242 6972 42252 7028
rect 42308 6972 43484 7028
rect 43540 6972 52332 7028
rect 52388 6972 52780 7028
rect 52836 6972 53564 7028
rect 53620 6972 53630 7028
rect 26450 6860 26460 6916
rect 26516 6860 27580 6916
rect 27636 6860 35308 6916
rect 35364 6860 35980 6916
rect 36036 6860 36046 6916
rect 43698 6860 43708 6916
rect 43764 6860 48972 6916
rect 49028 6860 49038 6916
rect 49634 6860 49644 6916
rect 49700 6860 50092 6916
rect 50148 6860 52668 6916
rect 52724 6860 53116 6916
rect 53172 6860 53182 6916
rect 53330 6860 53340 6916
rect 53396 6860 54236 6916
rect 54292 6860 54302 6916
rect 21970 6748 21980 6804
rect 22036 6748 22876 6804
rect 22932 6748 22942 6804
rect 34626 6748 34636 6804
rect 34692 6748 34702 6804
rect 42242 6748 42252 6804
rect 42308 6748 43148 6804
rect 43204 6748 45612 6804
rect 45668 6748 46228 6804
rect 49298 6748 49308 6804
rect 49364 6748 50204 6804
rect 50260 6748 50764 6804
rect 50820 6748 50830 6804
rect 52882 6748 52892 6804
rect 52948 6748 55244 6804
rect 55300 6748 55310 6804
rect 34636 6692 34692 6748
rect 46172 6692 46228 6748
rect 8866 6636 8876 6692
rect 8932 6636 11228 6692
rect 11284 6636 11294 6692
rect 17378 6636 17388 6692
rect 17444 6636 19516 6692
rect 19572 6636 19582 6692
rect 19954 6636 19964 6692
rect 20020 6636 22988 6692
rect 23044 6636 24108 6692
rect 24164 6636 24174 6692
rect 33506 6636 33516 6692
rect 33572 6636 34692 6692
rect 41122 6636 41132 6692
rect 41188 6636 42700 6692
rect 42756 6636 42766 6692
rect 44370 6636 44380 6692
rect 44436 6636 45052 6692
rect 45108 6636 45500 6692
rect 45556 6636 45566 6692
rect 46162 6636 46172 6692
rect 46228 6636 47180 6692
rect 47236 6636 52108 6692
rect 52164 6636 52174 6692
rect 56018 6636 56028 6692
rect 56084 6636 58044 6692
rect 58100 6636 58110 6692
rect 14242 6524 14252 6580
rect 14308 6524 16268 6580
rect 16324 6524 16334 6580
rect 22754 6524 22764 6580
rect 22820 6524 23548 6580
rect 23604 6524 23884 6580
rect 23940 6524 25228 6580
rect 25284 6524 25294 6580
rect 40226 6524 40236 6580
rect 40292 6524 45388 6580
rect 45444 6524 45454 6580
rect 46050 6524 46060 6580
rect 46116 6524 46956 6580
rect 47012 6524 47022 6580
rect 47394 6524 47404 6580
rect 47460 6524 51100 6580
rect 51156 6524 51166 6580
rect 16370 6412 16380 6468
rect 16436 6412 16940 6468
rect 16996 6412 17006 6468
rect 21746 6412 21756 6468
rect 21812 6412 24780 6468
rect 24836 6412 24846 6468
rect 44034 6412 44044 6468
rect 44100 6412 44828 6468
rect 44884 6412 45612 6468
rect 45668 6412 46620 6468
rect 46676 6412 46686 6468
rect 16818 6300 16828 6356
rect 16884 6300 17948 6356
rect 18004 6300 19292 6356
rect 19348 6300 19358 6356
rect 34626 6300 34636 6356
rect 34692 6300 34972 6356
rect 35028 6300 35196 6356
rect 35252 6300 35262 6356
rect 45378 6300 45388 6356
rect 45444 6300 46396 6356
rect 46452 6300 46462 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 36306 6188 36316 6244
rect 36372 6188 37212 6244
rect 37268 6188 37278 6244
rect 16818 6076 16828 6132
rect 16884 6076 19068 6132
rect 19124 6076 19134 6132
rect 19282 6076 19292 6132
rect 19348 6076 21308 6132
rect 21364 6076 21374 6132
rect 45490 6076 45500 6132
rect 45556 6076 49644 6132
rect 49700 6076 50092 6132
rect 50148 6076 50158 6132
rect 7858 5964 7868 6020
rect 7924 5964 8540 6020
rect 8596 5964 25116 6020
rect 25172 5964 25788 6020
rect 25844 5964 26236 6020
rect 26292 5964 26302 6020
rect 46946 5964 46956 6020
rect 47012 5964 47852 6020
rect 47908 5964 47918 6020
rect 14914 5852 14924 5908
rect 14980 5852 15708 5908
rect 15764 5852 16828 5908
rect 16884 5852 16894 5908
rect 24434 5852 24444 5908
rect 24500 5852 25452 5908
rect 25508 5852 25518 5908
rect 37538 5852 37548 5908
rect 37604 5852 38556 5908
rect 38612 5852 41132 5908
rect 41188 5852 41198 5908
rect 47394 5852 47404 5908
rect 47460 5852 49980 5908
rect 50036 5852 50316 5908
rect 50372 5852 50382 5908
rect 16258 5740 16268 5796
rect 16324 5740 17724 5796
rect 17780 5740 17790 5796
rect 46610 5740 46620 5796
rect 46676 5740 47964 5796
rect 48020 5740 49084 5796
rect 49140 5740 49150 5796
rect 25778 5628 25788 5684
rect 25844 5628 26684 5684
rect 26740 5628 26750 5684
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 16034 5292 16044 5348
rect 16100 5292 19404 5348
rect 19460 5292 22764 5348
rect 22820 5292 22830 5348
rect 14578 5180 14588 5236
rect 14644 5180 15932 5236
rect 15988 5180 15998 5236
rect 17602 5180 17612 5236
rect 17668 5180 18452 5236
rect 22866 5180 22876 5236
rect 22932 5180 24108 5236
rect 24164 5180 24174 5236
rect 41010 5180 41020 5236
rect 41076 5180 42700 5236
rect 42756 5180 42766 5236
rect 50372 5180 53452 5236
rect 53508 5180 54684 5236
rect 54740 5180 54750 5236
rect 18396 5124 18452 5180
rect 50372 5124 50428 5180
rect 16706 5068 16716 5124
rect 16772 5068 17836 5124
rect 17892 5068 18172 5124
rect 18228 5068 18238 5124
rect 18386 5068 18396 5124
rect 18452 5068 19740 5124
rect 19796 5068 20412 5124
rect 20468 5068 20478 5124
rect 20738 5068 20748 5124
rect 20804 5068 21644 5124
rect 21700 5068 23772 5124
rect 23828 5068 26572 5124
rect 26628 5068 26638 5124
rect 29698 5068 29708 5124
rect 29764 5068 30380 5124
rect 30436 5068 30446 5124
rect 41122 5068 41132 5124
rect 41188 5068 43596 5124
rect 43652 5068 43662 5124
rect 49298 5068 49308 5124
rect 49364 5068 50428 5124
rect 24210 4956 24220 5012
rect 24276 4956 25228 5012
rect 25284 4956 29260 5012
rect 29316 4956 29326 5012
rect 34514 4956 34524 5012
rect 34580 4956 39228 5012
rect 39284 4956 39294 5012
rect 44930 4956 44940 5012
rect 44996 4956 46508 5012
rect 46564 4956 46574 5012
rect 9538 4844 9548 4900
rect 9604 4844 10892 4900
rect 10948 4844 10958 4900
rect 17826 4844 17836 4900
rect 17892 4844 18620 4900
rect 18676 4844 21420 4900
rect 21476 4844 21486 4900
rect 21858 4844 21868 4900
rect 21924 4844 24332 4900
rect 24388 4844 24398 4900
rect 46050 4844 46060 4900
rect 46116 4844 47404 4900
rect 47460 4844 47470 4900
rect 51314 4844 51324 4900
rect 51380 4844 52668 4900
rect 52724 4844 52734 4900
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 33282 4508 33292 4564
rect 33348 4508 34412 4564
rect 34468 4508 34478 4564
rect 32162 4396 32172 4452
rect 32228 4396 33180 4452
rect 33236 4396 33246 4452
rect 39554 4396 39564 4452
rect 39620 4396 57820 4452
rect 57876 4396 57886 4452
rect 10210 4284 10220 4340
rect 10276 4284 11228 4340
rect 11284 4284 13356 4340
rect 13412 4284 13422 4340
rect 13010 4172 13020 4228
rect 13076 4172 23100 4228
rect 23156 4172 23166 4228
rect 26898 4172 26908 4228
rect 26964 4172 28140 4228
rect 28196 4172 28206 4228
rect 20290 4060 20300 4116
rect 20356 4060 25228 4116
rect 25284 4060 25294 4116
rect 43026 4060 43036 4116
rect 43092 4060 45388 4116
rect 45444 4060 45454 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 25666 3724 25676 3780
rect 25732 3724 43148 3780
rect 43204 3724 44492 3780
rect 44548 3724 44558 3780
rect 59200 3668 60000 3696
rect 20850 3612 20860 3668
rect 20916 3612 22092 3668
rect 22148 3612 22158 3668
rect 24882 3612 24892 3668
rect 24948 3612 26124 3668
rect 26180 3612 26190 3668
rect 28578 3612 28588 3668
rect 28644 3612 38668 3668
rect 38882 3612 38892 3668
rect 38948 3612 40796 3668
rect 40852 3612 40862 3668
rect 43474 3612 43484 3668
rect 43540 3612 44380 3668
rect 44436 3612 44446 3668
rect 58146 3612 58156 3668
rect 58212 3612 60000 3668
rect 38612 3556 38668 3612
rect 59200 3584 60000 3612
rect 12786 3500 12796 3556
rect 12852 3500 21084 3556
rect 21140 3500 21150 3556
rect 28130 3500 28140 3556
rect 28196 3500 36652 3556
rect 36708 3500 36718 3556
rect 38612 3500 47404 3556
rect 47460 3500 48860 3556
rect 48916 3500 48926 3556
rect 45042 3388 45052 3444
rect 45108 3388 48972 3444
rect 49028 3388 49038 3444
rect 4722 3276 4732 3332
rect 4788 3276 5516 3332
rect 5572 3276 5582 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
<< via3 >>
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 23100 55916 23156 55972
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 26348 50540 26404 50596
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 26348 49532 26404 49588
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 23100 47292 23156 47348
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 34636 44492 34692 44548
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 43484 42140 43540 42196
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 29036 41020 29092 41076
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 34636 37772 34692 37828
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 43484 36652 43540 36708
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 29036 35868 29092 35924
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 52108 33516 52164 33572
rect 34188 32956 34244 33012
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 34524 32844 34580 32900
rect 52332 32396 52388 32452
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 34188 29820 34244 29876
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 8652 29372 8708 29428
rect 34524 29260 34580 29316
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 8652 28476 8708 28532
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 54124 27692 54180 27748
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 50988 26796 51044 26852
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 54124 26236 54180 26292
rect 52108 26124 52164 26180
rect 52332 26012 52388 26068
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 50988 25452 51044 25508
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 8652 24108 8708 24164
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 38444 19180 38500 19236
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 38444 18284 38500 18340
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 31836 17836 31892 17892
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 54460 16940 54516 16996
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 54460 12460 54516 12516
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 31836 11116 31892 11172
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 54348 8540 54404 8596
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 54348 7196 54404 7252
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
<< metal4 >>
rect 4448 55692 4768 56508
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 19808 56476 20128 56508
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 23100 55972 23156 55982
rect 23100 47348 23156 55916
rect 35168 55692 35488 56508
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 26348 50596 26404 50606
rect 26348 49588 26404 50540
rect 26348 49522 26404 49532
rect 23100 47282 23156 47292
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 34636 44548 34692 44558
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 29036 41076 29092 41086
rect 29036 35924 29092 41020
rect 34636 37828 34692 44492
rect 34636 37762 34692 37772
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 50528 56476 50848 56508
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 29036 35858 29092 35868
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 35168 35308 35488 36820
rect 43484 42196 43540 42206
rect 43484 36708 43540 42140
rect 43484 36642 43540 36652
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 34188 33012 34244 33022
rect 34188 29876 34244 32956
rect 34188 29810 34244 29820
rect 34524 32900 34580 32910
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 8652 29428 8708 29438
rect 8652 28532 8708 29372
rect 8652 24164 8708 28476
rect 8652 24098 8708 24108
rect 19808 28252 20128 29764
rect 34524 29316 34580 32844
rect 34524 29250 34580 29260
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 52108 33572 52164 33582
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50988 26852 51044 26862
rect 50988 25508 51044 26796
rect 52108 26180 52164 33516
rect 52108 26114 52164 26124
rect 52332 32452 52388 32462
rect 52332 26068 52388 32396
rect 54124 27748 54180 27758
rect 54124 26292 54180 27692
rect 54124 26226 54180 26236
rect 52332 26002 52388 26012
rect 50988 25442 51044 25452
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 38444 19236 38500 19246
rect 38444 18340 38500 19180
rect 38444 18274 38500 18284
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 31836 17892 31892 17902
rect 31836 11172 31892 17836
rect 31836 11106 31892 11116
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 54460 16996 54516 17006
rect 54460 12516 54516 16940
rect 54460 12450 54516 12460
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 54348 8596 54404 8606
rect 54348 7252 54404 8540
rect 54348 7186 54404 7196
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _1024_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15008 0 -1 42336
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1025_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23744 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1026_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 35056 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1027_
timestamp 1698431365
transform 1 0 30128 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1028_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31248 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1029_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30128 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1030_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30128 0 1 26656
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1031_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24416 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1032_
timestamp 1698431365
transform 1 0 22288 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1033_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 25312 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1034_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 25088 0 1 28224
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1035_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20720 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1036_
timestamp 1698431365
transform 1 0 23744 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1037_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22736 0 -1 26656
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1038_
timestamp 1698431365
transform 1 0 22288 0 1 26656
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1039_
timestamp 1698431365
transform -1 0 23520 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1040_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22176 0 -1 23520
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1041_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 24640 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1042_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22176 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1043_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22288 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1044_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22400 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1045_
timestamp 1698431365
transform -1 0 22848 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1046_
timestamp 1698431365
transform 1 0 27552 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1047_
timestamp 1698431365
transform -1 0 37632 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1048_
timestamp 1698431365
transform -1 0 38304 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1049_
timestamp 1698431365
transform -1 0 39200 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1050_
timestamp 1698431365
transform 1 0 37856 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1051_
timestamp 1698431365
transform 1 0 33040 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1052_
timestamp 1698431365
transform 1 0 33936 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1053_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 36848 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1054_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34608 0 1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1055_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36288 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1056_
timestamp 1698431365
transform 1 0 37520 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1057_
timestamp 1698431365
transform -1 0 27440 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1058_
timestamp 1698431365
transform 1 0 26656 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1059_
timestamp 1698431365
transform -1 0 37856 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1060_
timestamp 1698431365
transform -1 0 37520 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1061_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37408 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1062_
timestamp 1698431365
transform -1 0 36400 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1063_
timestamp 1698431365
transform -1 0 42112 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1064_
timestamp 1698431365
transform 1 0 37856 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1065_
timestamp 1698431365
transform 1 0 38416 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1066_
timestamp 1698431365
transform -1 0 42448 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1067_
timestamp 1698431365
transform 1 0 37744 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1068_
timestamp 1698431365
transform 1 0 38304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1069_
timestamp 1698431365
transform 1 0 42224 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1070_
timestamp 1698431365
transform 1 0 35616 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1071_
timestamp 1698431365
transform -1 0 37296 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1072_
timestamp 1698431365
transform -1 0 57904 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1073_
timestamp 1698431365
transform 1 0 35056 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1074_
timestamp 1698431365
transform 1 0 36176 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1075_
timestamp 1698431365
transform -1 0 34832 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1076_
timestamp 1698431365
transform -1 0 33936 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1077_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33936 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1078_
timestamp 1698431365
transform -1 0 35392 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1079_
timestamp 1698431365
transform 1 0 37184 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1080_
timestamp 1698431365
transform 1 0 38192 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1081_
timestamp 1698431365
transform -1 0 26656 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1082_
timestamp 1698431365
transform 1 0 26432 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1083_
timestamp 1698431365
transform 1 0 38640 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1084_
timestamp 1698431365
transform -1 0 39872 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1085_
timestamp 1698431365
transform -1 0 38304 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1086_
timestamp 1698431365
transform -1 0 41664 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1087_
timestamp 1698431365
transform 1 0 41104 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1088_
timestamp 1698431365
transform -1 0 41776 0 -1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1089_
timestamp 1698431365
transform -1 0 42896 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1090_
timestamp 1698431365
transform -1 0 40432 0 -1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1091_
timestamp 1698431365
transform -1 0 39424 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1092_
timestamp 1698431365
transform -1 0 36848 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1093_
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1094_
timestamp 1698431365
transform -1 0 39760 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1095_
timestamp 1698431365
transform -1 0 28784 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1096_
timestamp 1698431365
transform -1 0 28224 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1097_
timestamp 1698431365
transform 1 0 27440 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1098_
timestamp 1698431365
transform 1 0 37184 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1099_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28224 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1100_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27328 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1101_
timestamp 1698431365
transform 1 0 25872 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1102_
timestamp 1698431365
transform 1 0 27216 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1103_
timestamp 1698431365
transform 1 0 27328 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1104_
timestamp 1698431365
transform -1 0 29456 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1105_
timestamp 1698431365
transform -1 0 45584 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1106_
timestamp 1698431365
transform 1 0 29568 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1107_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29904 0 -1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1108_
timestamp 1698431365
transform -1 0 23520 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1109_
timestamp 1698431365
transform -1 0 15008 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1110_
timestamp 1698431365
transform 1 0 14000 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1111_
timestamp 1698431365
transform 1 0 22736 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1112_
timestamp 1698431365
transform -1 0 44128 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1113_
timestamp 1698431365
transform -1 0 29232 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1114_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23296 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1115_
timestamp 1698431365
transform 1 0 22848 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1116_
timestamp 1698431365
transform -1 0 46592 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1117_
timestamp 1698431365
transform -1 0 29568 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1118_
timestamp 1698431365
transform 1 0 23408 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1119_
timestamp 1698431365
transform 1 0 26992 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1120_
timestamp 1698431365
transform 1 0 26544 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1121_
timestamp 1698431365
transform -1 0 24864 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1122_
timestamp 1698431365
transform -1 0 25536 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1123_
timestamp 1698431365
transform 1 0 23408 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1124_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22848 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1125_
timestamp 1698431365
transform 1 0 23968 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1126_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24640 0 -1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1127_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23408 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1128_
timestamp 1698431365
transform -1 0 24304 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1129_
timestamp 1698431365
transform 1 0 23968 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1130_
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1131_
timestamp 1698431365
transform -1 0 15568 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1132_
timestamp 1698431365
transform 1 0 15568 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1133_
timestamp 1698431365
transform -1 0 23968 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1134_
timestamp 1698431365
transform 1 0 22512 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1135_
timestamp 1698431365
transform 1 0 24528 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1136_
timestamp 1698431365
transform -1 0 21616 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1137_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24528 0 1 14112
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1138_
timestamp 1698431365
transform -1 0 16912 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1139_
timestamp 1698431365
transform 1 0 17248 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1140_
timestamp 1698431365
transform -1 0 20944 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1141_
timestamp 1698431365
transform 1 0 13440 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1142_
timestamp 1698431365
transform -1 0 14000 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1143_
timestamp 1698431365
transform -1 0 14224 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1144_
timestamp 1698431365
transform 1 0 13104 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1145_
timestamp 1698431365
transform -1 0 17808 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1146_
timestamp 1698431365
transform -1 0 16352 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1147_
timestamp 1698431365
transform -1 0 14784 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1148_
timestamp 1698431365
transform 1 0 15344 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1149_
timestamp 1698431365
transform 1 0 16016 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1150_
timestamp 1698431365
transform -1 0 15456 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1151_
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1152_
timestamp 1698431365
transform 1 0 12096 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1153_
timestamp 1698431365
transform 1 0 11424 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1154_
timestamp 1698431365
transform -1 0 14784 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1155_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 14672 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1156_
timestamp 1698431365
transform -1 0 13104 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1157_
timestamp 1698431365
transform -1 0 24640 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1158_
timestamp 1698431365
transform -1 0 15344 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1159_
timestamp 1698431365
transform 1 0 13888 0 -1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1160_
timestamp 1698431365
transform 1 0 15120 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1161_
timestamp 1698431365
transform 1 0 34496 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1162_
timestamp 1698431365
transform 1 0 34832 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1163_
timestamp 1698431365
transform 1 0 33040 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1164_
timestamp 1698431365
transform -1 0 34832 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1165_
timestamp 1698431365
transform -1 0 26656 0 -1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1166_
timestamp 1698431365
transform -1 0 26096 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1167_
timestamp 1698431365
transform 1 0 26320 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1168_
timestamp 1698431365
transform -1 0 25088 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1169_
timestamp 1698431365
transform -1 0 34496 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1170_
timestamp 1698431365
transform -1 0 28336 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1171_
timestamp 1698431365
transform -1 0 32032 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1172_
timestamp 1698431365
transform 1 0 26656 0 -1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1173_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26096 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1174_
timestamp 1698431365
transform 1 0 19824 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1175_
timestamp 1698431365
transform -1 0 19600 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1176_
timestamp 1698431365
transform 1 0 18928 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1177_
timestamp 1698431365
transform 1 0 26320 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1178_
timestamp 1698431365
transform -1 0 24080 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1179_
timestamp 1698431365
transform -1 0 24304 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1180_
timestamp 1698431365
transform -1 0 22400 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1181_
timestamp 1698431365
transform -1 0 23296 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1182_
timestamp 1698431365
transform -1 0 20496 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1183_
timestamp 1698431365
transform 1 0 22400 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1184_
timestamp 1698431365
transform -1 0 22176 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1185_
timestamp 1698431365
transform -1 0 21840 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1186_
timestamp 1698431365
transform -1 0 20944 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1187_
timestamp 1698431365
transform -1 0 20160 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1188_
timestamp 1698431365
transform 1 0 20496 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1189_
timestamp 1698431365
transform -1 0 17024 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1190_
timestamp 1698431365
transform -1 0 17584 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1191_
timestamp 1698431365
transform -1 0 16576 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1192_
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1193_
timestamp 1698431365
transform -1 0 16464 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1194_
timestamp 1698431365
transform 1 0 18032 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1195_
timestamp 1698431365
transform 1 0 19040 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1196_
timestamp 1698431365
transform 1 0 21280 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1197_
timestamp 1698431365
transform 1 0 22288 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1198_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22624 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1199_
timestamp 1698431365
transform -1 0 24416 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1200_
timestamp 1698431365
transform -1 0 20048 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1201_
timestamp 1698431365
transform -1 0 14224 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1202_
timestamp 1698431365
transform 1 0 13888 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1203_
timestamp 1698431365
transform -1 0 12880 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1204_
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1205_
timestamp 1698431365
transform -1 0 6832 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1206_
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1207_
timestamp 1698431365
transform -1 0 5264 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1208_
timestamp 1698431365
transform 1 0 7616 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1209_
timestamp 1698431365
transform -1 0 7952 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1210_
timestamp 1698431365
transform -1 0 7056 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1211_
timestamp 1698431365
transform -1 0 6832 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1212_
timestamp 1698431365
transform 1 0 7392 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1213_
timestamp 1698431365
transform 1 0 6720 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1214_
timestamp 1698431365
transform 1 0 7952 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1215_
timestamp 1698431365
transform 1 0 7616 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1216_
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1217_
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1218_
timestamp 1698431365
transform 1 0 8176 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1219_
timestamp 1698431365
transform -1 0 10528 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1220_
timestamp 1698431365
transform 1 0 9072 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1221_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 35840 0 -1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1222_
timestamp 1698431365
transform 1 0 38416 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1223_
timestamp 1698431365
transform -1 0 42784 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1224_
timestamp 1698431365
transform 1 0 27552 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1225_
timestamp 1698431365
transform -1 0 42560 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1226_
timestamp 1698431365
transform -1 0 43232 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1227_
timestamp 1698431365
transform -1 0 41776 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1228_
timestamp 1698431365
transform 1 0 39872 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1229_
timestamp 1698431365
transform -1 0 42112 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1230_
timestamp 1698431365
transform 1 0 40320 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1231_
timestamp 1698431365
transform -1 0 42672 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1232_
timestamp 1698431365
transform 1 0 42672 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1233_
timestamp 1698431365
transform 1 0 41776 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1234_
timestamp 1698431365
transform 1 0 42448 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1235_
timestamp 1698431365
transform 1 0 48608 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1236_
timestamp 1698431365
transform 1 0 47824 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1237_
timestamp 1698431365
transform 1 0 49168 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1238_
timestamp 1698431365
transform 1 0 50176 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1239_
timestamp 1698431365
transform 1 0 52528 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1240_
timestamp 1698431365
transform -1 0 53536 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1241_
timestamp 1698431365
transform -1 0 52304 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1242_
timestamp 1698431365
transform -1 0 55664 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1243_
timestamp 1698431365
transform 1 0 54096 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1244_
timestamp 1698431365
transform 1 0 55216 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1245_
timestamp 1698431365
transform -1 0 55104 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1246_
timestamp 1698431365
transform 1 0 54208 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1247_
timestamp 1698431365
transform 1 0 55328 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1248_
timestamp 1698431365
transform 1 0 35616 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1249_
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1250_
timestamp 1698431365
transform 1 0 38080 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1251_
timestamp 1698431365
transform 1 0 37632 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1252_
timestamp 1698431365
transform -1 0 40544 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1253_
timestamp 1698431365
transform -1 0 39872 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1254_
timestamp 1698431365
transform -1 0 41664 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1255_
timestamp 1698431365
transform -1 0 42112 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1256_
timestamp 1698431365
transform -1 0 41776 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1257_
timestamp 1698431365
transform 1 0 41776 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1258_
timestamp 1698431365
transform -1 0 39536 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1259_
timestamp 1698431365
transform -1 0 38752 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1260_
timestamp 1698431365
transform 1 0 38080 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1261_
timestamp 1698431365
transform 1 0 37408 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1262_
timestamp 1698431365
transform 1 0 41328 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1263_
timestamp 1698431365
transform 1 0 41104 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1264_
timestamp 1698431365
transform -1 0 42336 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1265_
timestamp 1698431365
transform -1 0 42784 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1266_
timestamp 1698431365
transform 1 0 43008 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1267_
timestamp 1698431365
transform -1 0 42336 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1268_
timestamp 1698431365
transform -1 0 43008 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1269_
timestamp 1698431365
transform -1 0 41104 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1270_
timestamp 1698431365
transform -1 0 43232 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1271_
timestamp 1698431365
transform 1 0 40992 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1272_
timestamp 1698431365
transform -1 0 39648 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1273_
timestamp 1698431365
transform -1 0 42784 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1274_
timestamp 1698431365
transform -1 0 42672 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1275_
timestamp 1698431365
transform 1 0 41216 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1276_
timestamp 1698431365
transform 1 0 46704 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1277_
timestamp 1698431365
transform 1 0 47376 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1278_
timestamp 1698431365
transform -1 0 50400 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1279_
timestamp 1698431365
transform -1 0 49952 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1280_
timestamp 1698431365
transform -1 0 53536 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1281_
timestamp 1698431365
transform -1 0 52304 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1282_
timestamp 1698431365
transform -1 0 55328 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1283_
timestamp 1698431365
transform 1 0 55328 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1284_
timestamp 1698431365
transform 1 0 53648 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1285_
timestamp 1698431365
transform -1 0 56896 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1286_
timestamp 1698431365
transform -1 0 30912 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1287_
timestamp 1698431365
transform 1 0 29008 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1288_
timestamp 1698431365
transform 1 0 30128 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1289_
timestamp 1698431365
transform -1 0 30240 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1290_
timestamp 1698431365
transform 1 0 24864 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1291_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30464 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1292_
timestamp 1698431365
transform -1 0 30464 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1293_
timestamp 1698431365
transform 1 0 30128 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1294_
timestamp 1698431365
transform -1 0 32144 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1295_
timestamp 1698431365
transform -1 0 30128 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1296_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33040 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1297_
timestamp 1698431365
transform 1 0 34832 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1298_
timestamp 1698431365
transform 1 0 33712 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1299_
timestamp 1698431365
transform 1 0 34608 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1300_
timestamp 1698431365
transform -1 0 4368 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1301_
timestamp 1698431365
transform 1 0 3696 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1302_
timestamp 1698431365
transform -1 0 3696 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1303_
timestamp 1698431365
transform -1 0 4032 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1304_
timestamp 1698431365
transform 1 0 3360 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1305_
timestamp 1698431365
transform -1 0 3360 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1306_
timestamp 1698431365
transform -1 0 4256 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1307_
timestamp 1698431365
transform 1 0 6832 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1308_
timestamp 1698431365
transform 1 0 3472 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1309_
timestamp 1698431365
transform -1 0 3472 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1310_
timestamp 1698431365
transform -1 0 4928 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1311_
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1312_
timestamp 1698431365
transform -1 0 4704 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1313_
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1314_
timestamp 1698431365
transform -1 0 7168 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1315_
timestamp 1698431365
transform 1 0 5376 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1316_
timestamp 1698431365
transform 1 0 5824 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1317_
timestamp 1698431365
transform 1 0 14896 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1318_
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1319_
timestamp 1698431365
transform 1 0 8288 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1320_
timestamp 1698431365
transform 1 0 24528 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1321_
timestamp 1698431365
transform 1 0 7056 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1322_
timestamp 1698431365
transform 1 0 7056 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1323_
timestamp 1698431365
transform -1 0 8288 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1324_
timestamp 1698431365
transform 1 0 8512 0 1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1325_
timestamp 1698431365
transform 1 0 9856 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1326_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 38864 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1327_
timestamp 1698431365
transform -1 0 38752 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1328_
timestamp 1698431365
transform -1 0 29568 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1329_
timestamp 1698431365
transform -1 0 27552 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1330_
timestamp 1698431365
transform 1 0 26320 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1331_
timestamp 1698431365
transform 1 0 26768 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1332_
timestamp 1698431365
transform 1 0 43344 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1333_
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1334_
timestamp 1698431365
transform 1 0 25872 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1335_
timestamp 1698431365
transform -1 0 29792 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1336_
timestamp 1698431365
transform -1 0 28000 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1337_
timestamp 1698431365
transform -1 0 29680 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1338_
timestamp 1698431365
transform -1 0 27440 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1339_
timestamp 1698431365
transform 1 0 23856 0 -1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1340_
timestamp 1698431365
transform -1 0 22624 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1341_
timestamp 1698431365
transform 1 0 23520 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1342_
timestamp 1698431365
transform -1 0 22288 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1343_
timestamp 1698431365
transform -1 0 26656 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1344_
timestamp 1698431365
transform -1 0 25872 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1345_
timestamp 1698431365
transform -1 0 26544 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1346_
timestamp 1698431365
transform 1 0 24640 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1347_
timestamp 1698431365
transform 1 0 30016 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1348_
timestamp 1698431365
transform 1 0 29456 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1349_
timestamp 1698431365
transform 1 0 31696 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1350_
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1351_
timestamp 1698431365
transform 1 0 30464 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1352_
timestamp 1698431365
transform -1 0 29456 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1353_
timestamp 1698431365
transform 1 0 31696 0 -1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1354_
timestamp 1698431365
transform 1 0 32928 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1355_
timestamp 1698431365
transform 1 0 30128 0 1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1356_
timestamp 1698431365
transform -1 0 30352 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1357_
timestamp 1698431365
transform 1 0 26544 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1358_
timestamp 1698431365
transform 1 0 28112 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1359_
timestamp 1698431365
transform 1 0 35840 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1360_
timestamp 1698431365
transform 1 0 24192 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1361_
timestamp 1698431365
transform 1 0 26432 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1362_
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1363_
timestamp 1698431365
transform -1 0 34832 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1364_
timestamp 1698431365
transform -1 0 9184 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1365_
timestamp 1698431365
transform -1 0 8176 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1366_
timestamp 1698431365
transform -1 0 36736 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1367_
timestamp 1698431365
transform -1 0 31360 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1368_
timestamp 1698431365
transform -1 0 34048 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1369_
timestamp 1698431365
transform -1 0 31248 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1370_
timestamp 1698431365
transform -1 0 24864 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1371_
timestamp 1698431365
transform -1 0 23856 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1372_
timestamp 1698431365
transform 1 0 21840 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1373_
timestamp 1698431365
transform -1 0 20608 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1374_
timestamp 1698431365
transform 1 0 30576 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1375_
timestamp 1698431365
transform -1 0 29456 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1376_
timestamp 1698431365
transform 1 0 21952 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1377_
timestamp 1698431365
transform -1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1378_
timestamp 1698431365
transform 1 0 34160 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1379_
timestamp 1698431365
transform -1 0 36512 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1380_
timestamp 1698431365
transform -1 0 32368 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1381_
timestamp 1698431365
transform 1 0 30016 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1382_
timestamp 1698431365
transform 1 0 39312 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1383_
timestamp 1698431365
transform -1 0 47152 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1384_
timestamp 1698431365
transform 1 0 48944 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1385_
timestamp 1698431365
transform 1 0 48608 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1386_
timestamp 1698431365
transform 1 0 45584 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1387_
timestamp 1698431365
transform 1 0 48944 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1388_
timestamp 1698431365
transform 1 0 43792 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1389_
timestamp 1698431365
transform 1 0 45024 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1390_
timestamp 1698431365
transform 1 0 46032 0 1 42336
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1391_
timestamp 1698431365
transform -1 0 47824 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1392_
timestamp 1698431365
transform 1 0 44688 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1393_
timestamp 1698431365
transform 1 0 45360 0 -1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1394_
timestamp 1698431365
transform -1 0 53536 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1395_
timestamp 1698431365
transform 1 0 49280 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1396_
timestamp 1698431365
transform 1 0 47824 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1397_
timestamp 1698431365
transform 1 0 48944 0 1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1398_
timestamp 1698431365
transform 1 0 48608 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1399_
timestamp 1698431365
transform 1 0 47488 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1400_
timestamp 1698431365
transform 1 0 51632 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1401_
timestamp 1698431365
transform -1 0 54768 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1402_
timestamp 1698431365
transform 1 0 51408 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1403_
timestamp 1698431365
transform 1 0 52528 0 -1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1404_
timestamp 1698431365
transform 1 0 56672 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1405_
timestamp 1698431365
transform 1 0 55664 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1406_
timestamp 1698431365
transform -1 0 56224 0 -1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1407_
timestamp 1698431365
transform -1 0 57232 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1408_
timestamp 1698431365
transform 1 0 54432 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1409_
timestamp 1698431365
transform 1 0 55216 0 1 42336
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1410_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34944 0 -1 34496
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1411_
timestamp 1698431365
transform -1 0 19264 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1412_
timestamp 1698431365
transform -1 0 11200 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1413_
timestamp 1698431365
transform -1 0 16464 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1414_
timestamp 1698431365
transform 1 0 14448 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1415_
timestamp 1698431365
transform -1 0 18256 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1416_
timestamp 1698431365
transform -1 0 15008 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1417_
timestamp 1698431365
transform -1 0 13552 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1418_
timestamp 1698431365
transform -1 0 11424 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1419_
timestamp 1698431365
transform 1 0 20272 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1420_
timestamp 1698431365
transform -1 0 18816 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1421_
timestamp 1698431365
transform 1 0 9856 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1422_
timestamp 1698431365
transform 1 0 8960 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1423_
timestamp 1698431365
transform -1 0 20272 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1424_
timestamp 1698431365
transform -1 0 14448 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1425_
timestamp 1698431365
transform -1 0 8960 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1426_
timestamp 1698431365
transform -1 0 10528 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1427_
timestamp 1698431365
transform -1 0 8064 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1428_
timestamp 1698431365
transform 1 0 8400 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1429_
timestamp 1698431365
transform -1 0 8736 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1430_
timestamp 1698431365
transform 1 0 7840 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1431_
timestamp 1698431365
transform 1 0 9408 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1432_
timestamp 1698431365
transform 1 0 6160 0 1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1433_
timestamp 1698431365
transform 1 0 7280 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1434_
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1435_
timestamp 1698431365
transform 1 0 11872 0 1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1436_
timestamp 1698431365
transform -1 0 11872 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1437_
timestamp 1698431365
transform 1 0 48496 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1438_
timestamp 1698431365
transform -1 0 45696 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1439_
timestamp 1698431365
transform 1 0 44016 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1440_
timestamp 1698431365
transform 1 0 45472 0 -1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1441_
timestamp 1698431365
transform 1 0 44800 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1442_
timestamp 1698431365
transform -1 0 43792 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1443_
timestamp 1698431365
transform 1 0 42336 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1444_
timestamp 1698431365
transform 1 0 41664 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1445_
timestamp 1698431365
transform -1 0 42560 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1446_
timestamp 1698431365
transform 1 0 41888 0 1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1447_
timestamp 1698431365
transform -1 0 41776 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1448_
timestamp 1698431365
transform 1 0 39760 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1449_
timestamp 1698431365
transform 1 0 37744 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1450_
timestamp 1698431365
transform 1 0 36400 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1451_
timestamp 1698431365
transform 1 0 38976 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1452_
timestamp 1698431365
transform 1 0 36400 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1453_
timestamp 1698431365
transform -1 0 37744 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1454_
timestamp 1698431365
transform -1 0 33824 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1455_
timestamp 1698431365
transform 1 0 36848 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1456_
timestamp 1698431365
transform 1 0 37968 0 1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1457_
timestamp 1698431365
transform -1 0 42112 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1458_
timestamp 1698431365
transform 1 0 40208 0 1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1459_
timestamp 1698431365
transform 1 0 40768 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1460_
timestamp 1698431365
transform -1 0 43568 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1461_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42448 0 -1 48608
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1462_
timestamp 1698431365
transform 1 0 45024 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1463_
timestamp 1698431365
transform -1 0 54544 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1464_
timestamp 1698431365
transform -1 0 53088 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1465_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 52528 0 1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1466_
timestamp 1698431365
transform 1 0 50176 0 1 42336
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1467_
timestamp 1698431365
transform -1 0 50624 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1468_
timestamp 1698431365
transform 1 0 49616 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1469_
timestamp 1698431365
transform -1 0 53648 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1470_
timestamp 1698431365
transform 1 0 50288 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1471_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 54320 0 -1 43904
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1472_
timestamp 1698431365
transform 1 0 56896 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1473_
timestamp 1698431365
transform -1 0 56896 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1474_
timestamp 1698431365
transform 1 0 56448 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1475_
timestamp 1698431365
transform 1 0 56112 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1476_
timestamp 1698431365
transform 1 0 54768 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1477_
timestamp 1698431365
transform 1 0 54320 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1478_
timestamp 1698431365
transform 1 0 53536 0 1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1479_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 52528 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1480_
timestamp 1698431365
transform -1 0 54880 0 -1 47040
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1481_
timestamp 1698431365
transform -1 0 48272 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1482_
timestamp 1698431365
transform -1 0 47376 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1483_
timestamp 1698431365
transform 1 0 49504 0 -1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1484_
timestamp 1698431365
transform -1 0 52304 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1485_
timestamp 1698431365
transform 1 0 52640 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1486_
timestamp 1698431365
transform 1 0 54208 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1487_
timestamp 1698431365
transform 1 0 54880 0 -1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1488_
timestamp 1698431365
transform 1 0 45920 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1489_
timestamp 1698431365
transform 1 0 41216 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1490_
timestamp 1698431365
transform -1 0 39536 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1491_
timestamp 1698431365
transform 1 0 36176 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1492_
timestamp 1698431365
transform 1 0 36400 0 -1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1493_
timestamp 1698431365
transform 1 0 43680 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1494_
timestamp 1698431365
transform 1 0 37744 0 1 47040
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1495_
timestamp 1698431365
transform -1 0 45472 0 -1 48608
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1496_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 40544 0 -1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1497_
timestamp 1698431365
transform -1 0 41888 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1498_
timestamp 1698431365
transform 1 0 40544 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1499_
timestamp 1698431365
transform -1 0 57792 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1500_
timestamp 1698431365
transform -1 0 17584 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1501_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34384 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1502_
timestamp 1698431365
transform 1 0 16576 0 1 29792
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1503_
timestamp 1698431365
transform 1 0 33712 0 1 48608
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1504_
timestamp 1698431365
transform -1 0 34944 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1505_
timestamp 1698431365
transform 1 0 40656 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1506_
timestamp 1698431365
transform -1 0 41440 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1507_
timestamp 1698431365
transform -1 0 42448 0 -1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1508_
timestamp 1698431365
transform -1 0 18368 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1509_
timestamp 1698431365
transform -1 0 15456 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1510_
timestamp 1698431365
transform 1 0 14784 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1511_
timestamp 1698431365
transform -1 0 17248 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1512_
timestamp 1698431365
transform 1 0 15680 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1513_
timestamp 1698431365
transform 1 0 41440 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1514_
timestamp 1698431365
transform -1 0 32704 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1515_
timestamp 1698431365
transform -1 0 32368 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1516_
timestamp 1698431365
transform 1 0 32928 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1517_
timestamp 1698431365
transform 1 0 37296 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1518_
timestamp 1698431365
transform 1 0 41328 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1519_
timestamp 1698431365
transform -1 0 36624 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1520_
timestamp 1698431365
transform 1 0 35728 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1521_
timestamp 1698431365
transform 1 0 34944 0 -1 48608
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1522_
timestamp 1698431365
transform -1 0 36512 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1523_
timestamp 1698431365
transform 1 0 36848 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1524_
timestamp 1698431365
transform 1 0 35728 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1525_
timestamp 1698431365
transform -1 0 37744 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1526_
timestamp 1698431365
transform -1 0 43008 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1527_
timestamp 1698431365
transform 1 0 38976 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1528_
timestamp 1698431365
transform 1 0 39648 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1529_
timestamp 1698431365
transform 1 0 40768 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1530_
timestamp 1698431365
transform -1 0 40544 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1531_
timestamp 1698431365
transform 1 0 40768 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1532_
timestamp 1698431365
transform -1 0 41440 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1533_
timestamp 1698431365
transform 1 0 42224 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1534_
timestamp 1698431365
transform 1 0 40992 0 1 53312
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1535_
timestamp 1698431365
transform 1 0 42784 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1536_
timestamp 1698431365
transform 1 0 45584 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1537_
timestamp 1698431365
transform -1 0 47264 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1538_
timestamp 1698431365
transform 1 0 43568 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1539_
timestamp 1698431365
transform 1 0 44688 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1540_
timestamp 1698431365
transform 1 0 46368 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1541_
timestamp 1698431365
transform 1 0 55776 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1542_
timestamp 1698431365
transform 1 0 45808 0 -1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1543_
timestamp 1698431365
transform 1 0 47152 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1544_
timestamp 1698431365
transform -1 0 50512 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1545_
timestamp 1698431365
transform 1 0 47936 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1546_
timestamp 1698431365
transform 1 0 49392 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1547_
timestamp 1698431365
transform 1 0 48496 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1548_
timestamp 1698431365
transform 1 0 48608 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1549_
timestamp 1698431365
transform 1 0 50400 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1550_
timestamp 1698431365
transform -1 0 49952 0 -1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1551_
timestamp 1698431365
transform -1 0 48720 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1552_
timestamp 1698431365
transform -1 0 51408 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1553_
timestamp 1698431365
transform 1 0 50064 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1554_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 49504 0 -1 51744
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1555_
timestamp 1698431365
transform 1 0 50848 0 1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1556_
timestamp 1698431365
transform 1 0 51184 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1557_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 49280 0 1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1558_
timestamp 1698431365
transform 1 0 49728 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1559_
timestamp 1698431365
transform -1 0 51184 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1560_
timestamp 1698431365
transform 1 0 52528 0 1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1561_
timestamp 1698431365
transform 1 0 54208 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1562_
timestamp 1698431365
transform 1 0 54880 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1563_
timestamp 1698431365
transform 1 0 54544 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1564_
timestamp 1698431365
transform 1 0 56448 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1565_
timestamp 1698431365
transform 1 0 54880 0 -1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1566_
timestamp 1698431365
transform -1 0 56224 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1567_
timestamp 1698431365
transform 1 0 56448 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1568_
timestamp 1698431365
transform -1 0 57344 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1569_
timestamp 1698431365
transform 1 0 15344 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1570_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16912 0 1 43904
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1571_
timestamp 1698431365
transform -1 0 17024 0 -1 45472
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1572_
timestamp 1698431365
transform -1 0 15008 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1573_
timestamp 1698431365
transform -1 0 16128 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1574_
timestamp 1698431365
transform 1 0 13664 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1575_
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1576_
timestamp 1698431365
transform -1 0 9408 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1577_
timestamp 1698431365
transform 1 0 8512 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1578_
timestamp 1698431365
transform 1 0 11648 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1579_
timestamp 1698431365
transform -1 0 9968 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1580_
timestamp 1698431365
transform -1 0 8736 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1581_
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1582_
timestamp 1698431365
transform 1 0 10416 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1583_
timestamp 1698431365
transform 1 0 10864 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1584_
timestamp 1698431365
transform 1 0 11872 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1585_
timestamp 1698431365
transform -1 0 11872 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1586_
timestamp 1698431365
transform 1 0 10976 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1587_
timestamp 1698431365
transform 1 0 10976 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1588_
timestamp 1698431365
transform 1 0 10528 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1589_
timestamp 1698431365
transform 1 0 10304 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1590_
timestamp 1698431365
transform 1 0 10864 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1591_
timestamp 1698431365
transform -1 0 8176 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1592_
timestamp 1698431365
transform -1 0 7056 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1593_
timestamp 1698431365
transform 1 0 7168 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1594_
timestamp 1698431365
transform -1 0 9296 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1595_
timestamp 1698431365
transform -1 0 7728 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1596_
timestamp 1698431365
transform -1 0 8736 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1597_
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1598_
timestamp 1698431365
transform -1 0 6160 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1599_
timestamp 1698431365
transform 1 0 6384 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1600_
timestamp 1698431365
transform -1 0 6384 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1601_
timestamp 1698431365
transform -1 0 5152 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1602_
timestamp 1698431365
transform 1 0 3024 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1603_
timestamp 1698431365
transform 1 0 3584 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1604_
timestamp 1698431365
transform -1 0 4704 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1605_
timestamp 1698431365
transform -1 0 5376 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1606_
timestamp 1698431365
transform 1 0 3696 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1607_
timestamp 1698431365
transform -1 0 6608 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1608_
timestamp 1698431365
transform 1 0 4032 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1609_
timestamp 1698431365
transform -1 0 6048 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1610_
timestamp 1698431365
transform -1 0 6720 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1611_
timestamp 1698431365
transform -1 0 5264 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1612_
timestamp 1698431365
transform -1 0 6272 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1613_
timestamp 1698431365
transform -1 0 6160 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1614_
timestamp 1698431365
transform 1 0 4592 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1615_
timestamp 1698431365
transform 1 0 4816 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1616_
timestamp 1698431365
transform 1 0 4704 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1617_
timestamp 1698431365
transform 1 0 4144 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1618_
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1619_
timestamp 1698431365
transform -1 0 6048 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1620_
timestamp 1698431365
transform -1 0 5264 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1621_
timestamp 1698431365
transform 1 0 4256 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1622_
timestamp 1698431365
transform -1 0 7728 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1623_
timestamp 1698431365
transform -1 0 7056 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1624_
timestamp 1698431365
transform 1 0 5264 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1625_
timestamp 1698431365
transform -1 0 11536 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1626_
timestamp 1698431365
transform 1 0 5600 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1627_
timestamp 1698431365
transform 1 0 5488 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1628_
timestamp 1698431365
transform -1 0 9072 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1629_
timestamp 1698431365
transform -1 0 5488 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1630_
timestamp 1698431365
transform 1 0 6048 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1631_
timestamp 1698431365
transform -1 0 9856 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1632_
timestamp 1698431365
transform 1 0 7392 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1633_
timestamp 1698431365
transform -1 0 7840 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1634_
timestamp 1698431365
transform -1 0 9072 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1635_
timestamp 1698431365
transform 1 0 8736 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1636_
timestamp 1698431365
transform -1 0 9184 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1637_
timestamp 1698431365
transform 1 0 8624 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1638_
timestamp 1698431365
transform 1 0 8064 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1639_
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1640_
timestamp 1698431365
transform -1 0 6272 0 -1 29792
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1641_
timestamp 1698431365
transform 1 0 5152 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1642_
timestamp 1698431365
transform -1 0 8960 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1643_
timestamp 1698431365
transform -1 0 8064 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1644_
timestamp 1698431365
transform -1 0 9072 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1645_
timestamp 1698431365
transform 1 0 8176 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1646_
timestamp 1698431365
transform -1 0 10192 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1647_
timestamp 1698431365
transform -1 0 8064 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1648_
timestamp 1698431365
transform -1 0 8960 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1649_
timestamp 1698431365
transform -1 0 8064 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1650_
timestamp 1698431365
transform 1 0 33376 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1651_
timestamp 1698431365
transform -1 0 34944 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1652_
timestamp 1698431365
transform 1 0 33488 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1653_
timestamp 1698431365
transform -1 0 35728 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1654_
timestamp 1698431365
transform 1 0 33040 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1655_
timestamp 1698431365
transform 1 0 34048 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1656_
timestamp 1698431365
transform -1 0 33936 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1657_
timestamp 1698431365
transform -1 0 34608 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1658_
timestamp 1698431365
transform -1 0 38528 0 -1 14112
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1659_
timestamp 1698431365
transform -1 0 34160 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1660_
timestamp 1698431365
transform 1 0 34496 0 1 12544
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1661_
timestamp 1698431365
transform 1 0 35056 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1662_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34608 0 -1 15680
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1663_
timestamp 1698431365
transform -1 0 28560 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1664_
timestamp 1698431365
transform 1 0 27664 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1665_
timestamp 1698431365
transform 1 0 28784 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1666_
timestamp 1698431365
transform -1 0 32704 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1667_
timestamp 1698431365
transform 1 0 29456 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1668_
timestamp 1698431365
transform -1 0 31024 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1669_
timestamp 1698431365
transform -1 0 32592 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1670_
timestamp 1698431365
transform 1 0 41216 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1671_
timestamp 1698431365
transform 1 0 31472 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1672_
timestamp 1698431365
transform -1 0 31472 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1673_
timestamp 1698431365
transform -1 0 31696 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1674_
timestamp 1698431365
transform 1 0 31472 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1675_
timestamp 1698431365
transform -1 0 31472 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1676_
timestamp 1698431365
transform 1 0 30576 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1677_
timestamp 1698431365
transform -1 0 30576 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1678_
timestamp 1698431365
transform -1 0 28784 0 1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1679_
timestamp 1698431365
transform 1 0 26880 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1680_
timestamp 1698431365
transform -1 0 32032 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1681_
timestamp 1698431365
transform -1 0 19936 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1682_
timestamp 1698431365
transform 1 0 16576 0 1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1683_
timestamp 1698431365
transform -1 0 15008 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1684_
timestamp 1698431365
transform 1 0 18368 0 -1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1685_
timestamp 1698431365
transform 1 0 18480 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1686_
timestamp 1698431365
transform 1 0 16016 0 -1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1687_
timestamp 1698431365
transform -1 0 12992 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1688_
timestamp 1698431365
transform 1 0 18368 0 -1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1689_
timestamp 1698431365
transform -1 0 18256 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1690_
timestamp 1698431365
transform -1 0 47152 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1691_
timestamp 1698431365
transform -1 0 46032 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1692_
timestamp 1698431365
transform 1 0 40992 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1693_
timestamp 1698431365
transform -1 0 45136 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1694_
timestamp 1698431365
transform -1 0 48160 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1695_
timestamp 1698431365
transform -1 0 46256 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1696_
timestamp 1698431365
transform 1 0 45808 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1697_
timestamp 1698431365
transform 1 0 46032 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1698_
timestamp 1698431365
transform 1 0 46256 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1699_
timestamp 1698431365
transform -1 0 47488 0 -1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1700_
timestamp 1698431365
transform 1 0 47376 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1701_
timestamp 1698431365
transform -1 0 47712 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1702_
timestamp 1698431365
transform 1 0 45360 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1703_
timestamp 1698431365
transform -1 0 54656 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1704_
timestamp 1698431365
transform 1 0 39984 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1705_
timestamp 1698431365
transform 1 0 50848 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1706_
timestamp 1698431365
transform -1 0 49056 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1707_
timestamp 1698431365
transform -1 0 50400 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1708_
timestamp 1698431365
transform -1 0 50848 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1709_
timestamp 1698431365
transform -1 0 49952 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1710_
timestamp 1698431365
transform -1 0 48384 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1711_
timestamp 1698431365
transform 1 0 47936 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1712_
timestamp 1698431365
transform -1 0 49616 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1713_
timestamp 1698431365
transform -1 0 48384 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1714_
timestamp 1698431365
transform 1 0 47040 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1715_
timestamp 1698431365
transform -1 0 54208 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1716_
timestamp 1698431365
transform 1 0 51744 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1717_
timestamp 1698431365
transform 1 0 50512 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1718_
timestamp 1698431365
transform -1 0 54208 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1719_
timestamp 1698431365
transform 1 0 51856 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1720_
timestamp 1698431365
transform 1 0 52528 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1721_
timestamp 1698431365
transform 1 0 46816 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1722_
timestamp 1698431365
transform -1 0 48160 0 -1 12544
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1723_
timestamp 1698431365
transform -1 0 51296 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1724_
timestamp 1698431365
transform -1 0 50512 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1725_
timestamp 1698431365
transform 1 0 52640 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1726_
timestamp 1698431365
transform -1 0 53648 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1727_
timestamp 1698431365
transform -1 0 50176 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1728_
timestamp 1698431365
transform -1 0 51184 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1729_
timestamp 1698431365
transform 1 0 47936 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1730_
timestamp 1698431365
transform -1 0 51184 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1731_
timestamp 1698431365
transform 1 0 45024 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1732_
timestamp 1698431365
transform 1 0 46144 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1733_
timestamp 1698431365
transform 1 0 49616 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1734_
timestamp 1698431365
transform -1 0 51632 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1735_
timestamp 1698431365
transform 1 0 49616 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1736_
timestamp 1698431365
transform 1 0 49728 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1737_
timestamp 1698431365
transform -1 0 49504 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1738_
timestamp 1698431365
transform 1 0 46704 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1739_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 49728 0 1 9408
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1740_
timestamp 1698431365
transform -1 0 43792 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1741_
timestamp 1698431365
transform 1 0 43792 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1742_
timestamp 1698431365
transform 1 0 44912 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1743_
timestamp 1698431365
transform 1 0 43680 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1744_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 46144 0 -1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1745_
timestamp 1698431365
transform 1 0 39088 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1746_
timestamp 1698431365
transform 1 0 44128 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1747_
timestamp 1698431365
transform -1 0 44464 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1748_
timestamp 1698431365
transform -1 0 47040 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1749_
timestamp 1698431365
transform 1 0 47040 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1750_
timestamp 1698431365
transform 1 0 48608 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1751_
timestamp 1698431365
transform 1 0 49168 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1752_
timestamp 1698431365
transform 1 0 51632 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1753_
timestamp 1698431365
transform 1 0 47152 0 -1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1754_
timestamp 1698431365
transform 1 0 52304 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1755_
timestamp 1698431365
transform 1 0 53200 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1756_
timestamp 1698431365
transform 1 0 52864 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1757_
timestamp 1698431365
transform 1 0 54432 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1758_
timestamp 1698431365
transform 1 0 52864 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1759_
timestamp 1698431365
transform 1 0 54208 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1760_
timestamp 1698431365
transform 1 0 55552 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1761_
timestamp 1698431365
transform -1 0 42784 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1762_
timestamp 1698431365
transform 1 0 37520 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1763_
timestamp 1698431365
transform 1 0 52304 0 -1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1764_
timestamp 1698431365
transform 1 0 52640 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1765_
timestamp 1698431365
transform 1 0 52528 0 1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1766_
timestamp 1698431365
transform 1 0 53648 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1767_
timestamp 1698431365
transform 1 0 55216 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1768_
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1769_
timestamp 1698431365
transform -1 0 55664 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1770_
timestamp 1698431365
transform -1 0 53984 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1771_
timestamp 1698431365
transform 1 0 53648 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1772_
timestamp 1698431365
transform 1 0 56448 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1773_
timestamp 1698431365
transform 1 0 53312 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1774_
timestamp 1698431365
transform 1 0 54656 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1775_
timestamp 1698431365
transform 1 0 56448 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1776_
timestamp 1698431365
transform -1 0 54544 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1777_
timestamp 1698431365
transform -1 0 53648 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1778_
timestamp 1698431365
transform 1 0 52976 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1779_
timestamp 1698431365
transform 1 0 53648 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1780_
timestamp 1698431365
transform 1 0 49728 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1781_
timestamp 1698431365
transform -1 0 50288 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1782_
timestamp 1698431365
transform 1 0 49840 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1783_
timestamp 1698431365
transform 1 0 50848 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1784_
timestamp 1698431365
transform -1 0 47712 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1785_
timestamp 1698431365
transform 1 0 45360 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1786_
timestamp 1698431365
transform 1 0 47264 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1787_
timestamp 1698431365
transform -1 0 49728 0 1 6272
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1788_
timestamp 1698431365
transform -1 0 44128 0 1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1789_
timestamp 1698431365
transform -1 0 32256 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1790_
timestamp 1698431365
transform 1 0 31136 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1791_
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1792_
timestamp 1698431365
transform -1 0 47712 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1793_
timestamp 1698431365
transform 1 0 43120 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1794_
timestamp 1698431365
transform -1 0 54096 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1795_
timestamp 1698431365
transform -1 0 52976 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1796_
timestamp 1698431365
transform -1 0 51968 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1797_
timestamp 1698431365
transform -1 0 51296 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1798_
timestamp 1698431365
transform -1 0 54320 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1799_
timestamp 1698431365
transform -1 0 55104 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1800_
timestamp 1698431365
transform -1 0 54656 0 1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1801_
timestamp 1698431365
transform -1 0 53200 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1802_
timestamp 1698431365
transform 1 0 51632 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1803_
timestamp 1698431365
transform -1 0 52864 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1804_
timestamp 1698431365
transform 1 0 51408 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1805_
timestamp 1698431365
transform 1 0 50848 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1806_
timestamp 1698431365
transform -1 0 49392 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1807_
timestamp 1698431365
transform 1 0 47264 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1808_
timestamp 1698431365
transform 1 0 48048 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1809_
timestamp 1698431365
transform 1 0 43568 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1810_
timestamp 1698431365
transform 1 0 44352 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1811_
timestamp 1698431365
transform 1 0 45920 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1812_
timestamp 1698431365
transform 1 0 46256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1813_
timestamp 1698431365
transform 1 0 43120 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1814_
timestamp 1698431365
transform -1 0 47936 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1815_
timestamp 1698431365
transform 1 0 48608 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1816_
timestamp 1698431365
transform -1 0 48832 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1817_
timestamp 1698431365
transform 1 0 50624 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1818_
timestamp 1698431365
transform 1 0 49504 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1819_
timestamp 1698431365
transform 1 0 49840 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1820_
timestamp 1698431365
transform 1 0 50176 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1821_
timestamp 1698431365
transform -1 0 50624 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1822_
timestamp 1698431365
transform 1 0 49280 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1823_
timestamp 1698431365
transform -1 0 54656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1824_
timestamp 1698431365
transform 1 0 53200 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1825_
timestamp 1698431365
transform 1 0 53200 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1826_
timestamp 1698431365
transform 1 0 51408 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1827_
timestamp 1698431365
transform 1 0 52080 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1828_
timestamp 1698431365
transform -1 0 53648 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1829_
timestamp 1698431365
transform -1 0 53536 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1830_
timestamp 1698431365
transform -1 0 52976 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1831_
timestamp 1698431365
transform 1 0 50848 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1832_
timestamp 1698431365
transform 1 0 49280 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1833_
timestamp 1698431365
transform -1 0 52304 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1834_
timestamp 1698431365
transform -1 0 49616 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1835_
timestamp 1698431365
transform 1 0 49616 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1836_
timestamp 1698431365
transform 1 0 48608 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1837_
timestamp 1698431365
transform 1 0 49616 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1838_
timestamp 1698431365
transform 1 0 48944 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1839_
timestamp 1698431365
transform 1 0 49056 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1840_
timestamp 1698431365
transform -1 0 50848 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1841_
timestamp 1698431365
transform 1 0 48720 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1842_
timestamp 1698431365
transform 1 0 47376 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1843_
timestamp 1698431365
transform -1 0 52304 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1844_
timestamp 1698431365
transform -1 0 51632 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1845_
timestamp 1698431365
transform -1 0 51408 0 -1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1846_
timestamp 1698431365
transform 1 0 49504 0 1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1847_
timestamp 1698431365
transform -1 0 50960 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1848_
timestamp 1698431365
transform -1 0 38416 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1849_
timestamp 1698431365
transform -1 0 45584 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1850_
timestamp 1698431365
transform 1 0 44576 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1851_
timestamp 1698431365
transform 1 0 45136 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1852_
timestamp 1698431365
transform -1 0 46256 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1853_
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1854_
timestamp 1698431365
transform 1 0 44016 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1855_
timestamp 1698431365
transform 1 0 44912 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1856_
timestamp 1698431365
transform 1 0 46816 0 -1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1857_
timestamp 1698431365
transform 1 0 49056 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1858_
timestamp 1698431365
transform 1 0 45248 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1859_
timestamp 1698431365
transform -1 0 46256 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1860_
timestamp 1698431365
transform 1 0 46256 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1861_
timestamp 1698431365
transform 1 0 47040 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1862_
timestamp 1698431365
transform -1 0 48160 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1863_
timestamp 1698431365
transform 1 0 52528 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1864_
timestamp 1698431365
transform 1 0 53088 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1865_
timestamp 1698431365
transform 1 0 54432 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1866_
timestamp 1698431365
transform -1 0 54656 0 -1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1867_
timestamp 1698431365
transform 1 0 52976 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1868_
timestamp 1698431365
transform 1 0 52528 0 1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1869_
timestamp 1698431365
transform 1 0 54096 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1870_
timestamp 1698431365
transform 1 0 54096 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1871_
timestamp 1698431365
transform 1 0 55440 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1872_
timestamp 1698431365
transform 1 0 53872 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1873_
timestamp 1698431365
transform 1 0 54992 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1874_
timestamp 1698431365
transform -1 0 55104 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1875_
timestamp 1698431365
transform 1 0 54432 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1876_
timestamp 1698431365
transform 1 0 56448 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1877_
timestamp 1698431365
transform -1 0 56224 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1878_
timestamp 1698431365
transform -1 0 56112 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1879_
timestamp 1698431365
transform -1 0 55440 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1880_
timestamp 1698431365
transform 1 0 55104 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1881_
timestamp 1698431365
transform 1 0 51296 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1882_
timestamp 1698431365
transform 1 0 52640 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1883_
timestamp 1698431365
transform -1 0 53088 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1884_
timestamp 1698431365
transform -1 0 48384 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1885_
timestamp 1698431365
transform 1 0 35392 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1886_
timestamp 1698431365
transform -1 0 36400 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1887_
timestamp 1698431365
transform -1 0 37632 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1888_
timestamp 1698431365
transform 1 0 28112 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1889_
timestamp 1698431365
transform -1 0 30688 0 1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1890_
timestamp 1698431365
transform -1 0 21840 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1891_
timestamp 1698431365
transform -1 0 27552 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1892_
timestamp 1698431365
transform -1 0 23968 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1893_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20496 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1894_
timestamp 1698431365
transform 1 0 28336 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1895_
timestamp 1698431365
transform -1 0 30128 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1896_
timestamp 1698431365
transform 1 0 26656 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1897_
timestamp 1698431365
transform 1 0 25088 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1898_
timestamp 1698431365
transform 1 0 26544 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1899_
timestamp 1698431365
transform 1 0 24304 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1900_
timestamp 1698431365
transform -1 0 26544 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1901_
timestamp 1698431365
transform 1 0 26208 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1902_
timestamp 1698431365
transform -1 0 26544 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1903_
timestamp 1698431365
transform -1 0 28336 0 1 47040
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1904_
timestamp 1698431365
transform 1 0 26432 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1905_
timestamp 1698431365
transform 1 0 26992 0 -1 48608
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1906_
timestamp 1698431365
transform -1 0 30128 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1907_
timestamp 1698431365
transform -1 0 28560 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1908_
timestamp 1698431365
transform -1 0 30800 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1909_
timestamp 1698431365
transform -1 0 29680 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1910_
timestamp 1698431365
transform -1 0 32032 0 -1 47040
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1911_
timestamp 1698431365
transform 1 0 22736 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1912_
timestamp 1698431365
transform -1 0 27328 0 -1 47040
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1913_
timestamp 1698431365
transform 1 0 26656 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1914_
timestamp 1698431365
transform -1 0 29904 0 -1 45472
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1915_
timestamp 1698431365
transform -1 0 22176 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1916_
timestamp 1698431365
transform -1 0 26656 0 1 45472
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1917_
timestamp 1698431365
transform -1 0 24416 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1918_
timestamp 1698431365
transform -1 0 24416 0 -1 45472
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1919_
timestamp 1698431365
transform -1 0 23184 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1920_
timestamp 1698431365
transform 1 0 23184 0 1 43904
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1921_
timestamp 1698431365
transform 1 0 25536 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1922_
timestamp 1698431365
transform -1 0 24192 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1923_
timestamp 1698431365
transform 1 0 22624 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1924_
timestamp 1698431365
transform -1 0 24192 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1925_
timestamp 1698431365
transform 1 0 25984 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1926_
timestamp 1698431365
transform 1 0 30352 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1927_
timestamp 1698431365
transform -1 0 32368 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1928_
timestamp 1698431365
transform -1 0 32032 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1929_
timestamp 1698431365
transform 1 0 31360 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1930_
timestamp 1698431365
transform -1 0 31584 0 -1 50176
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1931_
timestamp 1698431365
transform 1 0 30464 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1932_
timestamp 1698431365
transform 1 0 31248 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1933_
timestamp 1698431365
transform 1 0 22848 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1934_
timestamp 1698431365
transform -1 0 26432 0 1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1935_
timestamp 1698431365
transform -1 0 24080 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1936_
timestamp 1698431365
transform 1 0 26656 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1937_
timestamp 1698431365
transform -1 0 27888 0 1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1938_
timestamp 1698431365
transform -1 0 27552 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1939_
timestamp 1698431365
transform -1 0 28784 0 1 53312
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1940_
timestamp 1698431365
transform 1 0 27888 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1941_
timestamp 1698431365
transform 1 0 29120 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1942_
timestamp 1698431365
transform 1 0 21168 0 -1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1943_
timestamp 1698431365
transform 1 0 22512 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1944_
timestamp 1698431365
transform -1 0 22288 0 1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1945_
timestamp 1698431365
transform -1 0 22064 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1946_
timestamp 1698431365
transform -1 0 20944 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1947_
timestamp 1698431365
transform 1 0 21168 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1948_
timestamp 1698431365
transform 1 0 18704 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1949_
timestamp 1698431365
transform 1 0 20496 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1950_
timestamp 1698431365
transform 1 0 19600 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1951_
timestamp 1698431365
transform 1 0 19600 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1952_
timestamp 1698431365
transform 1 0 19600 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1953_
timestamp 1698431365
transform 1 0 19376 0 1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1954_
timestamp 1698431365
transform -1 0 20496 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1955_
timestamp 1698431365
transform 1 0 21840 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1956_
timestamp 1698431365
transform -1 0 22176 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1957_
timestamp 1698431365
transform 1 0 25312 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1958_
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1959_
timestamp 1698431365
transform -1 0 28896 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1960_
timestamp 1698431365
transform -1 0 27328 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1961_
timestamp 1698431365
transform 1 0 25312 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1962_
timestamp 1698431365
transform 1 0 25760 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1963_
timestamp 1698431365
transform 1 0 24192 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1964_
timestamp 1698431365
transform 1 0 25200 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1965_
timestamp 1698431365
transform -1 0 15904 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1966_
timestamp 1698431365
transform 1 0 12208 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1967_
timestamp 1698431365
transform -1 0 16240 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1968_
timestamp 1698431365
transform -1 0 14000 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1969_
timestamp 1698431365
transform -1 0 14224 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1970_
timestamp 1698431365
transform 1 0 15008 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1971_
timestamp 1698431365
transform 1 0 15904 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1972_
timestamp 1698431365
transform -1 0 16688 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1973_
timestamp 1698431365
transform -1 0 18144 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1974_
timestamp 1698431365
transform 1 0 15680 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1975_
timestamp 1698431365
transform 1 0 16576 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1976_
timestamp 1698431365
transform -1 0 16800 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1977_
timestamp 1698431365
transform -1 0 16576 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1978_
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1979_
timestamp 1698431365
transform -1 0 16576 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1980_
timestamp 1698431365
transform -1 0 16352 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1981_
timestamp 1698431365
transform 1 0 16352 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1982_
timestamp 1698431365
transform -1 0 16800 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1983_
timestamp 1698431365
transform -1 0 17024 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1984_
timestamp 1698431365
transform 1 0 15680 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1985_
timestamp 1698431365
transform 1 0 54208 0 1 37632
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1986_
timestamp 1698431365
transform -1 0 37632 0 -1 39200
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1987_
timestamp 1698431365
transform -1 0 36512 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1988_
timestamp 1698431365
transform -1 0 34272 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1989_
timestamp 1698431365
transform -1 0 33712 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1990_
timestamp 1698431365
transform -1 0 32368 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1991_
timestamp 1698431365
transform -1 0 35840 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1992_
timestamp 1698431365
transform -1 0 33712 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1993_
timestamp 1698431365
transform 1 0 33040 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1994_
timestamp 1698431365
transform -1 0 32816 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1995_
timestamp 1698431365
transform 1 0 31808 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1996_
timestamp 1698431365
transform -1 0 36064 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1997_
timestamp 1698431365
transform -1 0 36624 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1998_
timestamp 1698431365
transform -1 0 36400 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1999_
timestamp 1698431365
transform -1 0 37296 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2000_
timestamp 1698431365
transform 1 0 38304 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2001_
timestamp 1698431365
transform -1 0 39424 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2002_
timestamp 1698431365
transform -1 0 41440 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2003_
timestamp 1698431365
transform -1 0 40096 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2004_
timestamp 1698431365
transform 1 0 37408 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2005_
timestamp 1698431365
transform -1 0 37408 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2006_
timestamp 1698431365
transform -1 0 38752 0 -1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2007_
timestamp 1698431365
transform -1 0 36512 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2008_
timestamp 1698431365
transform 1 0 37296 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2009_
timestamp 1698431365
transform -1 0 35616 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2010_
timestamp 1698431365
transform -1 0 39760 0 -1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2011_
timestamp 1698431365
transform -1 0 40208 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2012_
timestamp 1698431365
transform 1 0 41440 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2013_
timestamp 1698431365
transform 1 0 40880 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2014_
timestamp 1698431365
transform 1 0 41776 0 1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2015_
timestamp 1698431365
transform 1 0 41776 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2016_
timestamp 1698431365
transform -1 0 44352 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2017_
timestamp 1698431365
transform -1 0 42560 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2018_
timestamp 1698431365
transform -1 0 43232 0 1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2019_
timestamp 1698431365
transform -1 0 42224 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2020_
timestamp 1698431365
transform -1 0 44240 0 1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2021_
timestamp 1698431365
transform 1 0 43904 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2022_
timestamp 1698431365
transform -1 0 18144 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2023_
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2024_
timestamp 1698431365
transform -1 0 17024 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2025_
timestamp 1698431365
transform -1 0 14896 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2026_
timestamp 1698431365
transform -1 0 14672 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2027_
timestamp 1698431365
transform 1 0 13104 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2028_
timestamp 1698431365
transform -1 0 13104 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2029_
timestamp 1698431365
transform 1 0 12768 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2030_
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2031_
timestamp 1698431365
transform 1 0 13664 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2032_
timestamp 1698431365
transform 1 0 13328 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2033_
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2034_
timestamp 1698431365
transform 1 0 14224 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2035_
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2036_
timestamp 1698431365
transform 1 0 18144 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2037_
timestamp 1698431365
transform -1 0 16912 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2038_
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2039_
timestamp 1698431365
transform 1 0 19264 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2040_
timestamp 1698431365
transform 1 0 18816 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2041_
timestamp 1698431365
transform 1 0 18816 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2042_
timestamp 1698431365
transform 1 0 18592 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2043_
timestamp 1698431365
transform 1 0 19936 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2044_
timestamp 1698431365
transform -1 0 18592 0 1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2045_
timestamp 1698431365
transform 1 0 17696 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2046_
timestamp 1698431365
transform -1 0 34608 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2047_
timestamp 1698431365
transform -1 0 31920 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2048_
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2049_
timestamp 1698431365
transform 1 0 30688 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2050_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34160 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2051_
timestamp 1698431365
transform -1 0 40432 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2052_
timestamp 1698431365
transform -1 0 40096 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2053_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34272 0 -1 10976
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2054_
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2055_
timestamp 1698431365
transform 1 0 36400 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2056_
timestamp 1698431365
transform 1 0 41216 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2057_
timestamp 1698431365
transform 1 0 40992 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2058_
timestamp 1698431365
transform 1 0 37296 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2059_
timestamp 1698431365
transform 1 0 24080 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2060_
timestamp 1698431365
transform 1 0 26656 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2061_
timestamp 1698431365
transform 1 0 19712 0 -1 36064
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2062_
timestamp 1698431365
transform 1 0 20272 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2063_
timestamp 1698431365
transform -1 0 28784 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2064_
timestamp 1698431365
transform 1 0 22512 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2065_
timestamp 1698431365
transform -1 0 26768 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2066_
timestamp 1698431365
transform 1 0 19040 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2067_
timestamp 1698431365
transform 1 0 10192 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2068_
timestamp 1698431365
transform 1 0 15232 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2069_
timestamp 1698431365
transform 1 0 9856 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2070_
timestamp 1698431365
transform 1 0 11088 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2071_
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2072_
timestamp 1698431365
transform 1 0 23968 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2073_
timestamp 1698431365
transform -1 0 28448 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2074_
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2075_
timestamp 1698431365
transform 1 0 18704 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2076_
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2077_
timestamp 1698431365
transform -1 0 20384 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2078_
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2079_
timestamp 1698431365
transform 1 0 13664 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2080_
timestamp 1698431365
transform -1 0 20944 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2081_
timestamp 1698431365
transform 1 0 21168 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2082_
timestamp 1698431365
transform 1 0 17696 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2083_
timestamp 1698431365
transform 1 0 10528 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2084_
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2085_
timestamp 1698431365
transform -1 0 7616 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2086_
timestamp 1698431365
transform 1 0 4592 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2087_
timestamp 1698431365
transform -1 0 11984 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2088_
timestamp 1698431365
transform 1 0 6160 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2089_
timestamp 1698431365
transform 1 0 9968 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2090_
timestamp 1698431365
transform -1 0 41104 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2091_
timestamp 1698431365
transform 1 0 40768 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2092_
timestamp 1698431365
transform 1 0 42784 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2093_
timestamp 1698431365
transform -1 0 44464 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2094_
timestamp 1698431365
transform -1 0 51744 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2095_
timestamp 1698431365
transform 1 0 50960 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2096_
timestamp 1698431365
transform 1 0 55104 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2097_
timestamp 1698431365
transform 1 0 55104 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2098_
timestamp 1698431365
transform 1 0 38416 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2099_
timestamp 1698431365
transform 1 0 40880 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2100_
timestamp 1698431365
transform 1 0 41216 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2101_
timestamp 1698431365
transform 1 0 37072 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2102_
timestamp 1698431365
transform 1 0 43008 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2103_
timestamp 1698431365
transform 1 0 38976 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2104_
timestamp 1698431365
transform 1 0 37296 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2105_
timestamp 1698431365
transform 1 0 41664 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2106_
timestamp 1698431365
transform 1 0 48496 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2107_
timestamp 1698431365
transform 1 0 51072 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2108_
timestamp 1698431365
transform 1 0 55104 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2109_
timestamp 1698431365
transform -1 0 56224 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2110_
timestamp 1698431365
transform 1 0 29120 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2111_
timestamp 1698431365
transform 1 0 29232 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2112_
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2113_
timestamp 1698431365
transform -1 0 36624 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2114_
timestamp 1698431365
transform -1 0 36400 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2115_
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2116_
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2117_
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2118_
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2119_
timestamp 1698431365
transform 1 0 2016 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2120_
timestamp 1698431365
transform -1 0 10416 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2121_
timestamp 1698431365
transform -1 0 9072 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2122_
timestamp 1698431365
transform 1 0 9744 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2123_
timestamp 1698431365
transform -1 0 29680 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2124_
timestamp 1698431365
transform 1 0 21168 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2125_
timestamp 1698431365
transform 1 0 20608 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2126_
timestamp 1698431365
transform 1 0 20272 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2127_
timestamp 1698431365
transform 1 0 24192 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2128_
timestamp 1698431365
transform 1 0 25088 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2129_
timestamp 1698431365
transform -1 0 34496 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2130_
timestamp 1698431365
transform 1 0 27776 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2131_
timestamp 1698431365
transform -1 0 34608 0 1 43904
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2132_
timestamp 1698431365
transform -1 0 30800 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2133_
timestamp 1698431365
transform 1 0 35952 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2134_
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2135_
timestamp 1698431365
transform 1 0 38304 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2136_
timestamp 1698431365
transform 1 0 6496 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2137_
timestamp 1698431365
transform 1 0 21616 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2138_
timestamp 1698431365
transform 1 0 18816 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2139_
timestamp 1698431365
transform 1 0 27328 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2140_
timestamp 1698431365
transform 1 0 18704 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2141_
timestamp 1698431365
transform -1 0 36960 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2142_
timestamp 1698431365
transform 1 0 29456 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2143_
timestamp 1698431365
transform 1 0 44688 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2144_
timestamp 1698431365
transform 1 0 45136 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2145_
timestamp 1698431365
transform 1 0 45024 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2146_
timestamp 1698431365
transform 1 0 48720 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2147_
timestamp 1698431365
transform -1 0 53088 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2148_
timestamp 1698431365
transform 1 0 51968 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2149_
timestamp 1698431365
transform 1 0 55104 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2150_
timestamp 1698431365
transform 1 0 55104 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2151_
timestamp 1698431365
transform 1 0 17248 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2152_
timestamp 1698431365
transform 1 0 8288 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2153_
timestamp 1698431365
transform -1 0 7840 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2154_
timestamp 1698431365
transform 1 0 5936 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2155_
timestamp 1698431365
transform -1 0 7280 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2156_
timestamp 1698431365
transform 1 0 9968 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2157_
timestamp 1698431365
transform 1 0 13776 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2158_
timestamp 1698431365
transform 1 0 30912 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2159_
timestamp 1698431365
transform 1 0 34048 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2160_
timestamp 1698431365
transform 1 0 33376 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2161_
timestamp 1698431365
transform 1 0 37856 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2162_
timestamp 1698431365
transform 1 0 37184 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2163_
timestamp 1698431365
transform -1 0 45696 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2164_
timestamp 1698431365
transform -1 0 46368 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2165_
timestamp 1698431365
transform 1 0 45808 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2166_
timestamp 1698431365
transform 1 0 50624 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2167_
timestamp 1698431365
transform 1 0 47040 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2168_
timestamp 1698431365
transform -1 0 54768 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2169_
timestamp 1698431365
transform 1 0 49056 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2170_
timestamp 1698431365
transform 1 0 52528 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2171_
timestamp 1698431365
transform -1 0 58352 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2172_
timestamp 1698431365
transform 1 0 55104 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2173_
timestamp 1698431365
transform -1 0 58352 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2174_
timestamp 1698431365
transform 1 0 11760 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2175_
timestamp 1698431365
transform 1 0 17472 0 1 28224
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2176_
timestamp 1698431365
transform -1 0 14000 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2177_
timestamp 1698431365
transform -1 0 13104 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2178_
timestamp 1698431365
transform 1 0 7840 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2179_
timestamp 1698431365
transform 1 0 4816 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2180_
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2181_
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2182_
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2183_
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2184_
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2185_
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2186_
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2187_
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2188_
timestamp 1698431365
transform -1 0 8736 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2189_
timestamp 1698431365
transform -1 0 12656 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2190_
timestamp 1698431365
transform -1 0 11536 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2191_
timestamp 1698431365
transform 1 0 6832 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2192_
timestamp 1698431365
transform -1 0 28896 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2193_
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2194_
timestamp 1698431365
transform 1 0 29120 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2195_
timestamp 1698431365
transform 1 0 29456 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2196_
timestamp 1698431365
transform 1 0 26656 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2197_
timestamp 1698431365
transform 1 0 30912 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2198_
timestamp 1698431365
transform -1 0 14448 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2199_
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2200_
timestamp 1698431365
transform -1 0 20608 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2201_
timestamp 1698431365
transform 1 0 11200 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2202_
timestamp 1698431365
transform 1 0 16128 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2203_
timestamp 1698431365
transform 1 0 44464 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2204_
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2205_
timestamp 1698431365
transform -1 0 51968 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2206_
timestamp 1698431365
transform 1 0 55104 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2207_
timestamp 1698431365
transform 1 0 55104 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2208_
timestamp 1698431365
transform -1 0 58352 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2209_
timestamp 1698431365
transform -1 0 58352 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2210_
timestamp 1698431365
transform -1 0 58352 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2211_
timestamp 1698431365
transform -1 0 56224 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2212_
timestamp 1698431365
transform -1 0 53648 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2213_
timestamp 1698431365
transform -1 0 49504 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2214_
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2215_
timestamp 1698431365
transform -1 0 32256 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2216_
timestamp 1698431365
transform 1 0 44800 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2217_
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2218_
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2219_
timestamp 1698431365
transform 1 0 46480 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2220_
timestamp 1698431365
transform 1 0 55104 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2221_
timestamp 1698431365
transform 1 0 55104 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2222_
timestamp 1698431365
transform 1 0 55104 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2223_
timestamp 1698431365
transform 1 0 55104 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2224_
timestamp 1698431365
transform 1 0 55104 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2225_
timestamp 1698431365
transform 1 0 55104 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2226_
timestamp 1698431365
transform -1 0 54096 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2227_
timestamp 1698431365
transform 1 0 45136 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2228_
timestamp 1698431365
transform -1 0 36288 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2229_
timestamp 1698431365
transform 1 0 22512 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2230_
timestamp 1698431365
transform -1 0 34272 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2231_
timestamp 1698431365
transform -1 0 34384 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2232_
timestamp 1698431365
transform 1 0 22736 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2233_
timestamp 1698431365
transform 1 0 25536 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2234_
timestamp 1698431365
transform -1 0 32256 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2235_
timestamp 1698431365
transform 1 0 17360 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2236_
timestamp 1698431365
transform 1 0 17248 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2237_
timestamp 1698431365
transform 1 0 15232 0 1 48608
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2238_
timestamp 1698431365
transform 1 0 15008 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2239_
timestamp 1698431365
transform 1 0 17696 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2240_
timestamp 1698431365
transform 1 0 21056 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2241_
timestamp 1698431365
transform 1 0 23184 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2242_
timestamp 1698431365
transform -1 0 28336 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2243_
timestamp 1698431365
transform 1 0 19152 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2244_
timestamp 1698431365
transform 1 0 11536 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2245_
timestamp 1698431365
transform 1 0 12320 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2246_
timestamp 1698431365
transform -1 0 20496 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2247_
timestamp 1698431365
transform 1 0 13776 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2248_
timestamp 1698431365
transform 1 0 12880 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2249_
timestamp 1698431365
transform 1 0 13776 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2250_
timestamp 1698431365
transform 1 0 13776 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2251_
timestamp 1698431365
transform 1 0 30464 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2252_
timestamp 1698431365
transform 1 0 31360 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2253_
timestamp 1698431365
transform 1 0 29568 0 1 34496
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2254_
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2255_
timestamp 1698431365
transform 1 0 36960 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2256_
timestamp 1698431365
transform 1 0 35504 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2257_
timestamp 1698431365
transform 1 0 34496 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2258_
timestamp 1698431365
transform 1 0 33376 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2259_
timestamp 1698431365
transform -1 0 40880 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2260_
timestamp 1698431365
transform -1 0 44016 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2261_
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2262_
timestamp 1698431365
transform 1 0 40768 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2263_
timestamp 1698431365
transform 1 0 44016 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2264_
timestamp 1698431365
transform 1 0 15120 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2265_
timestamp 1698431365
transform 1 0 9856 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2266_
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2267_
timestamp 1698431365
transform 1 0 10080 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2268_
timestamp 1698431365
transform -1 0 18032 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2269_
timestamp 1698431365
transform -1 0 20944 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2270_
timestamp 1698431365
transform -1 0 22512 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2271_
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2272_
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2273_
timestamp 1698431365
transform -1 0 31024 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1025__A2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22736 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1034__B1
timestamp 1698431365
transform 1 0 22288 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1038__A1
timestamp 1698431365
transform 1 0 21616 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1038__B1
timestamp 1698431365
transform 1 0 22064 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1040__A3
timestamp 1698431365
transform 1 0 25312 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1043__A2
timestamp 1698431365
transform 1 0 24528 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1047__I
timestamp 1698431365
transform -1 0 38864 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1048__I
timestamp 1698431365
transform 1 0 38976 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1052__I
timestamp 1698431365
transform -1 0 34832 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1053__A3
timestamp 1698431365
transform 1 0 37856 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1053__A4
timestamp 1698431365
transform 1 0 32480 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1057__I
timestamp 1698431365
transform 1 0 26768 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1059__A1
timestamp 1698431365
transform 1 0 38080 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1061__A1
timestamp 1698431365
transform 1 0 39088 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1063__I
timestamp 1698431365
transform 1 0 42336 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1066__I
timestamp 1698431365
transform 1 0 42672 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1069__I
timestamp 1698431365
transform 1 0 43344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1070__A1
timestamp 1698431365
transform -1 0 35056 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1073__I
timestamp 1698431365
transform -1 0 36400 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1074__A1
timestamp 1698431365
transform 1 0 35952 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1080__I
timestamp 1698431365
transform 1 0 37968 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1082__I
timestamp 1698431365
transform -1 0 26432 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1083__A1
timestamp 1698431365
transform 1 0 38192 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1083__A2
timestamp 1698431365
transform 1 0 39984 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1084__A1
timestamp 1698431365
transform -1 0 37744 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1090__A1
timestamp 1698431365
transform 1 0 40432 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1092__I
timestamp 1698431365
transform 1 0 38528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1097__I
timestamp 1698431365
transform 1 0 27216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1098__I
timestamp 1698431365
transform 1 0 36400 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1100__A1
timestamp 1698431365
transform 1 0 28448 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1101__A1
timestamp 1698431365
transform 1 0 26992 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1102__I
timestamp 1698431365
transform -1 0 28336 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1103__I
timestamp 1698431365
transform 1 0 28224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1105__I
timestamp 1698431365
transform 1 0 45584 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1106__A1
timestamp 1698431365
transform 1 0 30128 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1107__A1
timestamp 1698431365
transform 1 0 29680 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1108__I
timestamp 1698431365
transform -1 0 23968 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1111__A1
timestamp 1698431365
transform 1 0 22512 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1112__I
timestamp 1698431365
transform 1 0 44128 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1113__A1
timestamp 1698431365
transform 1 0 29456 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1115__A1
timestamp 1698431365
transform -1 0 22848 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1116__I
timestamp 1698431365
transform 1 0 46816 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1117__A1
timestamp 1698431365
transform -1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1119__A2
timestamp 1698431365
transform 1 0 26768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1119__B
timestamp 1698431365
transform -1 0 28336 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1120__A2
timestamp 1698431365
transform 1 0 26320 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1121__I
timestamp 1698431365
transform 1 0 25312 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1127__A1
timestamp 1698431365
transform 1 0 22288 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1139__A1
timestamp 1698431365
transform 1 0 17024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1153__I
timestamp 1698431365
transform 1 0 12320 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1156__A1
timestamp 1698431365
transform 1 0 12208 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1158__I
timestamp 1698431365
transform 1 0 15568 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1165__A1
timestamp 1698431365
transform 1 0 25424 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1166__A1
timestamp 1698431365
transform -1 0 25536 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1170__A1
timestamp 1698431365
transform 1 0 28560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1172__B
timestamp 1698431365
transform 1 0 26432 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1174__I
timestamp 1698431365
transform 1 0 21392 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1175__I
timestamp 1698431365
transform 1 0 19824 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1176__I
timestamp 1698431365
transform 1 0 20720 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1189__I
timestamp 1698431365
transform -1 0 16352 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1200__A1
timestamp 1698431365
transform 1 0 20272 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1202__B
timestamp 1698431365
transform 1 0 15008 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1216__A1
timestamp 1698431365
transform 1 0 10528 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1222__A2
timestamp 1698431365
transform -1 0 38416 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1223__I
timestamp 1698431365
transform -1 0 42112 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1225__A1
timestamp 1698431365
transform -1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1225__A2
timestamp 1698431365
transform 1 0 42448 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1227__A1
timestamp 1698431365
transform 1 0 40544 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1233__A1
timestamp 1698431365
transform 1 0 43008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1235__I
timestamp 1698431365
transform 1 0 48160 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1237__A1
timestamp 1698431365
transform -1 0 49168 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1239__I
timestamp 1698431365
transform 1 0 53648 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1240__A1
timestamp 1698431365
transform 1 0 53760 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1243__A1
timestamp 1698431365
transform -1 0 56112 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1246__A1
timestamp 1698431365
transform -1 0 56224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1251__A1
timestamp 1698431365
transform 1 0 37408 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1252__A1
timestamp 1698431365
transform 1 0 39312 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1258__A1
timestamp 1698431365
transform 1 0 39760 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1260__I
timestamp 1698431365
transform 1 0 38080 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1263__A1
timestamp 1698431365
transform 1 0 40880 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1265__A1
timestamp 1698431365
transform 1 0 40432 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1267__I
timestamp 1698431365
transform 1 0 42560 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1268__A1
timestamp 1698431365
transform -1 0 42000 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1270__I
timestamp 1698431365
transform 1 0 43232 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1271__A1
timestamp 1698431365
transform -1 0 42448 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1273__I
timestamp 1698431365
transform 1 0 43008 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1274__A1
timestamp 1698431365
transform 1 0 42896 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1278__A1
timestamp 1698431365
transform 1 0 49168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1280__A1
timestamp 1698431365
transform 1 0 54880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1282__A1
timestamp 1698431365
transform 1 0 56000 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1284__A1
timestamp 1698431365
transform 1 0 56672 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1287__A1
timestamp 1698431365
transform 1 0 28784 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1291__C
timestamp 1698431365
transform -1 0 30464 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1300__A2
timestamp 1698431365
transform -1 0 3472 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1301__A2
timestamp 1698431365
transform -1 0 5040 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1308__B
timestamp 1698431365
transform 1 0 4592 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1311__B
timestamp 1698431365
transform 1 0 6608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1315__B
timestamp 1698431365
transform -1 0 6720 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1318__B
timestamp 1698431365
transform -1 0 10752 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1320__I
timestamp 1698431365
transform 1 0 25648 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1323__A1
timestamp 1698431365
transform 1 0 8512 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1328__A1
timestamp 1698431365
transform 1 0 29792 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1329__A1
timestamp 1698431365
transform 1 0 26768 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1331__A1
timestamp 1698431365
transform 1 0 28112 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1332__I
timestamp 1698431365
transform 1 0 44240 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1334__A1
timestamp 1698431365
transform 1 0 27776 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1335__A2
timestamp 1698431365
transform 1 0 30016 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1337__A1
timestamp 1698431365
transform -1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1339__A1
timestamp 1698431365
transform -1 0 25088 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1341__A1
timestamp 1698431365
transform 1 0 25312 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1343__A1
timestamp 1698431365
transform -1 0 27888 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1345__A1
timestamp 1698431365
transform -1 0 26992 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1349__A1
timestamp 1698431365
transform 1 0 33600 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1351__A1
timestamp 1698431365
transform -1 0 31920 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1353__A1
timestamp 1698431365
transform 1 0 33152 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1355__A1
timestamp 1698431365
transform 1 0 31136 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1357__I
timestamp 1698431365
transform 1 0 28336 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1358__I
timestamp 1698431365
transform 1 0 27888 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1359__A1
timestamp 1698431365
transform 1 0 35616 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1362__C
timestamp 1698431365
transform 1 0 26208 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1364__A1
timestamp 1698431365
transform 1 0 9184 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1368__A1
timestamp 1698431365
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1370__A1
timestamp 1698431365
transform -1 0 26432 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1372__A1
timestamp 1698431365
transform 1 0 22960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1374__A1
timestamp 1698431365
transform 1 0 31808 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1376__A1
timestamp 1698431365
transform -1 0 23408 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1378__A1
timestamp 1698431365
transform -1 0 35616 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1380__A1
timestamp 1698431365
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1382__A3
timestamp 1698431365
transform -1 0 39312 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1385__A1
timestamp 1698431365
transform -1 0 48608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1386__A1
timestamp 1698431365
transform 1 0 45360 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1389__A1
timestamp 1698431365
transform 1 0 44800 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1390__A1
timestamp 1698431365
transform -1 0 46032 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1392__A1
timestamp 1698431365
transform 1 0 44912 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1393__A1
timestamp 1698431365
transform 1 0 45360 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1396__A1
timestamp 1698431365
transform 1 0 47152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1397__A1
timestamp 1698431365
transform 1 0 48720 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1398__A1
timestamp 1698431365
transform 1 0 48160 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1399__A1
timestamp 1698431365
transform -1 0 47488 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1400__I
timestamp 1698431365
transform 1 0 51408 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1402__A1
timestamp 1698431365
transform 1 0 51184 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1403__A1
timestamp 1698431365
transform 1 0 52304 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1406__A1
timestamp 1698431365
transform 1 0 54208 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1409__A1
timestamp 1698431365
transform -1 0 55216 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1411__I
timestamp 1698431365
transform -1 0 19712 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1419__A1
timestamp 1698431365
transform 1 0 21168 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1423__A1
timestamp 1698431365
transform -1 0 20496 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1501__A1
timestamp 1698431365
transform -1 0 36064 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1501__A2
timestamp 1698431365
transform -1 0 35616 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1501__B
timestamp 1698431365
transform 1 0 34160 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1503__A1
timestamp 1698431365
transform 1 0 37072 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1503__A2
timestamp 1698431365
transform -1 0 37744 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1503__A3
timestamp 1698431365
transform -1 0 33712 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1505__I
timestamp 1698431365
transform 1 0 40992 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1507__B
timestamp 1698431365
transform 1 0 42672 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1508__A2
timestamp 1698431365
transform 1 0 18592 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1511__A2
timestamp 1698431365
transform 1 0 17472 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1514__A2
timestamp 1698431365
transform -1 0 33824 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1516__A2
timestamp 1698431365
transform 1 0 33712 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1517__I
timestamp 1698431365
transform 1 0 38192 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1520__A2
timestamp 1698431365
transform 1 0 37072 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1522__A1
timestamp 1698431365
transform -1 0 35616 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1525__A1
timestamp 1698431365
transform 1 0 37968 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1526__I
timestamp 1698431365
transform -1 0 42336 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1540__I
timestamp 1698431365
transform 1 0 46144 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1555__C
timestamp 1698431365
transform -1 0 51072 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1566__A1
timestamp 1698431365
transform 1 0 55328 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1576__A1
timestamp 1698431365
transform -1 0 9856 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1579__A1
timestamp 1698431365
transform 1 0 10192 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1582__A1
timestamp 1698431365
transform -1 0 11200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1583__I
timestamp 1698431365
transform -1 0 11760 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1595__I
timestamp 1698431365
transform 1 0 7728 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1610__I
timestamp 1698431365
transform -1 0 7168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1625__I
timestamp 1698431365
transform -1 0 11984 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1639__B
timestamp 1698431365
transform 1 0 10528 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1645__C
timestamp 1698431365
transform 1 0 9632 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1646__A2
timestamp 1698431365
transform 1 0 10192 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1648__B
timestamp 1698431365
transform -1 0 7392 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1663__A1
timestamp 1698431365
transform 1 0 26992 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1664__A1
timestamp 1698431365
transform -1 0 27664 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1665__A1
timestamp 1698431365
transform 1 0 28560 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__A2
timestamp 1698431365
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1669__A3
timestamp 1698431365
transform -1 0 32816 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1671__A2
timestamp 1698431365
transform 1 0 32592 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1681__A1
timestamp 1698431365
transform -1 0 20832 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1681__A2
timestamp 1698431365
transform 1 0 20160 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1682__A1
timestamp 1698431365
transform 1 0 17808 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1684__A1
timestamp 1698431365
transform 1 0 19600 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1686__A1
timestamp 1698431365
transform 1 0 17472 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__A1
timestamp 1698431365
transform 1 0 20048 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__A2
timestamp 1698431365
transform 1 0 19600 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1691__A2
timestamp 1698431365
transform -1 0 44800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1740__A1
timestamp 1698431365
transform 1 0 42784 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1740__B
timestamp 1698431365
transform 1 0 42560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1742__A2
timestamp 1698431365
transform 1 0 45696 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1745__I
timestamp 1698431365
transform 1 0 39760 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1747__A1
timestamp 1698431365
transform 1 0 45248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1750__A1
timestamp 1698431365
transform 1 0 49728 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1753__A4
timestamp 1698431365
transform 1 0 46928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1756__A1
timestamp 1698431365
transform 1 0 52752 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1759__A1
timestamp 1698431365
transform 1 0 53984 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1762__A1
timestamp 1698431365
transform 1 0 38640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1762__A2
timestamp 1698431365
transform 1 0 39088 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1766__A1
timestamp 1698431365
transform 1 0 54992 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1766__A2
timestamp 1698431365
transform 1 0 54432 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1768__I
timestamp 1698431365
transform 1 0 36960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1771__A1
timestamp 1698431365
transform 1 0 52304 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1771__A2
timestamp 1698431365
transform 1 0 54880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1774__A1
timestamp 1698431365
transform -1 0 54656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1778__A1
timestamp 1698431365
transform -1 0 52976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1778__A2
timestamp 1698431365
transform -1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1782__A1
timestamp 1698431365
transform 1 0 49616 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1785__A1
timestamp 1698431365
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1788__A1
timestamp 1698431365
transform 1 0 43568 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1788__A2
timestamp 1698431365
transform 1 0 42672 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1788__C
timestamp 1698431365
transform 1 0 42224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__A1
timestamp 1698431365
transform 1 0 32480 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__A2
timestamp 1698431365
transform 1 0 32480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1790__A2
timestamp 1698431365
transform 1 0 32480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1790__A3
timestamp 1698431365
transform 1 0 33152 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1791__B
timestamp 1698431365
transform 1 0 32704 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1793__A2
timestamp 1698431365
transform 1 0 42896 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1848__B
timestamp 1698431365
transform -1 0 37520 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1853__A3
timestamp 1698431365
transform 1 0 45024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1854__A2
timestamp 1698431365
transform 1 0 43792 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1856__A4
timestamp 1698431365
transform 1 0 46592 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1862__A1
timestamp 1698431365
transform 1 0 47264 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1865__A1
timestamp 1698431365
transform 1 0 54544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1871__A1
timestamp 1698431365
transform 1 0 55216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1884__B
timestamp 1698431365
transform -1 0 47488 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1887__A1
timestamp 1698431365
transform -1 0 36848 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1889__A2
timestamp 1698431365
transform 1 0 30128 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1920__C
timestamp 1698431365
transform 1 0 27776 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1921__A1
timestamp 1698431365
transform -1 0 26544 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1922__I
timestamp 1698431365
transform -1 0 24640 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1925__I
timestamp 1698431365
transform 1 0 25760 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1926__A3
timestamp 1698431365
transform -1 0 32480 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1927__A2
timestamp 1698431365
transform 1 0 33152 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1930__A4
timestamp 1698431365
transform -1 0 32032 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1933__I
timestamp 1698431365
transform -1 0 22848 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1957__B
timestamp 1698431365
transform 1 0 26208 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1960__A1
timestamp 1698431365
transform 1 0 27552 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1962__A1
timestamp 1698431365
transform -1 0 27328 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1964__A1
timestamp 1698431365
transform -1 0 27440 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1968__B
timestamp 1698431365
transform 1 0 14224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1972__A1
timestamp 1698431365
transform -1 0 15792 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1984__A1
timestamp 1698431365
transform -1 0 16800 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1985__A4
timestamp 1698431365
transform 1 0 58128 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1986__A1
timestamp 1698431365
transform 1 0 38528 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1986__A2
timestamp 1698431365
transform 1 0 39200 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1986__A3
timestamp 1698431365
transform -1 0 37856 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1988__A1
timestamp 1698431365
transform 1 0 34496 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1988__A2
timestamp 1698431365
transform 1 0 34496 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1990__B
timestamp 1698431365
transform 1 0 31248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1992__A1
timestamp 1698431365
transform 1 0 33936 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1992__B
timestamp 1698431365
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1994__A1
timestamp 1698431365
transform 1 0 33152 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1994__B
timestamp 1698431365
transform -1 0 31920 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1996__A1
timestamp 1698431365
transform 1 0 36288 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1996__B
timestamp 1698431365
transform 1 0 34944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1998__A1
timestamp 1698431365
transform 1 0 37520 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1998__B
timestamp 1698431365
transform 1 0 35280 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2002__A1
timestamp 1698431365
transform 1 0 40320 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2004__A1
timestamp 1698431365
transform 1 0 37184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2006__A1
timestamp 1698431365
transform 1 0 38976 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2008__A1
timestamp 1698431365
transform -1 0 38752 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2010__A1
timestamp 1698431365
transform 1 0 39760 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2014__A1
timestamp 1698431365
transform -1 0 43232 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2016__A1
timestamp 1698431365
transform -1 0 44576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2018__A1
timestamp 1698431365
transform 1 0 43232 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2020__A1
timestamp 1698431365
transform 1 0 44240 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2039__B
timestamp 1698431365
transform -1 0 20608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2043__A1
timestamp 1698431365
transform 1 0 21392 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2047__A1
timestamp 1698431365
transform 1 0 32144 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2049__A1
timestamp 1698431365
transform -1 0 32256 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2194__CLK
timestamp 1698431365
transform 1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 30016 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_0__f_wb_clk_i_I
timestamp 1698431365
transform -1 0 22064 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_1__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 21392 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_2__f_wb_clk_i_I
timestamp 1698431365
transform -1 0 45136 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_3__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 44688 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 9856 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_1_wb_clk_i_I
timestamp 1698431365
transform 1 0 19152 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_2_wb_clk_i_I
timestamp 1698431365
transform 1 0 18032 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_3_wb_clk_i_I
timestamp 1698431365
transform -1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_4_wb_clk_i_I
timestamp 1698431365
transform 1 0 19152 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_5_wb_clk_i_I
timestamp 1698431365
transform 1 0 9632 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_6_wb_clk_i_I
timestamp 1698431365
transform 1 0 9632 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_7_wb_clk_i_I
timestamp 1698431365
transform 1 0 16352 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_8_wb_clk_i_I
timestamp 1698431365
transform 1 0 11312 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_9_wb_clk_i_I
timestamp 1698431365
transform 1 0 19600 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_10_wb_clk_i_I
timestamp 1698431365
transform 1 0 18704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_11_wb_clk_i_I
timestamp 1698431365
transform 1 0 19040 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_12_wb_clk_i_I
timestamp 1698431365
transform -1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_13_wb_clk_i_I
timestamp 1698431365
transform 1 0 25312 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_14_wb_clk_i_I
timestamp 1698431365
transform -1 0 29792 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_15_wb_clk_i_I
timestamp 1698431365
transform 1 0 43344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_16_wb_clk_i_I
timestamp 1698431365
transform 1 0 40544 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_17_wb_clk_i_I
timestamp 1698431365
transform 1 0 37072 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_18_wb_clk_i_I
timestamp 1698431365
transform 1 0 40768 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_19_wb_clk_i_I
timestamp 1698431365
transform 1 0 51072 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_20_wb_clk_i_I
timestamp 1698431365
transform -1 0 48384 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_21_wb_clk_i_I
timestamp 1698431365
transform 1 0 52528 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_22_wb_clk_i_I
timestamp 1698431365
transform 1 0 50512 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_23_wb_clk_i_I
timestamp 1698431365
transform 1 0 51856 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_24_wb_clk_i_I
timestamp 1698431365
transform 1 0 52080 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_25_wb_clk_i_I
timestamp 1698431365
transform 1 0 48384 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_26_wb_clk_i_I
timestamp 1698431365
transform 1 0 50512 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_27_wb_clk_i_I
timestamp 1698431365
transform -1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_28_wb_clk_i_I
timestamp 1698431365
transform 1 0 46592 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_29_wb_clk_i_I
timestamp 1698431365
transform 1 0 50848 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_30_wb_clk_i_I
timestamp 1698431365
transform 1 0 52080 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_31_wb_clk_i_I
timestamp 1698431365
transform 1 0 52080 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_32_wb_clk_i_I
timestamp 1698431365
transform 1 0 52080 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_33_wb_clk_i_I
timestamp 1698431365
transform 1 0 52080 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_34_wb_clk_i_I
timestamp 1698431365
transform -1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_35_wb_clk_i_I
timestamp 1698431365
transform 1 0 50512 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_36_wb_clk_i_I
timestamp 1698431365
transform 1 0 46816 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_37_wb_clk_i_I
timestamp 1698431365
transform 1 0 47152 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_38_wb_clk_i_I
timestamp 1698431365
transform 1 0 43120 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_39_wb_clk_i_I
timestamp 1698431365
transform 1 0 39872 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_40_wb_clk_i_I
timestamp 1698431365
transform 1 0 45920 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_41_wb_clk_i_I
timestamp 1698431365
transform 1 0 40208 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_42_wb_clk_i_I
timestamp 1698431365
transform 1 0 28560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_44_wb_clk_i_I
timestamp 1698431365
transform 1 0 21728 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_45_wb_clk_i_I
timestamp 1698431365
transform 1 0 26880 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_46_wb_clk_i_I
timestamp 1698431365
transform -1 0 27552 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_47_wb_clk_i_I
timestamp 1698431365
transform 1 0 19040 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_48_wb_clk_i_I
timestamp 1698431365
transform 1 0 18144 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_49_wb_clk_i_I
timestamp 1698431365
transform 1 0 18480 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_50_wb_clk_i_I
timestamp 1698431365
transform 1 0 16800 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_51_wb_clk_i_I
timestamp 1698431365
transform 1 0 9296 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_52_wb_clk_i_I
timestamp 1698431365
transform 1 0 15232 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_53_wb_clk_i_I
timestamp 1698431365
transform 1 0 8848 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 57456 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 57680 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 57680 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 57680 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 57680 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 57680 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 57680 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 57456 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 57680 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform 1 0 58128 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform -1 0 37520 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform -1 0 52528 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform -1 0 22512 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output19_I
timestamp 1698431365
transform -1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output20_I
timestamp 1698431365
transform 1 0 48832 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30464 0 1 29792
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_wb_clk_i
timestamp 1698431365
transform -1 0 20944 0 1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_wb_clk_i
timestamp 1698431365
transform -1 0 20944 0 1 42336
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_wb_clk_i
timestamp 1698431365
transform 1 0 45136 0 1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_wb_clk_i
timestamp 1698431365
transform 1 0 44688 0 1 43904
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_0_wb_clk_i
timestamp 1698431365
transform 1 0 3584 0 -1 26656
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_1_wb_clk_i
timestamp 1698431365
transform -1 0 18928 0 1 25088
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_2_wb_clk_i
timestamp 1698431365
transform -1 0 23856 0 -1 25088
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_3_wb_clk_i
timestamp 1698431365
transform -1 0 26768 0 1 32928
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_4_wb_clk_i
timestamp 1698431365
transform -1 0 18928 0 1 34496
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_5_wb_clk_i
timestamp 1698431365
transform -1 0 8400 0 -1 34496
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_6_wb_clk_i
timestamp 1698431365
transform 1 0 3584 0 -1 40768
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_7_wb_clk_i
timestamp 1698431365
transform -1 0 15232 0 -1 43904
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_8_wb_clk_i
timestamp 1698431365
transform -1 0 11088 0 1 47040
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_9_wb_clk_i
timestamp 1698431365
transform -1 0 19600 0 1 50176
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_10_wb_clk_i
timestamp 1698431365
transform -1 0 24528 0 -1 47040
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_11_wb_clk_i
timestamp 1698431365
transform -1 0 24864 0 -1 53312
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_12_wb_clk_i
timestamp 1698431365
transform -1 0 30688 0 -1 54880
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_13_wb_clk_i
timestamp 1698431365
transform -1 0 30688 0 -1 40768
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_14_wb_clk_i
timestamp 1698431365
transform 1 0 29792 0 1 32928
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_15_wb_clk_i
timestamp 1698431365
transform -1 0 43344 0 1 40768
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_16_wb_clk_i
timestamp 1698431365
transform 1 0 34944 0 -1 45472
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_17_wb_clk_i
timestamp 1698431365
transform -1 0 36400 0 1 45472
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_18_wb_clk_i
timestamp 1698431365
transform -1 0 40432 0 -1 53312
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_19_wb_clk_i
timestamp 1698431365
transform -1 0 50848 0 1 47040
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_20_wb_clk_i
timestamp 1698431365
transform -1 0 54208 0 -1 54880
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_21_wb_clk_i
timestamp 1698431365
transform 1 0 52752 0 1 50176
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_22_wb_clk_i
timestamp 1698431365
transform 1 0 50624 0 -1 45472
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_23_wb_clk_i
timestamp 1698431365
transform 1 0 52528 0 1 40768
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_24_wb_clk_i
timestamp 1698431365
transform 1 0 52752 0 1 34496
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_25_wb_clk_i
timestamp 1698431365
transform -1 0 54208 0 -1 36064
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_26_wb_clk_i
timestamp 1698431365
transform -1 0 50288 0 1 37632
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_27_wb_clk_i
timestamp 1698431365
transform -1 0 44016 0 1 31360
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_28_wb_clk_i
timestamp 1698431365
transform -1 0 46368 0 -1 26656
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_29_wb_clk_i
timestamp 1698431365
transform -1 0 50624 0 1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_30_wb_clk_i
timestamp 1698431365
transform 1 0 52752 0 1 26656
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_31_wb_clk_i
timestamp 1698431365
transform 1 0 52752 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_32_wb_clk_i
timestamp 1698431365
transform 1 0 52752 0 1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_33_wb_clk_i
timestamp 1698431365
transform 1 0 52752 0 1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_34_wb_clk_i
timestamp 1698431365
transform 1 0 52528 0 1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_35_wb_clk_i
timestamp 1698431365
transform -1 0 50288 0 1 14112
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_36_wb_clk_i
timestamp 1698431365
transform -1 0 46592 0 -1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_37_wb_clk_i
timestamp 1698431365
transform -1 0 46368 0 -1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_38_wb_clk_i
timestamp 1698431365
transform -1 0 42448 0 1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_39_wb_clk_i
timestamp 1698431365
transform -1 0 39872 0 -1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_40_wb_clk_i
timestamp 1698431365
transform -1 0 46368 0 -1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_41_wb_clk_i
timestamp 1698431365
transform -1 0 39984 0 -1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_42_wb_clk_i
timestamp 1698431365
transform 1 0 29232 0 1 25088
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_44_wb_clk_i
timestamp 1698431365
transform -1 0 27552 0 1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_45_wb_clk_i
timestamp 1698431365
transform 1 0 27104 0 -1 14112
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_46_wb_clk_i
timestamp 1698431365
transform 1 0 26992 0 -1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_47_wb_clk_i
timestamp 1698431365
transform -1 0 24864 0 -1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_48_wb_clk_i
timestamp 1698431365
transform -1 0 23968 0 -1 14112
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_49_wb_clk_i
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_50_wb_clk_i
timestamp 1698431365
transform -1 0 15904 0 -1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_51_wb_clk_i
timestamp 1698431365
transform -1 0 8960 0 -1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_52_wb_clk_i
timestamp 1698431365
transform -1 0 15008 0 -1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_53_wb_clk_i
timestamp 1698431365
transform -1 0 8624 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_10 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_12 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2688 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_17 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3248 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_33
timestamp 1698431365
transform 1 0 5040 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_40
timestamp 1698431365
transform 1 0 5824 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_48
timestamp 1698431365
transform 1 0 6720 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_53
timestamp 1698431365
transform 1 0 7280 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_61 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8176 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_65
timestamp 1698431365
transform 1 0 8624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_67
timestamp 1698431365
transform 1 0 8848 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_74
timestamp 1698431365
transform 1 0 9632 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_82
timestamp 1698431365
transform 1 0 10528 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_84
timestamp 1698431365
transform 1 0 10752 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_89
timestamp 1698431365
transform 1 0 11312 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_97
timestamp 1698431365
transform 1 0 12208 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_101
timestamp 1698431365
transform 1 0 12656 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_108
timestamp 1698431365
transform 1 0 13440 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_116
timestamp 1698431365
transform 1 0 14336 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_120
timestamp 1698431365
transform 1 0 14784 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_125
timestamp 1698431365
transform 1 0 15344 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_133
timestamp 1698431365
transform 1 0 16240 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_135
timestamp 1698431365
transform 1 0 16464 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_143
timestamp 1698431365
transform 1 0 17360 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_174
timestamp 1698431365
transform 1 0 20832 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698431365
transform 1 0 23856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698431365
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_210
timestamp 1698431365
transform 1 0 24864 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_237
timestamp 1698431365
transform 1 0 27888 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_244
timestamp 1698431365
transform 1 0 28672 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_246
timestamp 1698431365
transform 1 0 28896 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_251
timestamp 1698431365
transform 1 0 29456 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_259
timestamp 1698431365
transform 1 0 30352 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_263
timestamp 1698431365
transform 1 0 30800 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_269
timestamp 1698431365
transform 1 0 31472 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_271
timestamp 1698431365
transform 1 0 31696 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_282
timestamp 1698431365
transform 1 0 32928 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_287
timestamp 1698431365
transform 1 0 33488 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_295
timestamp 1698431365
transform 1 0 34384 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_299
timestamp 1698431365
transform 1 0 34832 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_305
timestamp 1698431365
transform 1 0 35504 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_308
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_312
timestamp 1698431365
transform 1 0 36288 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_368
timestamp 1698431365
transform 1 0 42560 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_405
timestamp 1698431365
transform 1 0 46704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_407
timestamp 1698431365
transform 1 0 46928 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_440
timestamp 1698431365
transform 1 0 50624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_444
timestamp 1698431365
transform 1 0 51072 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_449
timestamp 1698431365
transform 1 0 51632 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_457
timestamp 1698431365
transform 1 0 52528 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_461
timestamp 1698431365
transform 1 0 52976 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_467
timestamp 1698431365
transform 1 0 53648 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_475
timestamp 1698431365
transform 1 0 54544 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_478
timestamp 1698431365
transform 1 0 54880 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_480
timestamp 1698431365
transform 1 0 55104 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_485
timestamp 1698431365
transform 1 0 55664 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_493
timestamp 1698431365
transform 1 0 56560 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_497
timestamp 1698431365
transform 1 0 57008 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_503
timestamp 1698431365
transform 1 0 57680 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_507
timestamp 1698431365
transform 1 0 58128 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_76
timestamp 1698431365
transform 1 0 9856 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_106
timestamp 1698431365
transform 1 0 13216 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_139
timestamp 1698431365
transform 1 0 16912 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_175
timestamp 1698431365
transform 1 0 20944 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698431365
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_241
timestamp 1698431365
transform 1 0 28336 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_245
timestamp 1698431365
transform 1 0 28784 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_247
timestamp 1698431365
transform 1 0 29008 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_277
timestamp 1698431365
transform 1 0 32368 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698431365
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_287
timestamp 1698431365
transform 1 0 33488 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_291
timestamp 1698431365
transform 1 0 33936 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_299
timestamp 1698431365
transform 1 0 34832 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_307
timestamp 1698431365
transform 1 0 35728 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_338
timestamp 1698431365
transform 1 0 39200 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_346
timestamp 1698431365
transform 1 0 40096 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_352
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_409
timestamp 1698431365
transform 1 0 47152 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_422
timestamp 1698431365
transform 1 0 48608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_426
timestamp 1698431365
transform 1 0 49056 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_434
timestamp 1698431365
transform 1 0 49952 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_473
timestamp 1698431365
transform 1 0 54320 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_489
timestamp 1698431365
transform 1 0 56112 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_492
timestamp 1698431365
transform 1 0 56448 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_500
timestamp 1698431365
transform 1 0 57344 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_104
timestamp 1698431365
transform 1 0 12992 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_123
timestamp 1698431365
transform 1 0 15120 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_127
timestamp 1698431365
transform 1 0 15568 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_135
timestamp 1698431365
transform 1 0 16464 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_143
timestamp 1698431365
transform 1 0 17360 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_147
timestamp 1698431365
transform 1 0 17808 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_164
timestamp 1698431365
transform 1 0 19712 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_168
timestamp 1698431365
transform 1 0 20160 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_219
timestamp 1698431365
transform 1 0 25872 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_221
timestamp 1698431365
transform 1 0 26096 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_230
timestamp 1698431365
transform 1 0 27104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_234
timestamp 1698431365
transform 1 0 27552 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_242
timestamp 1698431365
transform 1 0 28448 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_244
timestamp 1698431365
transform 1 0 28672 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_251
timestamp 1698431365
transform 1 0 29456 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_264
timestamp 1698431365
transform 1 0 30912 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_274
timestamp 1698431365
transform 1 0 32032 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_282
timestamp 1698431365
transform 1 0 32928 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_325
timestamp 1698431365
transform 1 0 37744 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_329
timestamp 1698431365
transform 1 0 38192 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_391
timestamp 1698431365
transform 1 0 45136 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_430
timestamp 1698431365
transform 1 0 49504 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_438
timestamp 1698431365
transform 1 0 50400 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_448
timestamp 1698431365
transform 1 0 51520 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_452
timestamp 1698431365
transform 1 0 51968 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_507
timestamp 1698431365
transform 1 0 58128 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_34
timestamp 1698431365
transform 1 0 5152 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_50
timestamp 1698431365
transform 1 0 6944 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_54
timestamp 1698431365
transform 1 0 7392 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_62
timestamp 1698431365
transform 1 0 8288 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_151
timestamp 1698431365
transform 1 0 18256 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_167
timestamp 1698431365
transform 1 0 20048 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_175
timestamp 1698431365
transform 1 0 20944 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_183
timestamp 1698431365
transform 1 0 21840 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_191
timestamp 1698431365
transform 1 0 22736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_195
timestamp 1698431365
transform 1 0 23184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_203
timestamp 1698431365
transform 1 0 24080 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_208
timestamp 1698431365
transform 1 0 24640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_222
timestamp 1698431365
transform 1 0 26208 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_279
timestamp 1698431365
transform 1 0 32592 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_286
timestamp 1698431365
transform 1 0 33376 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_288
timestamp 1698431365
transform 1 0 33600 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_305
timestamp 1698431365
transform 1 0 35504 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_418
timestamp 1698431365
transform 1 0 48160 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_422
timestamp 1698431365
transform 1 0 48608 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_430
timestamp 1698431365
transform 1 0 49504 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_443
timestamp 1698431365
transform 1 0 50960 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_459
timestamp 1698431365
transform 1 0 52752 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_492
timestamp 1698431365
transform 1 0 56448 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_508
timestamp 1698431365
transform 1 0 58240 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_39
timestamp 1698431365
transform 1 0 5712 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_69
timestamp 1698431365
transform 1 0 9072 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_145
timestamp 1698431365
transform 1 0 17584 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_153
timestamp 1698431365
transform 1 0 18480 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_157
timestamp 1698431365
transform 1 0 18928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_168
timestamp 1698431365
transform 1 0 20160 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_172
timestamp 1698431365
transform 1 0 20608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_174
timestamp 1698431365
transform 1 0 20832 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_179
timestamp 1698431365
transform 1 0 21392 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_186
timestamp 1698431365
transform 1 0 22176 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_197
timestamp 1698431365
transform 1 0 23408 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_201
timestamp 1698431365
transform 1 0 23856 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_231
timestamp 1698431365
transform 1 0 27216 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_239
timestamp 1698431365
transform 1 0 28112 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_243
timestamp 1698431365
transform 1 0 28560 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_276
timestamp 1698431365
transform 1 0 32256 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_280
timestamp 1698431365
transform 1 0 32704 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_282
timestamp 1698431365
transform 1 0 32928 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_296
timestamp 1698431365
transform 1 0 34496 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_298
timestamp 1698431365
transform 1 0 34720 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_305
timestamp 1698431365
transform 1 0 35504 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_307
timestamp 1698431365
transform 1 0 35728 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_313
timestamp 1698431365
transform 1 0 36400 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_382
timestamp 1698431365
transform 1 0 44128 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_384
timestamp 1698431365
transform 1 0 44352 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_387
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_389
timestamp 1698431365
transform 1 0 44912 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_407
timestamp 1698431365
transform 1 0 46928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_411
timestamp 1698431365
transform 1 0 47376 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_419
timestamp 1698431365
transform 1 0 48272 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_423
timestamp 1698431365
transform 1 0 48720 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_446
timestamp 1698431365
transform 1 0 51296 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_450
timestamp 1698431365
transform 1 0 51744 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_452
timestamp 1698431365
transform 1 0 51968 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_457
timestamp 1698431365
transform 1 0 52528 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_471
timestamp 1698431365
transform 1 0 54096 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_473
timestamp 1698431365
transform 1 0 54320 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_476
timestamp 1698431365
transform 1 0 54656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_34
timestamp 1698431365
transform 1 0 5152 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_50
timestamp 1698431365
transform 1 0 6944 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_63
timestamp 1698431365
transform 1 0 8400 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_67
timestamp 1698431365
transform 1 0 8848 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_69
timestamp 1698431365
transform 1 0 9072 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_82
timestamp 1698431365
transform 1 0 10528 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_86
timestamp 1698431365
transform 1 0 10976 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_116
timestamp 1698431365
transform 1 0 14336 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_132
timestamp 1698431365
transform 1 0 16128 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_216
timestamp 1698431365
transform 1 0 25536 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_237
timestamp 1698431365
transform 1 0 27888 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_245
timestamp 1698431365
transform 1 0 28784 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_275
timestamp 1698431365
transform 1 0 32144 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_279
timestamp 1698431365
transform 1 0 32592 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_290
timestamp 1698431365
transform 1 0 33824 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_294
timestamp 1698431365
transform 1 0 34272 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_304
timestamp 1698431365
transform 1 0 35392 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_308
timestamp 1698431365
transform 1 0 35840 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_324
timestamp 1698431365
transform 1 0 37632 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_332
timestamp 1698431365
transform 1 0 38528 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_349
timestamp 1698431365
transform 1 0 40432 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_361
timestamp 1698431365
transform 1 0 41776 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_367
timestamp 1698431365
transform 1 0 42448 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_371
timestamp 1698431365
transform 1 0 42896 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_375
timestamp 1698431365
transform 1 0 43344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_379
timestamp 1698431365
transform 1 0 43792 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_395
timestamp 1698431365
transform 1 0 45584 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_412
timestamp 1698431365
transform 1 0 47488 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_422
timestamp 1698431365
transform 1 0 48608 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_430
timestamp 1698431365
transform 1 0 49504 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_437
timestamp 1698431365
transform 1 0 50288 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_453
timestamp 1698431365
transform 1 0 52080 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_475
timestamp 1698431365
transform 1 0 54544 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_484
timestamp 1698431365
transform 1 0 55552 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_488
timestamp 1698431365
transform 1 0 56000 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_498
timestamp 1698431365
transform 1 0 57120 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_506
timestamp 1698431365
transform 1 0 58016 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_508
timestamp 1698431365
transform 1 0 58240 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_53
timestamp 1698431365
transform 1 0 7280 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_61
timestamp 1698431365
transform 1 0 8176 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_63
timestamp 1698431365
transform 1 0 8400 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_75
timestamp 1698431365
transform 1 0 9744 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_91
timestamp 1698431365
transform 1 0 11536 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_99
timestamp 1698431365
transform 1 0 12432 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_103
timestamp 1698431365
transform 1 0 12880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_139
timestamp 1698431365
transform 1 0 16912 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_170
timestamp 1698431365
transform 1 0 20384 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_174
timestamp 1698431365
transform 1 0 20832 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_212
timestamp 1698431365
transform 1 0 25088 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_214
timestamp 1698431365
transform 1 0 25312 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_221
timestamp 1698431365
transform 1 0 26096 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_223
timestamp 1698431365
transform 1 0 26320 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_226
timestamp 1698431365
transform 1 0 26656 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_242
timestamp 1698431365
transform 1 0 28448 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_244
timestamp 1698431365
transform 1 0 28672 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_255
timestamp 1698431365
transform 1 0 29904 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_263
timestamp 1698431365
transform 1 0 30800 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_279
timestamp 1698431365
transform 1 0 32592 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_287
timestamp 1698431365
transform 1 0 33488 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_303
timestamp 1698431365
transform 1 0 35280 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698431365
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_325
timestamp 1698431365
transform 1 0 37744 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_330
timestamp 1698431365
transform 1 0 38304 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_346
timestamp 1698431365
transform 1 0 40096 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_348
timestamp 1698431365
transform 1 0 40320 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_351
timestamp 1698431365
transform 1 0 40656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_355
timestamp 1698431365
transform 1 0 41104 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_387
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_403
timestamp 1698431365
transform 1 0 46480 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_416
timestamp 1698431365
transform 1 0 47936 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_424
timestamp 1698431365
transform 1 0 48832 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_428
timestamp 1698431365
transform 1 0 49280 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_439
timestamp 1698431365
transform 1 0 50512 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_457
timestamp 1698431365
transform 1 0 52528 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_476
timestamp 1698431365
transform 1 0 54656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_34
timestamp 1698431365
transform 1 0 5152 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_38
timestamp 1698431365
transform 1 0 5600 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_46
timestamp 1698431365
transform 1 0 6496 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_50
timestamp 1698431365
transform 1 0 6944 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_56
timestamp 1698431365
transform 1 0 7616 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_60
timestamp 1698431365
transform 1 0 8064 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_80
timestamp 1698431365
transform 1 0 10304 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_84
timestamp 1698431365
transform 1 0 10752 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_92
timestamp 1698431365
transform 1 0 11648 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_96
timestamp 1698431365
transform 1 0 12096 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_105
timestamp 1698431365
transform 1 0 13104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_125
timestamp 1698431365
transform 1 0 15344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_129
timestamp 1698431365
transform 1 0 15792 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_131
timestamp 1698431365
transform 1 0 16016 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_177
timestamp 1698431365
transform 1 0 21168 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_209
timestamp 1698431365
transform 1 0 24752 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_214
timestamp 1698431365
transform 1 0 25312 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_217
timestamp 1698431365
transform 1 0 25648 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_233
timestamp 1698431365
transform 1 0 27440 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_241
timestamp 1698431365
transform 1 0 28336 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_252
timestamp 1698431365
transform 1 0 29568 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_256
timestamp 1698431365
transform 1 0 30016 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_260
timestamp 1698431365
transform 1 0 30464 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698431365
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_342
timestamp 1698431365
transform 1 0 39648 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_344
timestamp 1698431365
transform 1 0 39872 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_349
timestamp 1698431365
transform 1 0 40432 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_352
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_354
timestamp 1698431365
transform 1 0 40992 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_359
timestamp 1698431365
transform 1 0 41552 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_367
timestamp 1698431365
transform 1 0 42448 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_369
timestamp 1698431365
transform 1 0 42672 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_403
timestamp 1698431365
transform 1 0 46480 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_411
timestamp 1698431365
transform 1 0 47376 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_415
timestamp 1698431365
transform 1 0 47824 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_436
timestamp 1698431365
transform 1 0 50176 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_440
timestamp 1698431365
transform 1 0 50624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_451
timestamp 1698431365
transform 1 0 51856 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_485
timestamp 1698431365
transform 1 0 55664 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_489
timestamp 1698431365
transform 1 0 56112 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_498
timestamp 1698431365
transform 1 0 57120 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_500
timestamp 1698431365
transform 1 0 57344 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_45
timestamp 1698431365
transform 1 0 6384 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_81
timestamp 1698431365
transform 1 0 10416 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_97
timestamp 1698431365
transform 1 0 12208 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_163
timestamp 1698431365
transform 1 0 19600 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_171
timestamp 1698431365
transform 1 0 20496 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_181
timestamp 1698431365
transform 1 0 21616 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_188
timestamp 1698431365
transform 1 0 22400 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_220
timestamp 1698431365
transform 1 0 25984 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_231
timestamp 1698431365
transform 1 0 27216 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_241
timestamp 1698431365
transform 1 0 28336 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_251
timestamp 1698431365
transform 1 0 29456 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_270
timestamp 1698431365
transform 1 0 31584 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_286
timestamp 1698431365
transform 1 0 33376 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_290
timestamp 1698431365
transform 1 0 33824 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_296
timestamp 1698431365
transform 1 0 34496 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_312
timestamp 1698431365
transform 1 0 36288 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_314
timestamp 1698431365
transform 1 0 36512 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_321
timestamp 1698431365
transform 1 0 37296 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_325
timestamp 1698431365
transform 1 0 37744 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_344
timestamp 1698431365
transform 1 0 39872 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_348
timestamp 1698431365
transform 1 0 40320 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_350
timestamp 1698431365
transform 1 0 40544 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_360
timestamp 1698431365
transform 1 0 41664 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_370
timestamp 1698431365
transform 1 0 42784 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_378
timestamp 1698431365
transform 1 0 43680 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_382
timestamp 1698431365
transform 1 0 44128 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_384
timestamp 1698431365
transform 1 0 44352 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_387
timestamp 1698431365
transform 1 0 44688 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_403
timestamp 1698431365
transform 1 0 46480 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_407
timestamp 1698431365
transform 1 0 46928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_440
timestamp 1698431365
transform 1 0 50624 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_448
timestamp 1698431365
transform 1 0 51520 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_452
timestamp 1698431365
transform 1 0 51968 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_457
timestamp 1698431365
transform 1 0 52528 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_18
timestamp 1698431365
transform 1 0 3360 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_22
timestamp 1698431365
transform 1 0 3808 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_32
timestamp 1698431365
transform 1 0 4928 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_44
timestamp 1698431365
transform 1 0 6272 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_48
timestamp 1698431365
transform 1 0 6720 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_64
timestamp 1698431365
transform 1 0 8512 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_68
timestamp 1698431365
transform 1 0 8960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_104
timestamp 1698431365
transform 1 0 12992 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_129
timestamp 1698431365
transform 1 0 15792 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_137
timestamp 1698431365
transform 1 0 16688 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_139
timestamp 1698431365
transform 1 0 16912 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_150
timestamp 1698431365
transform 1 0 18144 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_152
timestamp 1698431365
transform 1 0 18368 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_184
timestamp 1698431365
transform 1 0 21952 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_186
timestamp 1698431365
transform 1 0 22176 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_205
timestamp 1698431365
transform 1 0 24304 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_209
timestamp 1698431365
transform 1 0 24752 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_242
timestamp 1698431365
transform 1 0 28448 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_246
timestamp 1698431365
transform 1 0 28896 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_248
timestamp 1698431365
transform 1 0 29120 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_278
timestamp 1698431365
transform 1 0 32480 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_290
timestamp 1698431365
transform 1 0 33824 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_325
timestamp 1698431365
transform 1 0 37744 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_331
timestamp 1698431365
transform 1 0 38416 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_343
timestamp 1698431365
transform 1 0 39760 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_347
timestamp 1698431365
transform 1 0 40208 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_349
timestamp 1698431365
transform 1 0 40432 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_404
timestamp 1698431365
transform 1 0 46592 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_418
timestamp 1698431365
transform 1 0 48160 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_426
timestamp 1698431365
transform 1 0 49056 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_430
timestamp 1698431365
transform 1 0 49504 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_439
timestamp 1698431365
transform 1 0 50512 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_455
timestamp 1698431365
transform 1 0 52304 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_463
timestamp 1698431365
transform 1 0 53200 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_470
timestamp 1698431365
transform 1 0 53984 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_486
timestamp 1698431365
transform 1 0 55776 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_492
timestamp 1698431365
transform 1 0 56448 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_508
timestamp 1698431365
transform 1 0 58240 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_31
timestamp 1698431365
transform 1 0 4816 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_45
timestamp 1698431365
transform 1 0 6384 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_49
timestamp 1698431365
transform 1 0 6832 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_57
timestamp 1698431365
transform 1 0 7728 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_69
timestamp 1698431365
transform 1 0 9072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_73
timestamp 1698431365
transform 1 0 9520 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_75
timestamp 1698431365
transform 1 0 9744 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_120
timestamp 1698431365
transform 1 0 14784 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_153
timestamp 1698431365
transform 1 0 18480 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_169
timestamp 1698431365
transform 1 0 20272 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_173
timestamp 1698431365
transform 1 0 20720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_206
timestamp 1698431365
transform 1 0 24416 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_215
timestamp 1698431365
transform 1 0 25424 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_219
timestamp 1698431365
transform 1 0 25872 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_227
timestamp 1698431365
transform 1 0 26768 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_243
timestamp 1698431365
transform 1 0 28560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_263
timestamp 1698431365
transform 1 0 30800 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_293
timestamp 1698431365
transform 1 0 34160 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_309
timestamp 1698431365
transform 1 0 35952 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_313
timestamp 1698431365
transform 1 0 36400 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_325
timestamp 1698431365
transform 1 0 37744 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_355
timestamp 1698431365
transform 1 0 41104 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_359
timestamp 1698431365
transform 1 0 41552 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_373
timestamp 1698431365
transform 1 0 43120 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_381
timestamp 1698431365
transform 1 0 44016 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_387
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_391
timestamp 1698431365
transform 1 0 45136 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_403
timestamp 1698431365
transform 1 0 46480 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_405
timestamp 1698431365
transform 1 0 46704 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_412
timestamp 1698431365
transform 1 0 47488 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_414
timestamp 1698431365
transform 1 0 47712 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_420
timestamp 1698431365
transform 1 0 48384 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_428
timestamp 1698431365
transform 1 0 49280 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_449
timestamp 1698431365
transform 1 0 51632 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_473
timestamp 1698431365
transform 1 0 54320 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_477
timestamp 1698431365
transform 1 0 54768 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_479
timestamp 1698431365
transform 1 0 54992 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_68
timestamp 1698431365
transform 1 0 8960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_80
timestamp 1698431365
transform 1 0 10304 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_104
timestamp 1698431365
transform 1 0 12992 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_112
timestamp 1698431365
transform 1 0 13888 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_134
timestamp 1698431365
transform 1 0 16352 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_138
timestamp 1698431365
transform 1 0 16800 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_147
timestamp 1698431365
transform 1 0 17808 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_155
timestamp 1698431365
transform 1 0 18704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_157
timestamp 1698431365
transform 1 0 18928 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_187
timestamp 1698431365
transform 1 0 22288 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_203
timestamp 1698431365
transform 1 0 24080 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_207
timestamp 1698431365
transform 1 0 24528 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_209
timestamp 1698431365
transform 1 0 24752 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_220
timestamp 1698431365
transform 1 0 25984 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_224
timestamp 1698431365
transform 1 0 26432 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_255
timestamp 1698431365
transform 1 0 29904 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_271
timestamp 1698431365
transform 1 0 31696 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_279
timestamp 1698431365
transform 1 0 32592 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_290
timestamp 1698431365
transform 1 0 33824 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_348
timestamp 1698431365
transform 1 0 40320 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_370
timestamp 1698431365
transform 1 0 42784 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_374
timestamp 1698431365
transform 1 0 43232 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_418
timestamp 1698431365
transform 1 0 48160 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_455
timestamp 1698431365
transform 1 0 52304 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_457
timestamp 1698431365
transform 1 0 52528 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_466
timestamp 1698431365
transform 1 0 53536 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_477
timestamp 1698431365
transform 1 0 54768 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_487
timestamp 1698431365
transform 1 0 55888 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_489
timestamp 1698431365
transform 1 0 56112 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_492
timestamp 1698431365
transform 1 0 56448 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_508
timestamp 1698431365
transform 1 0 58240 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_18
timestamp 1698431365
transform 1 0 3360 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_22
timestamp 1698431365
transform 1 0 3808 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_30
timestamp 1698431365
transform 1 0 4704 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_41
timestamp 1698431365
transform 1 0 5936 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_82
timestamp 1698431365
transform 1 0 10528 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_98
timestamp 1698431365
transform 1 0 12320 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_102
timestamp 1698431365
transform 1 0 12768 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_104
timestamp 1698431365
transform 1 0 12992 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_123
timestamp 1698431365
transform 1 0 15120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_181
timestamp 1698431365
transform 1 0 21616 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_185
timestamp 1698431365
transform 1 0 22064 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_194
timestamp 1698431365
transform 1 0 23072 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_227
timestamp 1698431365
transform 1 0 26768 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_251
timestamp 1698431365
transform 1 0 29456 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_274
timestamp 1698431365
transform 1 0 32032 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_282
timestamp 1698431365
transform 1 0 32928 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_286
timestamp 1698431365
transform 1 0 33376 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_288
timestamp 1698431365
transform 1 0 33600 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_293
timestamp 1698431365
transform 1 0 34160 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_295
timestamp 1698431365
transform 1 0 34384 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_321
timestamp 1698431365
transform 1 0 37296 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_331
timestamp 1698431365
transform 1 0 38416 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_335
timestamp 1698431365
transform 1 0 38864 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_339
timestamp 1698431365
transform 1 0 39312 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_343
timestamp 1698431365
transform 1 0 39760 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_346
timestamp 1698431365
transform 1 0 40096 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_352
timestamp 1698431365
transform 1 0 40768 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_387
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_445
timestamp 1698431365
transform 1 0 51184 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_453
timestamp 1698431365
transform 1 0 52080 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_472
timestamp 1698431365
transform 1 0 54208 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_476
timestamp 1698431365
transform 1 0 54656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_10
timestamp 1698431365
transform 1 0 2464 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_12
timestamp 1698431365
transform 1 0 2688 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_27
timestamp 1698431365
transform 1 0 4368 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_31
timestamp 1698431365
transform 1 0 4816 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_63
timestamp 1698431365
transform 1 0 8400 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_67
timestamp 1698431365
transform 1 0 8848 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_69
timestamp 1698431365
transform 1 0 9072 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_76
timestamp 1698431365
transform 1 0 9856 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_78
timestamp 1698431365
transform 1 0 10080 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_112
timestamp 1698431365
transform 1 0 13888 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_120
timestamp 1698431365
transform 1 0 14784 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_124
timestamp 1698431365
transform 1 0 15232 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_139
timestamp 1698431365
transform 1 0 16912 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_218
timestamp 1698431365
transform 1 0 25760 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_226
timestamp 1698431365
transform 1 0 26656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_332
timestamp 1698431365
transform 1 0 38528 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_348
timestamp 1698431365
transform 1 0 40320 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_354
timestamp 1698431365
transform 1 0 40992 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_364
timestamp 1698431365
transform 1 0 42112 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_366
timestamp 1698431365
transform 1 0 42336 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_371
timestamp 1698431365
transform 1 0 42896 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_387
timestamp 1698431365
transform 1 0 44688 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_395
timestamp 1698431365
transform 1 0 45584 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_397
timestamp 1698431365
transform 1 0 45808 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_414
timestamp 1698431365
transform 1 0 47712 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_422
timestamp 1698431365
transform 1 0 48608 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_424
timestamp 1698431365
transform 1 0 48832 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_442
timestamp 1698431365
transform 1 0 50848 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_454
timestamp 1698431365
transform 1 0 52192 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_462
timestamp 1698431365
transform 1 0 53088 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_472
timestamp 1698431365
transform 1 0 54208 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_480
timestamp 1698431365
transform 1 0 55104 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_492
timestamp 1698431365
transform 1 0 56448 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_508
timestamp 1698431365
transform 1 0 58240 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_31
timestamp 1698431365
transform 1 0 4816 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_53
timestamp 1698431365
transform 1 0 7280 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_62
timestamp 1698431365
transform 1 0 8288 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_94
timestamp 1698431365
transform 1 0 11872 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_102
timestamp 1698431365
transform 1 0 12768 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_104
timestamp 1698431365
transform 1 0 12992 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_115
timestamp 1698431365
transform 1 0 14224 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_136
timestamp 1698431365
transform 1 0 16576 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_147
timestamp 1698431365
transform 1 0 17808 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_163
timestamp 1698431365
transform 1 0 19600 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_185
timestamp 1698431365
transform 1 0 22064 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_213
timestamp 1698431365
transform 1 0 25200 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_271
timestamp 1698431365
transform 1 0 31696 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_287
timestamp 1698431365
transform 1 0 33488 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_295
timestamp 1698431365
transform 1 0 34384 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_346
timestamp 1698431365
transform 1 0 40096 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_381
timestamp 1698431365
transform 1 0 44016 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_437
timestamp 1698431365
transform 1 0 50288 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_441
timestamp 1698431365
transform 1 0 50736 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_449
timestamp 1698431365
transform 1 0 51632 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_453
timestamp 1698431365
transform 1 0 52080 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_457
timestamp 1698431365
transform 1 0 52528 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_459
timestamp 1698431365
transform 1 0 52752 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_26
timestamp 1698431365
transform 1 0 4256 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_28
timestamp 1698431365
transform 1 0 4480 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_58
timestamp 1698431365
transform 1 0 7840 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_67
timestamp 1698431365
transform 1 0 8848 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_69
timestamp 1698431365
transform 1 0 9072 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_80
timestamp 1698431365
transform 1 0 10304 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_84
timestamp 1698431365
transform 1 0 10752 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_100
timestamp 1698431365
transform 1 0 12544 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_104
timestamp 1698431365
transform 1 0 12992 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_113
timestamp 1698431365
transform 1 0 14000 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_115
timestamp 1698431365
transform 1 0 14224 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_122
timestamp 1698431365
transform 1 0 15008 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_138
timestamp 1698431365
transform 1 0 16800 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_171
timestamp 1698431365
transform 1 0 20496 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_187
timestamp 1698431365
transform 1 0 22288 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_195
timestamp 1698431365
transform 1 0 23184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_202
timestamp 1698431365
transform 1 0 23968 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_228
timestamp 1698431365
transform 1 0 26880 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_236
timestamp 1698431365
transform 1 0 27776 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_240
timestamp 1698431365
transform 1 0 28224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_242
timestamp 1698431365
transform 1 0 28448 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_250
timestamp 1698431365
transform 1 0 29344 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_334
timestamp 1698431365
transform 1 0 38752 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_430
timestamp 1698431365
transform 1 0 49504 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_434
timestamp 1698431365
transform 1 0 49952 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_442
timestamp 1698431365
transform 1 0 50848 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_446
timestamp 1698431365
transform 1 0 51296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_448
timestamp 1698431365
transform 1 0 51520 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_468
timestamp 1698431365
transform 1 0 53760 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_484
timestamp 1698431365
transform 1 0 55552 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_488
timestamp 1698431365
transform 1 0 56000 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_492
timestamp 1698431365
transform 1 0 56448 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_500
timestamp 1698431365
transform 1 0 57344 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_45
timestamp 1698431365
transform 1 0 6384 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_47
timestamp 1698431365
transform 1 0 6608 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_95
timestamp 1698431365
transform 1 0 11984 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_103
timestamp 1698431365
transform 1 0 12880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_129
timestamp 1698431365
transform 1 0 15792 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_145
timestamp 1698431365
transform 1 0 17584 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_152
timestamp 1698431365
transform 1 0 18368 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_168
timestamp 1698431365
transform 1 0 20160 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1698431365
transform 1 0 20608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698431365
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_193
timestamp 1698431365
transform 1 0 22960 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_197
timestamp 1698431365
transform 1 0 23408 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_199
timestamp 1698431365
transform 1 0 23632 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_208
timestamp 1698431365
transform 1 0 24640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_218
timestamp 1698431365
transform 1 0 25760 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_226
timestamp 1698431365
transform 1 0 26656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_228
timestamp 1698431365
transform 1 0 26880 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_243
timestamp 1698431365
transform 1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_255
timestamp 1698431365
transform 1 0 29904 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_259
timestamp 1698431365
transform 1 0 30352 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_275
timestamp 1698431365
transform 1 0 32144 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_334
timestamp 1698431365
transform 1 0 38752 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_350
timestamp 1698431365
transform 1 0 40544 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_358
timestamp 1698431365
transform 1 0 41440 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_364
timestamp 1698431365
transform 1 0 42112 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_372
timestamp 1698431365
transform 1 0 43008 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_374
timestamp 1698431365
transform 1 0 43232 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_420
timestamp 1698431365
transform 1 0 48384 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_422
timestamp 1698431365
transform 1 0 48608 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_452
timestamp 1698431365
transform 1 0 51968 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_454
timestamp 1698431365
transform 1 0 52192 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_457
timestamp 1698431365
transform 1 0 52528 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_459
timestamp 1698431365
transform 1 0 52752 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_470
timestamp 1698431365
transform 1 0 53984 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_10
timestamp 1698431365
transform 1 0 2464 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_14
timestamp 1698431365
transform 1 0 2912 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_24
timestamp 1698431365
transform 1 0 4032 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_56
timestamp 1698431365
transform 1 0 7616 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_64
timestamp 1698431365
transform 1 0 8512 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698431365
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_122
timestamp 1698431365
transform 1 0 15008 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_126
timestamp 1698431365
transform 1 0 15456 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_133
timestamp 1698431365
transform 1 0 16240 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_137
timestamp 1698431365
transform 1 0 16688 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698431365
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_158
timestamp 1698431365
transform 1 0 19040 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_189
timestamp 1698431365
transform 1 0 22512 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_191
timestamp 1698431365
transform 1 0 22736 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_198
timestamp 1698431365
transform 1 0 23520 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_216
timestamp 1698431365
transform 1 0 25536 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_246
timestamp 1698431365
transform 1 0 28896 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_254
timestamp 1698431365
transform 1 0 29792 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_258
timestamp 1698431365
transform 1 0 30240 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_260
timestamp 1698431365
transform 1 0 30464 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_269
timestamp 1698431365
transform 1 0 31472 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_277
timestamp 1698431365
transform 1 0 32368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698431365
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_346
timestamp 1698431365
transform 1 0 40096 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_370
timestamp 1698431365
transform 1 0 42784 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_378
timestamp 1698431365
transform 1 0 43680 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_390
timestamp 1698431365
transform 1 0 45024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_394
timestamp 1698431365
transform 1 0 45472 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_398
timestamp 1698431365
transform 1 0 45920 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_407
timestamp 1698431365
transform 1 0 46928 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_422
timestamp 1698431365
transform 1 0 48608 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_426
timestamp 1698431365
transform 1 0 49056 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_433
timestamp 1698431365
transform 1 0 49840 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_441
timestamp 1698431365
transform 1 0 50736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_445
timestamp 1698431365
transform 1 0 51184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_457
timestamp 1698431365
transform 1 0 52528 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_461
timestamp 1698431365
transform 1 0 52976 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_465
timestamp 1698431365
transform 1 0 53424 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_467
timestamp 1698431365
transform 1 0 53648 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_472
timestamp 1698431365
transform 1 0 54208 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_488
timestamp 1698431365
transform 1 0 56000 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_492
timestamp 1698431365
transform 1 0 56448 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_508
timestamp 1698431365
transform 1 0 58240 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_31
timestamp 1698431365
transform 1 0 4816 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_41
timestamp 1698431365
transform 1 0 5936 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_51
timestamp 1698431365
transform 1 0 7056 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_59
timestamp 1698431365
transform 1 0 7952 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_91
timestamp 1698431365
transform 1 0 11536 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_99
timestamp 1698431365
transform 1 0 12432 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_103
timestamp 1698431365
transform 1 0 12880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_111
timestamp 1698431365
transform 1 0 13776 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_119
timestamp 1698431365
transform 1 0 14672 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_127
timestamp 1698431365
transform 1 0 15568 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_172
timestamp 1698431365
transform 1 0 20608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698431365
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_181
timestamp 1698431365
transform 1 0 21616 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_218
timestamp 1698431365
transform 1 0 25760 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_226
timestamp 1698431365
transform 1 0 26656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_230
timestamp 1698431365
transform 1 0 27104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_232
timestamp 1698431365
transform 1 0 27328 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_240
timestamp 1698431365
transform 1 0 28224 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_242
timestamp 1698431365
transform 1 0 28448 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_277
timestamp 1698431365
transform 1 0 32368 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_281
timestamp 1698431365
transform 1 0 32816 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_285
timestamp 1698431365
transform 1 0 33264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_297
timestamp 1698431365
transform 1 0 34608 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_301
timestamp 1698431365
transform 1 0 35056 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_307
timestamp 1698431365
transform 1 0 35728 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_313
timestamp 1698431365
transform 1 0 36400 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_319
timestamp 1698431365
transform 1 0 37072 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_349
timestamp 1698431365
transform 1 0 40432 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_365
timestamp 1698431365
transform 1 0 42224 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_369
timestamp 1698431365
transform 1 0 42672 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_387
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_403
timestamp 1698431365
transform 1 0 46480 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_409
timestamp 1698431365
transform 1 0 47152 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_441
timestamp 1698431365
transform 1 0 50736 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_449
timestamp 1698431365
transform 1 0 51632 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_457
timestamp 1698431365
transform 1 0 52528 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_10
timestamp 1698431365
transform 1 0 2464 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_26
timestamp 1698431365
transform 1 0 4256 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_64
timestamp 1698431365
transform 1 0 8512 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698431365
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_76
timestamp 1698431365
transform 1 0 9856 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_121
timestamp 1698431365
transform 1 0 14896 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_129
timestamp 1698431365
transform 1 0 15792 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698431365
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_161
timestamp 1698431365
transform 1 0 19376 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_177
timestamp 1698431365
transform 1 0 21168 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_185
timestamp 1698431365
transform 1 0 22064 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_208
timestamp 1698431365
transform 1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_216
timestamp 1698431365
transform 1 0 25536 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_220
timestamp 1698431365
transform 1 0 25984 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_232
timestamp 1698431365
transform 1 0 27328 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_264
timestamp 1698431365
transform 1 0 30912 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_268
timestamp 1698431365
transform 1 0 31360 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698431365
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_335
timestamp 1698431365
transform 1 0 38864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_339
timestamp 1698431365
transform 1 0 39312 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_347
timestamp 1698431365
transform 1 0 40208 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_352
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_374
timestamp 1698431365
transform 1 0 43232 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_384
timestamp 1698431365
transform 1 0 44352 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_388
timestamp 1698431365
transform 1 0 44800 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_394
timestamp 1698431365
transform 1 0 45472 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_398
timestamp 1698431365
transform 1 0 45920 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_414
timestamp 1698431365
transform 1 0 47712 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_428
timestamp 1698431365
transform 1 0 49280 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_436
timestamp 1698431365
transform 1 0 50176 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_440
timestamp 1698431365
transform 1 0 50624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_442
timestamp 1698431365
transform 1 0 50848 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_476
timestamp 1698431365
transform 1 0 54656 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_480
timestamp 1698431365
transform 1 0 55104 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_485
timestamp 1698431365
transform 1 0 55664 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_489
timestamp 1698431365
transform 1 0 56112 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_492
timestamp 1698431365
transform 1 0 56448 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_508
timestamp 1698431365
transform 1 0 58240 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_41
timestamp 1698431365
transform 1 0 5936 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_49
timestamp 1698431365
transform 1 0 6832 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_65
timestamp 1698431365
transform 1 0 8624 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_69
timestamp 1698431365
transform 1 0 9072 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_72
timestamp 1698431365
transform 1 0 9408 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_104
timestamp 1698431365
transform 1 0 12992 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_115
timestamp 1698431365
transform 1 0 14224 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_119
timestamp 1698431365
transform 1 0 14672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_149
timestamp 1698431365
transform 1 0 18032 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_165
timestamp 1698431365
transform 1 0 19824 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_173
timestamp 1698431365
transform 1 0 20720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_181
timestamp 1698431365
transform 1 0 21616 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_242
timestamp 1698431365
transform 1 0 28448 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698431365
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_263
timestamp 1698431365
transform 1 0 30800 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_267
timestamp 1698431365
transform 1 0 31248 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_277
timestamp 1698431365
transform 1 0 32368 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_281
timestamp 1698431365
transform 1 0 32816 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_289
timestamp 1698431365
transform 1 0 33712 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_293
timestamp 1698431365
transform 1 0 34160 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_295
timestamp 1698431365
transform 1 0 34384 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_300
timestamp 1698431365
transform 1 0 34944 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_308
timestamp 1698431365
transform 1 0 35840 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_312
timestamp 1698431365
transform 1 0 36288 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698431365
transform 1 0 36512 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_325
timestamp 1698431365
transform 1 0 37744 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_335
timestamp 1698431365
transform 1 0 38864 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_343
timestamp 1698431365
transform 1 0 39760 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_347
timestamp 1698431365
transform 1 0 40208 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_349
timestamp 1698431365
transform 1 0 40432 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_366
timestamp 1698431365
transform 1 0 42336 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_370
timestamp 1698431365
transform 1 0 42784 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_399
timestamp 1698431365
transform 1 0 46032 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_409
timestamp 1698431365
transform 1 0 47152 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_413
timestamp 1698431365
transform 1 0 47600 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_450
timestamp 1698431365
transform 1 0 51744 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_466
timestamp 1698431365
transform 1 0 53536 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_470
timestamp 1698431365
transform 1 0 53984 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_10
timestamp 1698431365
transform 1 0 2464 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_14
timestamp 1698431365
transform 1 0 2912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_29
timestamp 1698431365
transform 1 0 4592 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_33
timestamp 1698431365
transform 1 0 5040 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_41
timestamp 1698431365
transform 1 0 5936 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_49
timestamp 1698431365
transform 1 0 6832 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_57
timestamp 1698431365
transform 1 0 7728 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_61
timestamp 1698431365
transform 1 0 8176 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_101
timestamp 1698431365
transform 1 0 12656 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_116
timestamp 1698431365
transform 1 0 14336 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_132
timestamp 1698431365
transform 1 0 16128 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_148
timestamp 1698431365
transform 1 0 17920 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_156
timestamp 1698431365
transform 1 0 18816 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_168
timestamp 1698431365
transform 1 0 20160 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_172
timestamp 1698431365
transform 1 0 20608 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_188
timestamp 1698431365
transform 1 0 22400 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_190
timestamp 1698431365
transform 1 0 22624 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_205
timestamp 1698431365
transform 1 0 24304 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698431365
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_216
timestamp 1698431365
transform 1 0 25536 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_242
timestamp 1698431365
transform 1 0 28448 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_250
timestamp 1698431365
transform 1 0 29344 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_265
timestamp 1698431365
transform 1 0 31024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_267
timestamp 1698431365
transform 1 0 31248 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_286
timestamp 1698431365
transform 1 0 33376 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_352
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_356
timestamp 1698431365
transform 1 0 41216 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_364
timestamp 1698431365
transform 1 0 42112 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_368
timestamp 1698431365
transform 1 0 42560 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_372
timestamp 1698431365
transform 1 0 43008 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_380
timestamp 1698431365
transform 1 0 43904 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_384
timestamp 1698431365
transform 1 0 44352 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_414
timestamp 1698431365
transform 1 0 47712 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_418
timestamp 1698431365
transform 1 0 48160 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_422
timestamp 1698431365
transform 1 0 48608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_424
timestamp 1698431365
transform 1 0 48832 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_440
timestamp 1698431365
transform 1 0 50624 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_481
timestamp 1698431365
transform 1 0 55216 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_486
timestamp 1698431365
transform 1 0 55776 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_492
timestamp 1698431365
transform 1 0 56448 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_508
timestamp 1698431365
transform 1 0 58240 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_31
timestamp 1698431365
transform 1 0 4816 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_45
timestamp 1698431365
transform 1 0 6384 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_61
timestamp 1698431365
transform 1 0 8176 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_93
timestamp 1698431365
transform 1 0 11760 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698431365
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_115
timestamp 1698431365
transform 1 0 14224 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_131
timestamp 1698431365
transform 1 0 16016 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_139
timestamp 1698431365
transform 1 0 16912 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_143
timestamp 1698431365
transform 1 0 17360 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_145
timestamp 1698431365
transform 1 0 17584 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_185
timestamp 1698431365
transform 1 0 22064 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_211
timestamp 1698431365
transform 1 0 24976 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_233
timestamp 1698431365
transform 1 0 27440 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_241
timestamp 1698431365
transform 1 0 28336 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_276
timestamp 1698431365
transform 1 0 32256 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_292
timestamp 1698431365
transform 1 0 34048 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_294
timestamp 1698431365
transform 1 0 34272 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_299
timestamp 1698431365
transform 1 0 34832 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_307
timestamp 1698431365
transform 1 0 35728 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698431365
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_329
timestamp 1698431365
transform 1 0 38192 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_341
timestamp 1698431365
transform 1 0 39536 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_345
timestamp 1698431365
transform 1 0 39984 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_367
timestamp 1698431365
transform 1 0 42448 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_371
timestamp 1698431365
transform 1 0 42896 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_379
timestamp 1698431365
transform 1 0 43792 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_383
timestamp 1698431365
transform 1 0 44240 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_387
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_451
timestamp 1698431365
transform 1 0 51856 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_457
timestamp 1698431365
transform 1 0 52528 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_10
timestamp 1698431365
transform 1 0 2464 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_14
timestamp 1698431365
transform 1 0 2912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_65
timestamp 1698431365
transform 1 0 8624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_69
timestamp 1698431365
transform 1 0 9072 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_88
timestamp 1698431365
transform 1 0 11200 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_96
timestamp 1698431365
transform 1 0 12096 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_98
timestamp 1698431365
transform 1 0 12320 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_121
timestamp 1698431365
transform 1 0 14896 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_125
timestamp 1698431365
transform 1 0 15344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_127
timestamp 1698431365
transform 1 0 15568 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_150
timestamp 1698431365
transform 1 0 18144 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_154
timestamp 1698431365
transform 1 0 18592 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_164
timestamp 1698431365
transform 1 0 19712 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_180
timestamp 1698431365
transform 1 0 21504 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_184
timestamp 1698431365
transform 1 0 21952 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_186
timestamp 1698431365
transform 1 0 22176 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_205
timestamp 1698431365
transform 1 0 24304 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698431365
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_220
timestamp 1698431365
transform 1 0 25984 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_224
timestamp 1698431365
transform 1 0 26432 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_226
timestamp 1698431365
transform 1 0 26656 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_237
timestamp 1698431365
transform 1 0 27888 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_241
timestamp 1698431365
transform 1 0 28336 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_273
timestamp 1698431365
transform 1 0 31920 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_277
timestamp 1698431365
transform 1 0 32368 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_326
timestamp 1698431365
transform 1 0 37856 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_330
timestamp 1698431365
transform 1 0 38304 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_341
timestamp 1698431365
transform 1 0 39536 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_345
timestamp 1698431365
transform 1 0 39984 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_349
timestamp 1698431365
transform 1 0 40432 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_361
timestamp 1698431365
transform 1 0 41776 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_373
timestamp 1698431365
transform 1 0 43120 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_377
timestamp 1698431365
transform 1 0 43568 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_385
timestamp 1698431365
transform 1 0 44464 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_389
timestamp 1698431365
transform 1 0 44912 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_432
timestamp 1698431365
transform 1 0 49728 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_440
timestamp 1698431365
transform 1 0 50624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_471
timestamp 1698431365
transform 1 0 54096 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_479
timestamp 1698431365
transform 1 0 54992 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_488
timestamp 1698431365
transform 1 0 56000 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_492
timestamp 1698431365
transform 1 0 56448 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_500
timestamp 1698431365
transform 1 0 57344 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_10
timestamp 1698431365
transform 1 0 2464 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_14
timestamp 1698431365
transform 1 0 2912 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_16
timestamp 1698431365
transform 1 0 3136 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_27
timestamp 1698431365
transform 1 0 4368 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_45
timestamp 1698431365
transform 1 0 6384 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_75
timestamp 1698431365
transform 1 0 9744 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_152
timestamp 1698431365
transform 1 0 18368 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_168
timestamp 1698431365
transform 1 0 20160 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_172
timestamp 1698431365
transform 1 0 20608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698431365
transform 1 0 20832 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_185
timestamp 1698431365
transform 1 0 22064 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_187
timestamp 1698431365
transform 1 0 22288 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_204
timestamp 1698431365
transform 1 0 24192 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_263
timestamp 1698431365
transform 1 0 30800 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_265
timestamp 1698431365
transform 1 0 31024 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_276
timestamp 1698431365
transform 1 0 32256 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_282
timestamp 1698431365
transform 1 0 32928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_286
timestamp 1698431365
transform 1 0 33376 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_302
timestamp 1698431365
transform 1 0 35168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_314
timestamp 1698431365
transform 1 0 36512 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_348
timestamp 1698431365
transform 1 0 40320 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_387
timestamp 1698431365
transform 1 0 44688 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_389
timestamp 1698431365
transform 1 0 44912 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_440
timestamp 1698431365
transform 1 0 50624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_444
timestamp 1698431365
transform 1 0 51072 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_448
timestamp 1698431365
transform 1 0 51520 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_450
timestamp 1698431365
transform 1 0 51744 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_462
timestamp 1698431365
transform 1 0 53088 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_478
timestamp 1698431365
transform 1 0 54880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_31
timestamp 1698431365
transform 1 0 4816 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_63
timestamp 1698431365
transform 1 0 8400 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_67
timestamp 1698431365
transform 1 0 8848 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_69
timestamp 1698431365
transform 1 0 9072 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_76
timestamp 1698431365
transform 1 0 9856 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_92
timestamp 1698431365
transform 1 0 11648 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_100
timestamp 1698431365
transform 1 0 12544 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_104
timestamp 1698431365
transform 1 0 12992 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_106
timestamp 1698431365
transform 1 0 13216 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_115
timestamp 1698431365
transform 1 0 14224 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_131
timestamp 1698431365
transform 1 0 16016 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698431365
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_150
timestamp 1698431365
transform 1 0 18144 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_158
timestamp 1698431365
transform 1 0 19040 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_167
timestamp 1698431365
transform 1 0 20048 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_171
timestamp 1698431365
transform 1 0 20496 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_179
timestamp 1698431365
transform 1 0 21392 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_216
timestamp 1698431365
transform 1 0 25536 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_220
timestamp 1698431365
transform 1 0 25984 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_222
timestamp 1698431365
transform 1 0 26208 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_233
timestamp 1698431365
transform 1 0 27440 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_276
timestamp 1698431365
transform 1 0 32256 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_290
timestamp 1698431365
transform 1 0 33824 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_294
timestamp 1698431365
transform 1 0 34272 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_345
timestamp 1698431365
transform 1 0 39984 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_349
timestamp 1698431365
transform 1 0 40432 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_352
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_360
timestamp 1698431365
transform 1 0 41664 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_365
timestamp 1698431365
transform 1 0 42224 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_397
timestamp 1698431365
transform 1 0 45808 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_405
timestamp 1698431365
transform 1 0 46704 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_409
timestamp 1698431365
transform 1 0 47152 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_437
timestamp 1698431365
transform 1 0 50288 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_445
timestamp 1698431365
transform 1 0 51184 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_464
timestamp 1698431365
transform 1 0 53312 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_472
timestamp 1698431365
transform 1 0 54208 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_474
timestamp 1698431365
transform 1 0 54432 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_489
timestamp 1698431365
transform 1 0 56112 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_492
timestamp 1698431365
transform 1 0 56448 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_508
timestamp 1698431365
transform 1 0 58240 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_53
timestamp 1698431365
transform 1 0 7280 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_61
timestamp 1698431365
transform 1 0 8176 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_63
timestamp 1698431365
transform 1 0 8400 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_77
timestamp 1698431365
transform 1 0 9968 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_81
timestamp 1698431365
transform 1 0 10416 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_103
timestamp 1698431365
transform 1 0 12880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_111
timestamp 1698431365
transform 1 0 13776 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_120
timestamp 1698431365
transform 1 0 14784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_124
timestamp 1698431365
transform 1 0 15232 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_134
timestamp 1698431365
transform 1 0 16352 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_138
timestamp 1698431365
transform 1 0 16800 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_179
timestamp 1698431365
transform 1 0 21392 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_206
timestamp 1698431365
transform 1 0 24416 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_238
timestamp 1698431365
transform 1 0 28000 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_242
timestamp 1698431365
transform 1 0 28448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698431365
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_247
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_263
timestamp 1698431365
transform 1 0 30800 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_267
timestamp 1698431365
transform 1 0 31248 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_276
timestamp 1698431365
transform 1 0 32256 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_280
timestamp 1698431365
transform 1 0 32704 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_282
timestamp 1698431365
transform 1 0 32928 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_312
timestamp 1698431365
transform 1 0 36288 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_314
timestamp 1698431365
transform 1 0 36512 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_324
timestamp 1698431365
transform 1 0 37632 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_328
timestamp 1698431365
transform 1 0 38080 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_334
timestamp 1698431365
transform 1 0 38752 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_350
timestamp 1698431365
transform 1 0 40544 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_364
timestamp 1698431365
transform 1 0 42112 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_380
timestamp 1698431365
transform 1 0 43904 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_384
timestamp 1698431365
transform 1 0 44352 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_387
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_407
timestamp 1698431365
transform 1 0 46928 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_437
timestamp 1698431365
transform 1 0 50288 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_453
timestamp 1698431365
transform 1 0 52080 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_457
timestamp 1698431365
transform 1 0 52528 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_465
timestamp 1698431365
transform 1 0 53424 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_471
timestamp 1698431365
transform 1 0 54096 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_479
timestamp 1698431365
transform 1 0 54992 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_60
timestamp 1698431365
transform 1 0 8064 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698431365
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_76
timestamp 1698431365
transform 1 0 9856 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_80
timestamp 1698431365
transform 1 0 10304 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_146
timestamp 1698431365
transform 1 0 17696 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_148
timestamp 1698431365
transform 1 0 17920 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_206
timestamp 1698431365
transform 1 0 24416 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_244
timestamp 1698431365
transform 1 0 28672 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_252
timestamp 1698431365
transform 1 0 29568 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_256
timestamp 1698431365
transform 1 0 30016 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_261
timestamp 1698431365
transform 1 0 30576 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_277
timestamp 1698431365
transform 1 0 32368 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698431365
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_298
timestamp 1698431365
transform 1 0 34720 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_302
timestamp 1698431365
transform 1 0 35168 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_304
timestamp 1698431365
transform 1 0 35392 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_313
timestamp 1698431365
transform 1 0 36400 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_317
timestamp 1698431365
transform 1 0 36848 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_331
timestamp 1698431365
transform 1 0 38416 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_352
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_382
timestamp 1698431365
transform 1 0 44128 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_394
timestamp 1698431365
transform 1 0 45472 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_410
timestamp 1698431365
transform 1 0 47264 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_418
timestamp 1698431365
transform 1 0 48160 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_422
timestamp 1698431365
transform 1 0 48608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_424
timestamp 1698431365
transform 1 0 48832 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_435
timestamp 1698431365
transform 1 0 50064 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_439
timestamp 1698431365
transform 1 0 50512 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_441
timestamp 1698431365
transform 1 0 50736 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_446
timestamp 1698431365
transform 1 0 51296 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_462
timestamp 1698431365
transform 1 0 53088 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_470
timestamp 1698431365
transform 1 0 53984 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_498
timestamp 1698431365
transform 1 0 57120 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_506
timestamp 1698431365
transform 1 0 58016 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_508
timestamp 1698431365
transform 1 0 58240 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_18
timestamp 1698431365
transform 1 0 3360 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698431365
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698431365
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_50
timestamp 1698431365
transform 1 0 6944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_57
timestamp 1698431365
transform 1 0 7728 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_87
timestamp 1698431365
transform 1 0 11088 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_103
timestamp 1698431365
transform 1 0 12880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_157
timestamp 1698431365
transform 1 0 18928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_161
timestamp 1698431365
transform 1 0 19376 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_169
timestamp 1698431365
transform 1 0 20272 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_173
timestamp 1698431365
transform 1 0 20720 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_185
timestamp 1698431365
transform 1 0 22064 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_200
timestamp 1698431365
transform 1 0 23744 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_208
timestamp 1698431365
transform 1 0 24640 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_241
timestamp 1698431365
transform 1 0 28336 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_299
timestamp 1698431365
transform 1 0 34832 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_307
timestamp 1698431365
transform 1 0 35728 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_311
timestamp 1698431365
transform 1 0 36176 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_319
timestamp 1698431365
transform 1 0 37072 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_328
timestamp 1698431365
transform 1 0 38080 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_330
timestamp 1698431365
transform 1 0 38304 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_360
timestamp 1698431365
transform 1 0 41664 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_368
timestamp 1698431365
transform 1 0 42560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_370
timestamp 1698431365
transform 1 0 42784 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_387
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_417
timestamp 1698431365
transform 1 0 48048 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_425
timestamp 1698431365
transform 1 0 48944 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_452
timestamp 1698431365
transform 1 0 51968 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_454
timestamp 1698431365
transform 1 0 52192 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_461
timestamp 1698431365
transform 1 0 52976 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_467
timestamp 1698431365
transform 1 0 53648 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_471
timestamp 1698431365
transform 1 0 54096 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_10
timestamp 1698431365
transform 1 0 2464 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_14
timestamp 1698431365
transform 1 0 2912 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_76
timestamp 1698431365
transform 1 0 9856 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_113
timestamp 1698431365
transform 1 0 14000 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_121
timestamp 1698431365
transform 1 0 14896 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_125
timestamp 1698431365
transform 1 0 15344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_158
timestamp 1698431365
transform 1 0 19040 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_188
timestamp 1698431365
transform 1 0 22400 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_190
timestamp 1698431365
transform 1 0 22624 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_228
timestamp 1698431365
transform 1 0 26880 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_232
timestamp 1698431365
transform 1 0 27328 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_265
timestamp 1698431365
transform 1 0 31024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_267
timestamp 1698431365
transform 1 0 31248 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_273
timestamp 1698431365
transform 1 0 31920 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_277
timestamp 1698431365
transform 1 0 32368 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698431365
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_311
timestamp 1698431365
transform 1 0 36176 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_317
timestamp 1698431365
transform 1 0 36848 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_330
timestamp 1698431365
transform 1 0 38304 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_334
timestamp 1698431365
transform 1 0 38752 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_338
timestamp 1698431365
transform 1 0 39200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_344
timestamp 1698431365
transform 1 0 39872 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_348
timestamp 1698431365
transform 1 0 40320 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_402
timestamp 1698431365
transform 1 0 46368 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_406
timestamp 1698431365
transform 1 0 46816 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_414
timestamp 1698431365
transform 1 0 47712 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_418
timestamp 1698431365
transform 1 0 48160 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_422
timestamp 1698431365
transform 1 0 48608 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_430
timestamp 1698431365
transform 1 0 49504 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_442
timestamp 1698431365
transform 1 0 50848 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_450
timestamp 1698431365
transform 1 0 51744 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_452
timestamp 1698431365
transform 1 0 51968 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_466
timestamp 1698431365
transform 1 0 53536 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_468
timestamp 1698431365
transform 1 0 53760 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_487
timestamp 1698431365
transform 1 0 55888 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_489
timestamp 1698431365
transform 1 0 56112 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_492
timestamp 1698431365
transform 1 0 56448 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_500
timestamp 1698431365
transform 1 0 57344 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_18
timestamp 1698431365
transform 1 0 3360 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_20
timestamp 1698431365
transform 1 0 3584 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_42
timestamp 1698431365
transform 1 0 6048 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_50
timestamp 1698431365
transform 1 0 6944 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_57
timestamp 1698431365
transform 1 0 7728 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_71
timestamp 1698431365
transform 1 0 9296 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_103
timestamp 1698431365
transform 1 0 12880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_123
timestamp 1698431365
transform 1 0 15120 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_131
timestamp 1698431365
transform 1 0 16016 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_138
timestamp 1698431365
transform 1 0 16800 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_170
timestamp 1698431365
transform 1 0 20384 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698431365
transform 1 0 20832 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_183
timestamp 1698431365
transform 1 0 21840 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_232
timestamp 1698431365
transform 1 0 27328 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_236
timestamp 1698431365
transform 1 0 27776 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698431365
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_301
timestamp 1698431365
transform 1 0 35056 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_309
timestamp 1698431365
transform 1 0 35952 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_313
timestamp 1698431365
transform 1 0 36400 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_325
timestamp 1698431365
transform 1 0 37744 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_331
timestamp 1698431365
transform 1 0 38416 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_335
timestamp 1698431365
transform 1 0 38864 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_367
timestamp 1698431365
transform 1 0 42448 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_375
timestamp 1698431365
transform 1 0 43344 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_381
timestamp 1698431365
transform 1 0 44016 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_387
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_397
timestamp 1698431365
transform 1 0 45808 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_405
timestamp 1698431365
transform 1 0 46704 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_407
timestamp 1698431365
transform 1 0 46928 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_414
timestamp 1698431365
transform 1 0 47712 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_449
timestamp 1698431365
transform 1 0 51632 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_457
timestamp 1698431365
transform 1 0 52528 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_36
timestamp 1698431365
transform 1 0 5376 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_52
timestamp 1698431365
transform 1 0 7168 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_56
timestamp 1698431365
transform 1 0 7616 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_69
timestamp 1698431365
transform 1 0 9072 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_76
timestamp 1698431365
transform 1 0 9856 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_78
timestamp 1698431365
transform 1 0 10080 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_81
timestamp 1698431365
transform 1 0 10416 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_85
timestamp 1698431365
transform 1 0 10864 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_91
timestamp 1698431365
transform 1 0 11536 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_97
timestamp 1698431365
transform 1 0 12208 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_105
timestamp 1698431365
transform 1 0 13104 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_109
timestamp 1698431365
transform 1 0 13552 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_158
timestamp 1698431365
transform 1 0 19040 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_166
timestamp 1698431365
transform 1 0 19936 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_170
timestamp 1698431365
transform 1 0 20384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_172
timestamp 1698431365
transform 1 0 20608 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_181
timestamp 1698431365
transform 1 0 21616 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_197
timestamp 1698431365
transform 1 0 23408 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_199
timestamp 1698431365
transform 1 0 23632 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_208
timestamp 1698431365
transform 1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_223
timestamp 1698431365
transform 1 0 26320 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_229
timestamp 1698431365
transform 1 0 26992 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_233
timestamp 1698431365
transform 1 0 27440 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_246
timestamp 1698431365
transform 1 0 28896 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_272
timestamp 1698431365
transform 1 0 31808 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698431365
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_297
timestamp 1698431365
transform 1 0 34608 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_305
timestamp 1698431365
transform 1 0 35504 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_309
timestamp 1698431365
transform 1 0 35952 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_311
timestamp 1698431365
transform 1 0 36176 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_328
timestamp 1698431365
transform 1 0 38080 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_330
timestamp 1698431365
transform 1 0 38304 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_339
timestamp 1698431365
transform 1 0 39312 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_347
timestamp 1698431365
transform 1 0 40208 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_349
timestamp 1698431365
transform 1 0 40432 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_397
timestamp 1698431365
transform 1 0 45808 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_405
timestamp 1698431365
transform 1 0 46704 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_409
timestamp 1698431365
transform 1 0 47152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_419
timestamp 1698431365
transform 1 0 48272 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_422
timestamp 1698431365
transform 1 0 48608 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_454
timestamp 1698431365
transform 1 0 52192 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_462
timestamp 1698431365
transform 1 0 53088 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_466
timestamp 1698431365
transform 1 0 53536 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_468
timestamp 1698431365
transform 1 0 53760 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_473
timestamp 1698431365
transform 1 0 54320 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_489
timestamp 1698431365
transform 1 0 56112 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_492
timestamp 1698431365
transform 1 0 56448 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_508
timestamp 1698431365
transform 1 0 58240 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_18
timestamp 1698431365
transform 1 0 3360 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_22
timestamp 1698431365
transform 1 0 3808 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_24
timestamp 1698431365
transform 1 0 4032 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_30
timestamp 1698431365
transform 1 0 4704 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_51
timestamp 1698431365
transform 1 0 7056 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_79
timestamp 1698431365
transform 1 0 10192 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_102
timestamp 1698431365
transform 1 0 12768 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_104
timestamp 1698431365
transform 1 0 12992 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_123
timestamp 1698431365
transform 1 0 15120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_125
timestamp 1698431365
transform 1 0 15344 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_142
timestamp 1698431365
transform 1 0 17248 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_185
timestamp 1698431365
transform 1 0 22064 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_212
timestamp 1698431365
transform 1 0 25088 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_216
timestamp 1698431365
transform 1 0 25536 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_218
timestamp 1698431365
transform 1 0 25760 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_234
timestamp 1698431365
transform 1 0 27552 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_238
timestamp 1698431365
transform 1 0 28000 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_242
timestamp 1698431365
transform 1 0 28448 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_244
timestamp 1698431365
transform 1 0 28672 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_252
timestamp 1698431365
transform 1 0 29568 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_256
timestamp 1698431365
transform 1 0 30016 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_260
timestamp 1698431365
transform 1 0 30464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_262
timestamp 1698431365
transform 1 0 30688 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_267
timestamp 1698431365
transform 1 0 31248 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_299
timestamp 1698431365
transform 1 0 34832 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_325
timestamp 1698431365
transform 1 0 37744 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_327
timestamp 1698431365
transform 1 0 37968 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_334
timestamp 1698431365
transform 1 0 38752 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_365
timestamp 1698431365
transform 1 0 42224 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_397
timestamp 1698431365
transform 1 0 45808 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_404
timestamp 1698431365
transform 1 0 46592 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_424
timestamp 1698431365
transform 1 0 48832 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_432
timestamp 1698431365
transform 1 0 49728 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_440
timestamp 1698431365
transform 1 0 50624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_461
timestamp 1698431365
transform 1 0 52976 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_465
timestamp 1698431365
transform 1 0 53424 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_18
timestamp 1698431365
transform 1 0 3360 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_44
timestamp 1698431365
transform 1 0 6272 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_60
timestamp 1698431365
transform 1 0 8064 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_80
timestamp 1698431365
transform 1 0 10304 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_84
timestamp 1698431365
transform 1 0 10752 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_88
timestamp 1698431365
transform 1 0 11200 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_94
timestamp 1698431365
transform 1 0 11872 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_126
timestamp 1698431365
transform 1 0 15456 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698431365
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_150
timestamp 1698431365
transform 1 0 18144 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_154
timestamp 1698431365
transform 1 0 18592 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_156
timestamp 1698431365
transform 1 0 18816 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_163
timestamp 1698431365
transform 1 0 19600 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_167
timestamp 1698431365
transform 1 0 20048 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_175
timestamp 1698431365
transform 1 0 20944 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698431365
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_216
timestamp 1698431365
transform 1 0 25536 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_220
timestamp 1698431365
transform 1 0 25984 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_222
timestamp 1698431365
transform 1 0 26208 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_237
timestamp 1698431365
transform 1 0 27888 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_241
timestamp 1698431365
transform 1 0 28336 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_249
timestamp 1698431365
transform 1 0 29232 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_286
timestamp 1698431365
transform 1 0 33376 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_288
timestamp 1698431365
transform 1 0 33600 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_318
timestamp 1698431365
transform 1 0 36960 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_334
timestamp 1698431365
transform 1 0 38752 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_352
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_368
timestamp 1698431365
transform 1 0 42560 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_376
timestamp 1698431365
transform 1 0 43456 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_383
timestamp 1698431365
transform 1 0 44240 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_388
timestamp 1698431365
transform 1 0 44800 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_392
timestamp 1698431365
transform 1 0 45248 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_400
timestamp 1698431365
transform 1 0 46144 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_417
timestamp 1698431365
transform 1 0 48048 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_419
timestamp 1698431365
transform 1 0 48272 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_422
timestamp 1698431365
transform 1 0 48608 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_426
timestamp 1698431365
transform 1 0 49056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_455
timestamp 1698431365
transform 1 0 52304 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_489
timestamp 1698431365
transform 1 0 56112 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_492
timestamp 1698431365
transform 1 0 56448 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_508
timestamp 1698431365
transform 1 0 58240 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_31
timestamp 1698431365
transform 1 0 4816 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_48
timestamp 1698431365
transform 1 0 6720 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_52
timestamp 1698431365
transform 1 0 7168 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_68
timestamp 1698431365
transform 1 0 8960 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_76
timestamp 1698431365
transform 1 0 9856 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_80
timestamp 1698431365
transform 1 0 10304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_87
timestamp 1698431365
transform 1 0 11088 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_103
timestamp 1698431365
transform 1 0 12880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_123
timestamp 1698431365
transform 1 0 15120 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_127
timestamp 1698431365
transform 1 0 15568 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_173
timestamp 1698431365
transform 1 0 20720 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_193
timestamp 1698431365
transform 1 0 22960 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_201
timestamp 1698431365
transform 1 0 23856 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_203
timestamp 1698431365
transform 1 0 24080 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_214
timestamp 1698431365
transform 1 0 25312 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_224
timestamp 1698431365
transform 1 0 26432 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_240
timestamp 1698431365
transform 1 0 28224 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_244
timestamp 1698431365
transform 1 0 28672 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_251
timestamp 1698431365
transform 1 0 29456 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_253
timestamp 1698431365
transform 1 0 29680 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_314
timestamp 1698431365
transform 1 0 36512 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_325
timestamp 1698431365
transform 1 0 37744 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_333
timestamp 1698431365
transform 1 0 38640 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_337
timestamp 1698431365
transform 1 0 39088 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_342
timestamp 1698431365
transform 1 0 39648 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_350
timestamp 1698431365
transform 1 0 40544 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_355
timestamp 1698431365
transform 1 0 41104 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_359
timestamp 1698431365
transform 1 0 41552 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_363
timestamp 1698431365
transform 1 0 42000 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_367
timestamp 1698431365
transform 1 0 42448 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_383
timestamp 1698431365
transform 1 0 44240 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_387
timestamp 1698431365
transform 1 0 44688 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_391
timestamp 1698431365
transform 1 0 45136 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_398
timestamp 1698431365
transform 1 0 45920 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_430
timestamp 1698431365
transform 1 0 49504 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_438
timestamp 1698431365
transform 1 0 50400 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_446
timestamp 1698431365
transform 1 0 51296 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_454
timestamp 1698431365
transform 1 0 52192 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_457
timestamp 1698431365
transform 1 0 52528 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_461
timestamp 1698431365
transform 1 0 52976 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_476
timestamp 1698431365
transform 1 0 54656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_480
timestamp 1698431365
transform 1 0 55104 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_483
timestamp 1698431365
transform 1 0 55440 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_499
timestamp 1698431365
transform 1 0 57232 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_507
timestamp 1698431365
transform 1 0 58128 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_18
timestamp 1698431365
transform 1 0 3360 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_26
timestamp 1698431365
transform 1 0 4256 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_35
timestamp 1698431365
transform 1 0 5264 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_43
timestamp 1698431365
transform 1 0 6160 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_51
timestamp 1698431365
transform 1 0 7056 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_53
timestamp 1698431365
transform 1 0 7280 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698431365
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_78
timestamp 1698431365
transform 1 0 10080 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_93
timestamp 1698431365
transform 1 0 11760 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_101
timestamp 1698431365
transform 1 0 12656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_132
timestamp 1698431365
transform 1 0 16128 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_150
timestamp 1698431365
transform 1 0 18144 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_154
timestamp 1698431365
transform 1 0 18592 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_185
timestamp 1698431365
transform 1 0 22064 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_191
timestamp 1698431365
transform 1 0 22736 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_195
timestamp 1698431365
transform 1 0 23184 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_203
timestamp 1698431365
transform 1 0 24080 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_207
timestamp 1698431365
transform 1 0 24528 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_209
timestamp 1698431365
transform 1 0 24752 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_222
timestamp 1698431365
transform 1 0 26208 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_253
timestamp 1698431365
transform 1 0 29680 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_267
timestamp 1698431365
transform 1 0 31248 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_277
timestamp 1698431365
transform 1 0 32368 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_279
timestamp 1698431365
transform 1 0 32592 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_292
timestamp 1698431365
transform 1 0 34048 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_302
timestamp 1698431365
transform 1 0 35168 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_306
timestamp 1698431365
transform 1 0 35616 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_316
timestamp 1698431365
transform 1 0 36736 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_320
timestamp 1698431365
transform 1 0 37184 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_352
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_372
timestamp 1698431365
transform 1 0 43008 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_388
timestamp 1698431365
transform 1 0 44800 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_392
timestamp 1698431365
transform 1 0 45248 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_401
timestamp 1698431365
transform 1 0 46256 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_409
timestamp 1698431365
transform 1 0 47152 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_414
timestamp 1698431365
transform 1 0 47712 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_418
timestamp 1698431365
transform 1 0 48160 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_430
timestamp 1698431365
transform 1 0 49504 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_446
timestamp 1698431365
transform 1 0 51296 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_454
timestamp 1698431365
transform 1 0 52192 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_458
timestamp 1698431365
transform 1 0 52640 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_467
timestamp 1698431365
transform 1 0 53648 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_483
timestamp 1698431365
transform 1 0 55440 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_487
timestamp 1698431365
transform 1 0 55888 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_489
timestamp 1698431365
transform 1 0 56112 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_492
timestamp 1698431365
transform 1 0 56448 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_508
timestamp 1698431365
transform 1 0 58240 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_18
timestamp 1698431365
transform 1 0 3360 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_22
timestamp 1698431365
transform 1 0 3808 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_43
timestamp 1698431365
transform 1 0 6160 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_51
timestamp 1698431365
transform 1 0 7056 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_68
timestamp 1698431365
transform 1 0 8960 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_123
timestamp 1698431365
transform 1 0 15120 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_131
timestamp 1698431365
transform 1 0 16016 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_135
timestamp 1698431365
transform 1 0 16464 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_144
timestamp 1698431365
transform 1 0 17472 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_160
timestamp 1698431365
transform 1 0 19264 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_172
timestamp 1698431365
transform 1 0 20608 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_174
timestamp 1698431365
transform 1 0 20832 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_181
timestamp 1698431365
transform 1 0 21616 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_192
timestamp 1698431365
transform 1 0 22848 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_194
timestamp 1698431365
transform 1 0 23072 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_224
timestamp 1698431365
transform 1 0 26432 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_240
timestamp 1698431365
transform 1 0 28224 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_244
timestamp 1698431365
transform 1 0 28672 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_251
timestamp 1698431365
transform 1 0 29456 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_259
timestamp 1698431365
transform 1 0 30352 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_261
timestamp 1698431365
transform 1 0 30576 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698431365
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_325
timestamp 1698431365
transform 1 0 37744 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_329
timestamp 1698431365
transform 1 0 38192 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_381
timestamp 1698431365
transform 1 0 44016 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_416
timestamp 1698431365
transform 1 0 47936 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_432
timestamp 1698431365
transform 1 0 49728 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_448
timestamp 1698431365
transform 1 0 51520 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_452
timestamp 1698431365
transform 1 0 51968 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_454
timestamp 1698431365
transform 1 0 52192 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_468
timestamp 1698431365
transform 1 0 53760 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_470
timestamp 1698431365
transform 1 0 53984 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_479
timestamp 1698431365
transform 1 0 54992 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_44
timestamp 1698431365
transform 1 0 6272 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_60
timestamp 1698431365
transform 1 0 8064 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_68
timestamp 1698431365
transform 1 0 8960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_104
timestamp 1698431365
transform 1 0 12992 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_108
timestamp 1698431365
transform 1 0 13440 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_110
timestamp 1698431365
transform 1 0 13664 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_150
timestamp 1698431365
transform 1 0 18144 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_154
timestamp 1698431365
transform 1 0 18592 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_193
timestamp 1698431365
transform 1 0 22960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_220
timestamp 1698431365
transform 1 0 25984 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_224
timestamp 1698431365
transform 1 0 26432 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_270
timestamp 1698431365
transform 1 0 31584 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_274
timestamp 1698431365
transform 1 0 32032 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_278
timestamp 1698431365
transform 1 0 32480 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_308
timestamp 1698431365
transform 1 0 35840 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_340
timestamp 1698431365
transform 1 0 39424 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_348
timestamp 1698431365
transform 1 0 40320 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_389
timestamp 1698431365
transform 1 0 44912 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_405
timestamp 1698431365
transform 1 0 46704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_407
timestamp 1698431365
transform 1 0 46928 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_422
timestamp 1698431365
transform 1 0 48608 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_424
timestamp 1698431365
transform 1 0 48832 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_429
timestamp 1698431365
transform 1 0 49392 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_434
timestamp 1698431365
transform 1 0 49952 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_445
timestamp 1698431365
transform 1 0 51184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_460
timestamp 1698431365
transform 1 0 52864 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_476
timestamp 1698431365
transform 1 0 54656 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_484
timestamp 1698431365
transform 1 0 55552 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_488
timestamp 1698431365
transform 1 0 56000 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_492
timestamp 1698431365
transform 1 0 56448 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_496
timestamp 1698431365
transform 1 0 56896 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_498
timestamp 1698431365
transform 1 0 57120 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_31
timestamp 1698431365
transform 1 0 4816 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_47
timestamp 1698431365
transform 1 0 6608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_78
timestamp 1698431365
transform 1 0 10080 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_86
timestamp 1698431365
transform 1 0 10976 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_90
timestamp 1698431365
transform 1 0 11424 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_93
timestamp 1698431365
transform 1 0 11760 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_103
timestamp 1698431365
transform 1 0 12880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_123
timestamp 1698431365
transform 1 0 15120 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_131
timestamp 1698431365
transform 1 0 16016 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_138
timestamp 1698431365
transform 1 0 16800 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_154
timestamp 1698431365
transform 1 0 18592 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_162
timestamp 1698431365
transform 1 0 19488 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_166
timestamp 1698431365
transform 1 0 19936 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_171
timestamp 1698431365
transform 1 0 20496 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_227
timestamp 1698431365
transform 1 0 26768 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_237
timestamp 1698431365
transform 1 0 27888 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698431365
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_251
timestamp 1698431365
transform 1 0 29456 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_304
timestamp 1698431365
transform 1 0 35392 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_312
timestamp 1698431365
transform 1 0 36288 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_314
timestamp 1698431365
transform 1 0 36512 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_321
timestamp 1698431365
transform 1 0 37296 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_338
timestamp 1698431365
transform 1 0 39200 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_354
timestamp 1698431365
transform 1 0 40992 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_358
timestamp 1698431365
transform 1 0 41440 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_369
timestamp 1698431365
transform 1 0 42672 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_373
timestamp 1698431365
transform 1 0 43120 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_381
timestamp 1698431365
transform 1 0 44016 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_387
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_432
timestamp 1698431365
transform 1 0 49728 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_439
timestamp 1698431365
transform 1 0 50512 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_444
timestamp 1698431365
transform 1 0 51072 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_448
timestamp 1698431365
transform 1 0 51520 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_10
timestamp 1698431365
transform 1 0 2464 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_12
timestamp 1698431365
transform 1 0 2688 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_69
timestamp 1698431365
transform 1 0 9072 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_76
timestamp 1698431365
transform 1 0 9856 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_84
timestamp 1698431365
transform 1 0 10752 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_120
timestamp 1698431365
transform 1 0 14784 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_124
timestamp 1698431365
transform 1 0 15232 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_126
timestamp 1698431365
transform 1 0 15456 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_137
timestamp 1698431365
transform 1 0 16688 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_139
timestamp 1698431365
transform 1 0 16912 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_171
timestamp 1698431365
transform 1 0 20496 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_179
timestamp 1698431365
transform 1 0 21392 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_220
timestamp 1698431365
transform 1 0 25984 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_224
timestamp 1698431365
transform 1 0 26432 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_239
timestamp 1698431365
transform 1 0 28112 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_243
timestamp 1698431365
transform 1 0 28560 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_275
timestamp 1698431365
transform 1 0 32144 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_279
timestamp 1698431365
transform 1 0 32592 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_299
timestamp 1698431365
transform 1 0 34832 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_343
timestamp 1698431365
transform 1 0 39760 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_347
timestamp 1698431365
transform 1 0 40208 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_349
timestamp 1698431365
transform 1 0 40432 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_352
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_356
timestamp 1698431365
transform 1 0 41216 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_363
timestamp 1698431365
transform 1 0 42000 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_371
timestamp 1698431365
transform 1 0 42896 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_405
timestamp 1698431365
transform 1 0 46704 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_409
timestamp 1698431365
transform 1 0 47152 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_418
timestamp 1698431365
transform 1 0 48160 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_422
timestamp 1698431365
transform 1 0 48608 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_438
timestamp 1698431365
transform 1 0 50400 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_442
timestamp 1698431365
transform 1 0 50848 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_473
timestamp 1698431365
transform 1 0 54320 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_477
timestamp 1698431365
transform 1 0 54768 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_485
timestamp 1698431365
transform 1 0 55664 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_489
timestamp 1698431365
transform 1 0 56112 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_492
timestamp 1698431365
transform 1 0 56448 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_508
timestamp 1698431365
transform 1 0 58240 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_18
timestamp 1698431365
transform 1 0 3360 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_22
timestamp 1698431365
transform 1 0 3808 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_24
timestamp 1698431365
transform 1 0 4032 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_45
timestamp 1698431365
transform 1 0 6384 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_61
timestamp 1698431365
transform 1 0 8176 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_91
timestamp 1698431365
transform 1 0 11536 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_99
timestamp 1698431365
transform 1 0 12432 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_103
timestamp 1698431365
transform 1 0 12880 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_157
timestamp 1698431365
transform 1 0 18928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_161
timestamp 1698431365
transform 1 0 19376 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_169
timestamp 1698431365
transform 1 0 20272 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_173
timestamp 1698431365
transform 1 0 20720 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_209
timestamp 1698431365
transform 1 0 24752 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_213
timestamp 1698431365
transform 1 0 25200 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_215
timestamp 1698431365
transform 1 0 25424 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_221
timestamp 1698431365
transform 1 0 26096 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_225
timestamp 1698431365
transform 1 0 26544 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_229
timestamp 1698431365
transform 1 0 26992 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_233
timestamp 1698431365
transform 1 0 27440 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_251
timestamp 1698431365
transform 1 0 29456 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_291
timestamp 1698431365
transform 1 0 33936 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_293
timestamp 1698431365
transform 1 0 34160 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_304
timestamp 1698431365
transform 1 0 35392 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_312
timestamp 1698431365
transform 1 0 36288 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_314
timestamp 1698431365
transform 1 0 36512 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_346
timestamp 1698431365
transform 1 0 40096 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_348
timestamp 1698431365
transform 1 0 40320 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_351
timestamp 1698431365
transform 1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_370
timestamp 1698431365
transform 1 0 42784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_376
timestamp 1698431365
transform 1 0 43456 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_384
timestamp 1698431365
transform 1 0 44352 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_387
timestamp 1698431365
transform 1 0 44688 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_419
timestamp 1698431365
transform 1 0 48272 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_422
timestamp 1698431365
transform 1 0 48608 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_426
timestamp 1698431365
transform 1 0 49056 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_438
timestamp 1698431365
transform 1 0 50400 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_446
timestamp 1698431365
transform 1 0 51296 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_450
timestamp 1698431365
transform 1 0 51744 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_452
timestamp 1698431365
transform 1 0 51968 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_457
timestamp 1698431365
transform 1 0 52528 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_18
timestamp 1698431365
transform 1 0 3360 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_44
timestamp 1698431365
transform 1 0 6272 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_52
timestamp 1698431365
transform 1 0 7168 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_54
timestamp 1698431365
transform 1 0 7392 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_80
timestamp 1698431365
transform 1 0 10304 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_84
timestamp 1698431365
transform 1 0 10752 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_100
timestamp 1698431365
transform 1 0 12544 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_104
timestamp 1698431365
transform 1 0 12992 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_113
timestamp 1698431365
transform 1 0 14000 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_117
timestamp 1698431365
transform 1 0 14448 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_121
timestamp 1698431365
transform 1 0 14896 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_158
timestamp 1698431365
transform 1 0 19040 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_162
timestamp 1698431365
transform 1 0 19488 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_195
timestamp 1698431365
transform 1 0 23184 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_203
timestamp 1698431365
transform 1 0 24080 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_207
timestamp 1698431365
transform 1 0 24528 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_209
timestamp 1698431365
transform 1 0 24752 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_216
timestamp 1698431365
transform 1 0 25536 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_218
timestamp 1698431365
transform 1 0 25760 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_227
timestamp 1698431365
transform 1 0 26768 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_231
timestamp 1698431365
transform 1 0 27216 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_233
timestamp 1698431365
transform 1 0 27440 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_254
timestamp 1698431365
transform 1 0 29792 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_258
timestamp 1698431365
transform 1 0 30240 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_266
timestamp 1698431365
transform 1 0 31136 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_270
timestamp 1698431365
transform 1 0 31584 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_286
timestamp 1698431365
transform 1 0 33376 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_302
timestamp 1698431365
transform 1 0 35168 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_306
timestamp 1698431365
transform 1 0 35616 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_315
timestamp 1698431365
transform 1 0 36624 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_323
timestamp 1698431365
transform 1 0 37520 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_338
timestamp 1698431365
transform 1 0 39200 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_349
timestamp 1698431365
transform 1 0 40432 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_366
timestamp 1698431365
transform 1 0 42336 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_370
timestamp 1698431365
transform 1 0 42784 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_376
timestamp 1698431365
transform 1 0 43456 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_380
timestamp 1698431365
transform 1 0 43904 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_384
timestamp 1698431365
transform 1 0 44352 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_392
timestamp 1698431365
transform 1 0 45248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_394
timestamp 1698431365
transform 1 0 45472 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_397
timestamp 1698431365
transform 1 0 45808 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_417
timestamp 1698431365
transform 1 0 48048 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_419
timestamp 1698431365
transform 1 0 48272 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_472
timestamp 1698431365
transform 1 0 54208 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_486
timestamp 1698431365
transform 1 0 55776 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_492
timestamp 1698431365
transform 1 0 56448 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_496
timestamp 1698431365
transform 1 0 56896 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_504
timestamp 1698431365
transform 1 0 57792 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_508
timestamp 1698431365
transform 1 0 58240 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_31
timestamp 1698431365
transform 1 0 4816 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_42
timestamp 1698431365
transform 1 0 6048 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_74
timestamp 1698431365
transform 1 0 9632 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_90
timestamp 1698431365
transform 1 0 11424 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_100
timestamp 1698431365
transform 1 0 12544 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_104
timestamp 1698431365
transform 1 0 12992 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_115
timestamp 1698431365
transform 1 0 14224 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_123
timestamp 1698431365
transform 1 0 15120 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_130
timestamp 1698431365
transform 1 0 15904 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_145
timestamp 1698431365
transform 1 0 17584 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_161
timestamp 1698431365
transform 1 0 19376 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_173
timestamp 1698431365
transform 1 0 20720 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_181
timestamp 1698431365
transform 1 0 21616 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_197
timestamp 1698431365
transform 1 0 23408 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_201
timestamp 1698431365
transform 1 0 23856 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_240
timestamp 1698431365
transform 1 0 28224 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_244
timestamp 1698431365
transform 1 0 28672 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_263
timestamp 1698431365
transform 1 0 30800 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_289
timestamp 1698431365
transform 1 0 33712 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_293
timestamp 1698431365
transform 1 0 34160 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_297
timestamp 1698431365
transform 1 0 34608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_299
timestamp 1698431365
transform 1 0 34832 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_310
timestamp 1698431365
transform 1 0 36064 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_314
timestamp 1698431365
transform 1 0 36512 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_325
timestamp 1698431365
transform 1 0 37744 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_332
timestamp 1698431365
transform 1 0 38528 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_336
timestamp 1698431365
transform 1 0 38976 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_339
timestamp 1698431365
transform 1 0 39312 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_355
timestamp 1698431365
transform 1 0 41104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_357
timestamp 1698431365
transform 1 0 41328 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_382
timestamp 1698431365
transform 1 0 44128 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_384
timestamp 1698431365
transform 1 0 44352 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_395
timestamp 1698431365
transform 1 0 45584 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_404
timestamp 1698431365
transform 1 0 46592 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_408
timestamp 1698431365
transform 1 0 47040 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_416
timestamp 1698431365
transform 1 0 47936 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_420
timestamp 1698431365
transform 1 0 48384 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_450
timestamp 1698431365
transform 1 0 51744 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_466
timestamp 1698431365
transform 1 0 53536 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_476
timestamp 1698431365
transform 1 0 54656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_18
timestamp 1698431365
transform 1 0 3360 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_26
timestamp 1698431365
transform 1 0 4256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_40
timestamp 1698431365
transform 1 0 5824 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_48
timestamp 1698431365
transform 1 0 6720 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_50
timestamp 1698431365
transform 1 0 6944 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_57
timestamp 1698431365
transform 1 0 7728 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_68
timestamp 1698431365
transform 1 0 8960 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_88
timestamp 1698431365
transform 1 0 11200 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_133
timestamp 1698431365
transform 1 0 16240 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_137
timestamp 1698431365
transform 1 0 16688 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_139
timestamp 1698431365
transform 1 0 16912 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_150
timestamp 1698431365
transform 1 0 18144 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_154
timestamp 1698431365
transform 1 0 18592 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_166
timestamp 1698431365
transform 1 0 19936 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_170
timestamp 1698431365
transform 1 0 20384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_174
timestamp 1698431365
transform 1 0 20832 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_182
timestamp 1698431365
transform 1 0 21728 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_186
timestamp 1698431365
transform 1 0 22176 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_188
timestamp 1698431365
transform 1 0 22400 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_204
timestamp 1698431365
transform 1 0 24192 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_208
timestamp 1698431365
transform 1 0 24640 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_228
timestamp 1698431365
transform 1 0 26880 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_236
timestamp 1698431365
transform 1 0 27776 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_242
timestamp 1698431365
transform 1 0 28448 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_249
timestamp 1698431365
transform 1 0 29232 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_253
timestamp 1698431365
transform 1 0 29680 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_259
timestamp 1698431365
transform 1 0 30352 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_277
timestamp 1698431365
transform 1 0 32368 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698431365
transform 1 0 32592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_286
timestamp 1698431365
transform 1 0 33376 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_302
timestamp 1698431365
transform 1 0 35168 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_321
timestamp 1698431365
transform 1 0 37296 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_325
timestamp 1698431365
transform 1 0 37744 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_335
timestamp 1698431365
transform 1 0 38864 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_343
timestamp 1698431365
transform 1 0 39760 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_347
timestamp 1698431365
transform 1 0 40208 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_349
timestamp 1698431365
transform 1 0 40432 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_360
timestamp 1698431365
transform 1 0 41664 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_370
timestamp 1698431365
transform 1 0 42784 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_374
timestamp 1698431365
transform 1 0 43232 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_382
timestamp 1698431365
transform 1 0 44128 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_386
timestamp 1698431365
transform 1 0 44576 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_416
timestamp 1698431365
transform 1 0 47936 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_434
timestamp 1698431365
transform 1 0 49952 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_450
timestamp 1698431365
transform 1 0 51744 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_458
timestamp 1698431365
transform 1 0 52640 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_460
timestamp 1698431365
transform 1 0 52864 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_496
timestamp 1698431365
transform 1 0 56896 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_504
timestamp 1698431365
transform 1 0 57792 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_506
timestamp 1698431365
transform 1 0 58016 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_51
timestamp 1698431365
transform 1 0 7056 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_53
timestamp 1698431365
transform 1 0 7280 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_59
timestamp 1698431365
transform 1 0 7952 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_63
timestamp 1698431365
transform 1 0 8400 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_69
timestamp 1698431365
transform 1 0 9072 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_91
timestamp 1698431365
transform 1 0 11536 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_95
timestamp 1698431365
transform 1 0 11984 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_103
timestamp 1698431365
transform 1 0 12880 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_123
timestamp 1698431365
transform 1 0 15120 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_131
timestamp 1698431365
transform 1 0 16016 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_161
timestamp 1698431365
transform 1 0 19376 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_169
timestamp 1698431365
transform 1 0 20272 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_173
timestamp 1698431365
transform 1 0 20720 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_185
timestamp 1698431365
transform 1 0 22064 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_189
timestamp 1698431365
transform 1 0 22512 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_205
timestamp 1698431365
transform 1 0 24304 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_221
timestamp 1698431365
transform 1 0 26096 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_229
timestamp 1698431365
transform 1 0 26992 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_231
timestamp 1698431365
transform 1 0 27216 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_240
timestamp 1698431365
transform 1 0 28224 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_242
timestamp 1698431365
transform 1 0 28448 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_257
timestamp 1698431365
transform 1 0 30128 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_259
timestamp 1698431365
transform 1 0 30352 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_289
timestamp 1698431365
transform 1 0 33712 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_295
timestamp 1698431365
transform 1 0 34384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_299
timestamp 1698431365
transform 1 0 34832 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_301
timestamp 1698431365
transform 1 0 35056 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_314
timestamp 1698431365
transform 1 0 36512 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_347
timestamp 1698431365
transform 1 0 40208 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_355
timestamp 1698431365
transform 1 0 41104 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_359
timestamp 1698431365
transform 1 0 41552 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_365
timestamp 1698431365
transform 1 0 42224 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_373
timestamp 1698431365
transform 1 0 43120 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_381
timestamp 1698431365
transform 1 0 44016 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_437
timestamp 1698431365
transform 1 0 50288 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_441
timestamp 1698431365
transform 1 0 50736 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_449
timestamp 1698431365
transform 1 0 51632 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_453
timestamp 1698431365
transform 1 0 52080 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_457
timestamp 1698431365
transform 1 0 52528 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_465
timestamp 1698431365
transform 1 0 53424 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_469
timestamp 1698431365
transform 1 0 53872 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_471
timestamp 1698431365
transform 1 0 54096 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_31
timestamp 1698431365
transform 1 0 4816 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_58
timestamp 1698431365
transform 1 0 7840 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_101
timestamp 1698431365
transform 1 0 12656 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_117
timestamp 1698431365
transform 1 0 14448 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_122
timestamp 1698431365
transform 1 0 15008 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_138
timestamp 1698431365
transform 1 0 16800 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_146
timestamp 1698431365
transform 1 0 17696 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_151
timestamp 1698431365
transform 1 0 18256 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_161
timestamp 1698431365
transform 1 0 19376 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_165
timestamp 1698431365
transform 1 0 19824 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_198
timestamp 1698431365
transform 1 0 23520 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_206
timestamp 1698431365
transform 1 0 24416 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_220
timestamp 1698431365
transform 1 0 25984 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_224
timestamp 1698431365
transform 1 0 26432 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_266
timestamp 1698431365
transform 1 0 31136 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_274
timestamp 1698431365
transform 1 0 32032 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_284
timestamp 1698431365
transform 1 0 33152 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_324
timestamp 1698431365
transform 1 0 37632 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_336
timestamp 1698431365
transform 1 0 38976 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_340
timestamp 1698431365
transform 1 0 39424 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_348
timestamp 1698431365
transform 1 0 40320 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_381
timestamp 1698431365
transform 1 0 44016 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_389
timestamp 1698431365
transform 1 0 44912 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_409
timestamp 1698431365
transform 1 0 47152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_411
timestamp 1698431365
transform 1 0 47376 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_430
timestamp 1698431365
transform 1 0 49504 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_432
timestamp 1698431365
transform 1 0 49728 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_462
timestamp 1698431365
transform 1 0 53088 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_470
timestamp 1698431365
transform 1 0 53984 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_474
timestamp 1698431365
transform 1 0 54432 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_476
timestamp 1698431365
transform 1 0 54656 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_492
timestamp 1698431365
transform 1 0 56448 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_496
timestamp 1698431365
transform 1 0 56896 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_505
timestamp 1698431365
transform 1 0 57904 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_31
timestamp 1698431365
transform 1 0 4816 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_76
timestamp 1698431365
transform 1 0 9856 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_92
timestamp 1698431365
transform 1 0 11648 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_100
timestamp 1698431365
transform 1 0 12544 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_104
timestamp 1698431365
transform 1 0 12992 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_145
timestamp 1698431365
transform 1 0 17584 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_149
timestamp 1698431365
transform 1 0 18032 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_153
timestamp 1698431365
transform 1 0 18480 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_160
timestamp 1698431365
transform 1 0 19264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_164
timestamp 1698431365
transform 1 0 19712 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_172
timestamp 1698431365
transform 1 0 20608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_174
timestamp 1698431365
transform 1 0 20832 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_185
timestamp 1698431365
transform 1 0 22064 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_190
timestamp 1698431365
transform 1 0 22624 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_206
timestamp 1698431365
transform 1 0 24416 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_241
timestamp 1698431365
transform 1 0 28336 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_251
timestamp 1698431365
transform 1 0 29456 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_255
timestamp 1698431365
transform 1 0 29904 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_271
timestamp 1698431365
transform 1 0 31696 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_279
timestamp 1698431365
transform 1 0 32592 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_283
timestamp 1698431365
transform 1 0 33040 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_294
timestamp 1698431365
transform 1 0 34272 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_298
timestamp 1698431365
transform 1 0 34720 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_300
timestamp 1698431365
transform 1 0 34944 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_309
timestamp 1698431365
transform 1 0 35952 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_313
timestamp 1698431365
transform 1 0 36400 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_321
timestamp 1698431365
transform 1 0 37296 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_323
timestamp 1698431365
transform 1 0 37520 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_326
timestamp 1698431365
transform 1 0 37856 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_330
timestamp 1698431365
transform 1 0 38304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_334
timestamp 1698431365
transform 1 0 38752 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_350
timestamp 1698431365
transform 1 0 40544 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_352
timestamp 1698431365
transform 1 0 40768 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_359
timestamp 1698431365
transform 1 0 41552 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_370
timestamp 1698431365
transform 1 0 42784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_374
timestamp 1698431365
transform 1 0 43232 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_382
timestamp 1698431365
transform 1 0 44128 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_384
timestamp 1698431365
transform 1 0 44352 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_387
timestamp 1698431365
transform 1 0 44688 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_391
timestamp 1698431365
transform 1 0 45136 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_395
timestamp 1698431365
transform 1 0 45584 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_403
timestamp 1698431365
transform 1 0 46480 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_407
timestamp 1698431365
transform 1 0 46928 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_409
timestamp 1698431365
transform 1 0 47152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_412
timestamp 1698431365
transform 1 0 47488 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_422
timestamp 1698431365
transform 1 0 48608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_424
timestamp 1698431365
transform 1 0 48832 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_431
timestamp 1698431365
transform 1 0 49616 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_447
timestamp 1698431365
transform 1 0 51408 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_465
timestamp 1698431365
transform 1 0 53424 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_469
timestamp 1698431365
transform 1 0 53872 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_471
timestamp 1698431365
transform 1 0 54096 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_18
timestamp 1698431365
transform 1 0 3360 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_76
timestamp 1698431365
transform 1 0 9856 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_84
timestamp 1698431365
transform 1 0 10752 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_117
timestamp 1698431365
transform 1 0 14448 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_125
timestamp 1698431365
transform 1 0 15344 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_129
timestamp 1698431365
transform 1 0 15792 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_146
timestamp 1698431365
transform 1 0 17696 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_150
timestamp 1698431365
transform 1 0 18144 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_161
timestamp 1698431365
transform 1 0 19376 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_165
timestamp 1698431365
transform 1 0 19824 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_169
timestamp 1698431365
transform 1 0 20272 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_171
timestamp 1698431365
transform 1 0 20496 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_262
timestamp 1698431365
transform 1 0 30688 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_278
timestamp 1698431365
transform 1 0 32480 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_290
timestamp 1698431365
transform 1 0 33824 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_294
timestamp 1698431365
transform 1 0 34272 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_298
timestamp 1698431365
transform 1 0 34720 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_302
timestamp 1698431365
transform 1 0 35168 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_304
timestamp 1698431365
transform 1 0 35392 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_346
timestamp 1698431365
transform 1 0 40096 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_368
timestamp 1698431365
transform 1 0 42560 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_372
timestamp 1698431365
transform 1 0 43008 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_374
timestamp 1698431365
transform 1 0 43232 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_377
timestamp 1698431365
transform 1 0 43568 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_385
timestamp 1698431365
transform 1 0 44464 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_392
timestamp 1698431365
transform 1 0 45248 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_404
timestamp 1698431365
transform 1 0 46592 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_422
timestamp 1698431365
transform 1 0 48608 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_426
timestamp 1698431365
transform 1 0 49056 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_434
timestamp 1698431365
transform 1 0 49952 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_450
timestamp 1698431365
transform 1 0 51744 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_453
timestamp 1698431365
transform 1 0 52080 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_468
timestamp 1698431365
transform 1 0 53760 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_492
timestamp 1698431365
transform 1 0 56448 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_500
timestamp 1698431365
transform 1 0 57344 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_53
timestamp 1698431365
transform 1 0 7280 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_61
timestamp 1698431365
transform 1 0 8176 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_91
timestamp 1698431365
transform 1 0 11536 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_99
timestamp 1698431365
transform 1 0 12432 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_104
timestamp 1698431365
transform 1 0 12992 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_123
timestamp 1698431365
transform 1 0 15120 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_137
timestamp 1698431365
transform 1 0 16688 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_141
timestamp 1698431365
transform 1 0 17136 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_172
timestamp 1698431365
transform 1 0 20608 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_174
timestamp 1698431365
transform 1 0 20832 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_209
timestamp 1698431365
transform 1 0 24752 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_212
timestamp 1698431365
transform 1 0 25088 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_225
timestamp 1698431365
transform 1 0 26544 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_229
timestamp 1698431365
transform 1 0 26992 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_231
timestamp 1698431365
transform 1 0 27216 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_238
timestamp 1698431365
transform 1 0 28000 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_242
timestamp 1698431365
transform 1 0 28448 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_253
timestamp 1698431365
transform 1 0 29680 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_255
timestamp 1698431365
transform 1 0 29904 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_262
timestamp 1698431365
transform 1 0 30688 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_266
timestamp 1698431365
transform 1 0 31136 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_296
timestamp 1698431365
transform 1 0 34496 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_312
timestamp 1698431365
transform 1 0 36288 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_314
timestamp 1698431365
transform 1 0 36512 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_322
timestamp 1698431365
transform 1 0 37408 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_324
timestamp 1698431365
transform 1 0 37632 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_384
timestamp 1698431365
transform 1 0 44352 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_387
timestamp 1698431365
transform 1 0 44688 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_389
timestamp 1698431365
transform 1 0 44912 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_419
timestamp 1698431365
transform 1 0 48272 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_436
timestamp 1698431365
transform 1 0 50176 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_444
timestamp 1698431365
transform 1 0 51072 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_452
timestamp 1698431365
transform 1 0 51968 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_454
timestamp 1698431365
transform 1 0 52192 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_507
timestamp 1698431365
transform 1 0 58128 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_66
timestamp 1698431365
transform 1 0 8736 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_88
timestamp 1698431365
transform 1 0 11200 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_92
timestamp 1698431365
transform 1 0 11648 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_139
timestamp 1698431365
transform 1 0 16912 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_142
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_150
timestamp 1698431365
transform 1 0 18144 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_152
timestamp 1698431365
transform 1 0 18368 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_157
timestamp 1698431365
transform 1 0 18928 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_165
timestamp 1698431365
transform 1 0 19824 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_207
timestamp 1698431365
transform 1 0 24528 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_209
timestamp 1698431365
transform 1 0 24752 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_212
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_216
timestamp 1698431365
transform 1 0 25536 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_226
timestamp 1698431365
transform 1 0 26656 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_233
timestamp 1698431365
transform 1 0 27440 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_235
timestamp 1698431365
transform 1 0 27664 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_265
timestamp 1698431365
transform 1 0 31024 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_269
timestamp 1698431365
transform 1 0 31472 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_286
timestamp 1698431365
transform 1 0 33376 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_290
timestamp 1698431365
transform 1 0 33824 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_298
timestamp 1698431365
transform 1 0 34720 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_306
timestamp 1698431365
transform 1 0 35616 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_314
timestamp 1698431365
transform 1 0 36512 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_318
timestamp 1698431365
transform 1 0 36960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_331
timestamp 1698431365
transform 1 0 38416 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_347
timestamp 1698431365
transform 1 0 40208 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_349
timestamp 1698431365
transform 1 0 40432 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_381
timestamp 1698431365
transform 1 0 44016 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_383
timestamp 1698431365
transform 1 0 44240 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_386
timestamp 1698431365
transform 1 0 44576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_395
timestamp 1698431365
transform 1 0 45584 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_403
timestamp 1698431365
transform 1 0 46480 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_407
timestamp 1698431365
transform 1 0 46928 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_422
timestamp 1698431365
transform 1 0 48608 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_481
timestamp 1698431365
transform 1 0 55216 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_489
timestamp 1698431365
transform 1 0 56112 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_492
timestamp 1698431365
transform 1 0 56448 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_508
timestamp 1698431365
transform 1 0 58240 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_2
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698431365
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_37
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_69
timestamp 1698431365
transform 1 0 9072 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_71
timestamp 1698431365
transform 1 0 9296 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_88
timestamp 1698431365
transform 1 0 11200 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_104
timestamp 1698431365
transform 1 0 12992 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_107
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_109
timestamp 1698431365
transform 1 0 13552 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_118
timestamp 1698431365
transform 1 0 14560 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_122
timestamp 1698431365
transform 1 0 15008 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_124
timestamp 1698431365
transform 1 0 15232 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_177
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_181
timestamp 1698431365
transform 1 0 21616 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_187
timestamp 1698431365
transform 1 0 22288 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_203
timestamp 1698431365
transform 1 0 24080 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_233
timestamp 1698431365
transform 1 0 27440 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_237
timestamp 1698431365
transform 1 0 27888 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_257
timestamp 1698431365
transform 1 0 30128 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_259
timestamp 1698431365
transform 1 0 30352 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_269
timestamp 1698431365
transform 1 0 31472 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_273
timestamp 1698431365
transform 1 0 31920 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_281
timestamp 1698431365
transform 1 0 32816 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_285
timestamp 1698431365
transform 1 0 33264 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_317
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_330
timestamp 1698431365
transform 1 0 38304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_334
timestamp 1698431365
transform 1 0 38752 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_338
timestamp 1698431365
transform 1 0 39200 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_342
timestamp 1698431365
transform 1 0 39648 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_345
timestamp 1698431365
transform 1 0 39984 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_377
timestamp 1698431365
transform 1 0 43568 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_387
timestamp 1698431365
transform 1 0 44688 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_395
timestamp 1698431365
transform 1 0 45584 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_410
timestamp 1698431365
transform 1 0 47264 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_426
timestamp 1698431365
transform 1 0 49056 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_434
timestamp 1698431365
transform 1 0 49952 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_466
timestamp 1698431365
transform 1 0 53536 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_474
timestamp 1698431365
transform 1 0 54432 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_478
timestamp 1698431365
transform 1 0 54880 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_492
timestamp 1698431365
transform 1 0 56448 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_498
timestamp 1698431365
transform 1 0 57120 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_506
timestamp 1698431365
transform 1 0 58016 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_508
timestamp 1698431365
transform 1 0 58240 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_2
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_18
timestamp 1698431365
transform 1 0 3360 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_26
timestamp 1698431365
transform 1 0 4256 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_28
timestamp 1698431365
transform 1 0 4480 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_58
timestamp 1698431365
transform 1 0 7840 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_66
timestamp 1698431365
transform 1 0 8736 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_72
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_132
timestamp 1698431365
transform 1 0 16128 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_136
timestamp 1698431365
transform 1 0 16576 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_142
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_146
timestamp 1698431365
transform 1 0 17696 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_151
timestamp 1698431365
transform 1 0 18256 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_183
timestamp 1698431365
transform 1 0 21840 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_199
timestamp 1698431365
transform 1 0 23632 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_207
timestamp 1698431365
transform 1 0 24528 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_209
timestamp 1698431365
transform 1 0 24752 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_212
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_214
timestamp 1698431365
transform 1 0 25312 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_219
timestamp 1698431365
transform 1 0 25872 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_227
timestamp 1698431365
transform 1 0 26768 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_231
timestamp 1698431365
transform 1 0 27216 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_233
timestamp 1698431365
transform 1 0 27440 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_263
timestamp 1698431365
transform 1 0 30800 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_265
timestamp 1698431365
transform 1 0 31024 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_268
timestamp 1698431365
transform 1 0 31360 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_270
timestamp 1698431365
transform 1 0 31584 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_282
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_286
timestamp 1698431365
transform 1 0 33376 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_294
timestamp 1698431365
transform 1 0 34272 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_347
timestamp 1698431365
transform 1 0 40208 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_349
timestamp 1698431365
transform 1 0 40432 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_352
timestamp 1698431365
transform 1 0 40768 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_368
timestamp 1698431365
transform 1 0 42560 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_372
timestamp 1698431365
transform 1 0 43008 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_376
timestamp 1698431365
transform 1 0 43456 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_380
timestamp 1698431365
transform 1 0 43904 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_382
timestamp 1698431365
transform 1 0 44128 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_385
timestamp 1698431365
transform 1 0 44464 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_389
timestamp 1698431365
transform 1 0 44912 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_422
timestamp 1698431365
transform 1 0 48608 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_481
timestamp 1698431365
transform 1 0 55216 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_489
timestamp 1698431365
transform 1 0 56112 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_492
timestamp 1698431365
transform 1 0 56448 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_494
timestamp 1698431365
transform 1 0 56672 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_499
timestamp 1698431365
transform 1 0 57232 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_507
timestamp 1698431365
transform 1 0 58128 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_2
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698431365
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_37
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_45
timestamp 1698431365
transform 1 0 6384 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_49
timestamp 1698431365
transform 1 0 6832 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_51
timestamp 1698431365
transform 1 0 7056 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_84
timestamp 1698431365
transform 1 0 10752 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_100
timestamp 1698431365
transform 1 0 12544 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_104
timestamp 1698431365
transform 1 0 12992 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_107
timestamp 1698431365
transform 1 0 13328 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_111
timestamp 1698431365
transform 1 0 13776 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_113
timestamp 1698431365
transform 1 0 14000 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_139
timestamp 1698431365
transform 1 0 16912 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_141
timestamp 1698431365
transform 1 0 17136 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_171
timestamp 1698431365
transform 1 0 20496 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_177
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_185
timestamp 1698431365
transform 1 0 22064 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_189
timestamp 1698431365
transform 1 0 22512 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_234
timestamp 1698431365
transform 1 0 27552 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_238
timestamp 1698431365
transform 1 0 28000 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_242
timestamp 1698431365
transform 1 0 28448 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_244
timestamp 1698431365
transform 1 0 28672 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_247
timestamp 1698431365
transform 1 0 29008 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_255
timestamp 1698431365
transform 1 0 29904 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_297
timestamp 1698431365
transform 1 0 34608 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_305
timestamp 1698431365
transform 1 0 35504 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_309
timestamp 1698431365
transform 1 0 35952 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_314
timestamp 1698431365
transform 1 0 36512 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_317
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_321
timestamp 1698431365
transform 1 0 37296 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_323
timestamp 1698431365
transform 1 0 37520 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_353
timestamp 1698431365
transform 1 0 40880 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_383
timestamp 1698431365
transform 1 0 44240 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_437
timestamp 1698431365
transform 1 0 50288 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_441
timestamp 1698431365
transform 1 0 50736 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_445
timestamp 1698431365
transform 1 0 51184 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_477
timestamp 1698431365
transform 1 0 54768 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_479
timestamp 1698431365
transform 1 0 54992 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_2
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_66
timestamp 1698431365
transform 1 0 8736 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_83
timestamp 1698431365
transform 1 0 10640 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_85
timestamp 1698431365
transform 1 0 10864 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_90
timestamp 1698431365
transform 1 0 11424 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_98
timestamp 1698431365
transform 1 0 12320 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_102
timestamp 1698431365
transform 1 0 12768 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_109
timestamp 1698431365
transform 1 0 13552 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_113
timestamp 1698431365
transform 1 0 14000 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_142
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_158
timestamp 1698431365
transform 1 0 19040 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_160
timestamp 1698431365
transform 1 0 19264 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_175
timestamp 1698431365
transform 1 0 20944 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_179
timestamp 1698431365
transform 1 0 21392 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_206
timestamp 1698431365
transform 1 0 24416 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_259
timestamp 1698431365
transform 1 0 30352 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_267
timestamp 1698431365
transform 1 0 31248 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_286
timestamp 1698431365
transform 1 0 33376 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_290
timestamp 1698431365
transform 1 0 33824 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_298
timestamp 1698431365
transform 1 0 34720 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_410
timestamp 1698431365
transform 1 0 47264 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_418
timestamp 1698431365
transform 1 0 48160 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_422
timestamp 1698431365
transform 1 0 48608 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_424
timestamp 1698431365
transform 1 0 48832 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_437
timestamp 1698431365
transform 1 0 50288 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_439
timestamp 1698431365
transform 1 0 50512 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_508
timestamp 1698431365
transform 1 0 58240 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_2
timestamp 1698431365
transform 1 0 1568 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_34
timestamp 1698431365
transform 1 0 5152 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_37
timestamp 1698431365
transform 1 0 5488 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_41
timestamp 1698431365
transform 1 0 5936 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_55
timestamp 1698431365
transform 1 0 7504 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_59
timestamp 1698431365
transform 1 0 7952 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_66
timestamp 1698431365
transform 1 0 8736 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_82
timestamp 1698431365
transform 1 0 10528 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_86
timestamp 1698431365
transform 1 0 10976 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_104
timestamp 1698431365
transform 1 0 12992 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_107
timestamp 1698431365
transform 1 0 13328 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_123
timestamp 1698431365
transform 1 0 15120 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_139
timestamp 1698431365
transform 1 0 16912 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_147
timestamp 1698431365
transform 1 0 17808 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_149
timestamp 1698431365
transform 1 0 18032 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_156
timestamp 1698431365
transform 1 0 18816 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_164
timestamp 1698431365
transform 1 0 19712 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_168
timestamp 1698431365
transform 1 0 20160 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_171
timestamp 1698431365
transform 1 0 20496 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_177
timestamp 1698431365
transform 1 0 21168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_179
timestamp 1698431365
transform 1 0 21392 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_231
timestamp 1698431365
transform 1 0 27216 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_239
timestamp 1698431365
transform 1 0 28112 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_243
timestamp 1698431365
transform 1 0 28560 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_257
timestamp 1698431365
transform 1 0 30128 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_261
timestamp 1698431365
transform 1 0 30576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_313
timestamp 1698431365
transform 1 0 36400 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_317
timestamp 1698431365
transform 1 0 36848 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_321
timestamp 1698431365
transform 1 0 37296 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_329
timestamp 1698431365
transform 1 0 38192 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_337
timestamp 1698431365
transform 1 0 39088 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_341
timestamp 1698431365
transform 1 0 39536 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_347
timestamp 1698431365
transform 1 0 40208 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_349
timestamp 1698431365
transform 1 0 40432 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_352
timestamp 1698431365
transform 1 0 40768 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_368
timestamp 1698431365
transform 1 0 42560 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_376
timestamp 1698431365
transform 1 0 43456 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_384
timestamp 1698431365
transform 1 0 44352 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_387
timestamp 1698431365
transform 1 0 44688 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_403
timestamp 1698431365
transform 1 0 46480 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_407
timestamp 1698431365
transform 1 0 46928 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_453
timestamp 1698431365
transform 1 0 52080 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_505
timestamp 1698431365
transform 1 0 57904 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_2
timestamp 1698431365
transform 1 0 1568 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_18
timestamp 1698431365
transform 1 0 3360 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_22
timestamp 1698431365
transform 1 0 3808 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_59
timestamp 1698431365
transform 1 0 7952 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_69
timestamp 1698431365
transform 1 0 9072 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_72
timestamp 1698431365
transform 1 0 9408 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_76
timestamp 1698431365
transform 1 0 9856 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_106
timestamp 1698431365
transform 1 0 13216 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_114
timestamp 1698431365
transform 1 0 14112 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_118
timestamp 1698431365
transform 1 0 14560 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_126
timestamp 1698431365
transform 1 0 15456 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_130
timestamp 1698431365
transform 1 0 15904 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_135
timestamp 1698431365
transform 1 0 16464 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_139
timestamp 1698431365
transform 1 0 16912 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_142
timestamp 1698431365
transform 1 0 17248 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_146
timestamp 1698431365
transform 1 0 17696 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_154
timestamp 1698431365
transform 1 0 18592 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_207
timestamp 1698431365
transform 1 0 24528 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_209
timestamp 1698431365
transform 1 0 24752 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_212
timestamp 1698431365
transform 1 0 25088 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_232
timestamp 1698431365
transform 1 0 27328 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_274
timestamp 1698431365
transform 1 0 32032 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_278
timestamp 1698431365
transform 1 0 32480 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_287
timestamp 1698431365
transform 1 0 33488 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_291
timestamp 1698431365
transform 1 0 33936 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_295
timestamp 1698431365
transform 1 0 34384 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_303
timestamp 1698431365
transform 1 0 35280 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_306
timestamp 1698431365
transform 1 0 35616 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_310
timestamp 1698431365
transform 1 0 36064 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_312
timestamp 1698431365
transform 1 0 36288 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_322
timestamp 1698431365
transform 1 0 37408 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_338
timestamp 1698431365
transform 1 0 39200 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_346
timestamp 1698431365
transform 1 0 40096 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_367
timestamp 1698431365
transform 1 0 42448 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_371
timestamp 1698431365
transform 1 0 42896 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_387
timestamp 1698431365
transform 1 0 44688 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_395
timestamp 1698431365
transform 1 0 45584 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_397
timestamp 1698431365
transform 1 0 45808 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_406
timestamp 1698431365
transform 1 0 46816 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_414
timestamp 1698431365
transform 1 0 47712 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_418
timestamp 1698431365
transform 1 0 48160 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_422
timestamp 1698431365
transform 1 0 48608 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_440
timestamp 1698431365
transform 1 0 50624 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_487
timestamp 1698431365
transform 1 0 55888 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_489
timestamp 1698431365
transform 1 0 56112 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_500
timestamp 1698431365
transform 1 0 57344 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_2
timestamp 1698431365
transform 1 0 1568 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_34
timestamp 1698431365
transform 1 0 5152 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_87
timestamp 1698431365
transform 1 0 11088 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_91
timestamp 1698431365
transform 1 0 11536 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_99
timestamp 1698431365
transform 1 0 12432 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_103
timestamp 1698431365
transform 1 0 12880 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_107
timestamp 1698431365
transform 1 0 13328 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_115
timestamp 1698431365
transform 1 0 14224 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_119
timestamp 1698431365
transform 1 0 14672 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_126
timestamp 1698431365
transform 1 0 15456 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_136
timestamp 1698431365
transform 1 0 16576 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_142
timestamp 1698431365
transform 1 0 17248 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_152
timestamp 1698431365
transform 1 0 18368 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_156
timestamp 1698431365
transform 1 0 18816 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_160
timestamp 1698431365
transform 1 0 19264 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_173
timestamp 1698431365
transform 1 0 20720 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_177
timestamp 1698431365
transform 1 0 21168 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_206
timestamp 1698431365
transform 1 0 24416 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_263
timestamp 1698431365
transform 1 0 30800 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_293
timestamp 1698431365
transform 1 0 34160 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_308
timestamp 1698431365
transform 1 0 35840 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_310
timestamp 1698431365
transform 1 0 36064 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_317
timestamp 1698431365
transform 1 0 36848 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_319
timestamp 1698431365
transform 1 0 37072 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_336
timestamp 1698431365
transform 1 0 38976 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_344
timestamp 1698431365
transform 1 0 39872 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_348
timestamp 1698431365
transform 1 0 40320 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_354
timestamp 1698431365
transform 1 0 40992 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_370
timestamp 1698431365
transform 1 0 42784 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_374
timestamp 1698431365
transform 1 0 43232 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_379
timestamp 1698431365
transform 1 0 43792 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_383
timestamp 1698431365
transform 1 0 44240 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_387
timestamp 1698431365
transform 1 0 44688 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_442
timestamp 1698431365
transform 1 0 50848 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_446
timestamp 1698431365
transform 1 0 51296 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_454
timestamp 1698431365
transform 1 0 52192 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_457
timestamp 1698431365
transform 1 0 52528 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_475
timestamp 1698431365
transform 1 0 54544 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_479
timestamp 1698431365
transform 1 0 54992 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_2
timestamp 1698431365
transform 1 0 1568 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_34
timestamp 1698431365
transform 1 0 5152 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_38
timestamp 1698431365
transform 1 0 5600 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_40
timestamp 1698431365
transform 1 0 5824 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_78
timestamp 1698431365
transform 1 0 10080 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_110
timestamp 1698431365
transform 1 0 13664 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_142
timestamp 1698431365
transform 1 0 17248 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_175
timestamp 1698431365
transform 1 0 20944 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_209
timestamp 1698431365
transform 1 0 24752 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_216
timestamp 1698431365
transform 1 0 25536 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_277
timestamp 1698431365
transform 1 0 32368 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_279
timestamp 1698431365
transform 1 0 32592 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_282
timestamp 1698431365
transform 1 0 32928 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_362
timestamp 1698431365
transform 1 0 41888 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_366
timestamp 1698431365
transform 1 0 42336 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_419
timestamp 1698431365
transform 1 0 48272 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_422
timestamp 1698431365
transform 1 0 48608 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_430
timestamp 1698431365
transform 1 0 49504 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_469
timestamp 1698431365
transform 1 0 53872 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_485
timestamp 1698431365
transform 1 0 55664 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_489
timestamp 1698431365
transform 1 0 56112 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_500
timestamp 1698431365
transform 1 0 57344 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_508
timestamp 1698431365
transform 1 0 58240 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_2
timestamp 1698431365
transform 1 0 1568 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_34
timestamp 1698431365
transform 1 0 5152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_37
timestamp 1698431365
transform 1 0 5488 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_53
timestamp 1698431365
transform 1 0 7280 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_57
timestamp 1698431365
transform 1 0 7728 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_63
timestamp 1698431365
transform 1 0 8400 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_95
timestamp 1698431365
transform 1 0 11984 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_103
timestamp 1698431365
transform 1 0 12880 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_107
timestamp 1698431365
transform 1 0 13328 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_123
timestamp 1698431365
transform 1 0 15120 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_155
timestamp 1698431365
transform 1 0 18704 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_163
timestamp 1698431365
transform 1 0 19600 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_171
timestamp 1698431365
transform 1 0 20496 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_188
timestamp 1698431365
transform 1 0 22400 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_220
timestamp 1698431365
transform 1 0 25984 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_238
timestamp 1698431365
transform 1 0 28000 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_242
timestamp 1698431365
transform 1 0 28448 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_244
timestamp 1698431365
transform 1 0 28672 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_247
timestamp 1698431365
transform 1 0 29008 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_251
timestamp 1698431365
transform 1 0 29456 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_257
timestamp 1698431365
transform 1 0 30128 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_273
timestamp 1698431365
transform 1 0 31920 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_281
timestamp 1698431365
transform 1 0 32816 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_285
timestamp 1698431365
transform 1 0 33264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_346
timestamp 1698431365
transform 1 0 40096 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_361
timestamp 1698431365
transform 1 0 41776 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_377
timestamp 1698431365
transform 1 0 43568 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_387
timestamp 1698431365
transform 1 0 44688 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_389
timestamp 1698431365
transform 1 0 44912 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_398
timestamp 1698431365
transform 1 0 45920 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_414
timestamp 1698431365
transform 1 0 47712 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_416
timestamp 1698431365
transform 1 0 47936 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_423
timestamp 1698431365
transform 1 0 48720 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_457
timestamp 1698431365
transform 1 0 52528 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_467
timestamp 1698431365
transform 1 0 53648 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_475
timestamp 1698431365
transform 1 0 54544 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_479
timestamp 1698431365
transform 1 0 54992 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_2
timestamp 1698431365
transform 1 0 1568 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_66
timestamp 1698431365
transform 1 0 8736 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_72
timestamp 1698431365
transform 1 0 9408 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_117
timestamp 1698431365
transform 1 0 14448 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_133
timestamp 1698431365
transform 1 0 16240 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_137
timestamp 1698431365
transform 1 0 16688 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_139
timestamp 1698431365
transform 1 0 16912 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_142
timestamp 1698431365
transform 1 0 17248 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_158
timestamp 1698431365
transform 1 0 19040 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_162
timestamp 1698431365
transform 1 0 19488 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_165
timestamp 1698431365
transform 1 0 19824 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_197
timestamp 1698431365
transform 1 0 23408 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_205
timestamp 1698431365
transform 1 0 24304 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_209
timestamp 1698431365
transform 1 0 24752 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_212
timestamp 1698431365
transform 1 0 25088 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_214
timestamp 1698431365
transform 1 0 25312 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_230
timestamp 1698431365
transform 1 0 27104 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_246
timestamp 1698431365
transform 1 0 28896 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_254
timestamp 1698431365
transform 1 0 29792 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_256
timestamp 1698431365
transform 1 0 30016 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_270
timestamp 1698431365
transform 1 0 31584 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_274
timestamp 1698431365
transform 1 0 32032 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_278
timestamp 1698431365
transform 1 0 32480 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_282
timestamp 1698431365
transform 1 0 32928 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_298
timestamp 1698431365
transform 1 0 34720 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_306
timestamp 1698431365
transform 1 0 35616 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_310
timestamp 1698431365
transform 1 0 36064 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_312
timestamp 1698431365
transform 1 0 36288 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_317
timestamp 1698431365
transform 1 0 36848 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_321
timestamp 1698431365
transform 1 0 37296 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_325
timestamp 1698431365
transform 1 0 37744 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_341
timestamp 1698431365
transform 1 0 39536 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_349
timestamp 1698431365
transform 1 0 40432 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_368
timestamp 1698431365
transform 1 0 42560 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_400
timestamp 1698431365
transform 1 0 46144 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_416
timestamp 1698431365
transform 1 0 47936 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_434
timestamp 1698431365
transform 1 0 49952 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_440
timestamp 1698431365
transform 1 0 50624 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_444
timestamp 1698431365
transform 1 0 51072 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_452
timestamp 1698431365
transform 1 0 51968 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_456
timestamp 1698431365
transform 1 0 52416 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_459
timestamp 1698431365
transform 1 0 52752 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_475
timestamp 1698431365
transform 1 0 54544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_477
timestamp 1698431365
transform 1 0 54768 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_497
timestamp 1698431365
transform 1 0 57008 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_2
timestamp 1698431365
transform 1 0 1568 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_34
timestamp 1698431365
transform 1 0 5152 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_37
timestamp 1698431365
transform 1 0 5488 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_101
timestamp 1698431365
transform 1 0 12656 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_107
timestamp 1698431365
transform 1 0 13328 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_111
timestamp 1698431365
transform 1 0 13776 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_171
timestamp 1698431365
transform 1 0 20496 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_183
timestamp 1698431365
transform 1 0 21840 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_187
timestamp 1698431365
transform 1 0 22288 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_218
timestamp 1698431365
transform 1 0 25760 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_232
timestamp 1698431365
transform 1 0 27328 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_236
timestamp 1698431365
transform 1 0 27776 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_238
timestamp 1698431365
transform 1 0 28000 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_247
timestamp 1698431365
transform 1 0 29008 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_249
timestamp 1698431365
transform 1 0 29232 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_262
timestamp 1698431365
transform 1 0 30688 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_264
timestamp 1698431365
transform 1 0 30912 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_294
timestamp 1698431365
transform 1 0 34272 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_302
timestamp 1698431365
transform 1 0 35168 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_306
timestamp 1698431365
transform 1 0 35616 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_317
timestamp 1698431365
transform 1 0 36848 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_321
timestamp 1698431365
transform 1 0 37296 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_387
timestamp 1698431365
transform 1 0 44688 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_389
timestamp 1698431365
transform 1 0 44912 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_396
timestamp 1698431365
transform 1 0 45696 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_402
timestamp 1698431365
transform 1 0 46368 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_418
timestamp 1698431365
transform 1 0 48160 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_426
timestamp 1698431365
transform 1 0 49056 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_452
timestamp 1698431365
transform 1 0 51968 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_454
timestamp 1698431365
transform 1 0 52192 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_457
timestamp 1698431365
transform 1 0 52528 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_2
timestamp 1698431365
transform 1 0 1568 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_66
timestamp 1698431365
transform 1 0 8736 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_72
timestamp 1698431365
transform 1 0 9408 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_136
timestamp 1698431365
transform 1 0 16576 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_142
timestamp 1698431365
transform 1 0 17248 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_150
timestamp 1698431365
transform 1 0 18144 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_154
timestamp 1698431365
transform 1 0 18592 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_179
timestamp 1698431365
transform 1 0 21392 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_187
timestamp 1698431365
transform 1 0 22288 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_189
timestamp 1698431365
transform 1 0 22512 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_204
timestamp 1698431365
transform 1 0 24192 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_208
timestamp 1698431365
transform 1 0 24640 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_212
timestamp 1698431365
transform 1 0 25088 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_216
timestamp 1698431365
transform 1 0 25536 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_226
timestamp 1698431365
transform 1 0 26656 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_234
timestamp 1698431365
transform 1 0 27552 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_236
timestamp 1698431365
transform 1 0 27776 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_243
timestamp 1698431365
transform 1 0 28560 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_277
timestamp 1698431365
transform 1 0 32368 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_279
timestamp 1698431365
transform 1 0 32592 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_282
timestamp 1698431365
transform 1 0 32928 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_286
timestamp 1698431365
transform 1 0 33376 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_290
timestamp 1698431365
transform 1 0 33824 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_327
timestamp 1698431365
transform 1 0 37968 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_331
timestamp 1698431365
transform 1 0 38416 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_347
timestamp 1698431365
transform 1 0 40208 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_349
timestamp 1698431365
transform 1 0 40432 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_352
timestamp 1698431365
transform 1 0 40768 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_360
timestamp 1698431365
transform 1 0 41664 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_364
timestamp 1698431365
transform 1 0 42112 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_370
timestamp 1698431365
transform 1 0 42784 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_372
timestamp 1698431365
transform 1 0 43008 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_408
timestamp 1698431365
transform 1 0 47040 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_416
timestamp 1698431365
transform 1 0 47936 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_477
timestamp 1698431365
transform 1 0 54768 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_481
timestamp 1698431365
transform 1 0 55216 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_492
timestamp 1698431365
transform 1 0 56448 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_508
timestamp 1698431365
transform 1 0 58240 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_2
timestamp 1698431365
transform 1 0 1568 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_34
timestamp 1698431365
transform 1 0 5152 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_37
timestamp 1698431365
transform 1 0 5488 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_101
timestamp 1698431365
transform 1 0 12656 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_107
timestamp 1698431365
transform 1 0 13328 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_115
timestamp 1698431365
transform 1 0 14224 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_119
timestamp 1698431365
transform 1 0 14672 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_121
timestamp 1698431365
transform 1 0 14896 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_151
timestamp 1698431365
transform 1 0 18256 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_159
timestamp 1698431365
transform 1 0 19152 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_169
timestamp 1698431365
transform 1 0 20272 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_173
timestamp 1698431365
transform 1 0 20720 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_177
timestamp 1698431365
transform 1 0 21168 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_185
timestamp 1698431365
transform 1 0 22064 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_189
timestamp 1698431365
transform 1 0 22512 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_204
timestamp 1698431365
transform 1 0 24192 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_208
timestamp 1698431365
transform 1 0 24640 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_247
timestamp 1698431365
transform 1 0 29008 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_263
timestamp 1698431365
transform 1 0 30800 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_265
timestamp 1698431365
transform 1 0 31024 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_274
timestamp 1698431365
transform 1 0 32032 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_278
timestamp 1698431365
transform 1 0 32480 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_294
timestamp 1698431365
transform 1 0 34272 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_302
timestamp 1698431365
transform 1 0 35168 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_314
timestamp 1698431365
transform 1 0 36512 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_323
timestamp 1698431365
transform 1 0 37520 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_325
timestamp 1698431365
transform 1 0 37744 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_361
timestamp 1698431365
transform 1 0 41776 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_363
timestamp 1698431365
transform 1 0 42000 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_372
timestamp 1698431365
transform 1 0 43008 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_376
timestamp 1698431365
transform 1 0 43456 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_383
timestamp 1698431365
transform 1 0 44240 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_403
timestamp 1698431365
transform 1 0 46480 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_411
timestamp 1698431365
transform 1 0 47376 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_415
timestamp 1698431365
transform 1 0 47824 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_439
timestamp 1698431365
transform 1 0 50512 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_447
timestamp 1698431365
transform 1 0 51408 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_457
timestamp 1698431365
transform 1 0 52528 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_473
timestamp 1698431365
transform 1 0 54320 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_477
timestamp 1698431365
transform 1 0 54768 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_479
timestamp 1698431365
transform 1 0 54992 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_2
timestamp 1698431365
transform 1 0 1568 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_66
timestamp 1698431365
transform 1 0 8736 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_72
timestamp 1698431365
transform 1 0 9408 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_136
timestamp 1698431365
transform 1 0 16576 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_142
timestamp 1698431365
transform 1 0 17248 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_212
timestamp 1698431365
transform 1 0 25088 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_220
timestamp 1698431365
transform 1 0 25984 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_225
timestamp 1698431365
transform 1 0 26544 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_233
timestamp 1698431365
transform 1 0 27440 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_243
timestamp 1698431365
transform 1 0 28560 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_259
timestamp 1698431365
transform 1 0 30352 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_267
timestamp 1698431365
transform 1 0 31248 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_274
timestamp 1698431365
transform 1 0 32032 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_278
timestamp 1698431365
transform 1 0 32480 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_282
timestamp 1698431365
transform 1 0 32928 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_298
timestamp 1698431365
transform 1 0 34720 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_349
timestamp 1698431365
transform 1 0 40432 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_360
timestamp 1698431365
transform 1 0 41664 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_392
timestamp 1698431365
transform 1 0 45248 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_400
timestamp 1698431365
transform 1 0 46144 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_410
timestamp 1698431365
transform 1 0 47264 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_418
timestamp 1698431365
transform 1 0 48160 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_422
timestamp 1698431365
transform 1 0 48608 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_430
timestamp 1698431365
transform 1 0 49504 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_442
timestamp 1698431365
transform 1 0 50848 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_474
timestamp 1698431365
transform 1 0 54432 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_485
timestamp 1698431365
transform 1 0 55664 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_489
timestamp 1698431365
transform 1 0 56112 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_500
timestamp 1698431365
transform 1 0 57344 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_508
timestamp 1698431365
transform 1 0 58240 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_2
timestamp 1698431365
transform 1 0 1568 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_34
timestamp 1698431365
transform 1 0 5152 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_37
timestamp 1698431365
transform 1 0 5488 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_101
timestamp 1698431365
transform 1 0 12656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_107
timestamp 1698431365
transform 1 0 13328 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_139
timestamp 1698431365
transform 1 0 16912 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_155
timestamp 1698431365
transform 1 0 18704 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_163
timestamp 1698431365
transform 1 0 19600 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_187
timestamp 1698431365
transform 1 0 22288 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_195
timestamp 1698431365
transform 1 0 23184 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_211
timestamp 1698431365
transform 1 0 24976 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_224
timestamp 1698431365
transform 1 0 26432 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_247
timestamp 1698431365
transform 1 0 29008 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_256
timestamp 1698431365
transform 1 0 30016 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_295
timestamp 1698431365
transform 1 0 34384 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_303
timestamp 1698431365
transform 1 0 35280 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_325
timestamp 1698431365
transform 1 0 37744 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_329
timestamp 1698431365
transform 1 0 38192 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_333
timestamp 1698431365
transform 1 0 38640 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_335
timestamp 1698431365
transform 1 0 38864 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_350
timestamp 1698431365
transform 1 0 40544 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_365
timestamp 1698431365
transform 1 0 42224 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_369
timestamp 1698431365
transform 1 0 42672 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_378
timestamp 1698431365
transform 1 0 43680 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_382
timestamp 1698431365
transform 1 0 44128 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_384
timestamp 1698431365
transform 1 0 44352 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_387
timestamp 1698431365
transform 1 0 44688 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_419
timestamp 1698431365
transform 1 0 48272 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_425
timestamp 1698431365
transform 1 0 48944 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_433
timestamp 1698431365
transform 1 0 49840 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_451
timestamp 1698431365
transform 1 0 51856 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_475
timestamp 1698431365
transform 1 0 54544 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_477
timestamp 1698431365
transform 1 0 54768 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_492
timestamp 1698431365
transform 1 0 56448 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_508
timestamp 1698431365
transform 1 0 58240 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_2
timestamp 1698431365
transform 1 0 1568 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_66
timestamp 1698431365
transform 1 0 8736 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_72
timestamp 1698431365
transform 1 0 9408 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_136
timestamp 1698431365
transform 1 0 16576 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_195
timestamp 1698431365
transform 1 0 23184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_203
timestamp 1698431365
transform 1 0 24080 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_207
timestamp 1698431365
transform 1 0 24528 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_262
timestamp 1698431365
transform 1 0 30688 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_266
timestamp 1698431365
transform 1 0 31136 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_275
timestamp 1698431365
transform 1 0 32144 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_279
timestamp 1698431365
transform 1 0 32592 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_282
timestamp 1698431365
transform 1 0 32928 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_298
timestamp 1698431365
transform 1 0 34720 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_306
timestamp 1698431365
transform 1 0 35616 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_310
timestamp 1698431365
transform 1 0 36064 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_312
timestamp 1698431365
transform 1 0 36288 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_319
timestamp 1698431365
transform 1 0 37072 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_335
timestamp 1698431365
transform 1 0 38864 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_343
timestamp 1698431365
transform 1 0 39760 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_366
timestamp 1698431365
transform 1 0 42336 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_396
timestamp 1698431365
transform 1 0 45696 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_415
timestamp 1698431365
transform 1 0 47824 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_417
timestamp 1698431365
transform 1 0 48048 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_478
timestamp 1698431365
transform 1 0 54880 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_486
timestamp 1698431365
transform 1 0 55776 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_492
timestamp 1698431365
transform 1 0 56448 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_508
timestamp 1698431365
transform 1 0 58240 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_2
timestamp 1698431365
transform 1 0 1568 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_34
timestamp 1698431365
transform 1 0 5152 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_37
timestamp 1698431365
transform 1 0 5488 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_101
timestamp 1698431365
transform 1 0 12656 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_107
timestamp 1698431365
transform 1 0 13328 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_139
timestamp 1698431365
transform 1 0 16912 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_172
timestamp 1698431365
transform 1 0 20608 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_174
timestamp 1698431365
transform 1 0 20832 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_185
timestamp 1698431365
transform 1 0 22064 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_189
timestamp 1698431365
transform 1 0 22512 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_220
timestamp 1698431365
transform 1 0 25984 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_224
timestamp 1698431365
transform 1 0 26432 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_226
timestamp 1698431365
transform 1 0 26656 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_237
timestamp 1698431365
transform 1 0 27888 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_276
timestamp 1698431365
transform 1 0 32256 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_284
timestamp 1698431365
transform 1 0 33152 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_317
timestamp 1698431365
transform 1 0 36848 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_319
timestamp 1698431365
transform 1 0 37072 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_349
timestamp 1698431365
transform 1 0 40432 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_358
timestamp 1698431365
transform 1 0 41440 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_362
timestamp 1698431365
transform 1 0 41888 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_364
timestamp 1698431365
transform 1 0 42112 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_371
timestamp 1698431365
transform 1 0 42896 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_379
timestamp 1698431365
transform 1 0 43792 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_383
timestamp 1698431365
transform 1 0 44240 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_387
timestamp 1698431365
transform 1 0 44688 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_395
timestamp 1698431365
transform 1 0 45584 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_486
timestamp 1698431365
transform 1 0 55776 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_494
timestamp 1698431365
transform 1 0 56672 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_504
timestamp 1698431365
transform 1 0 57792 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_508
timestamp 1698431365
transform 1 0 58240 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_2
timestamp 1698431365
transform 1 0 1568 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_36
timestamp 1698431365
transform 1 0 5376 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_70
timestamp 1698431365
transform 1 0 9184 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_104
timestamp 1698431365
transform 1 0 12992 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_138
timestamp 1698431365
transform 1 0 16800 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_172
timestamp 1698431365
transform 1 0 20608 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_180
timestamp 1698431365
transform 1 0 21504 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_184
timestamp 1698431365
transform 1 0 21952 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_186
timestamp 1698431365
transform 1 0 22176 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_197
timestamp 1698431365
transform 1 0 23408 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_201
timestamp 1698431365
transform 1 0 23856 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_203
timestamp 1698431365
transform 1 0 24080 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_206
timestamp 1698431365
transform 1 0 24416 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_222
timestamp 1698431365
transform 1 0 26208 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_234
timestamp 1698431365
transform 1 0 27552 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_240
timestamp 1698431365
transform 1 0 28224 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_274
timestamp 1698431365
transform 1 0 32032 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_308
timestamp 1698431365
transform 1 0 35840 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_316
timestamp 1698431365
transform 1 0 36736 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_320
timestamp 1698431365
transform 1 0 37184 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_331
timestamp 1698431365
transform 1 0 38416 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_339
timestamp 1698431365
transform 1 0 39312 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_342
timestamp 1698431365
transform 1 0 39648 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_376
timestamp 1698431365
transform 1 0 43456 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_410
timestamp 1698431365
transform 1 0 47264 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_444
timestamp 1698431365
transform 1 0 51072 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_452
timestamp 1698431365
transform 1 0 51968 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_454
timestamp 1698431365
transform 1 0 52192 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_463
timestamp 1698431365
transform 1 0 53200 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_471
timestamp 1698431365
transform 1 0 54096 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_475
timestamp 1698431365
transform 1 0 54544 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_478
timestamp 1698431365
transform 1 0 54880 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_494
timestamp 1698431365
transform 1 0 56672 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_498
timestamp 1698431365
transform 1 0 57120 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_500
timestamp 1698431365
transform 1 0 57344 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input1
timestamp 1698431365
transform -1 0 58352 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform -1 0 58352 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input3
timestamp 1698431365
transform -1 0 58352 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input4
timestamp 1698431365
transform -1 0 58352 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input5
timestamp 1698431365
transform -1 0 58352 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input6
timestamp 1698431365
transform -1 0 58352 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input7
timestamp 1698431365
transform -1 0 58352 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input8
timestamp 1698431365
transform -1 0 58352 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input9
timestamp 1698431365
transform -1 0 58352 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input10
timestamp 1698431365
transform -1 0 58352 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input11
timestamp 1698431365
transform 1 0 37520 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input12
timestamp 1698431365
transform -1 0 53200 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input13
timestamp 1698431365
transform 1 0 22512 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22960 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698431365
transform 1 0 24976 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698431365
transform 1 0 36512 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698431365
transform 1 0 41552 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698431365
transform 1 0 44240 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698431365
transform 1 0 47264 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698431365
transform -1 0 20384 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698431365
transform 1 0 20944 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_68 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 58576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_69
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 58576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_70
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 58576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_71
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 58576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_72
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 58576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_73
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 58576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_74
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 58576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_75
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 58576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_76
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 58576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_77
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 58576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_78
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 58576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_79
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 58576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_80
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 58576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_81
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 58576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_82
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 58576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_83
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 58576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_84
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 58576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_85
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 58576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_86
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 58576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_87
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 58576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_88
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 58576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_89
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 58576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_90
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 58576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_91
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 58576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_92
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 58576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_93
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 58576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_94
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 58576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_95
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 58576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_96
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 58576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_97
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 58576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_98
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 58576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_99
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 58576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_100
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 58576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_101
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 58576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_102
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 58576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_103
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 58576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_104
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 58576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_105
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 58576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_106
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 58576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_107
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 58576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_108
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 58576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_109
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 58576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_110
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 58576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_111
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 58576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_112
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 58576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_113
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 58576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_114
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 58576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_115
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 58576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_116
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 58576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_117
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 58576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_118
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 58576 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_119
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 58576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_120
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 58576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_121
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 58576 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_122
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 58576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_123
timestamp 1698431365
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698431365
transform -1 0 58576 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_124
timestamp 1698431365
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698431365
transform -1 0 58576 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_125
timestamp 1698431365
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698431365
transform -1 0 58576 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_126
timestamp 1698431365
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698431365
transform -1 0 58576 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_127
timestamp 1698431365
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698431365
transform -1 0 58576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_128
timestamp 1698431365
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698431365
transform -1 0 58576 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_129
timestamp 1698431365
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698431365
transform -1 0 58576 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_130
timestamp 1698431365
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1698431365
transform -1 0 58576 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_131
timestamp 1698431365
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1698431365
transform -1 0 58576 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_132
timestamp 1698431365
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1698431365
transform -1 0 58576 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_133
timestamp 1698431365
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1698431365
transform -1 0 58576 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_134
timestamp 1698431365
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1698431365
transform -1 0 58576 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_135
timestamp 1698431365
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1698431365
transform -1 0 58576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_136 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_137
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_138
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_139
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_140
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_141
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_142
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_143
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_144
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_145
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_146
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_147
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_148
timestamp 1698431365
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_149
timestamp 1698431365
transform 1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_150
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_151
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_152
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_153
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_154
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_155
timestamp 1698431365
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_156
timestamp 1698431365
transform 1 0 56224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_157
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_158
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_159
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_160
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_161
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_162
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_163
timestamp 1698431365
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_164
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_165
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_166
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_167
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_168
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_169
timestamp 1698431365
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_170
timestamp 1698431365
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_171
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_172
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_173
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_174
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_175
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_176
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_177
timestamp 1698431365
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_178
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_179
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_180
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_181
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_182
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_183
timestamp 1698431365
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_184
timestamp 1698431365
transform 1 0 56224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_185
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_186
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_187
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_188
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_189
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_190
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_191
timestamp 1698431365
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_192
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_193
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_194
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_195
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_196
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_197
timestamp 1698431365
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_198
timestamp 1698431365
transform 1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_199
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_200
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_201
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_202
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_203
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_204
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_205
timestamp 1698431365
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_206
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_207
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_208
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_209
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_210
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_211
timestamp 1698431365
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_212
timestamp 1698431365
transform 1 0 56224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_213
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_214
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_215
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_216
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_217
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_218
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_219
timestamp 1698431365
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_220
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_221
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_222
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_223
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_224
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_225
timestamp 1698431365
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_226
timestamp 1698431365
transform 1 0 56224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_227
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_228
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_229
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_230
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_231
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_232
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_233
timestamp 1698431365
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_234
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_235
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_236
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_237
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_238
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_239
timestamp 1698431365
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_240
timestamp 1698431365
transform 1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_241
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_242
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_243
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_244
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_245
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_246
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_247
timestamp 1698431365
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_248
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_249
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_250
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_251
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_252
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_253
timestamp 1698431365
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_254
timestamp 1698431365
transform 1 0 56224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_255
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_256
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_257
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_258
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_259
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_260
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_261
timestamp 1698431365
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_262
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_263
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_264
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_265
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_266
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_267
timestamp 1698431365
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_268
timestamp 1698431365
transform 1 0 56224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_269
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_270
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_271
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_272
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_273
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_274
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_275
timestamp 1698431365
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_276
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_277
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_278
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_279
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_280
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_281
timestamp 1698431365
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_282
timestamp 1698431365
transform 1 0 56224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_283
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_284
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_285
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_286
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_287
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_288
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_289
timestamp 1698431365
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_290
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_291
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_292
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_293
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_294
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_295
timestamp 1698431365
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_296
timestamp 1698431365
transform 1 0 56224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_297
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_298
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_299
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_300
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_301
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_302
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_303
timestamp 1698431365
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_304
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_305
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_306
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_307
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_308
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_309
timestamp 1698431365
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_310
timestamp 1698431365
transform 1 0 56224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_311
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_312
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_313
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_314
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_315
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_316
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_317
timestamp 1698431365
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_318
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_319
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_320
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_321
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_322
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_323
timestamp 1698431365
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_324
timestamp 1698431365
transform 1 0 56224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_325
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_326
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_327
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_328
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_329
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_330
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_331
timestamp 1698431365
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_332
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_333
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_334
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_335
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_336
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_337
timestamp 1698431365
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_338
timestamp 1698431365
transform 1 0 56224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_339
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_340
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_341
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_342
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_343
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_344
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_345
timestamp 1698431365
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_346
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_347
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_348
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_349
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_350
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_351
timestamp 1698431365
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_352
timestamp 1698431365
transform 1 0 56224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_353
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_354
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_355
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_356
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_357
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_358
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_359
timestamp 1698431365
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_360
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_361
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_362
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_363
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_364
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_365
timestamp 1698431365
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_366
timestamp 1698431365
transform 1 0 56224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_367
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_368
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_369
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_370
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_371
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_372
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_373
timestamp 1698431365
transform 1 0 52304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_374
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_375
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_376
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_377
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_378
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_379
timestamp 1698431365
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_380
timestamp 1698431365
transform 1 0 56224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_381
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_382
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_383
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_384
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_385
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_386
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_387
timestamp 1698431365
transform 1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_388
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_389
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_390
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_391
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_392
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_393
timestamp 1698431365
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_394
timestamp 1698431365
transform 1 0 56224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_395
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_396
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_397
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_398
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_399
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_400
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_401
timestamp 1698431365
transform 1 0 52304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_402
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_403
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_404
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_405
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_406
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_407
timestamp 1698431365
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_408
timestamp 1698431365
transform 1 0 56224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_409
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_410
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_411
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_412
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_413
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_414
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_415
timestamp 1698431365
transform 1 0 52304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_416
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_417
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_418
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_419
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_420
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_421
timestamp 1698431365
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_422
timestamp 1698431365
transform 1 0 56224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_423
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_424
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_425
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_426
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_427
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_428
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_429
timestamp 1698431365
transform 1 0 52304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_430
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_431
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_432
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_433
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_434
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_435
timestamp 1698431365
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_436
timestamp 1698431365
transform 1 0 56224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_437
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_438
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_439
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_440
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_441
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_442
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_443
timestamp 1698431365
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_444
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_445
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_446
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_447
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_448
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_449
timestamp 1698431365
transform 1 0 48384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_450
timestamp 1698431365
transform 1 0 56224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_451
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_452
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_453
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_454
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_455
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_456
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_457
timestamp 1698431365
transform 1 0 52304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_458
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_459
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_460
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_461
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_462
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_463
timestamp 1698431365
transform 1 0 48384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_464
timestamp 1698431365
transform 1 0 56224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_465
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_466
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_467
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_468
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_469
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_470
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_471
timestamp 1698431365
transform 1 0 52304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_472
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_473
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_474
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_475
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_476
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_477
timestamp 1698431365
transform 1 0 48384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_478
timestamp 1698431365
transform 1 0 56224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_479
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_480
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_481
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_482
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_483
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_484
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_485
timestamp 1698431365
transform 1 0 52304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_486
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_487
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_488
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_489
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_490
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_491
timestamp 1698431365
transform 1 0 48384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_492
timestamp 1698431365
transform 1 0 56224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_493
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_494
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_495
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_496
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_497
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_498
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_499
timestamp 1698431365
transform 1 0 52304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_500
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_501
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_502
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_503
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_504
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_505
timestamp 1698431365
transform 1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_506
timestamp 1698431365
transform 1 0 56224 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_507
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_508
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_509
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_510
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_511
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_512
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_513
timestamp 1698431365
transform 1 0 52304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_514
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_515
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_516
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_517
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_518
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_519
timestamp 1698431365
transform 1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_520
timestamp 1698431365
transform 1 0 56224 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_521
timestamp 1698431365
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_522
timestamp 1698431365
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_523
timestamp 1698431365
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_524
timestamp 1698431365
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_525
timestamp 1698431365
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_526
timestamp 1698431365
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_527
timestamp 1698431365
transform 1 0 52304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_528
timestamp 1698431365
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_529
timestamp 1698431365
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_530
timestamp 1698431365
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_531
timestamp 1698431365
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_532
timestamp 1698431365
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_533
timestamp 1698431365
transform 1 0 48384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_534
timestamp 1698431365
transform 1 0 56224 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_535
timestamp 1698431365
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_536
timestamp 1698431365
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_537
timestamp 1698431365
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_538
timestamp 1698431365
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_539
timestamp 1698431365
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_540
timestamp 1698431365
transform 1 0 44464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_541
timestamp 1698431365
transform 1 0 52304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_542
timestamp 1698431365
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_543
timestamp 1698431365
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_544
timestamp 1698431365
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_545
timestamp 1698431365
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_546
timestamp 1698431365
transform 1 0 40544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_547
timestamp 1698431365
transform 1 0 48384 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_548
timestamp 1698431365
transform 1 0 56224 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_549
timestamp 1698431365
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_550
timestamp 1698431365
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_551
timestamp 1698431365
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_552
timestamp 1698431365
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_553
timestamp 1698431365
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_554
timestamp 1698431365
transform 1 0 44464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_555
timestamp 1698431365
transform 1 0 52304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_556
timestamp 1698431365
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_557
timestamp 1698431365
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_558
timestamp 1698431365
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_559
timestamp 1698431365
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_560
timestamp 1698431365
transform 1 0 40544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_561
timestamp 1698431365
transform 1 0 48384 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_562
timestamp 1698431365
transform 1 0 56224 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_563
timestamp 1698431365
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_564
timestamp 1698431365
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_565
timestamp 1698431365
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_566
timestamp 1698431365
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_567
timestamp 1698431365
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_568
timestamp 1698431365
transform 1 0 44464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_569
timestamp 1698431365
transform 1 0 52304 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_570
timestamp 1698431365
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_571
timestamp 1698431365
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_572
timestamp 1698431365
transform 1 0 24864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_573
timestamp 1698431365
transform 1 0 32704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_574
timestamp 1698431365
transform 1 0 40544 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_575
timestamp 1698431365
transform 1 0 48384 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_576
timestamp 1698431365
transform 1 0 56224 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_577
timestamp 1698431365
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_578
timestamp 1698431365
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_579
timestamp 1698431365
transform 1 0 20944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_580
timestamp 1698431365
transform 1 0 28784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_581
timestamp 1698431365
transform 1 0 36624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_582
timestamp 1698431365
transform 1 0 44464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_583
timestamp 1698431365
transform 1 0 52304 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_584
timestamp 1698431365
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_585
timestamp 1698431365
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_586
timestamp 1698431365
transform 1 0 24864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_587
timestamp 1698431365
transform 1 0 32704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_588
timestamp 1698431365
transform 1 0 40544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_589
timestamp 1698431365
transform 1 0 48384 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_590
timestamp 1698431365
transform 1 0 56224 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_591
timestamp 1698431365
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_592
timestamp 1698431365
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_593
timestamp 1698431365
transform 1 0 20944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_594
timestamp 1698431365
transform 1 0 28784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_595
timestamp 1698431365
transform 1 0 36624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_596
timestamp 1698431365
transform 1 0 44464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_597
timestamp 1698431365
transform 1 0 52304 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_598
timestamp 1698431365
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_599
timestamp 1698431365
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_600
timestamp 1698431365
transform 1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_601
timestamp 1698431365
transform 1 0 32704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_602
timestamp 1698431365
transform 1 0 40544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_603
timestamp 1698431365
transform 1 0 48384 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_604
timestamp 1698431365
transform 1 0 56224 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_605
timestamp 1698431365
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_606
timestamp 1698431365
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_607
timestamp 1698431365
transform 1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_608
timestamp 1698431365
transform 1 0 28784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_609
timestamp 1698431365
transform 1 0 36624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_610
timestamp 1698431365
transform 1 0 44464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_611
timestamp 1698431365
transform 1 0 52304 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_612
timestamp 1698431365
transform 1 0 5152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_613
timestamp 1698431365
transform 1 0 8960 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_614
timestamp 1698431365
transform 1 0 12768 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_615
timestamp 1698431365
transform 1 0 16576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_616
timestamp 1698431365
transform 1 0 20384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_617
timestamp 1698431365
transform 1 0 24192 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_618
timestamp 1698431365
transform 1 0 28000 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_619
timestamp 1698431365
transform 1 0 31808 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_620
timestamp 1698431365
transform 1 0 35616 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_621
timestamp 1698431365
transform 1 0 39424 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_622
timestamp 1698431365
transform 1 0 43232 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_623
timestamp 1698431365
transform 1 0 47040 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_624
timestamp 1698431365
transform 1 0 50848 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_625
timestamp 1698431365
transform 1 0 54656 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_23 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 3248 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_24
timestamp 1698431365
transform -1 0 5824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_25
timestamp 1698431365
transform -1 0 7280 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_26
timestamp 1698431365
transform -1 0 9632 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_27
timestamp 1698431365
transform -1 0 11312 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_28
timestamp 1698431365
transform -1 0 13440 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_29
timestamp 1698431365
transform -1 0 15344 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_30
timestamp 1698431365
transform -1 0 17360 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_31
timestamp 1698431365
transform -1 0 28672 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_32
timestamp 1698431365
transform -1 0 29456 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_33
timestamp 1698431365
transform -1 0 31472 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_34
timestamp 1698431365
transform -1 0 33488 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_35
timestamp 1698431365
transform -1 0 35504 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_36
timestamp 1698431365
transform -1 0 50624 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_37
timestamp 1698431365
transform -1 0 51632 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_38
timestamp 1698431365
transform -1 0 53648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_39
timestamp 1698431365
transform -1 0 55664 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_40
timestamp 1698431365
transform -1 0 57680 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_41
timestamp 1698431365
transform -1 0 48384 0 -1 4704
box -86 -86 534 870
<< labels >>
flabel metal3 s 59200 50176 60000 50288 0 FreeSans 448 0 0 0 custom_settings[0]
port 0 nsew signal input
flabel metal3 s 59200 56000 60000 56112 0 FreeSans 448 0 0 0 custom_settings[1]
port 1 nsew signal input
flabel metal3 s 59200 3584 60000 3696 0 FreeSans 448 0 0 0 io_in_1[0]
port 2 nsew signal input
flabel metal3 s 59200 9408 60000 9520 0 FreeSans 448 0 0 0 io_in_1[1]
port 3 nsew signal input
flabel metal3 s 59200 15232 60000 15344 0 FreeSans 448 0 0 0 io_in_1[2]
port 4 nsew signal input
flabel metal3 s 59200 21056 60000 21168 0 FreeSans 448 0 0 0 io_in_1[3]
port 5 nsew signal input
flabel metal3 s 59200 26880 60000 26992 0 FreeSans 448 0 0 0 io_in_1[4]
port 6 nsew signal input
flabel metal3 s 59200 32704 60000 32816 0 FreeSans 448 0 0 0 io_in_1[5]
port 7 nsew signal input
flabel metal3 s 59200 38528 60000 38640 0 FreeSans 448 0 0 0 io_in_1[6]
port 8 nsew signal input
flabel metal3 s 59200 44352 60000 44464 0 FreeSans 448 0 0 0 io_in_1[7]
port 9 nsew signal input
flabel metal2 s 37408 59200 37520 60000 0 FreeSans 448 90 0 0 io_in_2[0]
port 10 nsew signal input
flabel metal2 s 52416 59200 52528 60000 0 FreeSans 448 90 0 0 io_in_2[1]
port 11 nsew signal input
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 io_out[0]
port 12 nsew signal tristate
flabel metal2 s 22848 0 22960 800 0 FreeSans 448 90 0 0 io_out[10]
port 13 nsew signal tristate
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 io_out[11]
port 14 nsew signal tristate
flabel metal2 s 26880 0 26992 800 0 FreeSans 448 90 0 0 io_out[12]
port 15 nsew signal tristate
flabel metal2 s 28896 0 29008 800 0 FreeSans 448 90 0 0 io_out[13]
port 16 nsew signal tristate
flabel metal2 s 30912 0 31024 800 0 FreeSans 448 90 0 0 io_out[14]
port 17 nsew signal tristate
flabel metal2 s 32928 0 33040 800 0 FreeSans 448 90 0 0 io_out[15]
port 18 nsew signal tristate
flabel metal2 s 34944 0 35056 800 0 FreeSans 448 90 0 0 io_out[16]
port 19 nsew signal tristate
flabel metal2 s 36960 0 37072 800 0 FreeSans 448 90 0 0 io_out[17]
port 20 nsew signal tristate
flabel metal2 s 38976 0 39088 800 0 FreeSans 448 90 0 0 io_out[18]
port 21 nsew signal tristate
flabel metal2 s 40992 0 41104 800 0 FreeSans 448 90 0 0 io_out[19]
port 22 nsew signal tristate
flabel metal2 s 4704 0 4816 800 0 FreeSans 448 90 0 0 io_out[1]
port 23 nsew signal tristate
flabel metal2 s 43008 0 43120 800 0 FreeSans 448 90 0 0 io_out[20]
port 24 nsew signal tristate
flabel metal2 s 45024 0 45136 800 0 FreeSans 448 90 0 0 io_out[21]
port 25 nsew signal tristate
flabel metal2 s 47040 0 47152 800 0 FreeSans 448 90 0 0 io_out[22]
port 26 nsew signal tristate
flabel metal2 s 49056 0 49168 800 0 FreeSans 448 90 0 0 io_out[23]
port 27 nsew signal tristate
flabel metal2 s 51072 0 51184 800 0 FreeSans 448 90 0 0 io_out[24]
port 28 nsew signal tristate
flabel metal2 s 53088 0 53200 800 0 FreeSans 448 90 0 0 io_out[25]
port 29 nsew signal tristate
flabel metal2 s 55104 0 55216 800 0 FreeSans 448 90 0 0 io_out[26]
port 30 nsew signal tristate
flabel metal2 s 57120 0 57232 800 0 FreeSans 448 90 0 0 io_out[27]
port 31 nsew signal tristate
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 io_out[2]
port 32 nsew signal tristate
flabel metal2 s 8736 0 8848 800 0 FreeSans 448 90 0 0 io_out[3]
port 33 nsew signal tristate
flabel metal2 s 10752 0 10864 800 0 FreeSans 448 90 0 0 io_out[4]
port 34 nsew signal tristate
flabel metal2 s 12768 0 12880 800 0 FreeSans 448 90 0 0 io_out[5]
port 35 nsew signal tristate
flabel metal2 s 14784 0 14896 800 0 FreeSans 448 90 0 0 io_out[6]
port 36 nsew signal tristate
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 io_out[7]
port 37 nsew signal tristate
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 io_out[8]
port 38 nsew signal tristate
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 io_out[9]
port 39 nsew signal tristate
flabel metal2 s 22400 59200 22512 60000 0 FreeSans 448 90 0 0 rst_n
port 40 nsew signal input
flabel metal4 s 4448 3076 4768 56508 0 FreeSans 1280 90 0 0 vdd
port 41 nsew power bidirectional
flabel metal4 s 35168 3076 35488 56508 0 FreeSans 1280 90 0 0 vdd
port 41 nsew power bidirectional
flabel metal4 s 19808 3076 20128 56508 0 FreeSans 1280 90 0 0 vss
port 42 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 56508 0 FreeSans 1280 90 0 0 vss
port 42 nsew ground bidirectional
flabel metal2 s 7392 59200 7504 60000 0 FreeSans 448 90 0 0 wb_clk_i
port 43 nsew signal input
rlabel metal1 29960 55664 29960 55664 0 vdd
rlabel metal1 29960 56448 29960 56448 0 vss
rlabel metal2 36120 18088 36120 18088 0 _0000_
rlabel metal2 39480 17864 39480 17864 0 _0001_
rlabel metal2 39144 14840 39144 14840 0 _0002_
rlabel metal2 35168 10696 35168 10696 0 _0003_
rlabel metal2 34552 21224 34552 21224 0 _0004_
rlabel metal2 38024 8680 38024 8680 0 _0005_
rlabel metal3 41776 8344 41776 8344 0 _0006_
rlabel metal2 41944 5432 41944 5432 0 _0007_
rlabel metal2 38248 6608 38248 6608 0 _0008_
rlabel metal2 26152 36120 26152 36120 0 _0009_
rlabel metal3 29008 38696 29008 38696 0 _0010_
rlabel metal2 20664 36456 20664 36456 0 _0011_
rlabel metal3 22456 38136 22456 38136 0 _0012_
rlabel metal2 27832 22736 27832 22736 0 _0013_
rlabel metal2 23464 17808 23464 17808 0 _0014_
rlabel metal3 25312 13048 25312 13048 0 _0015_
rlabel metal2 19992 12320 19992 12320 0 _0016_
rlabel metal3 12264 15176 12264 15176 0 _0017_
rlabel metal2 14952 11704 14952 11704 0 _0018_
rlabel metal2 10808 11760 10808 11760 0 _0019_
rlabel metal2 12040 7784 12040 7784 0 _0020_
rlabel metal3 16912 9128 16912 9128 0 _0021_
rlabel metal2 24920 7448 24920 7448 0 _0022_
rlabel metal2 26712 10024 26712 10024 0 _0023_
rlabel metal2 22120 10584 22120 10584 0 _0024_
rlabel metal2 19992 10248 19992 10248 0 _0025_
rlabel metal2 21896 7448 21896 7448 0 _0026_
rlabel metal2 19432 8624 19432 8624 0 _0027_
rlabel metal2 16296 6328 16296 6328 0 _0028_
rlabel metal2 14616 4816 14616 4816 0 _0029_
rlabel metal2 19992 4480 19992 4480 0 _0030_
rlabel metal2 22120 4480 22120 4480 0 _0031_
rlabel metal2 19320 23520 19320 23520 0 _0032_
rlabel metal2 12376 24360 12376 24360 0 _0033_
rlabel metal2 2520 22792 2520 22792 0 _0034_
rlabel metal2 6608 18536 6608 18536 0 _0035_
rlabel metal2 5544 15624 5544 15624 0 _0036_
rlabel metal2 10136 15456 10136 15456 0 _0037_
rlabel metal3 7784 11480 7784 11480 0 _0038_
rlabel metal2 10920 4648 10920 4648 0 _0039_
rlabel metal2 40152 11704 40152 11704 0 _0040_
rlabel metal2 41720 14336 41720 14336 0 _0041_
rlabel metal3 43400 9128 43400 9128 0 _0042_
rlabel metal2 43512 13216 43512 13216 0 _0043_
rlabel metal2 50792 19544 50792 19544 0 _0044_
rlabel metal2 51912 18760 51912 18760 0 _0045_
rlabel metal2 56000 16184 56000 16184 0 _0046_
rlabel metal2 56056 19544 56056 19544 0 _0047_
rlabel metal2 39368 25816 39368 25816 0 _0048_
rlabel metal2 41832 24360 41832 24360 0 _0049_
rlabel metal2 42168 22680 42168 22680 0 _0050_
rlabel metal2 38024 23072 38024 23072 0 _0051_
rlabel metal2 43960 34552 43960 34552 0 _0052_
rlabel metal2 39928 29344 39928 29344 0 _0053_
rlabel metal2 38248 30520 38248 30520 0 _0054_
rlabel metal3 42056 32424 42056 32424 0 _0055_
rlabel metal2 49448 36792 49448 36792 0 _0056_
rlabel metal2 52024 35224 52024 35224 0 _0057_
rlabel metal2 55608 36120 55608 36120 0 _0058_
rlabel metal3 55944 37128 55944 37128 0 _0059_
rlabel metal2 30016 4424 30016 4424 0 _0060_
rlabel metal2 30184 10192 30184 10192 0 _0061_
rlabel metal2 29960 7224 29960 7224 0 _0062_
rlabel metal2 35672 5432 35672 5432 0 _0063_
rlabel metal2 35112 8624 35112 8624 0 _0064_
rlabel metal2 2520 20412 2520 20412 0 _0065_
rlabel metal2 2520 17976 2520 17976 0 _0066_
rlabel metal2 2968 14000 2968 14000 0 _0067_
rlabel metal2 2520 12096 2520 12096 0 _0068_
rlabel metal2 2968 9464 2968 9464 0 _0069_
rlabel metal2 8680 9464 8680 9464 0 _0070_
rlabel metal2 8008 6328 8008 6328 0 _0071_
rlabel metal2 10696 6384 10696 6384 0 _0072_
rlabel metal2 27496 30240 27496 30240 0 _0073_
rlabel metal2 26600 28784 26600 28784 0 _0074_
rlabel metal3 21952 39816 21952 39816 0 _0075_
rlabel metal2 21224 42224 21224 42224 0 _0076_
rlabel metal2 25144 43064 25144 43064 0 _0077_
rlabel metal3 25480 39480 25480 39480 0 _0078_
rlabel metal2 33544 41496 33544 41496 0 _0079_
rlabel metal2 28728 42280 28728 42280 0 _0080_
rlabel metal2 33656 44632 33656 44632 0 _0081_
rlabel metal2 29960 43624 29960 43624 0 _0082_
rlabel metal2 36904 5432 36904 5432 0 _0083_
rlabel metal2 26040 5264 26040 5264 0 _0084_
rlabel metal2 34552 4760 34552 4760 0 _0085_
rlabel metal2 7672 21448 7672 21448 0 _0086_
rlabel metal3 23072 32760 23072 32760 0 _0087_
rlabel metal2 19768 31136 19768 31136 0 _0088_
rlabel metal3 28728 31864 28728 31864 0 _0089_
rlabel metal2 19656 32872 19656 32872 0 _0090_
rlabel metal2 36008 29736 36008 29736 0 _0091_
rlabel metal2 30352 29512 30352 29512 0 _0092_
rlabel metal2 45864 38668 45864 38668 0 _0093_
rlabel metal2 46312 43176 46312 43176 0 _0094_
rlabel metal2 45864 40768 45864 40768 0 _0095_
rlabel metal2 49448 41552 49448 41552 0 _0096_
rlabel metal3 49952 38696 49952 38696 0 _0097_
rlabel metal2 53032 41160 53032 41160 0 _0098_
rlabel metal2 56000 39704 56000 39704 0 _0099_
rlabel metal2 56056 43932 56056 43932 0 _0100_
rlabel metal2 19096 40320 19096 40320 0 _0101_
rlabel metal2 9240 42672 9240 42672 0 _0102_
rlabel metal2 7336 43932 7336 43932 0 _0103_
rlabel metal3 8288 48104 8288 48104 0 _0104_
rlabel metal3 7000 46536 7000 46536 0 _0105_
rlabel metal2 11368 46312 11368 46312 0 _0106_
rlabel metal2 15960 47824 15960 47824 0 _0107_
rlabel metal2 31864 47880 31864 47880 0 _0108_
rlabel metal2 35000 51744 35000 51744 0 _0109_
rlabel metal2 34328 54432 34328 54432 0 _0110_
rlabel metal2 38808 52472 38808 52472 0 _0111_
rlabel metal3 39424 55160 39424 55160 0 _0112_
rlabel metal2 43512 54040 43512 54040 0 _0113_
rlabel metal2 45416 51744 45416 51744 0 _0114_
rlabel metal3 47096 54712 47096 54712 0 _0115_
rlabel metal2 51576 48944 51576 48944 0 _0116_
rlabel metal2 47992 47544 47992 47544 0 _0117_
rlabel metal2 51800 50792 51800 50792 0 _0118_
rlabel metal2 50008 54432 50008 54432 0 _0119_
rlabel metal2 54488 54936 54488 54936 0 _0120_
rlabel metal2 57400 52472 57400 52472 0 _0121_
rlabel metal2 56000 49112 56000 49112 0 _0122_
rlabel metal2 57400 47656 57400 47656 0 _0123_
rlabel metal2 12712 42224 12712 42224 0 _0124_
rlabel metal3 15288 28728 15288 28728 0 _0125_
rlabel metal3 12208 28392 12208 28392 0 _0126_
rlabel metal2 11256 31416 11256 31416 0 _0127_
rlabel metal3 8624 25592 8624 25592 0 _0128_
rlabel metal2 5768 25032 5768 25032 0 _0129_
rlabel metal2 2520 25032 2520 25032 0 _0130_
rlabel metal2 3976 27440 3976 27440 0 _0131_
rlabel metal2 2520 30520 2520 30520 0 _0132_
rlabel metal3 3808 32424 3808 32424 0 _0133_
rlabel metal2 2520 34048 2520 34048 0 _0134_
rlabel metal2 4536 36120 4536 36120 0 _0135_
rlabel metal3 4200 38136 4200 38136 0 _0136_
rlabel metal3 6328 38864 6328 38864 0 _0137_
rlabel metal2 7560 39256 7560 39256 0 _0138_
rlabel metal3 10304 38696 10304 38696 0 _0139_
rlabel metal3 10136 35000 10136 35000 0 _0140_
rlabel metal2 7784 32536 7784 32536 0 _0141_
rlabel metal2 28000 16968 28000 16968 0 _0142_
rlabel metal2 30352 20104 30352 20104 0 _0143_
rlabel metal2 30744 17024 30744 17024 0 _0144_
rlabel metal2 30408 15680 30408 15680 0 _0145_
rlabel metal2 27608 12488 27608 12488 0 _0146_
rlabel metal2 31808 11480 31808 11480 0 _0147_
rlabel metal2 13496 48496 13496 48496 0 _0148_
rlabel metal2 14728 39256 14728 39256 0 _0149_
rlabel metal2 19656 41496 19656 41496 0 _0150_
rlabel metal2 12152 40712 12152 40712 0 _0151_
rlabel metal3 17528 38584 17528 38584 0 _0152_
rlabel metal2 45416 19264 45416 19264 0 _0153_
rlabel metal2 46536 15736 46536 15736 0 _0154_
rlabel metal2 49672 16576 49672 16576 0 _0155_
rlabel metal3 55496 14616 55496 14616 0 _0156_
rlabel metal2 56056 13440 56056 13440 0 _0157_
rlabel metal3 56560 11480 56560 11480 0 _0158_
rlabel metal2 57400 8372 57400 8372 0 _0159_
rlabel metal2 57232 6664 57232 6664 0 _0160_
rlabel metal2 54152 5152 54152 5152 0 _0161_
rlabel metal2 52696 4648 52696 4648 0 _0162_
rlabel metal2 47768 4760 47768 4760 0 _0163_
rlabel metal3 43960 3640 43960 3640 0 _0164_
rlabel metal3 32256 23016 32256 23016 0 _0165_
rlabel metal2 45752 26208 45752 26208 0 _0166_
rlabel metal3 43680 27720 43680 27720 0 _0167_
rlabel metal2 45528 31360 45528 31360 0 _0168_
rlabel metal2 47432 33656 47432 33656 0 _0169_
rlabel metal3 55440 33432 55440 33432 0 _0170_
rlabel metal3 55440 31640 55440 31640 0 _0171_
rlabel metal2 56000 28728 56000 28728 0 _0172_
rlabel metal2 56056 25312 56056 25312 0 _0173_
rlabel metal2 56000 24024 56000 24024 0 _0174_
rlabel metal2 55832 21952 55832 21952 0 _0175_
rlabel metal2 53144 22288 53144 22288 0 _0176_
rlabel metal2 46088 22344 46088 22344 0 _0177_
rlabel metal3 36120 23800 36120 23800 0 _0178_
rlabel metal2 23464 51072 23464 51072 0 _0179_
rlabel metal2 33320 51296 33320 51296 0 _0180_
rlabel metal2 33432 54040 33432 54040 0 _0181_
rlabel metal2 23800 54936 23800 54936 0 _0182_
rlabel metal2 26488 52864 26488 52864 0 _0183_
rlabel metal2 29848 54432 29848 54432 0 _0184_
rlabel metal2 22792 54936 22792 54936 0 _0185_
rlabel metal2 18200 54040 18200 54040 0 _0186_
rlabel metal3 18704 51128 18704 51128 0 _0187_
rlabel metal2 20328 51744 20328 51744 0 _0188_
rlabel metal2 18648 48720 18648 48720 0 _0189_
rlabel metal2 21896 47824 21896 47824 0 _0190_
rlabel metal2 24136 31920 24136 31920 0 _0191_
rlabel metal2 27384 25872 27384 25872 0 _0192_
rlabel metal3 22960 26376 22960 26376 0 _0193_
rlabel metal2 12488 33712 12488 33712 0 _0194_
rlabel metal3 13552 36232 13552 36232 0 _0195_
rlabel metal2 16408 34216 16408 34216 0 _0196_
rlabel metal2 14728 32872 14728 32872 0 _0197_
rlabel metal2 13832 30240 13832 30240 0 _0198_
rlabel metal2 16296 27496 16296 27496 0 _0199_
rlabel metal2 15960 24304 15960 24304 0 _0200_
rlabel metal3 31752 37464 31752 37464 0 _0201_
rlabel metal2 32312 33264 32312 33264 0 _0202_
rlabel metal2 30520 35280 30520 35280 0 _0203_
rlabel metal3 37072 35000 37072 35000 0 _0204_
rlabel metal2 37016 37520 37016 37520 0 _0205_
rlabel metal2 36456 40768 36456 40768 0 _0206_
rlabel metal2 35448 43848 35448 43848 0 _0207_
rlabel metal3 34832 41944 34832 41944 0 _0208_
rlabel metal2 39928 43960 39928 43960 0 _0209_
rlabel metal2 42560 38696 42560 38696 0 _0210_
rlabel metal2 42280 41216 42280 41216 0 _0211_
rlabel metal2 41944 44744 41944 44744 0 _0212_
rlabel metal2 44968 45416 44968 45416 0 _0213_
rlabel metal2 16520 21840 16520 21840 0 _0214_
rlabel metal3 11816 21784 11816 21784 0 _0215_
rlabel metal3 12152 19880 12152 19880 0 _0216_
rlabel metal3 12768 18312 12768 18312 0 _0217_
rlabel metal2 17080 19376 17080 19376 0 _0218_
rlabel metal2 19992 21336 19992 21336 0 _0219_
rlabel metal2 21560 17360 21560 17360 0 _0220_
rlabel metal2 18200 15624 18200 15624 0 _0221_
rlabel metal2 33880 26628 33880 26628 0 _0222_
rlabel metal3 30744 27720 30744 27720 0 _0223_
rlabel metal2 56056 50512 56056 50512 0 _0224_
rlabel metal2 57064 48328 57064 48328 0 _0225_
rlabel metal2 16520 43120 16520 43120 0 _0226_
rlabel metal2 15904 45080 15904 45080 0 _0227_
rlabel metal2 16072 44352 16072 44352 0 _0228_
rlabel metal2 14728 43848 14728 43848 0 _0229_
rlabel metal2 15848 43064 15848 43064 0 _0230_
rlabel metal2 9688 23912 9688 23912 0 _0231_
rlabel metal3 8344 28504 8344 28504 0 _0232_
rlabel metal2 9016 30576 9016 30576 0 _0233_
rlabel metal2 12208 28056 12208 28056 0 _0234_
rlabel metal2 8568 30576 8568 30576 0 _0235_
rlabel metal2 5992 31360 5992 31360 0 _0236_
rlabel metal2 11144 27440 11144 27440 0 _0237_
rlabel metal3 11480 28616 11480 28616 0 _0238_
rlabel metal2 11480 29792 11480 29792 0 _0239_
rlabel metal2 11368 29008 11368 29008 0 _0240_
rlabel metal2 11480 28112 11480 28112 0 _0241_
rlabel metal2 11144 30184 11144 30184 0 _0242_
rlabel metal2 10808 31024 10808 31024 0 _0243_
rlabel metal2 7672 28560 7672 28560 0 _0244_
rlabel metal3 6496 27048 6496 27048 0 _0245_
rlabel metal2 8176 26936 8176 26936 0 _0246_
rlabel metal2 8680 26936 8680 26936 0 _0247_
rlabel metal3 7616 26936 7616 26936 0 _0248_
rlabel metal2 5992 26152 5992 26152 0 _0249_
rlabel metal2 5768 30184 5768 30184 0 _0250_
rlabel metal2 6496 25704 6496 25704 0 _0251_
rlabel metal2 4648 26488 4648 26488 0 _0252_
rlabel metal2 3640 25872 3640 25872 0 _0253_
rlabel metal2 4200 27720 4200 27720 0 _0254_
rlabel metal2 3864 27440 3864 27440 0 _0255_
rlabel metal3 5152 32536 5152 32536 0 _0256_
rlabel metal2 4704 31080 4704 31080 0 _0257_
rlabel metal2 5544 30576 5544 30576 0 _0258_
rlabel metal3 5376 31080 5376 31080 0 _0259_
rlabel metal2 5600 32760 5600 32760 0 _0260_
rlabel metal2 4760 31556 4760 31556 0 _0261_
rlabel metal2 4872 32256 4872 32256 0 _0262_
rlabel metal2 5880 34944 5880 34944 0 _0263_
rlabel metal3 5152 34776 5152 34776 0 _0264_
rlabel metal2 4760 36008 4760 36008 0 _0265_
rlabel metal2 4312 36456 4312 36456 0 _0266_
rlabel metal3 6272 38024 6272 38024 0 _0267_
rlabel metal2 6104 38080 6104 38080 0 _0268_
rlabel metal2 5768 37688 5768 37688 0 _0269_
rlabel metal3 7000 38808 7000 38808 0 _0270_
rlabel metal2 6216 39032 6216 39032 0 _0271_
rlabel metal2 7560 38360 7560 38360 0 _0272_
rlabel metal2 6216 38640 6216 38640 0 _0273_
rlabel metal2 7336 39144 7336 39144 0 _0274_
rlabel metal2 7672 38528 7672 38528 0 _0275_
rlabel metal2 8792 38528 8792 38528 0 _0276_
rlabel metal2 9128 39088 9128 39088 0 _0277_
rlabel metal2 9240 35672 9240 35672 0 _0278_
rlabel metal2 9464 35840 9464 35840 0 _0279_
rlabel metal2 8624 28616 8624 28616 0 _0280_
rlabel metal3 6944 35784 6944 35784 0 _0281_
rlabel metal2 7952 35784 7952 35784 0 _0282_
rlabel metal2 7952 35448 7952 35448 0 _0283_
rlabel metal2 8344 28280 8344 28280 0 _0284_
rlabel metal2 9128 28448 9128 28448 0 _0285_
rlabel metal2 7896 29736 7896 29736 0 _0286_
rlabel metal2 7784 31360 7784 31360 0 _0287_
rlabel metal3 8288 31640 8288 31640 0 _0288_
rlabel metal2 34328 13888 34328 13888 0 _0289_
rlabel metal3 34048 18424 34048 18424 0 _0290_
rlabel metal2 34328 17360 34328 17360 0 _0291_
rlabel metal2 35224 17864 35224 17864 0 _0292_
rlabel metal2 34216 17808 34216 17808 0 _0293_
rlabel metal2 34496 15400 34496 15400 0 _0294_
rlabel metal2 33600 15064 33600 15064 0 _0295_
rlabel metal2 34328 15148 34328 15148 0 _0296_
rlabel metal2 36008 15204 36008 15204 0 _0297_
rlabel metal3 32760 12936 32760 12936 0 _0298_
rlabel metal2 36288 12824 36288 12824 0 _0299_
rlabel metal3 36120 15288 36120 15288 0 _0300_
rlabel metal3 32144 15400 32144 15400 0 _0301_
rlabel metal2 27384 16464 27384 16464 0 _0302_
rlabel metal3 30240 16744 30240 16744 0 _0303_
rlabel metal3 30688 19992 30688 19992 0 _0304_
rlabel metal2 30856 19936 30856 19936 0 _0305_
rlabel metal2 31080 17528 31080 17528 0 _0306_
rlabel metal3 43568 18088 43568 18088 0 _0307_
rlabel metal2 31304 17304 31304 17304 0 _0308_
rlabel metal2 31024 14728 31024 14728 0 _0309_
rlabel metal2 31304 16128 31304 16128 0 _0310_
rlabel metal3 29568 13160 29568 13160 0 _0311_
rlabel metal2 28056 12992 28056 12992 0 _0312_
rlabel metal2 27384 12936 27384 12936 0 _0313_
rlabel metal2 18760 38080 18760 38080 0 _0314_
rlabel metal2 14840 39144 14840 39144 0 _0315_
rlabel metal2 18760 40600 18760 40600 0 _0316_
rlabel metal2 12824 40656 12824 40656 0 _0317_
rlabel metal3 18480 38696 18480 38696 0 _0318_
rlabel metal3 46088 19208 46088 19208 0 _0319_
rlabel metal2 45024 18648 45024 18648 0 _0320_
rlabel metal2 43400 25424 43400 25424 0 _0321_
rlabel metal3 46144 6440 46144 6440 0 _0322_
rlabel metal2 46984 6216 46984 6216 0 _0323_
rlabel metal3 46424 8008 46424 8008 0 _0324_
rlabel metal2 46648 7560 46648 7560 0 _0325_
rlabel metal2 47208 7560 47208 7560 0 _0326_
rlabel metal2 46872 7784 46872 7784 0 _0327_
rlabel metal2 46984 7728 46984 7728 0 _0328_
rlabel metal2 48776 8736 48776 8736 0 _0329_
rlabel metal2 45080 16856 45080 16856 0 _0330_
rlabel metal2 46088 11648 46088 11648 0 _0331_
rlabel metal2 52808 9408 52808 9408 0 _0332_
rlabel metal2 50008 8512 50008 8512 0 _0333_
rlabel metal2 48888 10248 48888 10248 0 _0334_
rlabel metal3 48104 10360 48104 10360 0 _0335_
rlabel metal3 49672 13496 49672 13496 0 _0336_
rlabel metal3 50064 13720 50064 13720 0 _0337_
rlabel metal2 50232 12208 50232 12208 0 _0338_
rlabel metal2 47936 15848 47936 15848 0 _0339_
rlabel metal2 49336 12208 49336 12208 0 _0340_
rlabel metal2 49112 12656 49112 12656 0 _0341_
rlabel metal2 47656 10864 47656 10864 0 _0342_
rlabel metal2 48104 10248 48104 10248 0 _0343_
rlabel metal2 52808 12432 52808 12432 0 _0344_
rlabel metal2 52024 14224 52024 14224 0 _0345_
rlabel metal2 51016 11872 51016 11872 0 _0346_
rlabel metal2 53928 15876 53928 15876 0 _0347_
rlabel metal2 52472 11144 52472 11144 0 _0348_
rlabel metal3 50316 11368 50316 11368 0 _0349_
rlabel metal2 46760 12992 46760 12992 0 _0350_
rlabel metal2 48104 12040 48104 12040 0 _0351_
rlabel metal2 49336 6720 49336 6720 0 _0352_
rlabel metal2 49728 9240 49728 9240 0 _0353_
rlabel metal2 53144 8568 53144 8568 0 _0354_
rlabel metal2 50064 9128 50064 9128 0 _0355_
rlabel metal2 49896 9352 49896 9352 0 _0356_
rlabel metal2 49448 10584 49448 10584 0 _0357_
rlabel metal3 48608 9016 48608 9016 0 _0358_
rlabel metal2 50008 12544 50008 12544 0 _0359_
rlabel metal2 45528 13048 45528 13048 0 _0360_
rlabel metal2 49784 12600 49784 12600 0 _0361_
rlabel metal2 49840 10696 49840 10696 0 _0362_
rlabel metal2 50344 10920 50344 10920 0 _0363_
rlabel metal2 49896 10136 49896 10136 0 _0364_
rlabel metal2 49448 9240 49448 9240 0 _0365_
rlabel metal2 49112 9520 49112 9520 0 _0366_
rlabel metal2 47208 9128 47208 9128 0 _0367_
rlabel metal2 42616 9912 42616 9912 0 _0368_
rlabel metal3 43736 18984 43736 18984 0 _0369_
rlabel metal3 49280 15288 49280 15288 0 _0370_
rlabel metal2 45304 17304 45304 17304 0 _0371_
rlabel via2 46872 15960 46872 15960 0 _0372_
rlabel metal3 41776 20552 41776 20552 0 _0373_
rlabel metal2 43960 16184 43960 16184 0 _0374_
rlabel metal2 46760 15568 46760 15568 0 _0375_
rlabel metal3 48608 15176 48608 15176 0 _0376_
rlabel metal2 49336 16184 49336 16184 0 _0377_
rlabel metal2 52752 13720 52752 13720 0 _0378_
rlabel metal3 50512 16632 50512 16632 0 _0379_
rlabel metal2 53144 15512 53144 15512 0 _0380_
rlabel metal2 53704 15736 53704 15736 0 _0381_
rlabel metal3 54208 15960 54208 15960 0 _0382_
rlabel metal2 54320 14392 54320 14392 0 _0383_
rlabel metal2 55720 14056 55720 14056 0 _0384_
rlabel metal2 39144 13104 39144 13104 0 _0385_
rlabel metal2 38248 12264 38248 12264 0 _0386_
rlabel metal2 53088 12152 53088 12152 0 _0387_
rlabel metal3 53704 11928 53704 11928 0 _0388_
rlabel metal2 53816 10304 53816 10304 0 _0389_
rlabel metal3 54992 12152 54992 12152 0 _0390_
rlabel metal2 26264 30632 26264 30632 0 _0391_
rlabel metal3 54488 8344 54488 8344 0 _0392_
rlabel metal2 53760 9016 53760 9016 0 _0393_
rlabel metal3 55608 9016 55608 9016 0 _0394_
rlabel metal2 55048 7560 55048 7560 0 _0395_
rlabel metal3 56000 7448 56000 7448 0 _0396_
rlabel metal3 53816 6888 53816 6888 0 _0397_
rlabel metal3 49896 6888 49896 6888 0 _0398_
rlabel metal2 53760 4424 53760 4424 0 _0399_
rlabel metal2 50232 6216 50232 6216 0 _0400_
rlabel metal3 48888 5880 48888 5880 0 _0401_
rlabel metal2 50904 5096 50904 5096 0 _0402_
rlabel metal2 45752 5376 45752 5376 0 _0403_
rlabel metal2 47432 4648 47432 4648 0 _0404_
rlabel metal2 43736 6776 43736 6776 0 _0405_
rlabel metal2 33320 23520 33320 23520 0 _0406_
rlabel metal2 32088 22624 32088 22624 0 _0407_
rlabel metal3 44072 27832 44072 27832 0 _0408_
rlabel metal2 44744 25088 44744 25088 0 _0409_
rlabel metal3 49336 24752 49336 24752 0 _0410_
rlabel metal3 52248 25368 52248 25368 0 _0411_
rlabel metal2 51128 25200 51128 25200 0 _0412_
rlabel metal2 50456 25592 50456 25592 0 _0413_
rlabel metal2 54040 28224 54040 28224 0 _0414_
rlabel metal2 54824 29120 54824 29120 0 _0415_
rlabel metal2 52024 28616 52024 28616 0 _0416_
rlabel metal2 53144 32592 53144 32592 0 _0417_
rlabel metal2 52696 32704 52696 32704 0 _0418_
rlabel metal3 52136 32536 52136 32536 0 _0419_
rlabel metal2 51016 30408 51016 30408 0 _0420_
rlabel metal2 51800 29792 51800 29792 0 _0421_
rlabel metal3 48440 32536 48440 32536 0 _0422_
rlabel metal2 48216 31416 48216 31416 0 _0423_
rlabel metal2 49616 29400 49616 29400 0 _0424_
rlabel metal2 46424 29008 46424 29008 0 _0425_
rlabel metal2 46088 29008 46088 29008 0 _0426_
rlabel metal3 47320 28392 47320 28392 0 _0427_
rlabel metal2 47880 30352 47880 30352 0 _0428_
rlabel metal3 45752 28616 45752 28616 0 _0429_
rlabel metal2 48664 27664 48664 27664 0 _0430_
rlabel metal2 48216 29624 48216 29624 0 _0431_
rlabel metal2 48552 29064 48552 29064 0 _0432_
rlabel metal2 50904 32928 50904 32928 0 _0433_
rlabel metal3 50176 32536 50176 32536 0 _0434_
rlabel metal2 50344 32928 50344 32928 0 _0435_
rlabel metal2 50960 29512 50960 29512 0 _0436_
rlabel metal2 50344 29120 50344 29120 0 _0437_
rlabel metal3 50624 29624 50624 29624 0 _0438_
rlabel metal3 54208 30184 54208 30184 0 _0439_
rlabel metal2 53592 30464 53592 30464 0 _0440_
rlabel metal2 52248 29848 52248 29848 0 _0441_
rlabel metal2 51016 28728 51016 28728 0 _0442_
rlabel metal2 52528 26376 52528 26376 0 _0443_
rlabel metal2 53312 25704 53312 25704 0 _0444_
rlabel metal2 52808 29064 52808 29064 0 _0445_
rlabel metal3 52136 28616 52136 28616 0 _0446_
rlabel metal3 50904 26376 50904 26376 0 _0447_
rlabel metal2 49000 22904 49000 22904 0 _0448_
rlabel metal2 49448 22736 49448 22736 0 _0449_
rlabel metal2 48888 24192 48888 24192 0 _0450_
rlabel metal2 50008 23856 50008 23856 0 _0451_
rlabel metal2 49112 22008 49112 22008 0 _0452_
rlabel metal2 49896 24360 49896 24360 0 _0453_
rlabel metal2 49224 25200 49224 25200 0 _0454_
rlabel metal2 49336 26292 49336 26292 0 _0455_
rlabel metal2 50120 25536 50120 25536 0 _0456_
rlabel metal2 49504 24136 49504 24136 0 _0457_
rlabel metal2 51240 27496 51240 27496 0 _0458_
rlabel metal2 51632 27048 51632 27048 0 _0459_
rlabel metal3 50736 26936 50736 26936 0 _0460_
rlabel metal2 50232 28112 50232 28112 0 _0461_
rlabel metal3 50904 25480 50904 25480 0 _0462_
rlabel metal3 44184 24920 44184 24920 0 _0463_
rlabel metal3 45640 23912 45640 23912 0 _0464_
rlabel metal2 45080 24192 45080 24192 0 _0465_
rlabel metal2 45304 25900 45304 25900 0 _0466_
rlabel metal2 45640 23800 45640 23800 0 _0467_
rlabel metal2 45584 28840 45584 28840 0 _0468_
rlabel metal2 45080 27720 45080 27720 0 _0469_
rlabel metal3 48608 31528 48608 31528 0 _0470_
rlabel metal2 47320 32200 47320 32200 0 _0471_
rlabel metal2 45864 30408 45864 30408 0 _0472_
rlabel metal2 46760 24024 46760 24024 0 _0473_
rlabel metal2 48216 33264 48216 33264 0 _0474_
rlabel metal2 53200 33320 53200 33320 0 _0475_
rlabel metal2 54432 33208 54432 33208 0 _0476_
rlabel metal3 53648 32312 53648 32312 0 _0477_
rlabel metal3 54096 31864 54096 31864 0 _0478_
rlabel metal2 54264 31696 54264 31696 0 _0479_
rlabel metal2 55440 29288 55440 29288 0 _0480_
rlabel metal2 54824 24416 54824 24416 0 _0481_
rlabel metal2 54936 25592 54936 25592 0 _0482_
rlabel metal3 55496 24472 55496 24472 0 _0483_
rlabel metal2 56392 24696 56392 24696 0 _0484_
rlabel metal2 55552 21560 55552 21560 0 _0485_
rlabel metal2 52920 22568 52920 22568 0 _0486_
rlabel metal2 52640 23016 52640 23016 0 _0487_
rlabel metal2 48328 22848 48328 22848 0 _0488_
rlabel metal2 36456 23128 36456 23128 0 _0489_
rlabel metal3 36792 23912 36792 23912 0 _0490_
rlabel metal2 29960 50512 29960 50512 0 _0491_
rlabel metal2 22792 50960 22792 50960 0 _0492_
rlabel metal2 23240 45528 23240 45528 0 _0493_
rlabel metal2 26376 45136 26376 45136 0 _0494_
rlabel metal2 23464 46480 23464 46480 0 _0495_
rlabel metal2 26488 46760 26488 46760 0 _0496_
rlabel metal2 30408 47768 30408 47768 0 _0497_
rlabel metal3 28840 48888 28840 48888 0 _0498_
rlabel metal2 26824 50176 26824 50176 0 _0499_
rlabel metal3 25760 49672 25760 49672 0 _0500_
rlabel metal2 26824 49224 26824 49224 0 _0501_
rlabel metal2 24584 49112 24584 49112 0 _0502_
rlabel metal2 25816 49504 25816 49504 0 _0503_
rlabel metal2 27272 48496 27272 48496 0 _0504_
rlabel metal2 26264 53200 26264 53200 0 _0505_
rlabel metal2 27496 47936 27496 47936 0 _0506_
rlabel metal2 26768 47992 26768 47992 0 _0507_
rlabel metal2 30968 47376 30968 47376 0 _0508_
rlabel metal2 29848 46760 29848 46760 0 _0509_
rlabel metal3 29176 49000 29176 49000 0 _0510_
rlabel metal3 30632 46648 30632 46648 0 _0511_
rlabel metal2 29400 46312 29400 46312 0 _0512_
rlabel metal2 29624 45416 29624 45416 0 _0513_
rlabel metal2 25816 47656 25816 47656 0 _0514_
rlabel metal2 26488 45752 26488 45752 0 _0515_
rlabel metal2 27160 45360 27160 45360 0 _0516_
rlabel metal2 26152 45360 26152 45360 0 _0517_
rlabel metal2 21784 45920 21784 45920 0 _0518_
rlabel metal2 24584 45024 24584 45024 0 _0519_
rlabel metal2 21784 47320 21784 47320 0 _0520_
rlabel metal2 23464 44632 23464 44632 0 _0521_
rlabel metal2 22904 44408 22904 44408 0 _0522_
rlabel metal2 25312 32760 25312 32760 0 _0523_
rlabel metal2 26208 44520 26208 44520 0 _0524_
rlabel metal2 20328 51240 20328 51240 0 _0525_
rlabel metal2 24024 51296 24024 51296 0 _0526_
rlabel metal2 26544 51576 26544 51576 0 _0527_
rlabel metal2 31584 52360 31584 52360 0 _0528_
rlabel metal2 31920 51576 31920 51576 0 _0529_
rlabel metal2 31640 53704 31640 53704 0 _0530_
rlabel metal2 30408 50204 30408 50204 0 _0531_
rlabel metal2 26152 54488 26152 54488 0 _0532_
rlabel metal3 21504 48776 21504 48776 0 _0533_
rlabel metal3 24584 53704 24584 53704 0 _0534_
rlabel metal2 27160 54320 27160 54320 0 _0535_
rlabel metal2 27160 53704 27160 53704 0 _0536_
rlabel metal2 21728 53592 21728 53592 0 _0537_
rlabel metal2 28168 53480 28168 53480 0 _0538_
rlabel metal2 22512 54376 22512 54376 0 _0539_
rlabel metal3 20216 50680 20216 50680 0 _0540_
rlabel metal2 20720 53928 20720 53928 0 _0541_
rlabel metal2 21280 50456 21280 50456 0 _0542_
rlabel metal2 19432 51800 19432 51800 0 _0543_
rlabel metal2 19992 51464 19992 51464 0 _0544_
rlabel metal2 20160 50008 20160 50008 0 _0545_
rlabel metal2 20552 48216 20552 48216 0 _0546_
rlabel metal2 22176 47432 22176 47432 0 _0547_
rlabel metal2 25704 31920 25704 31920 0 _0548_
rlabel metal2 26600 27160 26600 27160 0 _0549_
rlabel metal3 25872 27720 25872 27720 0 _0550_
rlabel metal2 25760 26040 25760 26040 0 _0551_
rlabel metal3 24920 27608 24920 27608 0 _0552_
rlabel metal3 13160 35672 13160 35672 0 _0553_
rlabel metal2 14168 36400 14168 36400 0 _0554_
rlabel metal2 13664 35896 13664 35896 0 _0555_
rlabel metal2 16296 34384 16296 34384 0 _0556_
rlabel metal2 16408 33824 16408 33824 0 _0557_
rlabel metal3 16912 32760 16912 32760 0 _0558_
rlabel metal3 17360 23128 17360 23128 0 _0559_
rlabel metal3 16688 31864 16688 31864 0 _0560_
rlabel metal2 16072 29680 16072 29680 0 _0561_
rlabel metal2 16464 29512 16464 29512 0 _0562_
rlabel metal2 15904 28392 15904 28392 0 _0563_
rlabel metal2 16632 27832 16632 27832 0 _0564_
rlabel metal2 15848 25088 15848 25088 0 _0565_
rlabel metal2 37688 39368 37688 39368 0 _0566_
rlabel metal3 36624 38024 36624 38024 0 _0567_
rlabel metal2 35896 37128 35896 37128 0 _0568_
rlabel metal2 33656 39480 33656 39480 0 _0569_
rlabel metal2 32312 37912 32312 37912 0 _0570_
rlabel metal2 33096 35280 33096 35280 0 _0571_
rlabel metal2 33656 35056 33656 35056 0 _0572_
rlabel metal2 32536 36008 32536 36008 0 _0573_
rlabel metal2 35840 35784 35840 35784 0 _0574_
rlabel metal2 36568 37408 36568 37408 0 _0575_
rlabel metal3 40208 40152 40208 40152 0 _0576_
rlabel metal2 38808 41272 38808 41272 0 _0577_
rlabel metal3 40432 40264 40432 40264 0 _0578_
rlabel metal2 39592 41440 39592 41440 0 _0579_
rlabel metal2 37240 41384 37240 41384 0 _0580_
rlabel metal3 37296 43624 37296 43624 0 _0581_
rlabel metal2 35448 42056 35448 42056 0 _0582_
rlabel metal2 39256 43344 39256 43344 0 _0583_
rlabel metal2 43344 44296 43344 44296 0 _0584_
rlabel metal2 43848 44184 43848 44184 0 _0585_
rlabel metal2 42112 38920 42112 38920 0 _0586_
rlabel metal2 42392 40712 42392 40712 0 _0587_
rlabel metal2 42280 44408 42280 44408 0 _0588_
rlabel metal2 43512 45080 43512 45080 0 _0589_
rlabel metal2 16632 21616 16632 21616 0 _0590_
rlabel metal2 16856 21896 16856 21896 0 _0591_
rlabel metal3 13832 20776 13832 20776 0 _0592_
rlabel metal2 16072 18312 16072 18312 0 _0593_
rlabel metal2 13160 21336 13160 21336 0 _0594_
rlabel metal2 13552 19992 13552 19992 0 _0595_
rlabel metal2 13832 20440 13832 20440 0 _0596_
rlabel metal2 16744 18480 16744 18480 0 _0597_
rlabel metal2 14392 18760 14392 18760 0 _0598_
rlabel metal2 18424 18480 18424 18480 0 _0599_
rlabel metal2 18648 18088 18648 18088 0 _0600_
rlabel metal2 16632 19096 16632 19096 0 _0601_
rlabel metal2 19544 20888 19544 20888 0 _0602_
rlabel metal2 19320 18088 19320 18088 0 _0603_
rlabel metal2 19936 17528 19936 17528 0 _0604_
rlabel metal2 17864 16744 17864 16744 0 _0605_
rlabel metal2 31640 27832 31640 27832 0 _0606_
rlabel metal2 31752 26040 31752 26040 0 _0607_
rlabel metal2 23016 25536 23016 25536 0 _0608_
rlabel metal2 23856 23800 23856 23800 0 _0609_
rlabel metal2 33040 27048 33040 27048 0 _0610_
rlabel metal2 30408 25900 30408 25900 0 _0611_
rlabel metal2 30968 27664 30968 27664 0 _0612_
rlabel metal3 30912 27048 30912 27048 0 _0613_
rlabel metal2 24248 24976 24248 24976 0 _0614_
rlabel metal2 22904 23800 22904 23800 0 _0615_
rlabel metal2 22792 29624 22792 29624 0 _0616_
rlabel metal2 23800 29344 23800 29344 0 _0617_
rlabel metal2 23240 24024 23240 24024 0 _0618_
rlabel metal2 10248 27664 10248 27664 0 _0619_
rlabel metal2 24024 27328 24024 27328 0 _0620_
rlabel metal2 24136 26712 24136 26712 0 _0621_
rlabel metal2 23352 24528 23352 24528 0 _0622_
rlabel metal2 22456 22008 22456 22008 0 _0623_
rlabel metal2 24808 22680 24808 22680 0 _0624_
rlabel metal2 21672 22792 21672 22792 0 _0625_
rlabel metal2 23240 21224 23240 21224 0 _0626_
rlabel metal2 23520 21784 23520 21784 0 _0627_
rlabel metal2 22568 20048 22568 20048 0 _0628_
rlabel metal3 37632 26488 37632 26488 0 _0629_
rlabel metal3 39648 24696 39648 24696 0 _0630_
rlabel metal2 38920 34776 38920 34776 0 _0631_
rlabel metal2 36568 32200 36568 32200 0 _0632_
rlabel metal2 33320 33712 33320 33712 0 _0633_
rlabel metal2 34328 38248 34328 38248 0 _0634_
rlabel metal3 35056 36568 35056 36568 0 _0635_
rlabel metal3 36400 31976 36400 31976 0 _0636_
rlabel metal2 37072 21560 37072 21560 0 _0637_
rlabel metal2 38472 15792 38472 15792 0 _0638_
rlabel metal2 27160 20272 27160 20272 0 _0639_
rlabel metal2 42616 19544 42616 19544 0 _0640_
rlabel metal2 37352 21504 37352 21504 0 _0641_
rlabel metal3 37128 15848 37128 15848 0 _0642_
rlabel metal3 37072 17752 37072 17752 0 _0643_
rlabel metal2 41608 20216 41608 20216 0 _0644_
rlabel metal3 38472 18536 38472 18536 0 _0645_
rlabel metal2 41888 20552 41888 20552 0 _0646_
rlabel metal2 38416 15400 38416 15400 0 _0647_
rlabel metal2 42952 20720 42952 20720 0 _0648_
rlabel metal3 36624 13048 36624 13048 0 _0649_
rlabel metal3 42784 39368 42784 39368 0 _0650_
rlabel metal2 49784 20216 49784 20216 0 _0651_
rlabel metal2 34664 21168 34664 21168 0 _0652_
rlabel metal2 33600 34328 33600 34328 0 _0653_
rlabel metal2 34664 34608 34664 34608 0 _0654_
rlabel metal2 28616 27720 28616 27720 0 _0655_
rlabel metal3 39704 10584 39704 10584 0 _0656_
rlabel metal3 40320 7448 40320 7448 0 _0657_
rlabel metal3 23576 19992 23576 19992 0 _0658_
rlabel metal2 25368 17584 25368 17584 0 _0659_
rlabel metal2 39480 10080 39480 10080 0 _0660_
rlabel metal2 38136 8960 38136 8960 0 _0661_
rlabel metal2 41216 9128 41216 9128 0 _0662_
rlabel metal3 41944 6664 41944 6664 0 _0663_
rlabel metal2 39256 7616 39256 7616 0 _0664_
rlabel metal3 35056 27832 35056 27832 0 _0665_
rlabel metal2 45696 39032 45696 39032 0 _0666_
rlabel metal2 29624 35336 29624 35336 0 _0667_
rlabel metal2 28056 35392 28056 35392 0 _0668_
rlabel metal2 26040 35560 26040 35560 0 _0669_
rlabel metal2 26712 34048 26712 34048 0 _0670_
rlabel metal2 48552 39424 48552 39424 0 _0671_
rlabel metal2 29568 37912 29568 37912 0 _0672_
rlabel metal2 26600 36008 26600 36008 0 _0673_
rlabel metal2 11704 37352 11704 37352 0 _0674_
rlabel metal2 45416 39760 45416 39760 0 _0675_
rlabel metal2 21952 45752 21952 45752 0 _0676_
rlabel metal3 45080 42168 45080 42168 0 _0677_
rlabel metal2 30072 38304 30072 38304 0 _0678_
rlabel metal2 23016 16800 23016 16800 0 _0679_
rlabel metal2 14280 16856 14280 16856 0 _0680_
rlabel metal2 17528 14504 17528 14504 0 _0681_
rlabel metal2 23352 37240 23352 37240 0 _0682_
rlabel metal2 44968 39312 44968 39312 0 _0683_
rlabel metal3 26432 37240 26432 37240 0 _0684_
rlabel metal2 23464 37800 23464 37800 0 _0685_
rlabel metal2 48104 42224 48104 42224 0 _0686_
rlabel metal3 26544 37800 26544 37800 0 _0687_
rlabel metal2 27272 22456 27272 22456 0 _0688_
rlabel metal2 20328 21588 20328 21588 0 _0689_
rlabel metal2 23016 21224 23016 21224 0 _0690_
rlabel metal2 24360 20832 24360 20832 0 _0691_
rlabel metal2 24024 20664 24024 20664 0 _0692_
rlabel metal2 23016 18816 23016 18816 0 _0693_
rlabel metal2 23520 18200 23520 18200 0 _0694_
rlabel metal2 24024 17444 24024 17444 0 _0695_
rlabel metal3 24248 13944 24248 13944 0 _0696_
rlabel metal2 25368 14224 25368 14224 0 _0697_
rlabel metal2 15848 21000 15848 21000 0 _0698_
rlabel metal2 16072 16408 16072 16408 0 _0699_
rlabel metal2 22736 12936 22736 12936 0 _0700_
rlabel metal2 23016 13664 23016 13664 0 _0701_
rlabel metal2 21336 13384 21336 13384 0 _0702_
rlabel metal2 16744 14280 16744 14280 0 _0703_
rlabel metal2 15512 14224 15512 14224 0 _0704_
rlabel metal3 18984 14392 18984 14392 0 _0705_
rlabel metal2 15736 12936 15736 12936 0 _0706_
rlabel metal2 10248 12376 10248 12376 0 _0707_
rlabel metal2 13888 14616 13888 14616 0 _0708_
rlabel metal2 15960 12992 15960 12992 0 _0709_
rlabel metal2 14616 11760 14616 11760 0 _0710_
rlabel metal2 13496 11760 13496 11760 0 _0711_
rlabel metal2 15624 14168 15624 14168 0 _0712_
rlabel metal2 15288 13272 15288 13272 0 _0713_
rlabel metal3 13216 11480 13216 11480 0 _0714_
rlabel metal2 11984 28280 11984 28280 0 _0715_
rlabel metal2 14224 8904 14224 8904 0 _0716_
rlabel metal2 13216 8904 13216 8904 0 _0717_
rlabel metal2 23912 15624 23912 15624 0 _0718_
rlabel metal2 10192 15736 10192 15736 0 _0719_
rlabel metal2 15176 10584 15176 10584 0 _0720_
rlabel metal2 35112 6944 35112 6944 0 _0721_
rlabel metal2 26488 6328 26488 6328 0 _0722_
rlabel metal2 34440 5208 34440 5208 0 _0723_
rlabel metal2 21728 5880 21728 5880 0 _0724_
rlabel metal2 26152 7896 26152 7896 0 _0725_
rlabel metal2 26600 10472 26600 10472 0 _0726_
rlabel metal3 23912 8008 23912 8008 0 _0727_
rlabel metal3 32480 9688 32480 9688 0 _0728_
rlabel metal3 27328 10024 27328 10024 0 _0729_
rlabel metal2 26712 6552 26712 6552 0 _0730_
rlabel metal2 27104 9800 27104 9800 0 _0731_
rlabel metal3 19656 29624 19656 29624 0 _0732_
rlabel metal2 7112 29904 7112 29904 0 _0733_
rlabel metal2 21000 7840 21000 7840 0 _0734_
rlabel metal3 21224 5096 21224 5096 0 _0735_
rlabel metal3 23408 10584 23408 10584 0 _0736_
rlabel metal2 22232 10248 22232 10248 0 _0737_
rlabel metal2 20328 10080 20328 10080 0 _0738_
rlabel metal3 22456 6776 22456 6776 0 _0739_
rlabel metal2 17976 6216 17976 6216 0 _0740_
rlabel metal3 19432 5096 19432 5096 0 _0741_
rlabel metal2 19656 7784 19656 7784 0 _0742_
rlabel metal2 19432 5152 19432 5152 0 _0743_
rlabel metal2 16464 5992 16464 5992 0 _0744_
rlabel metal2 16296 5544 16296 5544 0 _0745_
rlabel metal2 18984 5208 18984 5208 0 _0746_
rlabel metal2 21784 4760 21784 4760 0 _0747_
rlabel metal2 21560 23408 21560 23408 0 _0748_
rlabel metal2 24024 23912 24024 23912 0 _0749_
rlabel metal2 5936 22344 5936 22344 0 _0750_
rlabel metal3 13440 23800 13440 23800 0 _0751_
rlabel metal3 5544 22120 5544 22120 0 _0752_
rlabel metal2 6328 18872 6328 18872 0 _0753_
rlabel metal2 5768 21112 5768 21112 0 _0754_
rlabel metal2 7784 17696 7784 17696 0 _0755_
rlabel metal3 6944 17528 6944 17528 0 _0756_
rlabel metal2 6776 18256 6776 18256 0 _0757_
rlabel metal2 7504 15960 7504 15960 0 _0758_
rlabel metal3 9016 15176 9016 15176 0 _0759_
rlabel metal2 9632 15736 9632 15736 0 _0760_
rlabel metal2 8960 11368 8960 11368 0 _0761_
rlabel metal2 9352 6944 9352 6944 0 _0762_
rlabel metal2 39928 35672 39928 35672 0 _0763_
rlabel metal2 42392 18984 42392 18984 0 _0764_
rlabel metal2 42280 16044 42280 16044 0 _0765_
rlabel metal2 40376 40712 40376 40712 0 _0766_
rlabel metal2 43064 18536 43064 18536 0 _0767_
rlabel metal3 42224 13944 42224 13944 0 _0768_
rlabel metal3 40656 12040 40656 12040 0 _0769_
rlabel metal2 41608 14056 41608 14056 0 _0770_
rlabel metal2 42616 11480 42616 11480 0 _0771_
rlabel metal2 42280 12992 42280 12992 0 _0772_
rlabel metal3 49560 19992 49560 19992 0 _0773_
rlabel metal2 49560 19544 49560 19544 0 _0774_
rlabel metal2 50344 19824 50344 19824 0 _0775_
rlabel metal2 53144 39368 53144 39368 0 _0776_
rlabel metal2 52752 19320 52752 19320 0 _0777_
rlabel metal2 54936 39144 54936 39144 0 _0778_
rlabel metal2 55328 18536 55328 18536 0 _0779_
rlabel metal2 54376 39872 54376 39872 0 _0780_
rlabel metal3 55104 19880 55104 19880 0 _0781_
rlabel metal2 36120 33376 36120 33376 0 _0782_
rlabel metal2 37744 29400 37744 29400 0 _0783_
rlabel metal2 39704 24808 39704 24808 0 _0784_
rlabel metal2 40152 24976 40152 24976 0 _0785_
rlabel metal2 40040 25536 40040 25536 0 _0786_
rlabel metal2 41832 23800 41832 23800 0 _0787_
rlabel metal2 41384 21784 41384 21784 0 _0788_
rlabel metal2 39032 22176 39032 22176 0 _0789_
rlabel metal2 38696 38920 38696 38920 0 _0790_
rlabel metal3 44072 35112 44072 35112 0 _0791_
rlabel metal2 41888 34328 41888 34328 0 _0792_
rlabel metal3 44856 35672 44856 35672 0 _0793_
rlabel metal3 42112 34776 42112 34776 0 _0794_
rlabel metal2 43176 34720 43176 34720 0 _0795_
rlabel metal2 25368 41496 25368 41496 0 _0796_
rlabel metal2 40936 30520 40936 30520 0 _0797_
rlabel metal2 17584 40600 17584 40600 0 _0798_
rlabel metal2 39480 30240 39480 30240 0 _0799_
rlabel metal3 21784 38696 21784 38696 0 _0800_
rlabel metal2 41384 33040 41384 33040 0 _0801_
rlabel metal2 49672 35560 49672 35560 0 _0802_
rlabel metal2 50008 35112 50008 35112 0 _0803_
rlabel metal2 49784 36064 49784 36064 0 _0804_
rlabel metal3 52472 36568 52472 36568 0 _0805_
rlabel metal3 55160 35560 55160 35560 0 _0806_
rlabel metal2 54376 36792 54376 36792 0 _0807_
rlabel metal3 30464 9800 30464 9800 0 _0808_
rlabel metal2 29512 8232 29512 8232 0 _0809_
rlabel metal2 30072 6608 30072 6608 0 _0810_
rlabel metal2 25984 25816 25984 25816 0 _0811_
rlabel metal2 29848 9744 29848 9744 0 _0812_
rlabel metal3 30072 7336 30072 7336 0 _0813_
rlabel metal2 33880 7448 33880 7448 0 _0814_
rlabel metal2 34944 5992 34944 5992 0 _0815_
rlabel metal3 34384 8232 34384 8232 0 _0816_
rlabel metal2 3528 21112 3528 21112 0 _0817_
rlabel metal2 3752 19768 3752 19768 0 _0818_
rlabel metal2 3192 17080 3192 17080 0 _0819_
rlabel metal3 3416 18312 3416 18312 0 _0820_
rlabel metal2 3080 14504 3080 14504 0 _0821_
rlabel metal3 7784 31752 7784 31752 0 _0822_
rlabel metal3 3528 13608 3528 13608 0 _0823_
rlabel metal2 4144 10808 4144 10808 0 _0824_
rlabel metal3 5320 11480 5320 11480 0 _0825_
rlabel metal2 6888 9744 6888 9744 0 _0826_
rlabel metal2 9576 8960 9576 8960 0 _0827_
rlabel metal2 5992 9856 5992 9856 0 _0828_
rlabel metal2 15344 16184 15344 16184 0 _0829_
rlabel metal2 9016 9184 9016 9184 0 _0830_
rlabel metal2 20328 17472 20328 17472 0 _0831_
rlabel metal2 7336 8120 7336 8120 0 _0832_
rlabel metal2 8176 5992 8176 5992 0 _0833_
rlabel metal2 10024 7784 10024 7784 0 _0834_
rlabel metal2 38248 34944 38248 34944 0 _0835_
rlabel metal3 38192 33544 38192 33544 0 _0836_
rlabel metal3 28224 28616 28224 28616 0 _0837_
rlabel metal2 26376 28672 26376 28672 0 _0838_
rlabel metal2 26768 29176 26768 29176 0 _0839_
rlabel metal3 26152 28392 26152 28392 0 _0840_
rlabel metal2 26040 29008 26040 29008 0 _0841_
rlabel metal3 29288 41048 29288 41048 0 _0842_
rlabel metal3 25032 41944 25032 41944 0 _0843_
rlabel metal2 29400 41888 29400 41888 0 _0844_
rlabel metal2 26152 41552 26152 41552 0 _0845_
rlabel metal3 23408 39704 23408 39704 0 _0846_
rlabel metal3 23072 41944 23072 41944 0 _0847_
rlabel metal2 25928 42616 25928 42616 0 _0848_
rlabel metal2 24808 40096 24808 40096 0 _0849_
rlabel metal3 31304 42672 31304 42672 0 _0850_
rlabel metal2 30856 43232 30856 43232 0 _0851_
rlabel metal3 32704 41832 32704 41832 0 _0852_
rlabel metal3 30128 42616 30128 42616 0 _0853_
rlabel metal2 32200 44184 32200 44184 0 _0854_
rlabel metal2 30632 44688 30632 44688 0 _0855_
rlabel metal3 20356 20104 20356 20104 0 _0856_
rlabel metal2 37016 23632 37016 23632 0 _0857_
rlabel metal3 24976 5880 24976 5880 0 _0858_
rlabel metal2 26712 5432 26712 5432 0 _0859_
rlabel metal2 8400 20104 8400 20104 0 _0860_
rlabel metal2 31528 31248 31528 31248 0 _0861_
rlabel metal2 22680 32816 22680 32816 0 _0862_
rlabel metal3 34160 30968 34160 30968 0 _0863_
rlabel metal3 23408 32648 23408 32648 0 _0864_
rlabel metal2 23688 32312 23688 32312 0 _0865_
rlabel metal3 21392 31640 21392 31640 0 _0866_
rlabel metal2 29288 32144 29288 32144 0 _0867_
rlabel metal2 22456 32984 22456 32984 0 _0868_
rlabel metal3 35616 30184 35616 30184 0 _0869_
rlabel metal2 30184 30520 30184 30520 0 _0870_
rlabel metal2 43960 39592 43960 39592 0 _0871_
rlabel via2 46648 40264 46648 40264 0 _0872_
rlabel metal2 54600 39760 54600 39760 0 _0873_
rlabel metal3 47600 38808 47600 38808 0 _0874_
rlabel metal3 50008 45640 50008 45640 0 _0875_
rlabel metal3 49784 42056 49784 42056 0 _0876_
rlabel metal2 45528 42392 45528 42392 0 _0877_
rlabel metal2 51128 43848 51128 43848 0 _0878_
rlabel metal2 45360 40376 45360 40376 0 _0879_
rlabel metal2 51352 42784 51352 42784 0 _0880_
rlabel metal2 49784 40880 49784 40880 0 _0881_
rlabel metal2 49112 41552 49112 41552 0 _0882_
rlabel metal3 48552 37464 48552 37464 0 _0883_
rlabel metal3 52584 40600 52584 40600 0 _0884_
rlabel metal3 54488 43904 54488 43904 0 _0885_
rlabel metal2 52640 40152 52640 40152 0 _0886_
rlabel metal2 57064 44408 57064 44408 0 _0887_
rlabel metal2 56168 39592 56168 39592 0 _0888_
rlabel metal2 54264 47096 54264 47096 0 _0889_
rlabel metal2 54936 40992 54936 40992 0 _0890_
rlabel metal2 19096 39200 19096 39200 0 _0891_
rlabel metal2 10248 44016 10248 44016 0 _0892_
rlabel metal2 15064 46312 15064 46312 0 _0893_
rlabel metal2 13272 45472 13272 45472 0 _0894_
rlabel metal2 16632 43960 16632 43960 0 _0895_
rlabel metal3 14056 45080 14056 45080 0 _0896_
rlabel metal2 12264 45472 12264 45472 0 _0897_
rlabel metal3 10584 44072 10584 44072 0 _0898_
rlabel metal2 21056 44968 21056 44968 0 _0899_
rlabel metal2 10696 45136 10696 45136 0 _0900_
rlabel metal2 9912 44296 9912 44296 0 _0901_
rlabel metal2 19544 45528 19544 45528 0 _0902_
rlabel metal2 7784 46088 7784 46088 0 _0903_
rlabel metal2 8568 44240 8568 44240 0 _0904_
rlabel metal2 8344 45080 8344 45080 0 _0905_
rlabel metal2 8904 46928 8904 46928 0 _0906_
rlabel metal2 8120 45864 8120 45864 0 _0907_
rlabel metal2 8344 48552 8344 48552 0 _0908_
rlabel metal2 7392 45976 7392 45976 0 _0909_
rlabel metal2 12040 45416 12040 45416 0 _0910_
rlabel metal3 12152 45752 12152 45752 0 _0911_
rlabel metal3 47656 53480 47656 53480 0 _0912_
rlabel metal2 45192 51184 45192 51184 0 _0913_
rlabel metal2 45640 48496 45640 48496 0 _0914_
rlabel metal3 45640 48104 45640 48104 0 _0915_
rlabel metal2 45136 47656 45136 47656 0 _0916_
rlabel metal2 43456 47656 43456 47656 0 _0917_
rlabel metal2 42504 50064 42504 50064 0 _0918_
rlabel metal2 42392 49336 42392 49336 0 _0919_
rlabel metal2 42168 49280 42168 49280 0 _0920_
rlabel metal2 42392 48664 42392 48664 0 _0921_
rlabel metal3 39984 49000 39984 49000 0 _0922_
rlabel metal2 39816 47432 39816 47432 0 _0923_
rlabel metal2 38696 48664 38696 48664 0 _0924_
rlabel metal2 38808 48048 38808 48048 0 _0925_
rlabel metal3 41160 49560 41160 49560 0 _0926_
rlabel metal2 37464 49280 37464 49280 0 _0927_
rlabel metal2 37240 47824 37240 47824 0 _0928_
rlabel metal3 32816 48104 32816 48104 0 _0929_
rlabel metal2 37856 49000 37856 49000 0 _0930_
rlabel metal2 38584 49448 38584 49448 0 _0931_
rlabel metal2 41048 49056 41048 49056 0 _0932_
rlabel metal2 41384 49448 41384 49448 0 _0933_
rlabel metal2 42504 48272 42504 48272 0 _0934_
rlabel metal2 43064 47936 43064 47936 0 _0935_
rlabel metal2 43624 48720 43624 48720 0 _0936_
rlabel metal2 46312 46536 46312 46536 0 _0937_
rlabel metal2 54488 45640 54488 45640 0 _0938_
rlabel metal2 52808 43624 52808 43624 0 _0939_
rlabel metal2 53032 45808 53032 45808 0 _0940_
rlabel metal2 51576 44800 51576 44800 0 _0941_
rlabel metal2 50120 46536 50120 46536 0 _0942_
rlabel metal2 49896 46984 49896 46984 0 _0943_
rlabel metal2 53088 49112 53088 49112 0 _0944_
rlabel metal2 52136 44408 52136 44408 0 _0945_
rlabel metal3 54096 45080 54096 45080 0 _0946_
rlabel metal2 57288 46872 57288 46872 0 _0947_
rlabel metal2 56616 47096 56616 47096 0 _0948_
rlabel metal2 52808 46256 52808 46256 0 _0949_
rlabel metal2 54488 44744 54488 44744 0 _0950_
rlabel metal2 55048 43848 55048 43848 0 _0951_
rlabel metal3 54376 45752 54376 45752 0 _0952_
rlabel metal2 54040 46536 54040 46536 0 _0953_
rlabel metal2 54152 46256 54152 46256 0 _0954_
rlabel metal2 47208 47936 47208 47936 0 _0955_
rlabel metal3 45976 48216 45976 48216 0 _0956_
rlabel metal2 46088 47376 46088 47376 0 _0957_
rlabel metal3 51016 44296 51016 44296 0 _0958_
rlabel metal2 52024 45808 52024 45808 0 _0959_
rlabel metal2 54376 44576 54376 44576 0 _0960_
rlabel metal2 54712 44800 54712 44800 0 _0961_
rlabel metal2 46648 46592 46648 46592 0 _0962_
rlabel metal3 43904 46648 43904 46648 0 _0963_
rlabel metal2 41552 48216 41552 48216 0 _0964_
rlabel metal2 39256 47432 39256 47432 0 _0965_
rlabel metal2 36792 47040 36792 47040 0 _0966_
rlabel metal2 39928 47600 39928 47600 0 _0967_
rlabel metal2 44632 48440 44632 48440 0 _0968_
rlabel metal2 44520 47936 44520 47936 0 _0969_
rlabel metal3 40376 48160 40376 48160 0 _0970_
rlabel metal3 40768 47992 40768 47992 0 _0971_
rlabel metal2 40712 47768 40712 47768 0 _0972_
rlabel metal2 40824 46928 40824 46928 0 _0973_
rlabel metal2 57512 52528 57512 52528 0 _0974_
rlabel metal2 17528 36008 17528 36008 0 _0975_
rlabel metal3 34776 48216 34776 48216 0 _0976_
rlabel metal2 20440 29904 20440 29904 0 _0977_
rlabel metal2 36232 48552 36232 48552 0 _0978_
rlabel metal2 46928 17752 46928 17752 0 _0979_
rlabel metal2 41440 18984 41440 18984 0 _0980_
rlabel metal2 42056 45976 42056 45976 0 _0981_
rlabel metal2 18648 46984 18648 46984 0 _0982_
rlabel metal2 16072 47544 16072 47544 0 _0983_
rlabel metal2 14952 46928 14952 46928 0 _0984_
rlabel metal2 16632 47432 16632 47432 0 _0985_
rlabel metal2 44968 19880 44968 19880 0 _0986_
rlabel metal2 31528 45472 31528 45472 0 _0987_
rlabel metal2 46200 50904 46200 50904 0 _0988_
rlabel metal2 51016 50120 51016 50120 0 _0989_
rlabel metal3 43848 16856 43848 16856 0 _0990_
rlabel metal2 36008 16128 36008 16128 0 _0991_
rlabel metal2 36008 51408 36008 51408 0 _0992_
rlabel metal2 37352 49420 37352 49420 0 _0993_
rlabel metal2 37352 53032 37352 53032 0 _0994_
rlabel metal3 40880 53816 40880 53816 0 _0995_
rlabel metal2 45304 52640 45304 52640 0 _0996_
rlabel metal3 40208 52920 40208 52920 0 _0997_
rlabel metal2 40376 54096 40376 54096 0 _0998_
rlabel metal3 40656 54712 40656 54712 0 _0999_
rlabel metal3 41832 55272 41832 55272 0 _1000_
rlabel metal2 43176 54656 43176 54656 0 _1001_
rlabel metal2 43064 53032 43064 53032 0 _1002_
rlabel metal3 48552 52920 48552 52920 0 _1003_
rlabel metal2 46760 53816 46760 53816 0 _1004_
rlabel metal2 44072 52192 44072 52192 0 _1005_
rlabel metal2 50568 53648 50568 53648 0 _1006_
rlabel metal2 47656 53144 47656 53144 0 _1007_
rlabel metal2 47152 54376 47152 54376 0 _1008_
rlabel metal2 50064 52136 50064 52136 0 _1009_
rlabel metal3 49000 52136 49000 52136 0 _1010_
rlabel metal2 49000 51856 49000 51856 0 _1011_
rlabel metal2 48888 51632 48888 51632 0 _1012_
rlabel metal2 50680 51072 50680 51072 0 _1013_
rlabel metal2 48552 49448 48552 49448 0 _1014_
rlabel metal2 51184 51464 51184 51464 0 _1015_
rlabel metal2 50736 50008 50736 50008 0 _1016_
rlabel metal2 51016 52416 51016 52416 0 _1017_
rlabel metal2 51128 53928 51128 53928 0 _1018_
rlabel metal2 50288 50792 50288 50792 0 _1019_
rlabel metal2 50904 53424 50904 53424 0 _1020_
rlabel metal2 53704 53760 53704 53760 0 _1021_
rlabel metal2 56840 53200 56840 53200 0 _1022_
rlabel metal3 56056 52920 56056 52920 0 _1023_
rlabel metal3 45136 43400 45136 43400 0 clknet_0_wb_clk_i
rlabel metal3 20216 25144 20216 25144 0 clknet_2_0__leaf_wb_clk_i
rlabel metal2 4984 40488 4984 40488 0 clknet_2_1__leaf_wb_clk_i
rlabel metal2 40152 23016 40152 23016 0 clknet_2_2__leaf_wb_clk_i
rlabel metal2 52920 52528 52920 52528 0 clknet_2_3__leaf_wb_clk_i
rlabel metal2 1848 26264 1848 26264 0 clknet_leaf_0_wb_clk_i
rlabel metal2 20216 46984 20216 46984 0 clknet_leaf_10_wb_clk_i
rlabel metal2 22680 51688 22680 51688 0 clknet_leaf_11_wb_clk_i
rlabel metal2 25480 54936 25480 54936 0 clknet_leaf_12_wb_clk_i
rlabel metal3 24808 39592 24808 39592 0 clknet_leaf_13_wb_clk_i
rlabel metal2 31528 32480 31528 32480 0 clknet_leaf_14_wb_clk_i
rlabel metal2 40712 43988 40712 43988 0 clknet_leaf_15_wb_clk_i
rlabel metal3 40544 45192 40544 45192 0 clknet_leaf_16_wb_clk_i
rlabel metal2 31192 46704 31192 46704 0 clknet_leaf_17_wb_clk_i
rlabel metal3 32816 55272 32816 55272 0 clknet_leaf_18_wb_clk_i
rlabel metal2 47096 48496 47096 48496 0 clknet_leaf_19_wb_clk_i
rlabel metal2 15288 23520 15288 23520 0 clknet_leaf_1_wb_clk_i
rlabel metal2 52024 54936 52024 54936 0 clknet_leaf_20_wb_clk_i
rlabel metal2 54600 50904 54600 50904 0 clknet_leaf_21_wb_clk_i
rlabel via2 51912 45192 51912 45192 0 clknet_leaf_22_wb_clk_i
rlabel metal2 52920 39480 52920 39480 0 clknet_leaf_23_wb_clk_i
rlabel metal2 55384 32536 55384 32536 0 clknet_leaf_24_wb_clk_i
rlabel metal2 46648 33264 46648 33264 0 clknet_leaf_25_wb_clk_i
rlabel metal2 45136 41160 45136 41160 0 clknet_leaf_26_wb_clk_i
rlabel metal2 41832 32200 41832 32200 0 clknet_leaf_27_wb_clk_i
rlabel metal2 41160 25536 41160 25536 0 clknet_leaf_28_wb_clk_i
rlabel metal2 45416 22960 45416 22960 0 clknet_leaf_29_wb_clk_i
rlabel metal2 17864 22512 17864 22512 0 clknet_leaf_2_wb_clk_i
rlabel metal2 55384 24696 55384 24696 0 clknet_leaf_30_wb_clk_i
rlabel metal2 55440 19208 55440 19208 0 clknet_leaf_31_wb_clk_i
rlabel metal2 51688 16464 51688 16464 0 clknet_leaf_32_wb_clk_i
rlabel metal2 55496 10808 55496 10808 0 clknet_leaf_33_wb_clk_i
rlabel metal3 49868 5096 49868 5096 0 clknet_leaf_34_wb_clk_i
rlabel metal2 44968 15596 44968 15596 0 clknet_leaf_35_wb_clk_i
rlabel metal2 40936 11032 40936 11032 0 clknet_leaf_36_wb_clk_i
rlabel metal2 41160 5824 41160 5824 0 clknet_leaf_37_wb_clk_i
rlabel metal2 36344 4704 36344 4704 0 clknet_leaf_38_wb_clk_i
rlabel metal2 34608 10584 34608 10584 0 clknet_leaf_39_wb_clk_i
rlabel metal2 21896 33768 21896 33768 0 clknet_leaf_3_wb_clk_i
rlabel metal2 41160 15148 41160 15148 0 clknet_leaf_40_wb_clk_i
rlabel metal2 32088 23240 32088 23240 0 clknet_leaf_41_wb_clk_i
rlabel metal2 30744 25928 30744 25928 0 clknet_leaf_42_wb_clk_i
rlabel metal2 22624 17640 22624 17640 0 clknet_leaf_44_wb_clk_i
rlabel metal2 26600 13160 26600 13160 0 clknet_leaf_45_wb_clk_i
rlabel metal2 25256 4648 25256 4648 0 clknet_leaf_46_wb_clk_i
rlabel metal2 20216 8344 20216 8344 0 clknet_leaf_47_wb_clk_i
rlabel metal2 17528 15204 17528 15204 0 clknet_leaf_48_wb_clk_i
rlabel metal2 17416 9352 17416 9352 0 clknet_leaf_49_wb_clk_i
rlabel metal2 12992 30968 12992 30968 0 clknet_leaf_4_wb_clk_i
rlabel metal2 13384 5040 13384 5040 0 clknet_leaf_50_wb_clk_i
rlabel metal2 1848 10584 1848 10584 0 clknet_leaf_51_wb_clk_i
rlabel metal3 8848 18424 8848 18424 0 clknet_leaf_52_wb_clk_i
rlabel metal2 1848 22400 1848 22400 0 clknet_leaf_53_wb_clk_i
rlabel metal2 4984 33656 4984 33656 0 clknet_leaf_5_wb_clk_i
rlabel metal2 1848 40040 1848 40040 0 clknet_leaf_6_wb_clk_i
rlabel metal2 10304 46648 10304 46648 0 clknet_leaf_7_wb_clk_i
rlabel metal2 6216 47880 6216 47880 0 clknet_leaf_8_wb_clk_i
rlabel metal2 14336 49784 14336 49784 0 clknet_leaf_9_wb_clk_i
rlabel metal2 58184 50120 58184 50120 0 custom_settings[0]
rlabel metal3 58730 56056 58730 56056 0 custom_settings[1]
rlabel metal2 58184 3976 58184 3976 0 io_in_1[0]
rlabel metal2 58184 9352 58184 9352 0 io_in_1[1]
rlabel metal3 58730 15288 58730 15288 0 io_in_1[2]
rlabel metal2 58184 21336 58184 21336 0 io_in_1[3]
rlabel metal2 58184 26656 58184 26656 0 io_in_1[4]
rlabel metal3 58730 32760 58730 32760 0 io_in_1[5]
rlabel metal2 58072 39536 58072 39536 0 io_in_1[6]
rlabel metal2 58240 45640 58240 45640 0 io_in_1[7]
rlabel metal2 37464 57778 37464 57778 0 io_in_2[0]
rlabel metal2 52472 57778 52472 57778 0 io_in_2[1]
rlabel metal3 23520 5208 23520 5208 0 io_out[10]
rlabel metal3 25536 3640 25536 3640 0 io_out[11]
rlabel metal2 37016 854 37016 854 0 io_out[17]
rlabel metal2 39032 1190 39032 1190 0 io_out[18]
rlabel metal3 41888 5208 41888 5208 0 io_out[19]
rlabel metal3 44240 4088 44240 4088 0 io_out[20]
rlabel metal3 47040 3416 47040 3416 0 io_out[21]
rlabel metal2 18872 2198 18872 2198 0 io_out[8]
rlabel metal3 21504 3640 21504 3640 0 io_out[9]
rlabel metal3 43680 49840 43680 49840 0 net1
rlabel metal2 54824 40040 54824 40040 0 net10
rlabel metal2 37240 39592 37240 39592 0 net11
rlabel metal2 52136 41048 52136 41048 0 net12
rlabel metal2 26488 20888 26488 20888 0 net13
rlabel metal2 23128 4648 23128 4648 0 net14
rlabel metal2 20328 6496 20328 6496 0 net15
rlabel metal2 28168 3864 28168 3864 0 net16
rlabel metal2 39032 3864 39032 3864 0 net17
rlabel metal2 41384 5152 41384 5152 0 net18
rlabel metal3 26432 21448 26432 21448 0 net19
rlabel metal2 57680 55384 57680 55384 0 net2
rlabel metal2 48888 3864 48888 3864 0 net20
rlabel metal2 20384 15176 20384 15176 0 net21
rlabel metal2 12824 4368 12824 4368 0 net22
rlabel metal2 2744 2030 2744 2030 0 net23
rlabel metal2 4760 2030 4760 2030 0 net24
rlabel metal2 6776 2030 6776 2030 0 net25
rlabel metal2 8792 854 8792 854 0 net26
rlabel metal2 10808 2030 10808 2030 0 net27
rlabel metal2 12824 2030 12824 2030 0 net28
rlabel metal2 14840 2030 14840 2030 0 net29
rlabel metal2 39648 10024 39648 10024 0 net3
rlabel metal2 16856 2030 16856 2030 0 net30
rlabel metal2 26936 1246 26936 1246 0 net31
rlabel metal2 28952 2030 28952 2030 0 net32
rlabel metal2 30968 2030 30968 2030 0 net33
rlabel metal2 32984 2030 32984 2030 0 net34
rlabel metal2 35000 2030 35000 2030 0 net35
rlabel metal2 49112 1246 49112 1246 0 net36
rlabel metal2 51128 2030 51128 2030 0 net37
rlabel metal2 53144 2030 53144 2030 0 net38
rlabel metal2 55160 2030 55160 2030 0 net39
rlabel metal3 42784 20104 42784 20104 0 net4
rlabel metal2 57176 2030 57176 2030 0 net40
rlabel metal2 47096 854 47096 854 0 net41
rlabel metal2 42728 20104 42728 20104 0 net5
rlabel metal2 42504 21616 42504 21616 0 net6
rlabel metal2 57848 26684 57848 26684 0 net7
rlabel metal3 44128 41160 44128 41160 0 net8
rlabel metal3 56896 39032 56896 39032 0 net9
rlabel metal2 22456 57778 22456 57778 0 rst_n
rlabel metal2 33432 39144 33432 39144 0 tt_um_rejunity_ay8913.active
rlabel metal2 26488 30184 26488 30184 0 tt_um_rejunity_ay8913.amplitude_A\[0\]
rlabel metal3 24920 26264 24920 26264 0 tt_um_rejunity_ay8913.amplitude_B\[0\]
rlabel metal3 35448 26712 35448 26712 0 tt_um_rejunity_ay8913.amplitude_C\[0\]
rlabel metal2 14616 34832 14616 34832 0 tt_um_rejunity_ay8913.clk_counter\[0\]
rlabel metal2 16072 36848 16072 36848 0 tt_um_rejunity_ay8913.clk_counter\[1\]
rlabel via2 16408 35224 16408 35224 0 tt_um_rejunity_ay8913.clk_counter\[2\]
rlabel metal2 17976 31248 17976 31248 0 tt_um_rejunity_ay8913.clk_counter\[3\]
rlabel metal3 16576 30184 16576 30184 0 tt_um_rejunity_ay8913.clk_counter\[4\]
rlabel metal3 17752 28504 17752 28504 0 tt_um_rejunity_ay8913.clk_counter\[5\]
rlabel metal2 16800 26264 16800 26264 0 tt_um_rejunity_ay8913.clk_counter\[6\]
rlabel metal2 24248 29624 24248 29624 0 tt_um_rejunity_ay8913.envelope_A
rlabel metal3 23520 26824 23520 26824 0 tt_um_rejunity_ay8913.envelope_B
rlabel metal2 27944 25760 27944 25760 0 tt_um_rejunity_ay8913.envelope_C
rlabel metal2 17528 41216 17528 41216 0 tt_um_rejunity_ay8913.envelope_alternate
rlabel metal2 14280 40320 14280 40320 0 tt_um_rejunity_ay8913.envelope_attack
rlabel metal2 18536 39480 18536 39480 0 tt_um_rejunity_ay8913.envelope_continue
rlabel metal2 11368 41496 11368 41496 0 tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[0\]
rlabel metal2 8232 44016 8232 44016 0 tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[1\]
rlabel metal2 8456 45416 8456 45416 0 tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[2\]
rlabel metal3 5488 45864 5488 45864 0 tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[3\]
rlabel metal2 14672 44408 14672 44408 0 tt_um_rejunity_ay8913.envelope_generator.hold
rlabel metal2 14840 44296 14840 44296 0 tt_um_rejunity_ay8913.envelope_generator.invert_output
rlabel metal2 37576 41832 37576 41832 0 tt_um_rejunity_ay8913.envelope_generator.period\[0\]
rlabel metal2 48104 41328 48104 41328 0 tt_um_rejunity_ay8913.envelope_generator.period\[10\]
rlabel metal3 52584 41832 52584 41832 0 tt_um_rejunity_ay8913.envelope_generator.period\[11\]
rlabel metal2 53704 45024 53704 45024 0 tt_um_rejunity_ay8913.envelope_generator.period\[12\]
rlabel metal3 54880 43736 54880 43736 0 tt_um_rejunity_ay8913.envelope_generator.period\[13\]
rlabel metal2 56840 44436 56840 44436 0 tt_um_rejunity_ay8913.envelope_generator.period\[14\]
rlabel metal3 57848 44408 57848 44408 0 tt_um_rejunity_ay8913.envelope_generator.period\[15\]
rlabel metal3 38080 43512 38080 43512 0 tt_um_rejunity_ay8913.envelope_generator.period\[1\]
rlabel metal2 37632 42728 37632 42728 0 tt_um_rejunity_ay8913.envelope_generator.period\[2\]
rlabel metal2 39760 45752 39760 45752 0 tt_um_rejunity_ay8913.envelope_generator.period\[3\]
rlabel metal2 42112 48776 42112 48776 0 tt_um_rejunity_ay8913.envelope_generator.period\[4\]
rlabel metal2 44072 48496 44072 48496 0 tt_um_rejunity_ay8913.envelope_generator.period\[5\]
rlabel metal2 45864 47880 45864 47880 0 tt_um_rejunity_ay8913.envelope_generator.period\[6\]
rlabel metal2 47096 44632 47096 44632 0 tt_um_rejunity_ay8913.envelope_generator.period\[7\]
rlabel metal2 49896 44968 49896 44968 0 tt_um_rejunity_ay8913.envelope_generator.period\[8\]
rlabel metal3 48664 44968 48664 44968 0 tt_um_rejunity_ay8913.envelope_generator.period\[9\]
rlabel metal2 14616 46760 14616 46760 0 tt_um_rejunity_ay8913.envelope_generator.signal_edge.previous_signal_state_0
rlabel metal3 16632 47208 16632 47208 0 tt_um_rejunity_ay8913.envelope_generator.signal_edge.signal
rlabel metal2 12488 45472 12488 45472 0 tt_um_rejunity_ay8913.envelope_generator.stop
rlabel metal2 36568 46872 36568 46872 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[0\]
rlabel metal2 51688 48496 51688 48496 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[10\]
rlabel metal2 51688 52584 51688 52584 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[11\]
rlabel metal2 55384 54544 55384 54544 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[12\]
rlabel metal2 55272 52696 55272 52696 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[13\]
rlabel metal2 58184 49168 58184 49168 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[14\]
rlabel metal2 55272 47488 55272 47488 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[15\]
rlabel metal2 36568 49280 36568 49280 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[1\]
rlabel metal2 36568 54432 36568 54432 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[2\]
rlabel metal2 41608 52864 41608 52864 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[3\]
rlabel metal2 41832 55048 41832 55048 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[4\]
rlabel metal2 42616 52920 42616 52920 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[5\]
rlabel metal2 45528 51352 45528 51352 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[6\]
rlabel metal2 48720 53704 48720 53704 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[7\]
rlabel metal2 53704 48440 53704 48440 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[8\]
rlabel metal2 50456 46368 50456 46368 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[9\]
rlabel metal2 34104 33264 34104 33264 0 tt_um_rejunity_ay8913.latched_register\[0\]
rlabel metal2 33208 34272 33208 34272 0 tt_um_rejunity_ay8913.latched_register\[1\]
rlabel metal2 39928 34608 39928 34608 0 tt_um_rejunity_ay8913.latched_register\[2\]
rlabel metal3 39368 36904 39368 36904 0 tt_um_rejunity_ay8913.latched_register\[3\]
rlabel metal2 22120 31808 22120 31808 0 tt_um_rejunity_ay8913.noise_disable_A
rlabel metal2 23912 28224 23912 28224 0 tt_um_rejunity_ay8913.noise_disable_B
rlabel metal2 32536 29008 32536 29008 0 tt_um_rejunity_ay8913.noise_disable_C
rlabel metal2 23128 28336 23128 28336 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[0\]
rlabel metal2 4760 36568 4760 36568 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[10\]
rlabel metal2 5544 37520 5544 37520 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[11\]
rlabel metal2 6776 37744 6776 37744 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[12\]
rlabel metal2 7672 37408 7672 37408 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[13\]
rlabel metal2 9576 37968 9576 37968 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[14\]
rlabel metal2 8344 37520 8344 37520 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[15\]
rlabel metal2 8120 36456 8120 36456 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[16\]
rlabel metal2 11256 27888 11256 27888 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[1\]
rlabel metal2 11592 29960 11592 29960 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[2\]
rlabel metal3 9352 28616 9352 28616 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[3\]
rlabel metal2 8288 27608 8288 27608 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[4\]
rlabel metal2 5768 26992 5768 26992 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[5\]
rlabel metal2 5096 28728 5096 28728 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[6\]
rlabel metal2 4984 29680 4984 29680 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[7\]
rlabel metal2 4312 30968 4312 30968 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[8\]
rlabel metal2 4648 33096 4648 33096 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[9\]
rlabel metal2 37240 18256 37240 18256 0 tt_um_rejunity_ay8913.noise_generator.period\[0\]
rlabel metal3 36400 19096 36400 19096 0 tt_um_rejunity_ay8913.noise_generator.period\[1\]
rlabel metal2 37856 13832 37856 13832 0 tt_um_rejunity_ay8913.noise_generator.period\[2\]
rlabel metal2 35896 11928 35896 11928 0 tt_um_rejunity_ay8913.noise_generator.period\[3\]
rlabel metal2 36008 21112 36008 21112 0 tt_um_rejunity_ay8913.noise_generator.period\[4\]
rlabel metal2 9576 22736 9576 22736 0 tt_um_rejunity_ay8913.noise_generator.signal_edge.previous_signal_state_0
rlabel metal2 25816 16632 25816 16632 0 tt_um_rejunity_ay8913.noise_generator.signal_edge.signal
rlabel metal3 32928 18536 32928 18536 0 tt_um_rejunity_ay8913.noise_generator.tone.counter\[0\]
rlabel metal2 33208 17808 33208 17808 0 tt_um_rejunity_ay8913.noise_generator.tone.counter\[1\]
rlabel metal3 32032 15176 32032 15176 0 tt_um_rejunity_ay8913.noise_generator.tone.counter\[2\]
rlabel metal3 32200 12824 32200 12824 0 tt_um_rejunity_ay8913.noise_generator.tone.counter\[3\]
rlabel metal2 33992 12152 33992 12152 0 tt_um_rejunity_ay8913.noise_generator.tone.counter\[4\]
rlabel metal2 18200 22512 18200 22512 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[2\]
rlabel metal2 13440 21784 13440 21784 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[3\]
rlabel metal2 12936 20272 12936 20272 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[4\]
rlabel metal3 13608 18424 13608 18424 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[5\]
rlabel metal2 16520 18984 16520 18984 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[6\]
rlabel metal2 17920 20888 17920 20888 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[7\]
rlabel metal2 19208 17192 19208 17192 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[8\]
rlabel metal2 4648 20944 4648 20944 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[2\]
rlabel metal2 4648 17808 4648 17808 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[3\]
rlabel metal2 4088 15148 4088 15148 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[4\]
rlabel metal2 4648 11424 4648 11424 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[5\]
rlabel metal2 5656 10080 5656 10080 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[6\]
rlabel metal2 7336 9576 7336 9576 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[7\]
rlabel metal2 7784 7784 7784 7784 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[8\]
rlabel metal2 22344 23968 22344 23968 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[2\]
rlabel metal2 14280 23968 14280 23968 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[3\]
rlabel metal2 5656 22176 5656 22176 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[4\]
rlabel metal2 6664 17976 6664 17976 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[5\]
rlabel metal2 7784 16128 7784 16128 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[6\]
rlabel metal2 8904 16128 8904 16128 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[7\]
rlabel via2 9240 12152 9240 12152 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[8\]
rlabel metal3 25200 22456 25200 22456 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[2\]
rlabel metal2 25592 18032 25592 18032 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[3\]
rlabel metal2 23632 15400 23632 15400 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[4\]
rlabel metal3 22176 13048 22176 13048 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[5\]
rlabel metal3 13440 13608 13440 13608 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[6\]
rlabel metal2 18312 11760 18312 11760 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[7\]
rlabel metal2 12936 11928 12936 11928 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[8\]
rlabel metal2 14056 8848 14056 8848 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[9\]
rlabel metal3 20160 44856 20160 44856 0 tt_um_rejunity_ay8913.restart_envelope
rlabel metal2 32200 4592 32200 4592 0 tt_um_rejunity_ay8913.spi_dac_i_2.counter\[0\]
rlabel metal2 30632 10136 30632 10136 0 tt_um_rejunity_ay8913.spi_dac_i_2.counter\[1\]
rlabel metal2 31640 7112 31640 7112 0 tt_um_rejunity_ay8913.spi_dac_i_2.counter\[2\]
rlabel metal2 33544 5936 33544 5936 0 tt_um_rejunity_ay8913.spi_dac_i_2.counter\[3\]
rlabel metal2 34440 8064 34440 8064 0 tt_um_rejunity_ay8913.spi_dac_i_2.counter\[4\]
rlabel metal3 20048 4872 20048 4872 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[10\]
rlabel metal2 24304 4200 24304 4200 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[11\]
rlabel metal2 26712 7504 26712 7504 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[2\]
rlabel metal2 25368 10864 25368 10864 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[3\]
rlabel metal2 23688 11144 23688 11144 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[4\]
rlabel metal2 22680 8568 22680 8568 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[5\]
rlabel metal3 23576 6664 23576 6664 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[6\]
rlabel metal3 18480 6664 18480 6664 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[7\]
rlabel metal2 16968 6216 16968 6216 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[8\]
rlabel metal3 17472 5096 17472 5096 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[9\]
rlabel via2 25480 30968 25480 30968 0 tt_um_rejunity_ay8913.tone_A
rlabel metal2 25592 50568 25592 50568 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[0\]
rlabel metal3 21224 48888 21224 48888 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[10\]
rlabel metal2 24192 47432 24192 47432 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[11\]
rlabel metal3 29064 50568 29064 50568 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[1\]
rlabel metal2 31416 49728 31416 49728 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[2\]
rlabel metal2 26376 53312 26376 53312 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[3\]
rlabel metal2 28392 51240 28392 51240 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[4\]
rlabel metal2 29120 45864 29120 45864 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[5\]
rlabel metal2 20664 54432 20664 54432 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[6\]
rlabel metal3 22512 53704 22512 53704 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[7\]
rlabel metal2 23408 45528 23408 45528 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[8\]
rlabel metal2 22568 47880 22568 47880 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[9\]
rlabel metal2 24136 40768 24136 40768 0 tt_um_rejunity_ay8913.tone_A_generator.period\[0\]
rlabel metal3 23240 45080 23240 45080 0 tt_um_rejunity_ay8913.tone_A_generator.period\[10\]
rlabel metal2 23016 44632 23016 44632 0 tt_um_rejunity_ay8913.tone_A_generator.period\[11\]
rlabel metal2 25368 48104 25368 48104 0 tt_um_rejunity_ay8913.tone_A_generator.period\[1\]
rlabel metal2 26488 42448 26488 42448 0 tt_um_rejunity_ay8913.tone_A_generator.period\[2\]
rlabel metal2 26712 44296 26712 44296 0 tt_um_rejunity_ay8913.tone_A_generator.period\[3\]
rlabel metal2 31864 41888 31864 41888 0 tt_um_rejunity_ay8913.tone_A_generator.period\[4\]
rlabel metal2 30520 42728 30520 42728 0 tt_um_rejunity_ay8913.tone_A_generator.period\[5\]
rlabel metal2 31528 44016 31528 44016 0 tt_um_rejunity_ay8913.tone_A_generator.period\[6\]
rlabel metal2 26824 46200 26824 46200 0 tt_um_rejunity_ay8913.tone_A_generator.period\[7\]
rlabel metal2 27272 36568 27272 36568 0 tt_um_rejunity_ay8913.tone_A_generator.period\[8\]
rlabel metal2 29680 38696 29680 38696 0 tt_um_rejunity_ay8913.tone_A_generator.period\[9\]
rlabel metal2 22904 25984 22904 25984 0 tt_um_rejunity_ay8913.tone_B
rlabel metal2 47544 26208 47544 26208 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[0\]
rlabel metal2 52136 22400 52136 22400 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[10\]
rlabel metal3 48832 21448 48832 21448 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[11\]
rlabel metal2 43848 28168 43848 28168 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[1\]
rlabel metal2 47432 31472 47432 31472 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[2\]
rlabel metal2 49560 33040 49560 33040 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[3\]
rlabel metal3 55048 33320 55048 33320 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[4\]
rlabel metal3 53088 31864 53088 31864 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[5\]
rlabel metal2 54936 29288 54936 29288 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[6\]
rlabel metal2 55720 25928 55720 25928 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[7\]
rlabel metal2 56952 24360 56952 24360 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[8\]
rlabel metal2 55720 22848 55720 22848 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[9\]
rlabel metal2 46088 34384 46088 34384 0 tt_um_rejunity_ay8913.tone_B_generator.period\[0\]
rlabel metal3 42952 22456 42952 22456 0 tt_um_rejunity_ay8913.tone_B_generator.period\[10\]
rlabel metal3 39760 22456 39760 22456 0 tt_um_rejunity_ay8913.tone_B_generator.period\[11\]
rlabel metal3 43176 28728 43176 28728 0 tt_um_rejunity_ay8913.tone_B_generator.period\[1\]
rlabel metal3 40768 30968 40768 30968 0 tt_um_rejunity_ay8913.tone_B_generator.period\[2\]
rlabel metal2 44744 32816 44744 32816 0 tt_um_rejunity_ay8913.tone_B_generator.period\[3\]
rlabel metal2 51576 35728 51576 35728 0 tt_um_rejunity_ay8913.tone_B_generator.period\[4\]
rlabel metal3 53760 33992 53760 33992 0 tt_um_rejunity_ay8913.tone_B_generator.period\[5\]
rlabel metal3 56672 35784 56672 35784 0 tt_um_rejunity_ay8913.tone_B_generator.period\[6\]
rlabel metal2 53480 26236 53480 26236 0 tt_um_rejunity_ay8913.tone_B_generator.period\[7\]
rlabel metal2 41496 25424 41496 25424 0 tt_um_rejunity_ay8913.tone_B_generator.period\[8\]
rlabel metal2 43960 24528 43960 24528 0 tt_um_rejunity_ay8913.tone_B_generator.period\[9\]
rlabel metal3 29456 23016 29456 23016 0 tt_um_rejunity_ay8913.tone_C
rlabel metal2 46984 19600 46984 19600 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[0\]
rlabel metal2 46424 5376 46424 5376 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[10\]
rlabel metal2 46536 4312 46536 4312 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[11\]
rlabel metal2 47712 16184 47712 16184 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[1\]
rlabel metal2 48216 16464 48216 16464 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[2\]
rlabel metal2 49336 14224 49336 14224 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[3\]
rlabel metal2 49784 13664 49784 13664 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[4\]
rlabel metal2 53144 11424 53144 11424 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[5\]
rlabel metal2 53648 10808 53648 10808 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[6\]
rlabel metal2 52920 7504 52920 7504 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[7\]
rlabel metal2 50344 8372 50344 8372 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[8\]
rlabel metal2 47432 7000 47432 7000 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[9\]
rlabel metal2 45864 12152 45864 12152 0 tt_um_rejunity_ay8913.tone_C_generator.period\[0\]
rlabel metal3 43792 7448 43792 7448 0 tt_um_rejunity_ay8913.tone_C_generator.period\[10\]
rlabel metal2 40320 5768 40320 5768 0 tt_um_rejunity_ay8913.tone_C_generator.period\[11\]
rlabel metal2 43848 14224 43848 14224 0 tt_um_rejunity_ay8913.tone_C_generator.period\[1\]
rlabel metal3 47880 11592 47880 11592 0 tt_um_rejunity_ay8913.tone_C_generator.period\[2\]
rlabel metal2 49224 12488 49224 12488 0 tt_um_rejunity_ay8913.tone_C_generator.period\[3\]
rlabel metal2 49448 19264 49448 19264 0 tt_um_rejunity_ay8913.tone_C_generator.period\[4\]
rlabel metal2 54040 17864 54040 17864 0 tt_um_rejunity_ay8913.tone_C_generator.period\[5\]
rlabel metal2 54040 16520 54040 16520 0 tt_um_rejunity_ay8913.tone_C_generator.period\[6\]
rlabel metal2 54488 19656 54488 19656 0 tt_um_rejunity_ay8913.tone_C_generator.period\[7\]
rlabel metal2 39536 8904 39536 8904 0 tt_um_rejunity_ay8913.tone_C_generator.period\[8\]
rlabel via2 44296 9016 44296 9016 0 tt_um_rejunity_ay8913.tone_C_generator.period\[9\]
rlabel metal2 24696 31416 24696 31416 0 tt_um_rejunity_ay8913.tone_disable_A
rlabel metal2 23072 26264 23072 26264 0 tt_um_rejunity_ay8913.tone_disable_B
rlabel metal2 30464 32424 30464 32424 0 tt_um_rejunity_ay8913.tone_disable_C
rlabel metal2 7504 43680 7504 43680 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
