magic
tech gf180mcuD
magscale 1 10
timestamp 1698874738
<< metal1 >>
rect 1344 32170 34608 32204
rect 1344 32118 5372 32170
rect 5424 32118 5476 32170
rect 5528 32118 5580 32170
rect 5632 32118 13688 32170
rect 13740 32118 13792 32170
rect 13844 32118 13896 32170
rect 13948 32118 22004 32170
rect 22056 32118 22108 32170
rect 22160 32118 22212 32170
rect 22264 32118 30320 32170
rect 30372 32118 30424 32170
rect 30476 32118 30528 32170
rect 30580 32118 34608 32170
rect 1344 32084 34608 32118
rect 1344 31386 34768 31420
rect 1344 31334 9530 31386
rect 9582 31334 9634 31386
rect 9686 31334 9738 31386
rect 9790 31334 17846 31386
rect 17898 31334 17950 31386
rect 18002 31334 18054 31386
rect 18106 31334 26162 31386
rect 26214 31334 26266 31386
rect 26318 31334 26370 31386
rect 26422 31334 34478 31386
rect 34530 31334 34582 31386
rect 34634 31334 34686 31386
rect 34738 31334 34768 31386
rect 1344 31300 34768 31334
rect 1344 30602 34608 30636
rect 1344 30550 5372 30602
rect 5424 30550 5476 30602
rect 5528 30550 5580 30602
rect 5632 30550 13688 30602
rect 13740 30550 13792 30602
rect 13844 30550 13896 30602
rect 13948 30550 22004 30602
rect 22056 30550 22108 30602
rect 22160 30550 22212 30602
rect 22264 30550 30320 30602
rect 30372 30550 30424 30602
rect 30476 30550 30528 30602
rect 30580 30550 34608 30602
rect 1344 30516 34608 30550
rect 1344 29818 34768 29852
rect 1344 29766 9530 29818
rect 9582 29766 9634 29818
rect 9686 29766 9738 29818
rect 9790 29766 17846 29818
rect 17898 29766 17950 29818
rect 18002 29766 18054 29818
rect 18106 29766 26162 29818
rect 26214 29766 26266 29818
rect 26318 29766 26370 29818
rect 26422 29766 34478 29818
rect 34530 29766 34582 29818
rect 34634 29766 34686 29818
rect 34738 29766 34768 29818
rect 1344 29732 34768 29766
rect 1344 29034 34608 29068
rect 1344 28982 5372 29034
rect 5424 28982 5476 29034
rect 5528 28982 5580 29034
rect 5632 28982 13688 29034
rect 13740 28982 13792 29034
rect 13844 28982 13896 29034
rect 13948 28982 22004 29034
rect 22056 28982 22108 29034
rect 22160 28982 22212 29034
rect 22264 28982 30320 29034
rect 30372 28982 30424 29034
rect 30476 28982 30528 29034
rect 30580 28982 34608 29034
rect 1344 28948 34608 28982
rect 11218 28702 11230 28754
rect 11282 28702 11294 28754
rect 8418 28590 8430 28642
rect 8482 28590 8494 28642
rect 9090 28478 9102 28530
rect 9154 28478 9166 28530
rect 1344 28250 34768 28284
rect 1344 28198 9530 28250
rect 9582 28198 9634 28250
rect 9686 28198 9738 28250
rect 9790 28198 17846 28250
rect 17898 28198 17950 28250
rect 18002 28198 18054 28250
rect 18106 28198 26162 28250
rect 26214 28198 26266 28250
rect 26318 28198 26370 28250
rect 26422 28198 34478 28250
rect 34530 28198 34582 28250
rect 34634 28198 34686 28250
rect 34738 28198 34768 28250
rect 1344 28164 34768 28198
rect 5070 27970 5122 27982
rect 5070 27906 5122 27918
rect 4510 27858 4562 27870
rect 4274 27806 4286 27858
rect 4338 27806 4350 27858
rect 4510 27794 4562 27806
rect 4846 27858 4898 27870
rect 4846 27794 4898 27806
rect 5182 27858 5234 27870
rect 20078 27858 20130 27870
rect 10210 27806 10222 27858
rect 10274 27806 10286 27858
rect 5182 27794 5234 27806
rect 20078 27794 20130 27806
rect 20302 27858 20354 27870
rect 20302 27794 20354 27806
rect 20638 27858 20690 27870
rect 20638 27794 20690 27806
rect 3614 27746 3666 27758
rect 20526 27746 20578 27758
rect 10994 27694 11006 27746
rect 11058 27694 11070 27746
rect 13122 27694 13134 27746
rect 13186 27694 13198 27746
rect 3614 27682 3666 27694
rect 20526 27682 20578 27694
rect 1344 27466 34608 27500
rect 1344 27414 5372 27466
rect 5424 27414 5476 27466
rect 5528 27414 5580 27466
rect 5632 27414 13688 27466
rect 13740 27414 13792 27466
rect 13844 27414 13896 27466
rect 13948 27414 22004 27466
rect 22056 27414 22108 27466
rect 22160 27414 22212 27466
rect 22264 27414 30320 27466
rect 30372 27414 30424 27466
rect 30476 27414 30528 27466
rect 30580 27414 34608 27466
rect 1344 27380 34608 27414
rect 5854 27298 5906 27310
rect 5854 27234 5906 27246
rect 4958 27186 5010 27198
rect 12238 27186 12290 27198
rect 4610 27134 4622 27186
rect 4674 27134 4686 27186
rect 10210 27134 10222 27186
rect 10274 27134 10286 27186
rect 17042 27134 17054 27186
rect 17106 27134 17118 27186
rect 20290 27134 20302 27186
rect 20354 27134 20366 27186
rect 4958 27122 5010 27134
rect 12238 27122 12290 27134
rect 5966 27074 6018 27086
rect 1810 27022 1822 27074
rect 1874 27022 1886 27074
rect 5966 27010 6018 27022
rect 6190 27074 6242 27086
rect 6190 27010 6242 27022
rect 6750 27074 6802 27086
rect 12014 27074 12066 27086
rect 7410 27022 7422 27074
rect 7474 27022 7486 27074
rect 14242 27022 14254 27074
rect 14306 27022 14318 27074
rect 17490 27022 17502 27074
rect 17554 27022 17566 27074
rect 6750 27010 6802 27022
rect 12014 27010 12066 27022
rect 5070 26962 5122 26974
rect 2482 26910 2494 26962
rect 2546 26910 2558 26962
rect 5070 26898 5122 26910
rect 6302 26962 6354 26974
rect 6302 26898 6354 26910
rect 6638 26962 6690 26974
rect 6638 26898 6690 26910
rect 6862 26962 6914 26974
rect 12462 26962 12514 26974
rect 8082 26910 8094 26962
rect 8146 26910 8158 26962
rect 6862 26898 6914 26910
rect 12462 26898 12514 26910
rect 12686 26962 12738 26974
rect 20638 26962 20690 26974
rect 14914 26910 14926 26962
rect 14978 26910 14990 26962
rect 18162 26910 18174 26962
rect 18226 26910 18238 26962
rect 12686 26898 12738 26910
rect 20638 26898 20690 26910
rect 20750 26962 20802 26974
rect 20750 26898 20802 26910
rect 1344 26682 34768 26716
rect 1344 26630 9530 26682
rect 9582 26630 9634 26682
rect 9686 26630 9738 26682
rect 9790 26630 17846 26682
rect 17898 26630 17950 26682
rect 18002 26630 18054 26682
rect 18106 26630 26162 26682
rect 26214 26630 26266 26682
rect 26318 26630 26370 26682
rect 26422 26630 34478 26682
rect 34530 26630 34582 26682
rect 34634 26630 34686 26682
rect 34738 26630 34768 26682
rect 1344 26596 34768 26630
rect 9886 26514 9938 26526
rect 9886 26450 9938 26462
rect 16382 26514 16434 26526
rect 16382 26450 16434 26462
rect 18174 26514 18226 26526
rect 18174 26450 18226 26462
rect 18958 26514 19010 26526
rect 18958 26450 19010 26462
rect 18286 26402 18338 26414
rect 7298 26350 7310 26402
rect 7362 26350 7374 26402
rect 18286 26338 18338 26350
rect 18510 26402 18562 26414
rect 18510 26338 18562 26350
rect 19070 26402 19122 26414
rect 25230 26402 25282 26414
rect 20514 26350 20526 26402
rect 20578 26350 20590 26402
rect 19070 26338 19122 26350
rect 25230 26338 25282 26350
rect 12350 26290 12402 26302
rect 16270 26290 16322 26302
rect 1810 26238 1822 26290
rect 1874 26238 1886 26290
rect 7970 26238 7982 26290
rect 8034 26238 8046 26290
rect 11778 26238 11790 26290
rect 11842 26238 11854 26290
rect 13122 26238 13134 26290
rect 13186 26238 13198 26290
rect 12350 26226 12402 26238
rect 16270 26226 16322 26238
rect 16494 26290 16546 26302
rect 16494 26226 16546 26238
rect 16942 26290 16994 26302
rect 16942 26226 16994 26238
rect 17838 26290 17890 26302
rect 17838 26226 17890 26238
rect 18846 26290 18898 26302
rect 18846 26226 18898 26238
rect 19518 26290 19570 26302
rect 23214 26290 23266 26302
rect 19730 26238 19742 26290
rect 19794 26238 19806 26290
rect 22978 26238 22990 26290
rect 23042 26238 23054 26290
rect 19518 26226 19570 26238
rect 23214 26226 23266 26238
rect 23326 26290 23378 26302
rect 23326 26226 23378 26238
rect 25566 26290 25618 26302
rect 25566 26226 25618 26238
rect 25678 26290 25730 26302
rect 25678 26226 25730 26238
rect 9998 26178 10050 26190
rect 2482 26126 2494 26178
rect 2546 26126 2558 26178
rect 4610 26126 4622 26178
rect 4674 26126 4686 26178
rect 5170 26126 5182 26178
rect 5234 26126 5246 26178
rect 9998 26114 10050 26126
rect 12462 26178 12514 26190
rect 25342 26178 25394 26190
rect 13794 26126 13806 26178
rect 13858 26126 13870 26178
rect 15922 26126 15934 26178
rect 15986 26126 15998 26178
rect 22642 26126 22654 26178
rect 22706 26126 22718 26178
rect 12462 26114 12514 26126
rect 25342 26114 25394 26126
rect 23762 26014 23774 26066
rect 23826 26014 23838 26066
rect 1344 25898 34608 25932
rect 1344 25846 5372 25898
rect 5424 25846 5476 25898
rect 5528 25846 5580 25898
rect 5632 25846 13688 25898
rect 13740 25846 13792 25898
rect 13844 25846 13896 25898
rect 13948 25846 22004 25898
rect 22056 25846 22108 25898
rect 22160 25846 22212 25898
rect 22264 25846 30320 25898
rect 30372 25846 30424 25898
rect 30476 25846 30528 25898
rect 30580 25846 34608 25898
rect 1344 25812 34608 25846
rect 2606 25730 2658 25742
rect 2606 25666 2658 25678
rect 2942 25730 2994 25742
rect 2942 25666 2994 25678
rect 3278 25730 3330 25742
rect 3278 25666 3330 25678
rect 18958 25730 19010 25742
rect 18958 25666 19010 25678
rect 12462 25618 12514 25630
rect 4946 25566 4958 25618
rect 5010 25566 5022 25618
rect 9874 25566 9886 25618
rect 9938 25566 9950 25618
rect 12462 25554 12514 25566
rect 13582 25618 13634 25630
rect 13582 25554 13634 25566
rect 14478 25618 14530 25630
rect 14478 25554 14530 25566
rect 15374 25618 15426 25630
rect 15374 25554 15426 25566
rect 19966 25618 20018 25630
rect 23090 25566 23102 25618
rect 23154 25566 23166 25618
rect 25218 25566 25230 25618
rect 25282 25566 25294 25618
rect 27346 25566 27358 25618
rect 27410 25566 27422 25618
rect 19966 25554 20018 25566
rect 12574 25506 12626 25518
rect 2594 25454 2606 25506
rect 2658 25454 2670 25506
rect 3266 25454 3278 25506
rect 3330 25454 3342 25506
rect 4610 25454 4622 25506
rect 4674 25454 4686 25506
rect 7074 25454 7086 25506
rect 7138 25454 7150 25506
rect 12574 25442 12626 25454
rect 13694 25506 13746 25518
rect 13694 25442 13746 25454
rect 14142 25506 14194 25518
rect 14142 25442 14194 25454
rect 14254 25506 14306 25518
rect 14254 25442 14306 25454
rect 14702 25506 14754 25518
rect 14702 25442 14754 25454
rect 15150 25506 15202 25518
rect 15150 25442 15202 25454
rect 15486 25506 15538 25518
rect 15486 25442 15538 25454
rect 15822 25506 15874 25518
rect 15822 25442 15874 25454
rect 16158 25506 16210 25518
rect 16158 25442 16210 25454
rect 19294 25506 19346 25518
rect 19294 25442 19346 25454
rect 19854 25506 19906 25518
rect 19854 25442 19906 25454
rect 20078 25506 20130 25518
rect 20078 25442 20130 25454
rect 20526 25506 20578 25518
rect 26350 25506 26402 25518
rect 21634 25454 21646 25506
rect 21698 25454 21710 25506
rect 22530 25454 22542 25506
rect 22594 25454 22606 25506
rect 26002 25454 26014 25506
rect 26066 25454 26078 25506
rect 20526 25442 20578 25454
rect 26350 25442 26402 25454
rect 3614 25394 3666 25406
rect 3614 25330 3666 25342
rect 4062 25394 4114 25406
rect 14926 25394 14978 25406
rect 7746 25342 7758 25394
rect 7810 25342 7822 25394
rect 4062 25330 4114 25342
rect 14926 25330 14978 25342
rect 16270 25394 16322 25406
rect 16270 25330 16322 25342
rect 19518 25394 19570 25406
rect 27022 25394 27074 25406
rect 22754 25342 22766 25394
rect 22818 25342 22830 25394
rect 26674 25342 26686 25394
rect 26738 25342 26750 25394
rect 19518 25330 19570 25342
rect 27022 25330 27074 25342
rect 12126 25282 12178 25294
rect 12126 25218 12178 25230
rect 12350 25282 12402 25294
rect 12350 25218 12402 25230
rect 13470 25282 13522 25294
rect 13470 25218 13522 25230
rect 16382 25282 16434 25294
rect 16382 25218 16434 25230
rect 16606 25282 16658 25294
rect 27246 25282 27298 25294
rect 21858 25230 21870 25282
rect 21922 25230 21934 25282
rect 16606 25218 16658 25230
rect 27246 25218 27298 25230
rect 1344 25114 34768 25148
rect 1344 25062 9530 25114
rect 9582 25062 9634 25114
rect 9686 25062 9738 25114
rect 9790 25062 17846 25114
rect 17898 25062 17950 25114
rect 18002 25062 18054 25114
rect 18106 25062 26162 25114
rect 26214 25062 26266 25114
rect 26318 25062 26370 25114
rect 26422 25062 34478 25114
rect 34530 25062 34582 25114
rect 34634 25062 34686 25114
rect 34738 25062 34768 25114
rect 1344 25028 34768 25062
rect 8878 24946 8930 24958
rect 4722 24894 4734 24946
rect 4786 24894 4798 24946
rect 6290 24894 6302 24946
rect 6354 24894 6366 24946
rect 8878 24882 8930 24894
rect 11006 24946 11058 24958
rect 11006 24882 11058 24894
rect 11118 24946 11170 24958
rect 11118 24882 11170 24894
rect 11230 24946 11282 24958
rect 11230 24882 11282 24894
rect 15150 24946 15202 24958
rect 23662 24946 23714 24958
rect 18834 24894 18846 24946
rect 18898 24894 18910 24946
rect 15150 24882 15202 24894
rect 23662 24882 23714 24894
rect 25678 24946 25730 24958
rect 25678 24882 25730 24894
rect 25790 24946 25842 24958
rect 25790 24882 25842 24894
rect 12350 24834 12402 24846
rect 4050 24782 4062 24834
rect 4114 24782 4126 24834
rect 5842 24782 5854 24834
rect 5906 24782 5918 24834
rect 6402 24782 6414 24834
rect 6466 24782 6478 24834
rect 12350 24770 12402 24782
rect 13246 24834 13298 24846
rect 13246 24770 13298 24782
rect 15710 24834 15762 24846
rect 18162 24782 18174 24834
rect 18226 24782 18238 24834
rect 28466 24782 28478 24834
rect 28530 24782 28542 24834
rect 15710 24770 15762 24782
rect 4398 24722 4450 24734
rect 4398 24658 4450 24670
rect 5070 24722 5122 24734
rect 5070 24658 5122 24670
rect 5294 24722 5346 24734
rect 12238 24722 12290 24734
rect 5618 24670 5630 24722
rect 5682 24670 5694 24722
rect 11442 24670 11454 24722
rect 11506 24670 11518 24722
rect 11666 24670 11678 24722
rect 11730 24670 11742 24722
rect 5294 24658 5346 24670
rect 12238 24658 12290 24670
rect 12574 24722 12626 24734
rect 12574 24658 12626 24670
rect 12686 24722 12738 24734
rect 12686 24658 12738 24670
rect 14590 24722 14642 24734
rect 14590 24658 14642 24670
rect 15038 24722 15090 24734
rect 15038 24658 15090 24670
rect 15262 24722 15314 24734
rect 15262 24658 15314 24670
rect 18510 24722 18562 24734
rect 20862 24722 20914 24734
rect 19058 24670 19070 24722
rect 19122 24670 19134 24722
rect 20178 24670 20190 24722
rect 20242 24670 20254 24722
rect 18510 24658 18562 24670
rect 20862 24658 20914 24670
rect 22878 24722 22930 24734
rect 22878 24658 22930 24670
rect 22990 24722 23042 24734
rect 22990 24658 23042 24670
rect 23886 24722 23938 24734
rect 23886 24658 23938 24670
rect 24334 24722 24386 24734
rect 24334 24658 24386 24670
rect 24446 24722 24498 24734
rect 24446 24658 24498 24670
rect 24558 24722 24610 24734
rect 24558 24658 24610 24670
rect 25118 24722 25170 24734
rect 25118 24658 25170 24670
rect 25566 24722 25618 24734
rect 29250 24670 29262 24722
rect 29314 24670 29326 24722
rect 25566 24658 25618 24670
rect 8990 24610 9042 24622
rect 8990 24546 9042 24558
rect 12462 24610 12514 24622
rect 12462 24546 12514 24558
rect 13358 24610 13410 24622
rect 13358 24546 13410 24558
rect 13470 24610 13522 24622
rect 13470 24546 13522 24558
rect 14142 24610 14194 24622
rect 20402 24558 20414 24610
rect 20466 24558 20478 24610
rect 26338 24558 26350 24610
rect 26402 24558 26414 24610
rect 14142 24546 14194 24558
rect 15598 24498 15650 24510
rect 15598 24434 15650 24446
rect 1344 24330 34608 24364
rect 1344 24278 5372 24330
rect 5424 24278 5476 24330
rect 5528 24278 5580 24330
rect 5632 24278 13688 24330
rect 13740 24278 13792 24330
rect 13844 24278 13896 24330
rect 13948 24278 22004 24330
rect 22056 24278 22108 24330
rect 22160 24278 22212 24330
rect 22264 24278 30320 24330
rect 30372 24278 30424 24330
rect 30476 24278 30528 24330
rect 30580 24278 34608 24330
rect 1344 24244 34608 24278
rect 12126 24162 12178 24174
rect 12126 24098 12178 24110
rect 13582 24162 13634 24174
rect 13582 24098 13634 24110
rect 11006 24050 11058 24062
rect 20302 24050 20354 24062
rect 9986 23998 9998 24050
rect 10050 23998 10062 24050
rect 15026 23998 15038 24050
rect 15090 23998 15102 24050
rect 11006 23986 11058 23998
rect 20302 23986 20354 23998
rect 26238 24050 26290 24062
rect 27010 23998 27022 24050
rect 27074 23998 27086 24050
rect 26238 23986 26290 23998
rect 10894 23938 10946 23950
rect 13470 23938 13522 23950
rect 7074 23886 7086 23938
rect 7138 23886 7150 23938
rect 11666 23886 11678 23938
rect 11730 23886 11742 23938
rect 10894 23874 10946 23886
rect 13470 23874 13522 23886
rect 14142 23938 14194 23950
rect 26126 23938 26178 23950
rect 17938 23886 17950 23938
rect 18002 23886 18014 23938
rect 19170 23886 19182 23938
rect 19234 23886 19246 23938
rect 14142 23874 14194 23886
rect 26126 23874 26178 23886
rect 5070 23826 5122 23838
rect 11118 23826 11170 23838
rect 7858 23774 7870 23826
rect 7922 23774 7934 23826
rect 5070 23762 5122 23774
rect 11118 23762 11170 23774
rect 11230 23826 11282 23838
rect 11230 23762 11282 23774
rect 12014 23826 12066 23838
rect 12014 23762 12066 23774
rect 14478 23826 14530 23838
rect 18846 23826 18898 23838
rect 17154 23774 17166 23826
rect 17218 23774 17230 23826
rect 14478 23762 14530 23774
rect 18846 23762 18898 23774
rect 26686 23826 26738 23838
rect 26686 23762 26738 23774
rect 4846 23714 4898 23726
rect 4846 23650 4898 23662
rect 4958 23714 5010 23726
rect 4958 23650 5010 23662
rect 12126 23714 12178 23726
rect 12126 23650 12178 23662
rect 13022 23714 13074 23726
rect 13022 23650 13074 23662
rect 13694 23714 13746 23726
rect 13694 23650 13746 23662
rect 13918 23714 13970 23726
rect 13918 23650 13970 23662
rect 14590 23714 14642 23726
rect 14590 23650 14642 23662
rect 14814 23714 14866 23726
rect 14814 23650 14866 23662
rect 18510 23714 18562 23726
rect 18510 23650 18562 23662
rect 18958 23714 19010 23726
rect 19854 23714 19906 23726
rect 19506 23662 19518 23714
rect 19570 23662 19582 23714
rect 18958 23650 19010 23662
rect 19854 23650 19906 23662
rect 25902 23714 25954 23726
rect 25902 23650 25954 23662
rect 26350 23714 26402 23726
rect 26350 23650 26402 23662
rect 26910 23714 26962 23726
rect 26910 23650 26962 23662
rect 1344 23546 34768 23580
rect 1344 23494 9530 23546
rect 9582 23494 9634 23546
rect 9686 23494 9738 23546
rect 9790 23494 17846 23546
rect 17898 23494 17950 23546
rect 18002 23494 18054 23546
rect 18106 23494 26162 23546
rect 26214 23494 26266 23546
rect 26318 23494 26370 23546
rect 26422 23494 34478 23546
rect 34530 23494 34582 23546
rect 34634 23494 34686 23546
rect 34738 23494 34768 23546
rect 1344 23460 34768 23494
rect 8430 23378 8482 23390
rect 5842 23326 5854 23378
rect 5906 23326 5918 23378
rect 8430 23314 8482 23326
rect 8878 23378 8930 23390
rect 8878 23314 8930 23326
rect 9998 23378 10050 23390
rect 9998 23314 10050 23326
rect 11006 23378 11058 23390
rect 11006 23314 11058 23326
rect 12910 23378 12962 23390
rect 15934 23378 15986 23390
rect 18846 23378 18898 23390
rect 14130 23326 14142 23378
rect 14194 23326 14206 23378
rect 17378 23326 17390 23378
rect 17442 23326 17454 23378
rect 12910 23314 12962 23326
rect 15934 23314 15986 23326
rect 18846 23314 18898 23326
rect 19070 23378 19122 23390
rect 25778 23326 25790 23378
rect 25842 23326 25854 23378
rect 19070 23314 19122 23326
rect 9886 23266 9938 23278
rect 9886 23202 9938 23214
rect 10222 23266 10274 23278
rect 10222 23202 10274 23214
rect 10894 23266 10946 23278
rect 10894 23202 10946 23214
rect 11790 23266 11842 23278
rect 11790 23202 11842 23214
rect 12686 23266 12738 23278
rect 12686 23202 12738 23214
rect 13694 23266 13746 23278
rect 13694 23202 13746 23214
rect 13806 23266 13858 23278
rect 15822 23266 15874 23278
rect 14802 23214 14814 23266
rect 14866 23214 14878 23266
rect 13806 23202 13858 23214
rect 15822 23202 15874 23214
rect 18622 23266 18674 23278
rect 22766 23266 22818 23278
rect 20290 23214 20302 23266
rect 20354 23214 20366 23266
rect 18622 23202 18674 23214
rect 22766 23202 22818 23214
rect 23102 23266 23154 23278
rect 24658 23214 24670 23266
rect 24722 23214 24734 23266
rect 29138 23214 29150 23266
rect 29202 23214 29214 23266
rect 23102 23202 23154 23214
rect 5518 23154 5570 23166
rect 6414 23154 6466 23166
rect 2034 23102 2046 23154
rect 2098 23102 2110 23154
rect 6178 23102 6190 23154
rect 6242 23102 6254 23154
rect 5518 23090 5570 23102
rect 6414 23090 6466 23102
rect 6638 23154 6690 23166
rect 6638 23090 6690 23102
rect 10334 23154 10386 23166
rect 11342 23154 11394 23166
rect 10658 23102 10670 23154
rect 10722 23102 10734 23154
rect 10334 23090 10386 23102
rect 11342 23090 11394 23102
rect 11678 23154 11730 23166
rect 13470 23154 13522 23166
rect 12114 23102 12126 23154
rect 12178 23102 12190 23154
rect 12450 23102 12462 23154
rect 12514 23102 12526 23154
rect 11678 23090 11730 23102
rect 13470 23090 13522 23102
rect 14478 23154 14530 23166
rect 15374 23154 15426 23166
rect 15026 23102 15038 23154
rect 15090 23102 15102 23154
rect 14478 23090 14530 23102
rect 15374 23090 15426 23102
rect 16046 23154 16098 23166
rect 19182 23154 19234 23166
rect 25230 23154 25282 23166
rect 26462 23154 26514 23166
rect 18386 23102 18398 23154
rect 18450 23102 18462 23154
rect 19506 23102 19518 23154
rect 19570 23102 19582 23154
rect 24434 23102 24446 23154
rect 24498 23102 24510 23154
rect 26114 23102 26126 23154
rect 26178 23102 26190 23154
rect 16046 23090 16098 23102
rect 19182 23090 19234 23102
rect 25230 23090 25282 23102
rect 26462 23090 26514 23102
rect 26686 23154 26738 23166
rect 29810 23102 29822 23154
rect 29874 23102 29886 23154
rect 26686 23090 26738 23102
rect 5294 23042 5346 23054
rect 2818 22990 2830 23042
rect 2882 22990 2894 23042
rect 4946 22990 4958 23042
rect 5010 22990 5022 23042
rect 5294 22978 5346 22990
rect 6750 23042 6802 23054
rect 6750 22978 6802 22990
rect 8542 23042 8594 23054
rect 8542 22978 8594 22990
rect 8990 23042 9042 23054
rect 17726 23042 17778 23054
rect 12562 22990 12574 23042
rect 12626 22990 12638 23042
rect 8990 22978 9042 22990
rect 17726 22978 17778 22990
rect 17950 23042 18002 23054
rect 22418 22990 22430 23042
rect 22482 22990 22494 23042
rect 27010 22990 27022 23042
rect 27074 22990 27086 23042
rect 17950 22978 18002 22990
rect 11454 22930 11506 22942
rect 11454 22866 11506 22878
rect 25454 22930 25506 22942
rect 25454 22866 25506 22878
rect 1344 22762 34608 22796
rect 1344 22710 5372 22762
rect 5424 22710 5476 22762
rect 5528 22710 5580 22762
rect 5632 22710 13688 22762
rect 13740 22710 13792 22762
rect 13844 22710 13896 22762
rect 13948 22710 22004 22762
rect 22056 22710 22108 22762
rect 22160 22710 22212 22762
rect 22264 22710 30320 22762
rect 30372 22710 30424 22762
rect 30476 22710 30528 22762
rect 30580 22710 34608 22762
rect 1344 22676 34608 22710
rect 5742 22594 5794 22606
rect 5742 22530 5794 22542
rect 5966 22594 6018 22606
rect 5966 22530 6018 22542
rect 19294 22594 19346 22606
rect 19294 22530 19346 22542
rect 19406 22482 19458 22494
rect 25342 22482 25394 22494
rect 4610 22430 4622 22482
rect 4674 22430 4686 22482
rect 7858 22430 7870 22482
rect 7922 22430 7934 22482
rect 24210 22430 24222 22482
rect 24274 22430 24286 22482
rect 19406 22418 19458 22430
rect 25342 22418 25394 22430
rect 6078 22370 6130 22382
rect 20302 22370 20354 22382
rect 25230 22370 25282 22382
rect 26910 22370 26962 22382
rect 1810 22318 1822 22370
rect 1874 22318 1886 22370
rect 12898 22318 12910 22370
rect 12962 22318 12974 22370
rect 15026 22318 15038 22370
rect 15090 22318 15102 22370
rect 19618 22318 19630 22370
rect 19682 22318 19694 22370
rect 19954 22318 19966 22370
rect 20018 22318 20030 22370
rect 21298 22318 21310 22370
rect 21362 22318 21374 22370
rect 26114 22318 26126 22370
rect 26178 22318 26190 22370
rect 26338 22318 26350 22370
rect 26402 22318 26414 22370
rect 6078 22306 6130 22318
rect 20302 22306 20354 22318
rect 25230 22306 25282 22318
rect 26910 22306 26962 22318
rect 5630 22258 5682 22270
rect 20638 22258 20690 22270
rect 2482 22206 2494 22258
rect 2546 22206 2558 22258
rect 18610 22206 18622 22258
rect 18674 22206 18686 22258
rect 20514 22206 20526 22258
rect 20578 22206 20590 22258
rect 5630 22194 5682 22206
rect 20638 22194 20690 22206
rect 20750 22258 20802 22270
rect 27022 22258 27074 22270
rect 22082 22206 22094 22258
rect 22146 22206 22158 22258
rect 20750 22194 20802 22206
rect 27022 22194 27074 22206
rect 27470 22258 27522 22270
rect 27470 22194 27522 22206
rect 25454 22146 25506 22158
rect 25454 22082 25506 22094
rect 25678 22146 25730 22158
rect 25678 22082 25730 22094
rect 26574 22146 26626 22158
rect 26574 22082 26626 22094
rect 26686 22146 26738 22158
rect 26686 22082 26738 22094
rect 27246 22146 27298 22158
rect 27246 22082 27298 22094
rect 27582 22146 27634 22158
rect 27582 22082 27634 22094
rect 1344 21978 34768 22012
rect 1344 21926 9530 21978
rect 9582 21926 9634 21978
rect 9686 21926 9738 21978
rect 9790 21926 17846 21978
rect 17898 21926 17950 21978
rect 18002 21926 18054 21978
rect 18106 21926 26162 21978
rect 26214 21926 26266 21978
rect 26318 21926 26370 21978
rect 26422 21926 34478 21978
rect 34530 21926 34582 21978
rect 34634 21926 34686 21978
rect 34738 21926 34768 21978
rect 1344 21892 34768 21926
rect 3614 21810 3666 21822
rect 3614 21746 3666 21758
rect 5518 21810 5570 21822
rect 5518 21746 5570 21758
rect 12686 21810 12738 21822
rect 12686 21746 12738 21758
rect 13582 21810 13634 21822
rect 13582 21746 13634 21758
rect 13694 21810 13746 21822
rect 13694 21746 13746 21758
rect 13806 21810 13858 21822
rect 13806 21746 13858 21758
rect 14702 21810 14754 21822
rect 14702 21746 14754 21758
rect 14926 21810 14978 21822
rect 14926 21746 14978 21758
rect 15710 21810 15762 21822
rect 15710 21746 15762 21758
rect 16830 21810 16882 21822
rect 19406 21810 19458 21822
rect 17938 21758 17950 21810
rect 18002 21758 18014 21810
rect 16830 21746 16882 21758
rect 19406 21746 19458 21758
rect 19966 21810 20018 21822
rect 19966 21746 20018 21758
rect 21086 21810 21138 21822
rect 21086 21746 21138 21758
rect 23662 21810 23714 21822
rect 23662 21746 23714 21758
rect 3950 21698 4002 21710
rect 3950 21634 4002 21646
rect 4622 21698 4674 21710
rect 4622 21634 4674 21646
rect 5406 21698 5458 21710
rect 5406 21634 5458 21646
rect 10782 21698 10834 21710
rect 10782 21634 10834 21646
rect 11342 21698 11394 21710
rect 13470 21698 13522 21710
rect 12338 21646 12350 21698
rect 12402 21646 12414 21698
rect 11342 21634 11394 21646
rect 13470 21634 13522 21646
rect 14814 21698 14866 21710
rect 19294 21698 19346 21710
rect 16482 21646 16494 21698
rect 16546 21646 16558 21698
rect 14814 21634 14866 21646
rect 19294 21634 19346 21646
rect 20638 21698 20690 21710
rect 20638 21634 20690 21646
rect 20862 21698 20914 21710
rect 20862 21634 20914 21646
rect 21758 21698 21810 21710
rect 21758 21634 21810 21646
rect 22542 21698 22594 21710
rect 26126 21698 26178 21710
rect 24210 21646 24222 21698
rect 24274 21646 24286 21698
rect 22542 21634 22594 21646
rect 26126 21634 26178 21646
rect 26238 21698 26290 21710
rect 26238 21634 26290 21646
rect 3390 21586 3442 21598
rect 3390 21522 3442 21534
rect 3614 21586 3666 21598
rect 3614 21522 3666 21534
rect 4398 21586 4450 21598
rect 4398 21522 4450 21534
rect 4510 21586 4562 21598
rect 4510 21522 4562 21534
rect 5742 21586 5794 21598
rect 5742 21522 5794 21534
rect 10670 21586 10722 21598
rect 11902 21586 11954 21598
rect 15150 21586 15202 21598
rect 20302 21586 20354 21598
rect 11554 21534 11566 21586
rect 11618 21534 11630 21586
rect 13010 21534 13022 21586
rect 13074 21534 13086 21586
rect 14130 21534 14142 21586
rect 14194 21534 14206 21586
rect 14466 21534 14478 21586
rect 14530 21534 14542 21586
rect 15474 21534 15486 21586
rect 15538 21534 15550 21586
rect 18162 21534 18174 21586
rect 18226 21534 18238 21586
rect 10670 21522 10722 21534
rect 11902 21522 11954 21534
rect 15150 21522 15202 21534
rect 20302 21522 20354 21534
rect 21310 21586 21362 21598
rect 21310 21522 21362 21534
rect 21870 21586 21922 21598
rect 21870 21522 21922 21534
rect 22094 21586 22146 21598
rect 22094 21522 22146 21534
rect 22430 21586 22482 21598
rect 24446 21586 24498 21598
rect 24098 21534 24110 21586
rect 24162 21534 24174 21586
rect 29474 21534 29486 21586
rect 29538 21534 29550 21586
rect 22430 21522 22482 21534
rect 24446 21522 24498 21534
rect 11678 21474 11730 21486
rect 5058 21422 5070 21474
rect 5122 21422 5134 21474
rect 11678 21410 11730 21422
rect 15374 21474 15426 21486
rect 15374 21410 15426 21422
rect 17614 21474 17666 21486
rect 17614 21410 17666 21422
rect 18958 21474 19010 21486
rect 24670 21474 24722 21486
rect 20738 21422 20750 21474
rect 20802 21422 20814 21474
rect 26562 21422 26574 21474
rect 26626 21422 26638 21474
rect 28690 21422 28702 21474
rect 28754 21422 28766 21474
rect 18958 21410 19010 21422
rect 24670 21410 24722 21422
rect 10782 21362 10834 21374
rect 10782 21298 10834 21310
rect 19406 21362 19458 21374
rect 19406 21298 19458 21310
rect 26126 21362 26178 21374
rect 26126 21298 26178 21310
rect 1344 21194 34608 21228
rect 1344 21142 5372 21194
rect 5424 21142 5476 21194
rect 5528 21142 5580 21194
rect 5632 21142 13688 21194
rect 13740 21142 13792 21194
rect 13844 21142 13896 21194
rect 13948 21142 22004 21194
rect 22056 21142 22108 21194
rect 22160 21142 22212 21194
rect 22264 21142 30320 21194
rect 30372 21142 30424 21194
rect 30476 21142 30528 21194
rect 30580 21142 34608 21194
rect 1344 21108 34608 21142
rect 2606 21026 2658 21038
rect 2606 20962 2658 20974
rect 11454 21026 11506 21038
rect 11454 20962 11506 20974
rect 12686 21026 12738 21038
rect 12686 20962 12738 20974
rect 15822 20914 15874 20926
rect 28030 20914 28082 20926
rect 10994 20862 11006 20914
rect 11058 20862 11070 20914
rect 25890 20862 25902 20914
rect 25954 20862 25966 20914
rect 15822 20850 15874 20862
rect 28030 20850 28082 20862
rect 3278 20802 3330 20814
rect 3278 20738 3330 20750
rect 4958 20802 5010 20814
rect 12574 20802 12626 20814
rect 5618 20750 5630 20802
rect 5682 20750 5694 20802
rect 7634 20750 7646 20802
rect 7698 20750 7710 20802
rect 4958 20738 5010 20750
rect 12574 20738 12626 20750
rect 13806 20802 13858 20814
rect 16046 20802 16098 20814
rect 27582 20802 27634 20814
rect 14130 20750 14142 20802
rect 14194 20750 14206 20802
rect 16930 20750 16942 20802
rect 16994 20750 17006 20802
rect 23090 20750 23102 20802
rect 23154 20750 23166 20802
rect 26450 20750 26462 20802
rect 26514 20750 26526 20802
rect 26674 20750 26686 20802
rect 26738 20750 26750 20802
rect 13806 20738 13858 20750
rect 16046 20738 16098 20750
rect 27582 20738 27634 20750
rect 27806 20802 27858 20814
rect 27806 20738 27858 20750
rect 3950 20690 4002 20702
rect 8206 20690 8258 20702
rect 5730 20638 5742 20690
rect 5794 20638 5806 20690
rect 3950 20626 4002 20638
rect 8206 20626 8258 20638
rect 10558 20690 10610 20702
rect 11342 20690 11394 20702
rect 10770 20638 10782 20690
rect 10834 20638 10846 20690
rect 10558 20626 10610 20638
rect 11342 20626 11394 20638
rect 11454 20690 11506 20702
rect 11454 20626 11506 20638
rect 12686 20690 12738 20702
rect 12686 20626 12738 20638
rect 13470 20690 13522 20702
rect 13470 20626 13522 20638
rect 14366 20690 14418 20702
rect 14366 20626 14418 20638
rect 16718 20690 16770 20702
rect 16718 20626 16770 20638
rect 17390 20690 17442 20702
rect 17390 20626 17442 20638
rect 17726 20690 17778 20702
rect 26238 20690 26290 20702
rect 23762 20638 23774 20690
rect 23826 20638 23838 20690
rect 17726 20626 17778 20638
rect 26238 20626 26290 20638
rect 28142 20690 28194 20702
rect 28142 20626 28194 20638
rect 2382 20578 2434 20590
rect 2382 20514 2434 20526
rect 2494 20578 2546 20590
rect 3614 20578 3666 20590
rect 2930 20526 2942 20578
rect 2994 20526 3006 20578
rect 2494 20514 2546 20526
rect 3614 20514 3666 20526
rect 4286 20578 4338 20590
rect 4286 20514 4338 20526
rect 4398 20578 4450 20590
rect 4398 20514 4450 20526
rect 4510 20578 4562 20590
rect 10222 20578 10274 20590
rect 7746 20526 7758 20578
rect 7810 20526 7822 20578
rect 4510 20514 4562 20526
rect 10222 20514 10274 20526
rect 10446 20578 10498 20590
rect 10446 20514 10498 20526
rect 13582 20578 13634 20590
rect 18398 20578 18450 20590
rect 16370 20526 16382 20578
rect 16434 20526 16446 20578
rect 18050 20526 18062 20578
rect 18114 20526 18126 20578
rect 13582 20514 13634 20526
rect 18398 20514 18450 20526
rect 1344 20410 34768 20444
rect 1344 20358 9530 20410
rect 9582 20358 9634 20410
rect 9686 20358 9738 20410
rect 9790 20358 17846 20410
rect 17898 20358 17950 20410
rect 18002 20358 18054 20410
rect 18106 20358 26162 20410
rect 26214 20358 26266 20410
rect 26318 20358 26370 20410
rect 26422 20358 34478 20410
rect 34530 20358 34582 20410
rect 34634 20358 34686 20410
rect 34738 20358 34768 20410
rect 1344 20324 34768 20358
rect 5070 20130 5122 20142
rect 5070 20066 5122 20078
rect 8206 20130 8258 20142
rect 8206 20066 8258 20078
rect 8878 20130 8930 20142
rect 8878 20066 8930 20078
rect 12014 20130 12066 20142
rect 12014 20066 12066 20078
rect 12574 20130 12626 20142
rect 14242 20078 14254 20130
rect 14306 20078 14318 20130
rect 14914 20078 14926 20130
rect 14978 20078 14990 20130
rect 15250 20078 15262 20130
rect 15314 20078 15326 20130
rect 16818 20078 16830 20130
rect 16882 20078 16894 20130
rect 12574 20066 12626 20078
rect 5294 20018 5346 20030
rect 1810 19966 1822 20018
rect 1874 19966 1886 20018
rect 5294 19954 5346 19966
rect 5518 20018 5570 20030
rect 10558 20018 10610 20030
rect 11454 20018 11506 20030
rect 7522 19966 7534 20018
rect 7586 19966 7598 20018
rect 9986 19966 9998 20018
rect 10050 19966 10062 20018
rect 10770 19966 10782 20018
rect 10834 19966 10846 20018
rect 5518 19954 5570 19966
rect 10558 19954 10610 19966
rect 11454 19954 11506 19966
rect 11902 20018 11954 20030
rect 11902 19954 11954 19966
rect 12126 20018 12178 20030
rect 12126 19954 12178 19966
rect 12686 20018 12738 20030
rect 17502 20018 17554 20030
rect 14018 19966 14030 20018
rect 14082 19966 14094 20018
rect 14690 19966 14702 20018
rect 14754 19966 14766 20018
rect 15474 19966 15486 20018
rect 15538 19966 15550 20018
rect 16594 19966 16606 20018
rect 16658 19966 16670 20018
rect 12686 19954 12738 19966
rect 17502 19954 17554 19966
rect 17950 20018 18002 20030
rect 17950 19954 18002 19966
rect 18174 20018 18226 20030
rect 18174 19954 18226 19966
rect 18510 20018 18562 20030
rect 18510 19954 18562 19966
rect 18846 20018 18898 20030
rect 18846 19954 18898 19966
rect 19070 20018 19122 20030
rect 19070 19954 19122 19966
rect 20302 20018 20354 20030
rect 20738 19966 20750 20018
rect 20802 19966 20814 20018
rect 21634 19966 21646 20018
rect 21698 19966 21710 20018
rect 25666 19966 25678 20018
rect 25730 19966 25742 20018
rect 20302 19954 20354 19966
rect 5182 19906 5234 19918
rect 16046 19906 16098 19918
rect 2594 19854 2606 19906
rect 2658 19854 2670 19906
rect 4722 19854 4734 19906
rect 4786 19854 4798 19906
rect 7410 19854 7422 19906
rect 7474 19854 7486 19906
rect 9650 19854 9662 19906
rect 9714 19854 9726 19906
rect 5182 19842 5234 19854
rect 16046 19842 16098 19854
rect 18062 19906 18114 19918
rect 18062 19842 18114 19854
rect 18958 19906 19010 19918
rect 18958 19842 19010 19854
rect 21198 19906 21250 19918
rect 22306 19854 22318 19906
rect 22370 19854 22382 19906
rect 24434 19854 24446 19906
rect 24498 19854 24510 19906
rect 26450 19854 26462 19906
rect 26514 19854 26526 19906
rect 28578 19854 28590 19906
rect 28642 19854 28654 19906
rect 21198 19842 21250 19854
rect 8654 19794 8706 19806
rect 8654 19730 8706 19742
rect 8990 19794 9042 19806
rect 12574 19794 12626 19806
rect 10210 19742 10222 19794
rect 10274 19742 10286 19794
rect 8990 19730 9042 19742
rect 12574 19730 12626 19742
rect 1344 19626 34608 19660
rect 1344 19574 5372 19626
rect 5424 19574 5476 19626
rect 5528 19574 5580 19626
rect 5632 19574 13688 19626
rect 13740 19574 13792 19626
rect 13844 19574 13896 19626
rect 13948 19574 22004 19626
rect 22056 19574 22108 19626
rect 22160 19574 22212 19626
rect 22264 19574 30320 19626
rect 30372 19574 30424 19626
rect 30476 19574 30528 19626
rect 30580 19574 34608 19626
rect 1344 19540 34608 19574
rect 9774 19458 9826 19470
rect 9774 19394 9826 19406
rect 12686 19458 12738 19470
rect 12686 19394 12738 19406
rect 17614 19458 17666 19470
rect 17614 19394 17666 19406
rect 21870 19458 21922 19470
rect 21870 19394 21922 19406
rect 22206 19458 22258 19470
rect 22206 19394 22258 19406
rect 7982 19346 8034 19358
rect 2482 19294 2494 19346
rect 2546 19294 2558 19346
rect 4610 19294 4622 19346
rect 4674 19294 4686 19346
rect 7982 19282 8034 19294
rect 8990 19346 9042 19358
rect 8990 19282 9042 19294
rect 9438 19346 9490 19358
rect 9438 19282 9490 19294
rect 11342 19346 11394 19358
rect 11342 19282 11394 19294
rect 12238 19346 12290 19358
rect 12238 19282 12290 19294
rect 17390 19346 17442 19358
rect 17390 19282 17442 19294
rect 18398 19346 18450 19358
rect 18398 19282 18450 19294
rect 22878 19346 22930 19358
rect 26002 19294 26014 19346
rect 26066 19294 26078 19346
rect 22878 19282 22930 19294
rect 7086 19234 7138 19246
rect 8654 19234 8706 19246
rect 1810 19182 1822 19234
rect 1874 19182 1886 19234
rect 7298 19182 7310 19234
rect 7362 19182 7374 19234
rect 7086 19170 7138 19182
rect 8654 19170 8706 19182
rect 8878 19234 8930 19246
rect 8878 19170 8930 19182
rect 9214 19234 9266 19246
rect 9214 19170 9266 19182
rect 10782 19234 10834 19246
rect 27234 19182 27246 19234
rect 27298 19182 27310 19234
rect 10782 19170 10834 19182
rect 9998 19122 10050 19134
rect 9998 19058 10050 19070
rect 10558 19122 10610 19134
rect 10558 19058 10610 19070
rect 11230 19122 11282 19134
rect 11230 19058 11282 19070
rect 12798 19122 12850 19134
rect 12798 19058 12850 19070
rect 11006 19010 11058 19022
rect 11006 18946 11058 18958
rect 11902 19010 11954 19022
rect 11902 18946 11954 18958
rect 12126 19010 12178 19022
rect 12126 18946 12178 18958
rect 12350 19010 12402 19022
rect 12350 18946 12402 18958
rect 14926 19010 14978 19022
rect 22094 19010 22146 19022
rect 17938 18958 17950 19010
rect 18002 18958 18014 19010
rect 14926 18946 14978 18958
rect 22094 18946 22146 18958
rect 1344 18842 34768 18876
rect 1344 18790 9530 18842
rect 9582 18790 9634 18842
rect 9686 18790 9738 18842
rect 9790 18790 17846 18842
rect 17898 18790 17950 18842
rect 18002 18790 18054 18842
rect 18106 18790 26162 18842
rect 26214 18790 26266 18842
rect 26318 18790 26370 18842
rect 26422 18790 34478 18842
rect 34530 18790 34582 18842
rect 34634 18790 34686 18842
rect 34738 18790 34768 18842
rect 1344 18756 34768 18790
rect 8206 18674 8258 18686
rect 7410 18622 7422 18674
rect 7474 18622 7486 18674
rect 8206 18610 8258 18622
rect 10782 18674 10834 18686
rect 22654 18674 22706 18686
rect 12674 18622 12686 18674
rect 12738 18622 12750 18674
rect 10782 18610 10834 18622
rect 22654 18610 22706 18622
rect 23326 18674 23378 18686
rect 23326 18610 23378 18622
rect 7982 18562 8034 18574
rect 5842 18510 5854 18562
rect 5906 18510 5918 18562
rect 6514 18510 6526 18562
rect 6578 18510 6590 18562
rect 7982 18498 8034 18510
rect 8766 18562 8818 18574
rect 8766 18498 8818 18510
rect 8878 18562 8930 18574
rect 8878 18498 8930 18510
rect 9550 18562 9602 18574
rect 9550 18498 9602 18510
rect 9662 18562 9714 18574
rect 9662 18498 9714 18510
rect 11454 18562 11506 18574
rect 26686 18562 26738 18574
rect 19506 18510 19518 18562
rect 19570 18510 19582 18562
rect 22978 18510 22990 18562
rect 23042 18510 23054 18562
rect 11454 18498 11506 18510
rect 26686 18498 26738 18510
rect 7870 18450 7922 18462
rect 5618 18398 5630 18450
rect 5682 18398 5694 18450
rect 6290 18398 6302 18450
rect 6354 18398 6366 18450
rect 7870 18386 7922 18398
rect 8318 18450 8370 18462
rect 8318 18386 8370 18398
rect 9886 18450 9938 18462
rect 9886 18386 9938 18398
rect 10558 18450 10610 18462
rect 10558 18386 10610 18398
rect 10670 18450 10722 18462
rect 10670 18386 10722 18398
rect 11342 18450 11394 18462
rect 11342 18386 11394 18398
rect 11678 18450 11730 18462
rect 11678 18386 11730 18398
rect 11790 18450 11842 18462
rect 17390 18450 17442 18462
rect 14018 18398 14030 18450
rect 14082 18398 14094 18450
rect 11790 18386 11842 18398
rect 17390 18386 17442 18398
rect 17614 18450 17666 18462
rect 17614 18386 17666 18398
rect 18062 18450 18114 18462
rect 23886 18450 23938 18462
rect 18722 18398 18734 18450
rect 18786 18398 18798 18450
rect 23650 18398 23662 18450
rect 23714 18398 23726 18450
rect 18062 18386 18114 18398
rect 23886 18386 23938 18398
rect 23998 18450 24050 18462
rect 23998 18386 24050 18398
rect 26238 18450 26290 18462
rect 27234 18398 27246 18450
rect 27298 18398 27310 18450
rect 26238 18386 26290 18398
rect 6862 18338 6914 18350
rect 6862 18274 6914 18286
rect 7086 18338 7138 18350
rect 7086 18274 7138 18286
rect 8094 18338 8146 18350
rect 8094 18274 8146 18286
rect 10334 18338 10386 18350
rect 10334 18274 10386 18286
rect 12126 18338 12178 18350
rect 12126 18274 12178 18286
rect 12350 18338 12402 18350
rect 17502 18338 17554 18350
rect 14690 18286 14702 18338
rect 14754 18286 14766 18338
rect 16818 18286 16830 18338
rect 16882 18286 16894 18338
rect 21634 18286 21646 18338
rect 21698 18286 21710 18338
rect 26562 18286 26574 18338
rect 26626 18286 26638 18338
rect 29250 18286 29262 18338
rect 29314 18286 29326 18338
rect 12350 18274 12402 18286
rect 17502 18274 17554 18286
rect 8878 18226 8930 18238
rect 8878 18162 8930 18174
rect 10110 18226 10162 18238
rect 10110 18162 10162 18174
rect 26910 18226 26962 18238
rect 26910 18162 26962 18174
rect 1344 18058 34608 18092
rect 1344 18006 5372 18058
rect 5424 18006 5476 18058
rect 5528 18006 5580 18058
rect 5632 18006 13688 18058
rect 13740 18006 13792 18058
rect 13844 18006 13896 18058
rect 13948 18006 22004 18058
rect 22056 18006 22108 18058
rect 22160 18006 22212 18058
rect 22264 18006 30320 18058
rect 30372 18006 30424 18058
rect 30476 18006 30528 18058
rect 30580 18006 34608 18058
rect 1344 17972 34608 18006
rect 6414 17890 6466 17902
rect 9550 17890 9602 17902
rect 6738 17838 6750 17890
rect 6802 17838 6814 17890
rect 6414 17826 6466 17838
rect 9550 17826 9602 17838
rect 9886 17890 9938 17902
rect 9886 17826 9938 17838
rect 26238 17890 26290 17902
rect 28466 17838 28478 17890
rect 28530 17838 28542 17890
rect 26238 17826 26290 17838
rect 8430 17778 8482 17790
rect 16046 17778 16098 17790
rect 27918 17778 27970 17790
rect 4610 17726 4622 17778
rect 4674 17726 4686 17778
rect 10434 17726 10446 17778
rect 10498 17726 10510 17778
rect 25890 17726 25902 17778
rect 25954 17726 25966 17778
rect 29138 17726 29150 17778
rect 29202 17726 29214 17778
rect 8430 17714 8482 17726
rect 16046 17714 16098 17726
rect 27918 17714 27970 17726
rect 6190 17666 6242 17678
rect 1810 17614 1822 17666
rect 1874 17614 1886 17666
rect 6190 17602 6242 17614
rect 7086 17666 7138 17678
rect 7086 17602 7138 17614
rect 7646 17666 7698 17678
rect 10894 17666 10946 17678
rect 7858 17614 7870 17666
rect 7922 17614 7934 17666
rect 9090 17614 9102 17666
rect 9154 17614 9166 17666
rect 10210 17614 10222 17666
rect 10274 17614 10286 17666
rect 7646 17602 7698 17614
rect 10894 17602 10946 17614
rect 11230 17666 11282 17678
rect 11230 17602 11282 17614
rect 15822 17666 15874 17678
rect 15822 17602 15874 17614
rect 16158 17666 16210 17678
rect 16158 17602 16210 17614
rect 16494 17666 16546 17678
rect 27470 17666 27522 17678
rect 27234 17614 27246 17666
rect 27298 17614 27310 17666
rect 16494 17602 16546 17614
rect 27470 17602 27522 17614
rect 28142 17666 28194 17678
rect 31938 17614 31950 17666
rect 32002 17614 32014 17666
rect 28142 17602 28194 17614
rect 10670 17554 10722 17566
rect 18958 17554 19010 17566
rect 2482 17502 2494 17554
rect 2546 17502 2558 17554
rect 17378 17502 17390 17554
rect 17442 17502 17454 17554
rect 18050 17502 18062 17554
rect 18114 17502 18126 17554
rect 10670 17490 10722 17502
rect 18958 17490 19010 17502
rect 26014 17554 26066 17566
rect 26014 17490 26066 17502
rect 26574 17554 26626 17566
rect 31266 17502 31278 17554
rect 31330 17502 31342 17554
rect 26574 17490 26626 17502
rect 5070 17442 5122 17454
rect 5070 17378 5122 17390
rect 7198 17442 7250 17454
rect 7198 17378 7250 17390
rect 7422 17442 7474 17454
rect 9774 17442 9826 17454
rect 8866 17390 8878 17442
rect 8930 17390 8942 17442
rect 7422 17378 7474 17390
rect 9774 17378 9826 17390
rect 10446 17442 10498 17454
rect 10446 17378 10498 17390
rect 11118 17442 11170 17454
rect 11118 17378 11170 17390
rect 17726 17442 17778 17454
rect 17726 17378 17778 17390
rect 18398 17442 18450 17454
rect 18398 17378 18450 17390
rect 19070 17442 19122 17454
rect 19070 17378 19122 17390
rect 1344 17274 34768 17308
rect 1344 17222 9530 17274
rect 9582 17222 9634 17274
rect 9686 17222 9738 17274
rect 9790 17222 17846 17274
rect 17898 17222 17950 17274
rect 18002 17222 18054 17274
rect 18106 17222 26162 17274
rect 26214 17222 26266 17274
rect 26318 17222 26370 17274
rect 26422 17222 34478 17274
rect 34530 17222 34582 17274
rect 34634 17222 34686 17274
rect 34738 17222 34768 17274
rect 1344 17188 34768 17222
rect 7422 17106 7474 17118
rect 7074 17054 7086 17106
rect 7138 17054 7150 17106
rect 7422 17042 7474 17054
rect 8206 17106 8258 17118
rect 8206 17042 8258 17054
rect 8430 17106 8482 17118
rect 14366 17106 14418 17118
rect 8642 17054 8654 17106
rect 8706 17054 8718 17106
rect 9874 17054 9886 17106
rect 9938 17054 9950 17106
rect 8430 17042 8482 17054
rect 14366 17042 14418 17054
rect 15822 17106 15874 17118
rect 15822 17042 15874 17054
rect 17390 17106 17442 17118
rect 17390 17042 17442 17054
rect 28926 17106 28978 17118
rect 28926 17042 28978 17054
rect 33070 17106 33122 17118
rect 33070 17042 33122 17054
rect 8094 16994 8146 17006
rect 8094 16930 8146 16942
rect 14142 16994 14194 17006
rect 14142 16930 14194 16942
rect 15262 16994 15314 17006
rect 15262 16930 15314 16942
rect 15934 16994 15986 17006
rect 15934 16930 15986 16942
rect 16718 16994 16770 17006
rect 16718 16930 16770 16942
rect 17614 16994 17666 17006
rect 17614 16930 17666 16942
rect 17726 16994 17778 17006
rect 29038 16994 29090 17006
rect 17938 16942 17950 16994
rect 18002 16942 18014 16994
rect 20626 16942 20638 16994
rect 20690 16942 20702 16994
rect 17726 16930 17778 16942
rect 29038 16930 29090 16942
rect 6750 16882 6802 16894
rect 3266 16830 3278 16882
rect 3330 16830 3342 16882
rect 3938 16830 3950 16882
rect 4002 16830 4014 16882
rect 6750 16818 6802 16830
rect 7534 16882 7586 16894
rect 9550 16882 9602 16894
rect 8866 16830 8878 16882
rect 8930 16830 8942 16882
rect 7534 16818 7586 16830
rect 9550 16818 9602 16830
rect 12126 16882 12178 16894
rect 12126 16818 12178 16830
rect 12238 16882 12290 16894
rect 15374 16882 15426 16894
rect 13570 16830 13582 16882
rect 13634 16830 13646 16882
rect 13906 16830 13918 16882
rect 13970 16830 13982 16882
rect 12238 16818 12290 16830
rect 15374 16818 15426 16830
rect 15710 16882 15762 16894
rect 15710 16818 15762 16830
rect 16382 16882 16434 16894
rect 16382 16818 16434 16830
rect 16830 16882 16882 16894
rect 28590 16882 28642 16894
rect 21410 16830 21422 16882
rect 21474 16830 21486 16882
rect 24546 16830 24558 16882
rect 24610 16830 24622 16882
rect 25330 16830 25342 16882
rect 25394 16830 25406 16882
rect 16830 16818 16882 16830
rect 28590 16818 28642 16830
rect 29262 16882 29314 16894
rect 33294 16882 33346 16894
rect 29586 16830 29598 16882
rect 29650 16830 29662 16882
rect 33618 16830 33630 16882
rect 33682 16830 33694 16882
rect 29262 16818 29314 16830
rect 33294 16818 33346 16830
rect 12798 16770 12850 16782
rect 33182 16770 33234 16782
rect 6066 16718 6078 16770
rect 6130 16718 6142 16770
rect 14018 16718 14030 16770
rect 14082 16718 14094 16770
rect 18162 16718 18174 16770
rect 18226 16718 18238 16770
rect 18498 16718 18510 16770
rect 18562 16718 18574 16770
rect 21746 16718 21758 16770
rect 21810 16718 21822 16770
rect 23874 16718 23886 16770
rect 23938 16718 23950 16770
rect 26002 16718 26014 16770
rect 26066 16718 26078 16770
rect 28130 16718 28142 16770
rect 28194 16718 28206 16770
rect 30370 16718 30382 16770
rect 30434 16718 30446 16770
rect 32498 16718 32510 16770
rect 32562 16718 32574 16770
rect 12798 16706 12850 16718
rect 33182 16706 33234 16718
rect 12686 16658 12738 16670
rect 12686 16594 12738 16606
rect 15262 16658 15314 16670
rect 15262 16594 15314 16606
rect 16718 16658 16770 16670
rect 16718 16594 16770 16606
rect 1344 16490 34608 16524
rect 1344 16438 5372 16490
rect 5424 16438 5476 16490
rect 5528 16438 5580 16490
rect 5632 16438 13688 16490
rect 13740 16438 13792 16490
rect 13844 16438 13896 16490
rect 13948 16438 22004 16490
rect 22056 16438 22108 16490
rect 22160 16438 22212 16490
rect 22264 16438 30320 16490
rect 30372 16438 30424 16490
rect 30476 16438 30528 16490
rect 30580 16438 34608 16490
rect 1344 16404 34608 16438
rect 17950 16322 18002 16334
rect 5730 16270 5742 16322
rect 5794 16319 5806 16322
rect 6290 16319 6302 16322
rect 5794 16273 6302 16319
rect 5794 16270 5806 16273
rect 6290 16270 6302 16273
rect 6354 16270 6366 16322
rect 17950 16258 18002 16270
rect 5742 16210 5794 16222
rect 5058 16158 5070 16210
rect 5122 16158 5134 16210
rect 5742 16146 5794 16158
rect 6302 16210 6354 16222
rect 17726 16210 17778 16222
rect 10770 16158 10782 16210
rect 10834 16158 10846 16210
rect 12898 16158 12910 16210
rect 12962 16158 12974 16210
rect 13682 16158 13694 16210
rect 13746 16158 13758 16210
rect 17378 16158 17390 16210
rect 17442 16158 17454 16210
rect 6302 16146 6354 16158
rect 17726 16146 17778 16158
rect 23438 16210 23490 16222
rect 23438 16146 23490 16158
rect 24446 16210 24498 16222
rect 24446 16146 24498 16158
rect 28030 16210 28082 16222
rect 28030 16146 28082 16158
rect 29262 16210 29314 16222
rect 34178 16158 34190 16210
rect 34242 16158 34254 16210
rect 29262 16146 29314 16158
rect 14814 16098 14866 16110
rect 2258 16046 2270 16098
rect 2322 16046 2334 16098
rect 10098 16046 10110 16098
rect 10162 16046 10174 16098
rect 13794 16046 13806 16098
rect 13858 16046 13870 16098
rect 14814 16034 14866 16046
rect 15486 16098 15538 16110
rect 15486 16034 15538 16046
rect 15710 16098 15762 16110
rect 15710 16034 15762 16046
rect 15934 16098 15986 16110
rect 15934 16034 15986 16046
rect 16606 16098 16658 16110
rect 22430 16098 22482 16110
rect 17266 16046 17278 16098
rect 17330 16046 17342 16098
rect 19058 16046 19070 16098
rect 19122 16046 19134 16098
rect 16606 16034 16658 16046
rect 22430 16034 22482 16046
rect 23662 16098 23714 16110
rect 27022 16098 27074 16110
rect 24658 16046 24670 16098
rect 24722 16046 24734 16098
rect 23662 16034 23714 16046
rect 27022 16034 27074 16046
rect 27918 16098 27970 16110
rect 27918 16034 27970 16046
rect 28142 16098 28194 16110
rect 28142 16034 28194 16046
rect 29150 16098 29202 16110
rect 29150 16034 29202 16046
rect 29374 16098 29426 16110
rect 29374 16034 29426 16046
rect 29822 16098 29874 16110
rect 29822 16034 29874 16046
rect 30046 16098 30098 16110
rect 31378 16046 31390 16098
rect 31442 16046 31454 16098
rect 30046 16034 30098 16046
rect 14142 15986 14194 15998
rect 2930 15934 2942 15986
rect 2994 15934 3006 15986
rect 14142 15922 14194 15934
rect 14478 15986 14530 15998
rect 14478 15922 14530 15934
rect 15038 15986 15090 15998
rect 15038 15922 15090 15934
rect 15150 15986 15202 15998
rect 15150 15922 15202 15934
rect 16046 15986 16098 15998
rect 16046 15922 16098 15934
rect 16158 15986 16210 15998
rect 16158 15922 16210 15934
rect 16942 15986 16994 15998
rect 16942 15922 16994 15934
rect 18510 15986 18562 15998
rect 18510 15922 18562 15934
rect 18622 15986 18674 15998
rect 18622 15922 18674 15934
rect 21422 15986 21474 15998
rect 21422 15922 21474 15934
rect 22206 15986 22258 15998
rect 22206 15922 22258 15934
rect 22654 15986 22706 15998
rect 22654 15922 22706 15934
rect 22766 15986 22818 15998
rect 22766 15922 22818 15934
rect 24334 15986 24386 15998
rect 24334 15922 24386 15934
rect 27582 15986 27634 15998
rect 27582 15922 27634 15934
rect 28366 15986 28418 15998
rect 32050 15934 32062 15986
rect 32114 15934 32126 15986
rect 28366 15922 28418 15934
rect 9662 15874 9714 15886
rect 9662 15810 9714 15822
rect 14254 15874 14306 15886
rect 14254 15810 14306 15822
rect 16830 15874 16882 15886
rect 18846 15874 18898 15886
rect 18274 15822 18286 15874
rect 18338 15822 18350 15874
rect 16830 15810 16882 15822
rect 18846 15810 18898 15822
rect 21534 15874 21586 15886
rect 21534 15810 21586 15822
rect 21646 15874 21698 15886
rect 27358 15874 27410 15886
rect 23986 15822 23998 15874
rect 24050 15822 24062 15874
rect 21646 15810 21698 15822
rect 27358 15810 27410 15822
rect 27694 15874 27746 15886
rect 30370 15822 30382 15874
rect 30434 15822 30446 15874
rect 27694 15810 27746 15822
rect 1344 15706 34768 15740
rect 1344 15654 9530 15706
rect 9582 15654 9634 15706
rect 9686 15654 9738 15706
rect 9790 15654 17846 15706
rect 17898 15654 17950 15706
rect 18002 15654 18054 15706
rect 18106 15654 26162 15706
rect 26214 15654 26266 15706
rect 26318 15654 26370 15706
rect 26422 15654 34478 15706
rect 34530 15654 34582 15706
rect 34634 15654 34686 15706
rect 34738 15654 34768 15706
rect 1344 15620 34768 15654
rect 14814 15538 14866 15550
rect 14814 15474 14866 15486
rect 15486 15538 15538 15550
rect 15486 15474 15538 15486
rect 15598 15538 15650 15550
rect 15598 15474 15650 15486
rect 27358 15538 27410 15550
rect 27358 15474 27410 15486
rect 27582 15538 27634 15550
rect 27582 15474 27634 15486
rect 29934 15538 29986 15550
rect 33058 15486 33070 15538
rect 33122 15486 33134 15538
rect 29934 15474 29986 15486
rect 14702 15426 14754 15438
rect 11890 15374 11902 15426
rect 11954 15374 11966 15426
rect 14702 15362 14754 15374
rect 16270 15426 16322 15438
rect 16270 15362 16322 15374
rect 16718 15426 16770 15438
rect 16718 15362 16770 15374
rect 16830 15426 16882 15438
rect 26126 15426 26178 15438
rect 22866 15374 22878 15426
rect 22930 15374 22942 15426
rect 16830 15362 16882 15374
rect 26126 15362 26178 15374
rect 26350 15426 26402 15438
rect 26350 15362 26402 15374
rect 27694 15426 27746 15438
rect 27694 15362 27746 15374
rect 28814 15426 28866 15438
rect 28814 15362 28866 15374
rect 29262 15426 29314 15438
rect 29262 15362 29314 15374
rect 29486 15426 29538 15438
rect 29486 15362 29538 15374
rect 30382 15426 30434 15438
rect 30382 15362 30434 15374
rect 30942 15426 30994 15438
rect 30942 15362 30994 15374
rect 32398 15426 32450 15438
rect 32398 15362 32450 15374
rect 8990 15314 9042 15326
rect 15262 15314 15314 15326
rect 5730 15262 5742 15314
rect 5794 15262 5806 15314
rect 11218 15262 11230 15314
rect 11282 15262 11294 15314
rect 8990 15250 9042 15262
rect 15262 15250 15314 15262
rect 15374 15314 15426 15326
rect 15374 15250 15426 15262
rect 15710 15314 15762 15326
rect 15710 15250 15762 15262
rect 17950 15314 18002 15326
rect 31054 15314 31106 15326
rect 18162 15262 18174 15314
rect 18226 15262 18238 15314
rect 28578 15262 28590 15314
rect 28642 15262 28654 15314
rect 17950 15250 18002 15262
rect 31054 15250 31106 15262
rect 31502 15314 31554 15326
rect 33630 15314 33682 15326
rect 31714 15262 31726 15314
rect 31778 15262 31790 15314
rect 32050 15262 32062 15314
rect 32114 15262 32126 15314
rect 31502 15250 31554 15262
rect 33630 15250 33682 15262
rect 16382 15202 16434 15214
rect 29822 15202 29874 15214
rect 6402 15150 6414 15202
rect 6466 15150 6478 15202
rect 8530 15150 8542 15202
rect 8594 15150 8606 15202
rect 14018 15150 14030 15202
rect 14082 15150 14094 15202
rect 26002 15150 26014 15202
rect 26066 15150 26078 15202
rect 29250 15150 29262 15202
rect 29314 15150 29326 15202
rect 16382 15138 16434 15150
rect 29822 15138 29874 15150
rect 30494 15202 30546 15214
rect 30494 15138 30546 15150
rect 30606 15202 30658 15214
rect 30606 15138 30658 15150
rect 33406 15202 33458 15214
rect 33406 15138 33458 15150
rect 31278 15090 31330 15102
rect 31278 15026 31330 15038
rect 32062 15090 32114 15102
rect 32062 15026 32114 15038
rect 1344 14922 34608 14956
rect 1344 14870 5372 14922
rect 5424 14870 5476 14922
rect 5528 14870 5580 14922
rect 5632 14870 13688 14922
rect 13740 14870 13792 14922
rect 13844 14870 13896 14922
rect 13948 14870 22004 14922
rect 22056 14870 22108 14922
rect 22160 14870 22212 14922
rect 22264 14870 30320 14922
rect 30372 14870 30424 14922
rect 30476 14870 30528 14922
rect 30580 14870 34608 14922
rect 1344 14836 34608 14870
rect 17950 14754 18002 14766
rect 17950 14690 18002 14702
rect 18174 14754 18226 14766
rect 18174 14690 18226 14702
rect 28254 14754 28306 14766
rect 28254 14690 28306 14702
rect 29262 14754 29314 14766
rect 29262 14690 29314 14702
rect 30830 14754 30882 14766
rect 30830 14690 30882 14702
rect 32174 14754 32226 14766
rect 32174 14690 32226 14702
rect 32622 14754 32674 14766
rect 32622 14690 32674 14702
rect 16494 14642 16546 14654
rect 29598 14642 29650 14654
rect 4610 14590 4622 14642
rect 4674 14590 4686 14642
rect 20626 14590 20638 14642
rect 20690 14590 20702 14642
rect 21298 14590 21310 14642
rect 21362 14590 21374 14642
rect 23426 14590 23438 14642
rect 23490 14590 23502 14642
rect 16494 14578 16546 14590
rect 29598 14578 29650 14590
rect 31166 14642 31218 14654
rect 31166 14578 31218 14590
rect 5630 14530 5682 14542
rect 16158 14530 16210 14542
rect 1810 14478 1822 14530
rect 1874 14478 1886 14530
rect 12674 14478 12686 14530
rect 12738 14478 12750 14530
rect 5630 14466 5682 14478
rect 16158 14466 16210 14478
rect 17054 14530 17106 14542
rect 17054 14466 17106 14478
rect 17390 14530 17442 14542
rect 17390 14466 17442 14478
rect 17502 14530 17554 14542
rect 27246 14530 27298 14542
rect 19618 14478 19630 14530
rect 19682 14478 19694 14530
rect 20738 14478 20750 14530
rect 20802 14478 20814 14530
rect 24210 14478 24222 14530
rect 24274 14478 24286 14530
rect 17502 14466 17554 14478
rect 27246 14466 27298 14478
rect 28030 14530 28082 14542
rect 28030 14466 28082 14478
rect 29374 14530 29426 14542
rect 32846 14530 32898 14542
rect 31826 14478 31838 14530
rect 31890 14478 31902 14530
rect 32386 14478 32398 14530
rect 32450 14478 32462 14530
rect 29374 14466 29426 14478
rect 32846 14466 32898 14478
rect 15822 14418 15874 14430
rect 2482 14366 2494 14418
rect 2546 14366 2558 14418
rect 8418 14366 8430 14418
rect 8482 14366 8494 14418
rect 15822 14354 15874 14366
rect 17726 14418 17778 14430
rect 20078 14418 20130 14430
rect 19394 14366 19406 14418
rect 19458 14366 19470 14418
rect 17726 14354 17778 14366
rect 20078 14354 20130 14366
rect 27470 14418 27522 14430
rect 27470 14354 27522 14366
rect 27582 14418 27634 14430
rect 27582 14354 27634 14366
rect 29710 14418 29762 14430
rect 29710 14354 29762 14366
rect 30718 14418 30770 14430
rect 31266 14366 31278 14418
rect 31330 14366 31342 14418
rect 31602 14366 31614 14418
rect 31666 14366 31678 14418
rect 30718 14354 30770 14366
rect 5070 14306 5122 14318
rect 13582 14306 13634 14318
rect 5954 14254 5966 14306
rect 6018 14254 6030 14306
rect 5070 14242 5122 14254
rect 13582 14242 13634 14254
rect 15934 14306 15986 14318
rect 15934 14242 15986 14254
rect 20302 14306 20354 14318
rect 20302 14242 20354 14254
rect 20526 14306 20578 14318
rect 20526 14242 20578 14254
rect 32510 14306 32562 14318
rect 32510 14242 32562 14254
rect 1344 14138 34768 14172
rect 1344 14086 9530 14138
rect 9582 14086 9634 14138
rect 9686 14086 9738 14138
rect 9790 14086 17846 14138
rect 17898 14086 17950 14138
rect 18002 14086 18054 14138
rect 18106 14086 26162 14138
rect 26214 14086 26266 14138
rect 26318 14086 26370 14138
rect 26422 14086 34478 14138
rect 34530 14086 34582 14138
rect 34634 14086 34686 14138
rect 34738 14086 34768 14138
rect 1344 14052 34768 14086
rect 6526 13970 6578 13982
rect 6526 13906 6578 13918
rect 10670 13970 10722 13982
rect 10670 13906 10722 13918
rect 11118 13970 11170 13982
rect 18398 13970 18450 13982
rect 17378 13918 17390 13970
rect 17442 13918 17454 13970
rect 11118 13906 11170 13918
rect 18398 13906 18450 13918
rect 18846 13970 18898 13982
rect 23662 13970 23714 13982
rect 22866 13918 22878 13970
rect 22930 13918 22942 13970
rect 18846 13906 18898 13918
rect 23662 13906 23714 13918
rect 24222 13970 24274 13982
rect 24222 13906 24274 13918
rect 25678 13970 25730 13982
rect 25678 13906 25730 13918
rect 31278 13970 31330 13982
rect 32274 13918 32286 13970
rect 32338 13918 32350 13970
rect 31278 13906 31330 13918
rect 10558 13858 10610 13870
rect 10558 13794 10610 13806
rect 10894 13858 10946 13870
rect 10894 13794 10946 13806
rect 11790 13858 11842 13870
rect 11790 13794 11842 13806
rect 15934 13858 15986 13870
rect 15934 13794 15986 13806
rect 19406 13858 19458 13870
rect 20402 13806 20414 13858
rect 20466 13806 20478 13858
rect 29922 13806 29934 13858
rect 29986 13806 29998 13858
rect 19406 13794 19458 13806
rect 6302 13746 6354 13758
rect 5394 13694 5406 13746
rect 5458 13694 5470 13746
rect 5618 13694 5630 13746
rect 5682 13694 5694 13746
rect 6302 13682 6354 13694
rect 6414 13746 6466 13758
rect 6414 13682 6466 13694
rect 6750 13746 6802 13758
rect 15822 13746 15874 13758
rect 10098 13694 10110 13746
rect 10162 13694 10174 13746
rect 10322 13694 10334 13746
rect 10386 13694 10398 13746
rect 11330 13694 11342 13746
rect 11394 13694 11406 13746
rect 15250 13694 15262 13746
rect 15314 13694 15326 13746
rect 6750 13682 6802 13694
rect 15822 13682 15874 13694
rect 17726 13746 17778 13758
rect 18734 13746 18786 13758
rect 18162 13694 18174 13746
rect 18226 13694 18238 13746
rect 17726 13682 17778 13694
rect 18734 13682 18786 13694
rect 19070 13746 19122 13758
rect 19070 13682 19122 13694
rect 20078 13746 20130 13758
rect 20078 13682 20130 13694
rect 22206 13746 22258 13758
rect 23550 13746 23602 13758
rect 22642 13694 22654 13746
rect 22706 13694 22718 13746
rect 22206 13682 22258 13694
rect 23550 13682 23602 13694
rect 23886 13746 23938 13758
rect 26126 13746 26178 13758
rect 25442 13694 25454 13746
rect 25506 13694 25518 13746
rect 23886 13682 23938 13694
rect 26126 13682 26178 13694
rect 26350 13746 26402 13758
rect 26350 13682 26402 13694
rect 26686 13746 26738 13758
rect 26686 13682 26738 13694
rect 27022 13746 27074 13758
rect 31726 13746 31778 13758
rect 30706 13694 30718 13746
rect 30770 13694 30782 13746
rect 27022 13682 27074 13694
rect 31726 13682 31778 13694
rect 33182 13746 33234 13758
rect 33182 13682 33234 13694
rect 33630 13746 33682 13758
rect 33630 13682 33682 13694
rect 5854 13634 5906 13646
rect 5854 13570 5906 13582
rect 7758 13634 7810 13646
rect 26462 13634 26514 13646
rect 10882 13582 10894 13634
rect 10946 13582 10958 13634
rect 7758 13570 7810 13582
rect 26462 13570 26514 13582
rect 27246 13634 27298 13646
rect 27794 13582 27806 13634
rect 27858 13582 27870 13634
rect 27246 13570 27298 13582
rect 7870 13522 7922 13534
rect 7870 13458 7922 13470
rect 11678 13522 11730 13534
rect 11678 13458 11730 13470
rect 21310 13522 21362 13534
rect 21310 13458 21362 13470
rect 21758 13522 21810 13534
rect 21758 13458 21810 13470
rect 21982 13522 22034 13534
rect 21982 13458 22034 13470
rect 26910 13522 26962 13534
rect 26910 13458 26962 13470
rect 27358 13522 27410 13534
rect 27358 13458 27410 13470
rect 31054 13522 31106 13534
rect 31054 13458 31106 13470
rect 31390 13522 31442 13534
rect 31390 13458 31442 13470
rect 31950 13522 32002 13534
rect 31950 13458 32002 13470
rect 33294 13522 33346 13534
rect 33294 13458 33346 13470
rect 33518 13522 33570 13534
rect 33518 13458 33570 13470
rect 1344 13354 34608 13388
rect 1344 13302 5372 13354
rect 5424 13302 5476 13354
rect 5528 13302 5580 13354
rect 5632 13302 13688 13354
rect 13740 13302 13792 13354
rect 13844 13302 13896 13354
rect 13948 13302 22004 13354
rect 22056 13302 22108 13354
rect 22160 13302 22212 13354
rect 22264 13302 30320 13354
rect 30372 13302 30424 13354
rect 30476 13302 30528 13354
rect 30580 13302 34608 13354
rect 1344 13268 34608 13302
rect 6526 13186 6578 13198
rect 6526 13122 6578 13134
rect 18622 13186 18674 13198
rect 18622 13122 18674 13134
rect 20302 13186 20354 13198
rect 20302 13122 20354 13134
rect 22094 13186 22146 13198
rect 29486 13186 29538 13198
rect 29138 13134 29150 13186
rect 29202 13134 29214 13186
rect 22094 13122 22146 13134
rect 29486 13122 29538 13134
rect 4622 13074 4674 13086
rect 4622 13010 4674 13022
rect 7422 13074 7474 13086
rect 11230 13074 11282 13086
rect 10770 13022 10782 13074
rect 10834 13022 10846 13074
rect 7422 13010 7474 13022
rect 11230 13010 11282 13022
rect 12126 13074 12178 13086
rect 12126 13010 12178 13022
rect 15374 13074 15426 13086
rect 15374 13010 15426 13022
rect 17054 13074 17106 13086
rect 17054 13010 17106 13022
rect 17950 13074 18002 13086
rect 17950 13010 18002 13022
rect 20078 13074 20130 13086
rect 20078 13010 20130 13022
rect 22318 13074 22370 13086
rect 22318 13010 22370 13022
rect 22990 13074 23042 13086
rect 29710 13074 29762 13086
rect 24770 13022 24782 13074
rect 24834 13022 24846 13074
rect 26898 13022 26910 13074
rect 26962 13022 26974 13074
rect 31266 13022 31278 13074
rect 31330 13022 31342 13074
rect 33394 13022 33406 13074
rect 33458 13022 33470 13074
rect 22990 13010 23042 13022
rect 29710 13010 29762 13022
rect 3614 12962 3666 12974
rect 3614 12898 3666 12910
rect 4286 12962 4338 12974
rect 5630 12962 5682 12974
rect 5058 12910 5070 12962
rect 5122 12910 5134 12962
rect 4286 12898 4338 12910
rect 5630 12898 5682 12910
rect 5854 12962 5906 12974
rect 5854 12898 5906 12910
rect 6078 12962 6130 12974
rect 6078 12898 6130 12910
rect 6750 12962 6802 12974
rect 6750 12898 6802 12910
rect 7086 12962 7138 12974
rect 12574 12962 12626 12974
rect 7970 12910 7982 12962
rect 8034 12910 8046 12962
rect 11666 12910 11678 12962
rect 11730 12910 11742 12962
rect 7086 12898 7138 12910
rect 12574 12898 12626 12910
rect 18846 12962 18898 12974
rect 18846 12898 18898 12910
rect 19518 12962 19570 12974
rect 20862 12962 20914 12974
rect 27470 12962 27522 12974
rect 20514 12910 20526 12962
rect 20578 12910 20590 12962
rect 21858 12910 21870 12962
rect 21922 12910 21934 12962
rect 24098 12910 24110 12962
rect 24162 12910 24174 12962
rect 34066 12910 34078 12962
rect 34130 12910 34142 12962
rect 19518 12898 19570 12910
rect 20862 12898 20914 12910
rect 27470 12898 27522 12910
rect 7534 12850 7586 12862
rect 13806 12850 13858 12862
rect 19294 12850 19346 12862
rect 8642 12798 8654 12850
rect 8706 12798 8718 12850
rect 14130 12798 14142 12850
rect 14194 12798 14206 12850
rect 7534 12786 7586 12798
rect 13806 12786 13858 12798
rect 19294 12786 19346 12798
rect 19854 12850 19906 12862
rect 19854 12786 19906 12798
rect 21646 12850 21698 12862
rect 21646 12786 21698 12798
rect 22542 12850 22594 12862
rect 22542 12786 22594 12798
rect 22878 12850 22930 12862
rect 22878 12786 22930 12798
rect 27358 12850 27410 12862
rect 27358 12786 27410 12798
rect 3726 12738 3778 12750
rect 3726 12674 3778 12686
rect 3838 12738 3890 12750
rect 3838 12674 3890 12686
rect 4510 12738 4562 12750
rect 4510 12674 4562 12686
rect 4734 12738 4786 12750
rect 4734 12674 4786 12686
rect 6862 12738 6914 12750
rect 6862 12674 6914 12686
rect 11118 12738 11170 12750
rect 11118 12674 11170 12686
rect 11342 12738 11394 12750
rect 11342 12674 11394 12686
rect 12014 12738 12066 12750
rect 12014 12674 12066 12686
rect 18398 12738 18450 12750
rect 18398 12674 18450 12686
rect 18510 12738 18562 12750
rect 18510 12674 18562 12686
rect 19406 12738 19458 12750
rect 19406 12674 19458 12686
rect 19742 12738 19794 12750
rect 19742 12674 19794 12686
rect 22430 12738 22482 12750
rect 22430 12674 22482 12686
rect 27134 12738 27186 12750
rect 27134 12674 27186 12686
rect 1344 12570 34768 12604
rect 1344 12518 9530 12570
rect 9582 12518 9634 12570
rect 9686 12518 9738 12570
rect 9790 12518 17846 12570
rect 17898 12518 17950 12570
rect 18002 12518 18054 12570
rect 18106 12518 26162 12570
rect 26214 12518 26266 12570
rect 26318 12518 26370 12570
rect 26422 12518 34478 12570
rect 34530 12518 34582 12570
rect 34634 12518 34686 12570
rect 34738 12518 34768 12570
rect 1344 12484 34768 12518
rect 4174 12402 4226 12414
rect 5630 12402 5682 12414
rect 5282 12350 5294 12402
rect 5346 12350 5358 12402
rect 4174 12338 4226 12350
rect 5630 12338 5682 12350
rect 6414 12402 6466 12414
rect 9886 12402 9938 12414
rect 7074 12350 7086 12402
rect 7138 12350 7150 12402
rect 6414 12338 6466 12350
rect 9886 12338 9938 12350
rect 20638 12402 20690 12414
rect 20962 12350 20974 12402
rect 21026 12350 21038 12402
rect 20638 12338 20690 12350
rect 3166 12290 3218 12302
rect 3166 12226 3218 12238
rect 3614 12290 3666 12302
rect 8654 12290 8706 12302
rect 6738 12238 6750 12290
rect 6802 12238 6814 12290
rect 7970 12238 7982 12290
rect 8034 12238 8046 12290
rect 3614 12226 3666 12238
rect 8654 12226 8706 12238
rect 8990 12290 9042 12302
rect 10558 12290 10610 12302
rect 9538 12238 9550 12290
rect 9602 12238 9614 12290
rect 18162 12238 18174 12290
rect 18226 12238 18238 12290
rect 23650 12238 23662 12290
rect 23714 12238 23726 12290
rect 8990 12226 9042 12238
rect 10558 12226 10610 12238
rect 2830 12178 2882 12190
rect 2830 12114 2882 12126
rect 3502 12178 3554 12190
rect 4510 12178 4562 12190
rect 4958 12178 5010 12190
rect 3826 12126 3838 12178
rect 3890 12126 3902 12178
rect 4386 12126 4398 12178
rect 4450 12126 4462 12178
rect 4722 12126 4734 12178
rect 4786 12126 4798 12178
rect 3502 12114 3554 12126
rect 4510 12114 4562 12126
rect 4958 12114 5010 12126
rect 7422 12178 7474 12190
rect 7422 12114 7474 12126
rect 8318 12178 8370 12190
rect 8318 12114 8370 12126
rect 10334 12178 10386 12190
rect 10334 12114 10386 12126
rect 11006 12178 11058 12190
rect 26014 12178 26066 12190
rect 31502 12178 31554 12190
rect 12674 12126 12686 12178
rect 12738 12126 12750 12178
rect 17490 12126 17502 12178
rect 17554 12126 17566 12178
rect 24322 12126 24334 12178
rect 24386 12126 24398 12178
rect 26562 12126 26574 12178
rect 26626 12126 26638 12178
rect 11006 12114 11058 12126
rect 26014 12114 26066 12126
rect 31502 12114 31554 12126
rect 6078 12066 6130 12078
rect 6078 12002 6130 12014
rect 10782 12066 10834 12078
rect 13570 12014 13582 12066
rect 13634 12014 13646 12066
rect 20290 12014 20302 12066
rect 20354 12014 20366 12066
rect 21522 12014 21534 12066
rect 21586 12014 21598 12066
rect 26674 12014 26686 12066
rect 26738 12014 26750 12066
rect 10782 12002 10834 12014
rect 31390 11954 31442 11966
rect 5842 11902 5854 11954
rect 5906 11951 5918 11954
rect 6178 11951 6190 11954
rect 5906 11905 6190 11951
rect 5906 11902 5918 11905
rect 6178 11902 6190 11905
rect 6242 11902 6254 11954
rect 31390 11890 31442 11902
rect 31726 11954 31778 11966
rect 31726 11890 31778 11902
rect 31838 11954 31890 11966
rect 31838 11890 31890 11902
rect 1344 11786 34608 11820
rect 1344 11734 5372 11786
rect 5424 11734 5476 11786
rect 5528 11734 5580 11786
rect 5632 11734 13688 11786
rect 13740 11734 13792 11786
rect 13844 11734 13896 11786
rect 13948 11734 22004 11786
rect 22056 11734 22108 11786
rect 22160 11734 22212 11786
rect 22264 11734 30320 11786
rect 30372 11734 30424 11786
rect 30476 11734 30528 11786
rect 30580 11734 34608 11786
rect 1344 11700 34608 11734
rect 6862 11618 6914 11630
rect 6862 11554 6914 11566
rect 8654 11618 8706 11630
rect 8654 11554 8706 11566
rect 8878 11618 8930 11630
rect 8878 11554 8930 11566
rect 17614 11618 17666 11630
rect 17614 11554 17666 11566
rect 20414 11618 20466 11630
rect 20414 11554 20466 11566
rect 22766 11618 22818 11630
rect 22766 11554 22818 11566
rect 2382 11506 2434 11518
rect 2382 11442 2434 11454
rect 3054 11506 3106 11518
rect 3054 11442 3106 11454
rect 4286 11506 4338 11518
rect 4286 11442 4338 11454
rect 6414 11506 6466 11518
rect 6414 11442 6466 11454
rect 9886 11506 9938 11518
rect 17838 11506 17890 11518
rect 10658 11454 10670 11506
rect 10722 11454 10734 11506
rect 14242 11454 14254 11506
rect 14306 11454 14318 11506
rect 16370 11454 16382 11506
rect 16434 11454 16446 11506
rect 9886 11442 9938 11454
rect 17838 11442 17890 11454
rect 18734 11506 18786 11518
rect 20526 11506 20578 11518
rect 19506 11454 19518 11506
rect 19570 11454 19582 11506
rect 18734 11442 18786 11454
rect 20526 11442 20578 11454
rect 21422 11506 21474 11518
rect 21422 11442 21474 11454
rect 22878 11506 22930 11518
rect 27346 11454 27358 11506
rect 27410 11454 27422 11506
rect 32050 11454 32062 11506
rect 32114 11454 32126 11506
rect 34178 11454 34190 11506
rect 34242 11454 34254 11506
rect 22878 11442 22930 11454
rect 2158 11394 2210 11406
rect 2158 11330 2210 11342
rect 3278 11394 3330 11406
rect 3278 11330 3330 11342
rect 3502 11394 3554 11406
rect 3502 11330 3554 11342
rect 3614 11394 3666 11406
rect 3614 11330 3666 11342
rect 4174 11394 4226 11406
rect 4174 11330 4226 11342
rect 5518 11394 5570 11406
rect 5518 11330 5570 11342
rect 6078 11394 6130 11406
rect 6078 11330 6130 11342
rect 6302 11394 6354 11406
rect 6302 11330 6354 11342
rect 6526 11394 6578 11406
rect 6526 11330 6578 11342
rect 7086 11394 7138 11406
rect 7086 11330 7138 11342
rect 7534 11394 7586 11406
rect 7534 11330 7586 11342
rect 8990 11394 9042 11406
rect 8990 11330 9042 11342
rect 9550 11394 9602 11406
rect 9550 11330 9602 11342
rect 10446 11394 10498 11406
rect 19630 11394 19682 11406
rect 13458 11342 13470 11394
rect 13522 11342 13534 11394
rect 19394 11342 19406 11394
rect 19458 11342 19470 11394
rect 10446 11330 10498 11342
rect 19630 11330 19682 11342
rect 19854 11394 19906 11406
rect 21534 11394 21586 11406
rect 29486 11394 29538 11406
rect 20066 11342 20078 11394
rect 20130 11342 20142 11394
rect 21858 11342 21870 11394
rect 21922 11342 21934 11394
rect 24434 11342 24446 11394
rect 24498 11342 24510 11394
rect 29138 11342 29150 11394
rect 29202 11342 29214 11394
rect 30258 11342 30270 11394
rect 30322 11342 30334 11394
rect 31266 11342 31278 11394
rect 31330 11342 31342 11394
rect 19854 11330 19906 11342
rect 21534 11330 21586 11342
rect 29486 11330 29538 11342
rect 4510 11282 4562 11294
rect 7422 11282 7474 11294
rect 4610 11230 4622 11282
rect 4674 11230 4686 11282
rect 5842 11230 5854 11282
rect 5906 11230 5918 11282
rect 4510 11218 4562 11230
rect 7422 11218 7474 11230
rect 7870 11282 7922 11294
rect 7870 11218 7922 11230
rect 8206 11282 8258 11294
rect 8206 11218 8258 11230
rect 8542 11282 8594 11294
rect 8542 11218 8594 11230
rect 9662 11282 9714 11294
rect 9662 11218 9714 11230
rect 9998 11282 10050 11294
rect 9998 11218 10050 11230
rect 16718 11282 16770 11294
rect 25218 11230 25230 11282
rect 25282 11230 25294 11282
rect 16718 11218 16770 11230
rect 2270 11170 2322 11182
rect 2270 11106 2322 11118
rect 2494 11170 2546 11182
rect 2494 11106 2546 11118
rect 2606 11170 2658 11182
rect 2606 11106 2658 11118
rect 3726 11170 3778 11182
rect 3726 11106 3778 11118
rect 4398 11170 4450 11182
rect 4398 11106 4450 11118
rect 7310 11170 7362 11182
rect 7310 11106 7362 11118
rect 8094 11170 8146 11182
rect 8094 11106 8146 11118
rect 10670 11170 10722 11182
rect 10670 11106 10722 11118
rect 16830 11170 16882 11182
rect 18286 11170 18338 11182
rect 17266 11118 17278 11170
rect 17330 11118 17342 11170
rect 16830 11106 16882 11118
rect 18286 11106 18338 11118
rect 29598 11170 29650 11182
rect 29598 11106 29650 11118
rect 29710 11170 29762 11182
rect 30034 11118 30046 11170
rect 30098 11118 30110 11170
rect 29710 11106 29762 11118
rect 1344 11002 34768 11036
rect 1344 10950 9530 11002
rect 9582 10950 9634 11002
rect 9686 10950 9738 11002
rect 9790 10950 17846 11002
rect 17898 10950 17950 11002
rect 18002 10950 18054 11002
rect 18106 10950 26162 11002
rect 26214 10950 26266 11002
rect 26318 10950 26370 11002
rect 26422 10950 34478 11002
rect 34530 10950 34582 11002
rect 34634 10950 34686 11002
rect 34738 10950 34768 11002
rect 1344 10916 34768 10950
rect 3278 10834 3330 10846
rect 3278 10770 3330 10782
rect 3726 10834 3778 10846
rect 3726 10770 3778 10782
rect 4734 10834 4786 10846
rect 4734 10770 4786 10782
rect 4958 10834 5010 10846
rect 4958 10770 5010 10782
rect 10334 10834 10386 10846
rect 10334 10770 10386 10782
rect 10894 10834 10946 10846
rect 10894 10770 10946 10782
rect 17390 10834 17442 10846
rect 17390 10770 17442 10782
rect 25790 10834 25842 10846
rect 25790 10770 25842 10782
rect 3838 10722 3890 10734
rect 3838 10658 3890 10670
rect 7982 10722 8034 10734
rect 7982 10658 8034 10670
rect 8990 10722 9042 10734
rect 8990 10658 9042 10670
rect 10446 10722 10498 10734
rect 10446 10658 10498 10670
rect 11118 10722 11170 10734
rect 26014 10722 26066 10734
rect 33294 10722 33346 10734
rect 13010 10670 13022 10722
rect 13074 10670 13086 10722
rect 30706 10670 30718 10722
rect 30770 10670 30782 10722
rect 11118 10658 11170 10670
rect 26014 10658 26066 10670
rect 33294 10658 33346 10670
rect 2718 10610 2770 10622
rect 5070 10610 5122 10622
rect 3042 10558 3054 10610
rect 3106 10558 3118 10610
rect 2718 10546 2770 10558
rect 5070 10546 5122 10558
rect 7870 10610 7922 10622
rect 7870 10546 7922 10558
rect 8206 10610 8258 10622
rect 8206 10546 8258 10558
rect 8542 10610 8594 10622
rect 8542 10546 8594 10558
rect 8878 10610 8930 10622
rect 9886 10610 9938 10622
rect 9538 10558 9550 10610
rect 9602 10558 9614 10610
rect 8878 10546 8930 10558
rect 9886 10546 9938 10558
rect 9998 10610 10050 10622
rect 9998 10546 10050 10558
rect 10670 10610 10722 10622
rect 10670 10546 10722 10558
rect 11342 10610 11394 10622
rect 16270 10610 16322 10622
rect 12338 10558 12350 10610
rect 12402 10558 12414 10610
rect 11342 10546 11394 10558
rect 16270 10546 16322 10558
rect 16494 10610 16546 10622
rect 16494 10546 16546 10558
rect 16606 10610 16658 10622
rect 16606 10546 16658 10558
rect 16830 10610 16882 10622
rect 22318 10610 22370 10622
rect 18498 10558 18510 10610
rect 18562 10558 18574 10610
rect 16830 10546 16882 10558
rect 22318 10546 22370 10558
rect 26910 10610 26962 10622
rect 27234 10558 27246 10610
rect 27298 10558 27310 10610
rect 26910 10546 26962 10558
rect 2942 10498 2994 10510
rect 2942 10434 2994 10446
rect 10222 10498 10274 10510
rect 15138 10446 15150 10498
rect 15202 10446 15214 10498
rect 17826 10446 17838 10498
rect 17890 10446 17902 10498
rect 19170 10446 19182 10498
rect 19234 10446 19246 10498
rect 21298 10446 21310 10498
rect 21362 10446 21374 10498
rect 25666 10446 25678 10498
rect 25730 10446 25742 10498
rect 10222 10434 10274 10446
rect 3614 10386 3666 10398
rect 3614 10322 3666 10334
rect 8654 10386 8706 10398
rect 33070 10386 33122 10398
rect 15810 10334 15822 10386
rect 15874 10334 15886 10386
rect 8654 10322 8706 10334
rect 33070 10322 33122 10334
rect 33406 10386 33458 10398
rect 33406 10322 33458 10334
rect 1344 10218 34608 10252
rect 1344 10166 5372 10218
rect 5424 10166 5476 10218
rect 5528 10166 5580 10218
rect 5632 10166 13688 10218
rect 13740 10166 13792 10218
rect 13844 10166 13896 10218
rect 13948 10166 22004 10218
rect 22056 10166 22108 10218
rect 22160 10166 22212 10218
rect 22264 10166 30320 10218
rect 30372 10166 30424 10218
rect 30476 10166 30528 10218
rect 30580 10166 34608 10218
rect 1344 10132 34608 10166
rect 2270 10050 2322 10062
rect 2270 9986 2322 9998
rect 2718 10050 2770 10062
rect 2718 9986 2770 9998
rect 9214 10050 9266 10062
rect 9214 9986 9266 9998
rect 19630 10050 19682 10062
rect 19630 9986 19682 9998
rect 31054 10050 31106 10062
rect 31054 9986 31106 9998
rect 6078 9938 6130 9950
rect 6078 9874 6130 9886
rect 8878 9938 8930 9950
rect 20414 9938 20466 9950
rect 30046 9938 30098 9950
rect 10546 9886 10558 9938
rect 10610 9886 10622 9938
rect 12450 9886 12462 9938
rect 12514 9886 12526 9938
rect 14466 9886 14478 9938
rect 14530 9886 14542 9938
rect 21746 9886 21758 9938
rect 21810 9886 21822 9938
rect 34178 9886 34190 9938
rect 34242 9886 34254 9938
rect 8878 9874 8930 9886
rect 20414 9874 20466 9886
rect 30046 9874 30098 9886
rect 2942 9826 2994 9838
rect 2942 9762 2994 9774
rect 3166 9826 3218 9838
rect 3166 9762 3218 9774
rect 5630 9826 5682 9838
rect 5630 9762 5682 9774
rect 9102 9826 9154 9838
rect 11454 9826 11506 9838
rect 9538 9774 9550 9826
rect 9602 9774 9614 9826
rect 9102 9762 9154 9774
rect 11454 9762 11506 9774
rect 11566 9826 11618 9838
rect 11566 9762 11618 9774
rect 12910 9826 12962 9838
rect 19742 9826 19794 9838
rect 29262 9826 29314 9838
rect 14018 9774 14030 9826
rect 14082 9774 14094 9826
rect 17826 9774 17838 9826
rect 17890 9774 17902 9826
rect 19282 9774 19294 9826
rect 19346 9774 19358 9826
rect 26898 9774 26910 9826
rect 26962 9774 26974 9826
rect 12910 9762 12962 9774
rect 19742 9762 19794 9774
rect 29262 9762 29314 9774
rect 29486 9826 29538 9838
rect 29486 9762 29538 9774
rect 29710 9826 29762 9838
rect 29710 9762 29762 9774
rect 30382 9826 30434 9838
rect 30382 9762 30434 9774
rect 30830 9826 30882 9838
rect 31266 9774 31278 9826
rect 31330 9774 31342 9826
rect 30830 9762 30882 9774
rect 3502 9714 3554 9726
rect 3502 9650 3554 9662
rect 3950 9714 4002 9726
rect 3950 9650 4002 9662
rect 5854 9714 5906 9726
rect 5854 9650 5906 9662
rect 6190 9714 6242 9726
rect 6190 9650 6242 9662
rect 8766 9714 8818 9726
rect 8766 9650 8818 9662
rect 9998 9714 10050 9726
rect 9998 9650 10050 9662
rect 10110 9714 10162 9726
rect 10110 9650 10162 9662
rect 10670 9714 10722 9726
rect 11230 9714 11282 9726
rect 10882 9662 10894 9714
rect 10946 9662 10958 9714
rect 10670 9650 10722 9662
rect 11230 9650 11282 9662
rect 13694 9714 13746 9726
rect 17278 9714 17330 9726
rect 19854 9714 19906 9726
rect 14130 9662 14142 9714
rect 14194 9662 14206 9714
rect 18610 9662 18622 9714
rect 18674 9662 18686 9714
rect 18946 9662 18958 9714
rect 19010 9662 19022 9714
rect 13694 9650 13746 9662
rect 17278 9650 17330 9662
rect 19854 9650 19906 9662
rect 21422 9714 21474 9726
rect 21422 9650 21474 9662
rect 22094 9714 22146 9726
rect 30270 9714 30322 9726
rect 22866 9662 22878 9714
rect 22930 9662 22942 9714
rect 32050 9662 32062 9714
rect 32114 9662 32126 9714
rect 22094 9650 22146 9662
rect 30270 9650 30322 9662
rect 3614 9602 3666 9614
rect 3614 9538 3666 9550
rect 3726 9602 3778 9614
rect 3726 9538 3778 9550
rect 10334 9602 10386 9614
rect 10334 9538 10386 9550
rect 12014 9602 12066 9614
rect 12014 9538 12066 9550
rect 13582 9602 13634 9614
rect 21870 9602 21922 9614
rect 18274 9550 18286 9602
rect 18338 9550 18350 9602
rect 13582 9538 13634 9550
rect 21870 9538 21922 9550
rect 28254 9602 28306 9614
rect 29486 9602 29538 9614
rect 28578 9550 28590 9602
rect 28642 9550 28654 9602
rect 28254 9538 28306 9550
rect 29486 9538 29538 9550
rect 1344 9434 34768 9468
rect 1344 9382 9530 9434
rect 9582 9382 9634 9434
rect 9686 9382 9738 9434
rect 9790 9382 17846 9434
rect 17898 9382 17950 9434
rect 18002 9382 18054 9434
rect 18106 9382 26162 9434
rect 26214 9382 26266 9434
rect 26318 9382 26370 9434
rect 26422 9382 34478 9434
rect 34530 9382 34582 9434
rect 34634 9382 34686 9434
rect 34738 9382 34768 9434
rect 1344 9348 34768 9382
rect 5294 9266 5346 9278
rect 3378 9214 3390 9266
rect 3442 9214 3454 9266
rect 5294 9202 5346 9214
rect 5406 9266 5458 9278
rect 5406 9202 5458 9214
rect 6862 9266 6914 9278
rect 6862 9202 6914 9214
rect 7870 9266 7922 9278
rect 26574 9266 26626 9278
rect 26226 9214 26238 9266
rect 26290 9214 26302 9266
rect 7870 9202 7922 9214
rect 26574 9202 26626 9214
rect 33182 9266 33234 9278
rect 33182 9202 33234 9214
rect 2494 9154 2546 9166
rect 2494 9090 2546 9102
rect 2830 9154 2882 9166
rect 2830 9090 2882 9102
rect 7758 9154 7810 9166
rect 16270 9154 16322 9166
rect 7758 9090 7810 9102
rect 9774 9098 9826 9110
rect 3166 9042 3218 9054
rect 3166 8978 3218 8990
rect 3502 9042 3554 9054
rect 4846 9042 4898 9054
rect 5518 9042 5570 9054
rect 3714 8990 3726 9042
rect 3778 8990 3790 9042
rect 5170 8990 5182 9042
rect 5234 8990 5246 9042
rect 3502 8978 3554 8990
rect 4846 8978 4898 8990
rect 5518 8978 5570 8990
rect 6414 9042 6466 9054
rect 6414 8978 6466 8990
rect 6638 9042 6690 9054
rect 6638 8978 6690 8990
rect 7646 9042 7698 9054
rect 7646 8978 7698 8990
rect 8318 9042 8370 9054
rect 8318 8978 8370 8990
rect 9550 9042 9602 9054
rect 9774 9034 9826 9046
rect 9886 9098 9938 9110
rect 10098 9102 10110 9154
rect 10162 9102 10174 9154
rect 16270 9090 16322 9102
rect 17278 9154 17330 9166
rect 33630 9154 33682 9166
rect 18834 9102 18846 9154
rect 18898 9102 18910 9154
rect 19730 9102 19742 9154
rect 19794 9102 19806 9154
rect 21746 9102 21758 9154
rect 21810 9102 21822 9154
rect 27794 9102 27806 9154
rect 27858 9102 27870 9154
rect 30370 9102 30382 9154
rect 30434 9102 30446 9154
rect 31826 9102 31838 9154
rect 31890 9102 31902 9154
rect 17278 9090 17330 9102
rect 33630 9090 33682 9102
rect 9886 9034 9938 9046
rect 11902 9042 11954 9054
rect 15038 9042 15090 9054
rect 9550 8978 9602 8990
rect 13234 8990 13246 9042
rect 13298 8990 13310 9042
rect 11902 8978 11954 8990
rect 15038 8978 15090 8990
rect 15374 9042 15426 9054
rect 24334 9042 24386 9054
rect 33070 9042 33122 9054
rect 18946 8990 18958 9042
rect 19010 8990 19022 9042
rect 19282 8990 19294 9042
rect 19346 8990 19358 9042
rect 20962 8990 20974 9042
rect 21026 8990 21038 9042
rect 24546 8990 24558 9042
rect 24610 8990 24622 9042
rect 27010 8990 27022 9042
rect 27074 8990 27086 9042
rect 30258 8990 30270 9042
rect 30322 8990 30334 9042
rect 31266 8990 31278 9042
rect 31330 8990 31342 9042
rect 15374 8978 15426 8990
rect 24334 8978 24386 8990
rect 33070 8978 33122 8990
rect 33294 9042 33346 9054
rect 33294 8978 33346 8990
rect 6526 8930 6578 8942
rect 14478 8930 14530 8942
rect 10322 8878 10334 8930
rect 10386 8878 10398 8930
rect 12226 8878 12238 8930
rect 12290 8878 12302 8930
rect 13122 8878 13134 8930
rect 13186 8878 13198 8930
rect 23874 8878 23886 8930
rect 23938 8878 23950 8930
rect 29922 8878 29934 8930
rect 29986 8878 29998 8930
rect 30594 8878 30606 8930
rect 30658 8878 30670 8930
rect 6526 8866 6578 8878
rect 14478 8866 14530 8878
rect 11678 8818 11730 8830
rect 3714 8766 3726 8818
rect 3778 8766 3790 8818
rect 11330 8766 11342 8818
rect 11394 8766 11406 8818
rect 11678 8754 11730 8766
rect 24222 8818 24274 8830
rect 24222 8754 24274 8766
rect 1344 8650 34608 8684
rect 1344 8598 5372 8650
rect 5424 8598 5476 8650
rect 5528 8598 5580 8650
rect 5632 8598 13688 8650
rect 13740 8598 13792 8650
rect 13844 8598 13896 8650
rect 13948 8598 22004 8650
rect 22056 8598 22108 8650
rect 22160 8598 22212 8650
rect 22264 8598 30320 8650
rect 30372 8598 30424 8650
rect 30476 8598 30528 8650
rect 30580 8598 34608 8650
rect 1344 8564 34608 8598
rect 12574 8482 12626 8494
rect 12574 8418 12626 8430
rect 19070 8482 19122 8494
rect 19070 8418 19122 8430
rect 2718 8370 2770 8382
rect 7198 8370 7250 8382
rect 9662 8370 9714 8382
rect 12798 8370 12850 8382
rect 22318 8370 22370 8382
rect 29934 8370 29986 8382
rect 3826 8318 3838 8370
rect 3890 8318 3902 8370
rect 9202 8318 9214 8370
rect 9266 8318 9278 8370
rect 12226 8318 12238 8370
rect 12290 8318 12302 8370
rect 13346 8318 13358 8370
rect 13410 8318 13422 8370
rect 18274 8318 18286 8370
rect 18338 8318 18350 8370
rect 23762 8318 23774 8370
rect 23826 8318 23838 8370
rect 25890 8318 25902 8370
rect 25954 8318 25966 8370
rect 28130 8318 28142 8370
rect 28194 8318 28206 8370
rect 2718 8306 2770 8318
rect 7198 8306 7250 8318
rect 9662 8306 9714 8318
rect 12798 8306 12850 8318
rect 22318 8306 22370 8318
rect 29934 8306 29986 8318
rect 30046 8370 30098 8382
rect 30046 8306 30098 8318
rect 30382 8370 30434 8382
rect 34178 8318 34190 8370
rect 34242 8318 34254 8370
rect 30382 8306 30434 8318
rect 3166 8258 3218 8270
rect 3166 8194 3218 8206
rect 3390 8258 3442 8270
rect 3390 8194 3442 8206
rect 3614 8258 3666 8270
rect 3614 8194 3666 8206
rect 4958 8258 5010 8270
rect 4958 8194 5010 8206
rect 5630 8258 5682 8270
rect 5630 8194 5682 8206
rect 5854 8258 5906 8270
rect 5854 8194 5906 8206
rect 6078 8258 6130 8270
rect 9438 8258 9490 8270
rect 6850 8206 6862 8258
rect 6914 8206 6926 8258
rect 6078 8194 6130 8206
rect 9438 8194 9490 8206
rect 9886 8258 9938 8270
rect 22094 8258 22146 8270
rect 26238 8258 26290 8270
rect 27694 8258 27746 8270
rect 30606 8258 30658 8270
rect 11666 8206 11678 8258
rect 11730 8206 11742 8258
rect 15138 8206 15150 8258
rect 15202 8206 15214 8258
rect 16706 8206 16718 8258
rect 16770 8206 16782 8258
rect 18050 8206 18062 8258
rect 18114 8206 18126 8258
rect 18946 8206 18958 8258
rect 19010 8206 19022 8258
rect 22978 8206 22990 8258
rect 23042 8206 23054 8258
rect 27122 8206 27134 8258
rect 27186 8206 27198 8258
rect 28018 8206 28030 8258
rect 28082 8206 28094 8258
rect 31266 8206 31278 8258
rect 31330 8206 31342 8258
rect 9886 8194 9938 8206
rect 22094 8194 22146 8206
rect 26238 8194 26290 8206
rect 27694 8194 27746 8206
rect 30606 8194 30658 8206
rect 2830 8146 2882 8158
rect 2830 8082 2882 8094
rect 3838 8146 3890 8158
rect 3838 8082 3890 8094
rect 4622 8146 4674 8158
rect 6526 8146 6578 8158
rect 6290 8094 6302 8146
rect 6354 8094 6366 8146
rect 4622 8082 4674 8094
rect 6526 8082 6578 8094
rect 7534 8146 7586 8158
rect 7534 8082 7586 8094
rect 8766 8146 8818 8158
rect 10110 8146 10162 8158
rect 8978 8094 8990 8146
rect 9042 8094 9054 8146
rect 8766 8082 8818 8094
rect 10110 8082 10162 8094
rect 10446 8146 10498 8158
rect 12014 8146 12066 8158
rect 11106 8094 11118 8146
rect 11170 8094 11182 8146
rect 11442 8094 11454 8146
rect 11506 8094 11518 8146
rect 10446 8082 10498 8094
rect 12014 8082 12066 8094
rect 12238 8146 12290 8158
rect 14914 8094 14926 8146
rect 14978 8094 14990 8146
rect 15810 8094 15822 8146
rect 15874 8094 15886 8146
rect 32050 8094 32062 8146
rect 32114 8094 32126 8146
rect 12238 8082 12290 8094
rect 2606 8034 2658 8046
rect 2606 7970 2658 7982
rect 4062 8034 4114 8046
rect 4062 7970 4114 7982
rect 4734 8034 4786 8046
rect 4734 7970 4786 7982
rect 5518 8034 5570 8046
rect 5518 7970 5570 7982
rect 7086 8034 7138 8046
rect 7086 7970 7138 7982
rect 7310 8034 7362 8046
rect 7310 7970 7362 7982
rect 8430 8034 8482 8046
rect 8430 7970 8482 7982
rect 8654 8034 8706 8046
rect 8654 7970 8706 7982
rect 17166 8034 17218 8046
rect 17166 7970 17218 7982
rect 21534 8034 21586 8046
rect 28254 8034 28306 8046
rect 21746 7982 21758 8034
rect 21810 7982 21822 8034
rect 26562 7982 26574 8034
rect 26626 7982 26638 8034
rect 26898 7982 26910 8034
rect 26962 7982 26974 8034
rect 30930 7982 30942 8034
rect 30994 7982 31006 8034
rect 21534 7970 21586 7982
rect 28254 7970 28306 7982
rect 1344 7866 34768 7900
rect 1344 7814 9530 7866
rect 9582 7814 9634 7866
rect 9686 7814 9738 7866
rect 9790 7814 17846 7866
rect 17898 7814 17950 7866
rect 18002 7814 18054 7866
rect 18106 7814 26162 7866
rect 26214 7814 26266 7866
rect 26318 7814 26370 7866
rect 26422 7814 34478 7866
rect 34530 7814 34582 7866
rect 34634 7814 34686 7866
rect 34738 7814 34768 7866
rect 1344 7780 34768 7814
rect 2942 7698 2994 7710
rect 6750 7698 6802 7710
rect 5170 7646 5182 7698
rect 5234 7646 5246 7698
rect 2942 7634 2994 7646
rect 6750 7634 6802 7646
rect 6862 7698 6914 7710
rect 6862 7634 6914 7646
rect 8094 7698 8146 7710
rect 8094 7634 8146 7646
rect 8878 7698 8930 7710
rect 8878 7634 8930 7646
rect 9662 7698 9714 7710
rect 11566 7698 11618 7710
rect 10546 7646 10558 7698
rect 10610 7646 10622 7698
rect 9662 7634 9714 7646
rect 11566 7634 11618 7646
rect 12574 7698 12626 7710
rect 12574 7634 12626 7646
rect 12910 7698 12962 7710
rect 12910 7634 12962 7646
rect 27470 7698 27522 7710
rect 27470 7634 27522 7646
rect 28142 7698 28194 7710
rect 28142 7634 28194 7646
rect 30270 7698 30322 7710
rect 30270 7634 30322 7646
rect 31726 7698 31778 7710
rect 31726 7634 31778 7646
rect 2158 7586 2210 7598
rect 2158 7522 2210 7534
rect 2494 7586 2546 7598
rect 2494 7522 2546 7534
rect 4510 7586 4562 7598
rect 4510 7522 4562 7534
rect 4846 7586 4898 7598
rect 23326 7586 23378 7598
rect 14354 7534 14366 7586
rect 14418 7534 14430 7586
rect 22418 7534 22430 7586
rect 22482 7534 22494 7586
rect 4846 7522 4898 7534
rect 23326 7522 23378 7534
rect 23550 7586 23602 7598
rect 23550 7522 23602 7534
rect 25902 7586 25954 7598
rect 25902 7522 25954 7534
rect 27918 7586 27970 7598
rect 27918 7522 27970 7534
rect 29486 7586 29538 7598
rect 29486 7522 29538 7534
rect 33070 7586 33122 7598
rect 33070 7522 33122 7534
rect 2830 7474 2882 7486
rect 2830 7410 2882 7422
rect 3054 7474 3106 7486
rect 3054 7410 3106 7422
rect 3502 7474 3554 7486
rect 3502 7410 3554 7422
rect 4398 7474 4450 7486
rect 4398 7410 4450 7422
rect 5182 7474 5234 7486
rect 5182 7410 5234 7422
rect 5294 7474 5346 7486
rect 5294 7410 5346 7422
rect 5518 7474 5570 7486
rect 5518 7410 5570 7422
rect 5742 7474 5794 7486
rect 5742 7410 5794 7422
rect 6638 7474 6690 7486
rect 7870 7474 7922 7486
rect 7186 7422 7198 7474
rect 7250 7422 7262 7474
rect 6638 7410 6690 7422
rect 7870 7410 7922 7422
rect 7982 7474 8034 7486
rect 7982 7410 8034 7422
rect 8206 7474 8258 7486
rect 8990 7474 9042 7486
rect 8418 7422 8430 7474
rect 8482 7422 8494 7474
rect 8206 7410 8258 7422
rect 8990 7410 9042 7422
rect 9550 7474 9602 7486
rect 9550 7410 9602 7422
rect 9774 7474 9826 7486
rect 9774 7410 9826 7422
rect 10222 7474 10274 7486
rect 10222 7410 10274 7422
rect 10894 7474 10946 7486
rect 10894 7410 10946 7422
rect 11454 7474 11506 7486
rect 11454 7410 11506 7422
rect 11678 7474 11730 7486
rect 11678 7410 11730 7422
rect 12014 7474 12066 7486
rect 15486 7474 15538 7486
rect 18286 7474 18338 7486
rect 21982 7474 22034 7486
rect 13122 7422 13134 7474
rect 13186 7422 13198 7474
rect 13346 7422 13358 7474
rect 13410 7422 13422 7474
rect 14130 7422 14142 7474
rect 14194 7422 14206 7474
rect 15250 7422 15262 7474
rect 15314 7422 15326 7474
rect 16258 7422 16270 7474
rect 16322 7422 16334 7474
rect 16482 7422 16494 7474
rect 16546 7422 16558 7474
rect 17826 7422 17838 7474
rect 17890 7422 17902 7474
rect 18722 7422 18734 7474
rect 18786 7422 18798 7474
rect 12014 7410 12066 7422
rect 15486 7410 15538 7422
rect 18286 7410 18338 7422
rect 21982 7410 22034 7422
rect 22206 7474 22258 7486
rect 22206 7410 22258 7422
rect 22766 7474 22818 7486
rect 22766 7410 22818 7422
rect 22990 7474 23042 7486
rect 22990 7410 23042 7422
rect 26014 7474 26066 7486
rect 29262 7474 29314 7486
rect 26226 7422 26238 7474
rect 26290 7422 26302 7474
rect 27570 7422 27582 7474
rect 27634 7422 27646 7474
rect 26014 7410 26066 7422
rect 29262 7410 29314 7422
rect 29598 7474 29650 7486
rect 31614 7474 31666 7486
rect 32286 7474 32338 7486
rect 33406 7474 33458 7486
rect 29810 7422 29822 7474
rect 29874 7422 29886 7474
rect 31826 7422 31838 7474
rect 31890 7422 31902 7474
rect 32498 7422 32510 7474
rect 32562 7422 32574 7474
rect 29598 7410 29650 7422
rect 31614 7410 31666 7422
rect 32286 7410 32338 7422
rect 33406 7410 33458 7422
rect 33518 7474 33570 7486
rect 33518 7410 33570 7422
rect 4174 7362 4226 7374
rect 4174 7298 4226 7310
rect 13918 7362 13970 7374
rect 17390 7362 17442 7374
rect 23438 7362 23490 7374
rect 14242 7310 14254 7362
rect 14306 7310 14318 7362
rect 16594 7310 16606 7362
rect 16658 7310 16670 7362
rect 19506 7310 19518 7362
rect 19570 7310 19582 7362
rect 21634 7310 21646 7362
rect 21698 7310 21710 7362
rect 13918 7298 13970 7310
rect 17390 7298 17442 7310
rect 23438 7298 23490 7310
rect 25678 7362 25730 7374
rect 25678 7298 25730 7310
rect 28030 7362 28082 7374
rect 28030 7298 28082 7310
rect 3838 7250 3890 7262
rect 3838 7186 3890 7198
rect 3950 7250 4002 7262
rect 3950 7186 4002 7198
rect 8878 7250 8930 7262
rect 8878 7186 8930 7198
rect 12798 7250 12850 7262
rect 12798 7186 12850 7198
rect 26686 7250 26738 7262
rect 26686 7186 26738 7198
rect 27134 7250 27186 7262
rect 27134 7186 27186 7198
rect 27358 7250 27410 7262
rect 27358 7186 27410 7198
rect 31390 7250 31442 7262
rect 31390 7186 31442 7198
rect 32174 7250 32226 7262
rect 32174 7186 32226 7198
rect 33182 7250 33234 7262
rect 33182 7186 33234 7198
rect 1344 7082 34608 7116
rect 1344 7030 5372 7082
rect 5424 7030 5476 7082
rect 5528 7030 5580 7082
rect 5632 7030 13688 7082
rect 13740 7030 13792 7082
rect 13844 7030 13896 7082
rect 13948 7030 22004 7082
rect 22056 7030 22108 7082
rect 22160 7030 22212 7082
rect 22264 7030 30320 7082
rect 30372 7030 30424 7082
rect 30476 7030 30528 7082
rect 30580 7030 34608 7082
rect 1344 6996 34608 7030
rect 9998 6914 10050 6926
rect 9998 6850 10050 6862
rect 27134 6914 27186 6926
rect 27134 6850 27186 6862
rect 29374 6914 29426 6926
rect 29374 6850 29426 6862
rect 5742 6802 5794 6814
rect 18174 6802 18226 6814
rect 29150 6802 29202 6814
rect 30382 6802 30434 6814
rect 7746 6750 7758 6802
rect 7810 6750 7822 6802
rect 23762 6750 23774 6802
rect 23826 6750 23838 6802
rect 29698 6750 29710 6802
rect 29762 6750 29774 6802
rect 33954 6750 33966 6802
rect 34018 6750 34030 6802
rect 5742 6738 5794 6750
rect 18174 6738 18226 6750
rect 29150 6738 29202 6750
rect 30382 6738 30434 6750
rect 4958 6690 5010 6702
rect 4958 6626 5010 6638
rect 5630 6690 5682 6702
rect 5630 6626 5682 6638
rect 6414 6690 6466 6702
rect 10222 6690 10274 6702
rect 7634 6638 7646 6690
rect 7698 6638 7710 6690
rect 8642 6638 8654 6690
rect 8706 6638 8718 6690
rect 6414 6626 6466 6638
rect 10222 6626 10274 6638
rect 10894 6690 10946 6702
rect 10894 6626 10946 6638
rect 12910 6690 12962 6702
rect 12910 6626 12962 6638
rect 13358 6690 13410 6702
rect 22094 6690 22146 6702
rect 27246 6690 27298 6702
rect 14578 6638 14590 6690
rect 14642 6638 14654 6690
rect 15250 6638 15262 6690
rect 15314 6638 15326 6690
rect 21746 6638 21758 6690
rect 21810 6638 21822 6690
rect 22306 6638 22318 6690
rect 22370 6638 22382 6690
rect 23202 6638 23214 6690
rect 23266 6638 23278 6690
rect 26450 6638 26462 6690
rect 26514 6638 26526 6690
rect 13358 6626 13410 6638
rect 22094 6626 22146 6638
rect 27246 6626 27298 6638
rect 27470 6690 27522 6702
rect 30158 6690 30210 6702
rect 28130 6638 28142 6690
rect 28194 6638 28206 6690
rect 30706 6638 30718 6690
rect 30770 6638 30782 6690
rect 31042 6638 31054 6690
rect 31106 6638 31118 6690
rect 27470 6626 27522 6638
rect 30158 6626 30210 6638
rect 5070 6578 5122 6590
rect 5070 6514 5122 6526
rect 6078 6578 6130 6590
rect 6078 6514 6130 6526
rect 6638 6578 6690 6590
rect 6638 6514 6690 6526
rect 6750 6578 6802 6590
rect 22990 6578 23042 6590
rect 27582 6578 27634 6590
rect 7970 6526 7982 6578
rect 8034 6526 8046 6578
rect 10546 6526 10558 6578
rect 10610 6526 10622 6578
rect 11218 6526 11230 6578
rect 11282 6526 11294 6578
rect 12562 6526 12574 6578
rect 12626 6526 12638 6578
rect 13794 6526 13806 6578
rect 13858 6526 13870 6578
rect 14242 6526 14254 6578
rect 14306 6526 14318 6578
rect 16034 6526 16046 6578
rect 16098 6526 16110 6578
rect 19058 6526 19070 6578
rect 19122 6526 19134 6578
rect 24098 6526 24110 6578
rect 24162 6526 24174 6578
rect 24770 6526 24782 6578
rect 24834 6526 24846 6578
rect 31826 6526 31838 6578
rect 31890 6526 31902 6578
rect 6750 6514 6802 6526
rect 22990 6514 23042 6526
rect 27582 6514 27634 6526
rect 5854 6466 5906 6478
rect 5854 6402 5906 6414
rect 8878 6466 8930 6478
rect 11566 6466 11618 6478
rect 9650 6414 9662 6466
rect 9714 6414 9726 6466
rect 8878 6402 8930 6414
rect 11566 6402 11618 6414
rect 18734 6466 18786 6478
rect 27906 6414 27918 6466
rect 27970 6414 27982 6466
rect 18734 6402 18786 6414
rect 1344 6298 34768 6332
rect 1344 6246 9530 6298
rect 9582 6246 9634 6298
rect 9686 6246 9738 6298
rect 9790 6246 17846 6298
rect 17898 6246 17950 6298
rect 18002 6246 18054 6298
rect 18106 6246 26162 6298
rect 26214 6246 26266 6298
rect 26318 6246 26370 6298
rect 26422 6246 34478 6298
rect 34530 6246 34582 6298
rect 34634 6246 34686 6298
rect 34738 6246 34768 6298
rect 1344 6212 34768 6246
rect 7646 6130 7698 6142
rect 3042 6078 3054 6130
rect 3106 6078 3118 6130
rect 4610 6078 4622 6130
rect 4674 6078 4686 6130
rect 5506 6078 5518 6130
rect 5570 6078 5582 6130
rect 6178 6078 6190 6130
rect 6242 6078 6254 6130
rect 7186 6078 7198 6130
rect 7250 6078 7262 6130
rect 3502 6018 3554 6030
rect 3502 5954 3554 5966
rect 5854 6018 5906 6030
rect 5854 5954 5906 5966
rect 6750 6018 6802 6030
rect 6750 5954 6802 5966
rect 6862 6018 6914 6030
rect 6862 5954 6914 5966
rect 5182 5906 5234 5918
rect 2818 5854 2830 5906
rect 2882 5854 2894 5906
rect 4386 5854 4398 5906
rect 4450 5854 4462 5906
rect 5182 5842 5234 5854
rect 6526 5906 6578 5918
rect 6526 5842 6578 5854
rect 3390 5682 3442 5694
rect 7201 5682 7247 6078
rect 7646 6066 7698 6078
rect 7982 6130 8034 6142
rect 7982 6066 8034 6078
rect 8206 6130 8258 6142
rect 8206 6066 8258 6078
rect 13694 6130 13746 6142
rect 13694 6066 13746 6078
rect 20974 6130 21026 6142
rect 20974 6066 21026 6078
rect 33294 6130 33346 6142
rect 33294 6066 33346 6078
rect 7870 6018 7922 6030
rect 7870 5954 7922 5966
rect 8430 6018 8482 6030
rect 8430 5954 8482 5966
rect 12014 6018 12066 6030
rect 16606 6018 16658 6030
rect 12674 5966 12686 6018
rect 12738 5966 12750 6018
rect 13010 5966 13022 6018
rect 13074 5966 13086 6018
rect 12014 5954 12066 5966
rect 16606 5954 16658 5966
rect 21310 6018 21362 6030
rect 21310 5954 21362 5966
rect 22990 6018 23042 6030
rect 22990 5954 23042 5966
rect 25678 6018 25730 6030
rect 25678 5954 25730 5966
rect 26686 6018 26738 6030
rect 26686 5954 26738 5966
rect 28702 6018 28754 6030
rect 28702 5954 28754 5966
rect 29822 6018 29874 6030
rect 29822 5954 29874 5966
rect 30942 6018 30994 6030
rect 30942 5954 30994 5966
rect 14142 5906 14194 5918
rect 7410 5854 7422 5906
rect 7474 5854 7486 5906
rect 8642 5854 8654 5906
rect 8706 5854 8718 5906
rect 8866 5854 8878 5906
rect 8930 5854 8942 5906
rect 13234 5854 13246 5906
rect 13298 5854 13310 5906
rect 14142 5842 14194 5854
rect 14366 5906 14418 5918
rect 14366 5842 14418 5854
rect 15710 5906 15762 5918
rect 17390 5906 17442 5918
rect 19294 5906 19346 5918
rect 15922 5854 15934 5906
rect 15986 5854 15998 5906
rect 17826 5854 17838 5906
rect 17890 5854 17902 5906
rect 18834 5854 18846 5906
rect 18898 5854 18910 5906
rect 15710 5842 15762 5854
rect 17390 5842 17442 5854
rect 19294 5842 19346 5854
rect 21646 5906 21698 5918
rect 21646 5842 21698 5854
rect 21758 5906 21810 5918
rect 21758 5842 21810 5854
rect 22654 5906 22706 5918
rect 25566 5906 25618 5918
rect 26462 5906 26514 5918
rect 24434 5854 24446 5906
rect 24498 5854 24510 5906
rect 25330 5854 25342 5906
rect 25394 5854 25406 5906
rect 26114 5854 26126 5906
rect 26178 5854 26190 5906
rect 22654 5842 22706 5854
rect 25566 5842 25618 5854
rect 26462 5842 26514 5854
rect 27022 5906 27074 5918
rect 27022 5842 27074 5854
rect 27694 5906 27746 5918
rect 30606 5906 30658 5918
rect 29026 5854 29038 5906
rect 29090 5854 29102 5906
rect 30034 5854 30046 5906
rect 30098 5854 30110 5906
rect 27694 5842 27746 5854
rect 30606 5842 30658 5854
rect 31166 5906 31218 5918
rect 31950 5906 32002 5918
rect 31490 5854 31502 5906
rect 31554 5854 31566 5906
rect 31166 5842 31218 5854
rect 31950 5842 32002 5854
rect 33070 5906 33122 5918
rect 33618 5854 33630 5906
rect 33682 5854 33694 5906
rect 33070 5842 33122 5854
rect 14590 5794 14642 5806
rect 8978 5742 8990 5794
rect 9042 5742 9054 5794
rect 14590 5730 14642 5742
rect 18398 5794 18450 5806
rect 18398 5730 18450 5742
rect 21422 5794 21474 5806
rect 26910 5794 26962 5806
rect 22530 5742 22542 5794
rect 22594 5742 22606 5794
rect 24322 5742 24334 5794
rect 24386 5742 24398 5794
rect 21422 5730 21474 5742
rect 26910 5730 26962 5742
rect 27806 5794 27858 5806
rect 27806 5730 27858 5742
rect 30718 5794 30770 5806
rect 30718 5730 30770 5742
rect 31726 5794 31778 5806
rect 31726 5730 31778 5742
rect 33182 5794 33234 5806
rect 33182 5730 33234 5742
rect 27358 5682 27410 5694
rect 7186 5630 7198 5682
rect 7250 5630 7262 5682
rect 24098 5630 24110 5682
rect 24162 5630 24174 5682
rect 3390 5618 3442 5630
rect 27358 5618 27410 5630
rect 27470 5682 27522 5694
rect 27470 5618 27522 5630
rect 29038 5682 29090 5694
rect 29038 5618 29090 5630
rect 32062 5682 32114 5694
rect 32062 5618 32114 5630
rect 1344 5514 34608 5548
rect 1344 5462 5372 5514
rect 5424 5462 5476 5514
rect 5528 5462 5580 5514
rect 5632 5462 13688 5514
rect 13740 5462 13792 5514
rect 13844 5462 13896 5514
rect 13948 5462 22004 5514
rect 22056 5462 22108 5514
rect 22160 5462 22212 5514
rect 22264 5462 30320 5514
rect 30372 5462 30424 5514
rect 30476 5462 30528 5514
rect 30580 5462 34608 5514
rect 1344 5428 34608 5462
rect 13582 5346 13634 5358
rect 3938 5294 3950 5346
rect 4002 5294 4014 5346
rect 4498 5294 4510 5346
rect 4562 5294 4574 5346
rect 13582 5282 13634 5294
rect 21982 5346 22034 5358
rect 21982 5282 22034 5294
rect 27358 5346 27410 5358
rect 27358 5282 27410 5294
rect 27694 5346 27746 5358
rect 27694 5282 27746 5294
rect 29262 5346 29314 5358
rect 29262 5282 29314 5294
rect 3390 5234 3442 5246
rect 3390 5170 3442 5182
rect 10782 5234 10834 5246
rect 10782 5170 10834 5182
rect 10894 5234 10946 5246
rect 19182 5234 19234 5246
rect 12114 5182 12126 5234
rect 12178 5182 12190 5234
rect 10894 5170 10946 5182
rect 19182 5170 19234 5182
rect 21646 5234 21698 5246
rect 30494 5234 30546 5246
rect 24098 5182 24110 5234
rect 24162 5182 24174 5234
rect 26226 5182 26238 5234
rect 26290 5182 26302 5234
rect 32050 5182 32062 5234
rect 32114 5182 32126 5234
rect 34178 5182 34190 5234
rect 34242 5182 34254 5234
rect 21646 5170 21698 5182
rect 30494 5170 30546 5182
rect 2718 5122 2770 5134
rect 2146 5070 2158 5122
rect 2210 5070 2222 5122
rect 2718 5058 2770 5070
rect 3614 5122 3666 5134
rect 10110 5122 10162 5134
rect 4274 5070 4286 5122
rect 4338 5070 4350 5122
rect 4834 5070 4846 5122
rect 4898 5070 4910 5122
rect 5954 5070 5966 5122
rect 6018 5070 6030 5122
rect 7410 5070 7422 5122
rect 7474 5070 7486 5122
rect 8082 5070 8094 5122
rect 8146 5070 8158 5122
rect 8866 5070 8878 5122
rect 8930 5070 8942 5122
rect 9090 5070 9102 5122
rect 9154 5070 9166 5122
rect 3614 5058 3666 5070
rect 10110 5058 10162 5070
rect 11230 5122 11282 5134
rect 11230 5058 11282 5070
rect 11790 5122 11842 5134
rect 13470 5122 13522 5134
rect 21870 5122 21922 5134
rect 12786 5070 12798 5122
rect 12850 5070 12862 5122
rect 13906 5070 13918 5122
rect 13970 5070 13982 5122
rect 15922 5070 15934 5122
rect 15986 5070 15998 5122
rect 18162 5070 18174 5122
rect 18226 5070 18238 5122
rect 11790 5058 11842 5070
rect 13470 5058 13522 5070
rect 21870 5058 21922 5070
rect 22766 5122 22818 5134
rect 22766 5058 22818 5070
rect 23326 5122 23378 5134
rect 29486 5122 29538 5134
rect 30270 5122 30322 5134
rect 27010 5070 27022 5122
rect 27074 5070 27086 5122
rect 27346 5070 27358 5122
rect 27410 5070 27422 5122
rect 29698 5070 29710 5122
rect 29762 5070 29774 5122
rect 23326 5058 23378 5070
rect 29486 5058 29538 5070
rect 30270 5058 30322 5070
rect 30718 5122 30770 5134
rect 30718 5058 30770 5070
rect 30942 5122 30994 5134
rect 31266 5070 31278 5122
rect 31330 5070 31342 5122
rect 30942 5058 30994 5070
rect 2382 5010 2434 5022
rect 5070 5010 5122 5022
rect 21534 5010 21586 5022
rect 3042 4958 3054 5010
rect 3106 4958 3118 5010
rect 7186 4958 7198 5010
rect 7250 4958 7262 5010
rect 7858 4958 7870 5010
rect 7922 4958 7934 5010
rect 9426 4958 9438 5010
rect 9490 4958 9502 5010
rect 9650 4958 9662 5010
rect 9714 4958 9726 5010
rect 12674 4958 12686 5010
rect 12738 4958 12750 5010
rect 14018 4958 14030 5010
rect 14082 4958 14094 5010
rect 17714 4958 17726 5010
rect 17778 4958 17790 5010
rect 2382 4946 2434 4958
rect 5070 4946 5122 4958
rect 21534 4946 21586 4958
rect 4286 4898 4338 4910
rect 4286 4834 4338 4846
rect 6190 4898 6242 4910
rect 29598 4898 29650 4910
rect 6290 4846 6302 4898
rect 6354 4846 6366 4898
rect 14130 4846 14142 4898
rect 14194 4846 14206 4898
rect 6190 4834 6242 4846
rect 29598 4834 29650 4846
rect 1344 4730 34768 4764
rect 1344 4678 9530 4730
rect 9582 4678 9634 4730
rect 9686 4678 9738 4730
rect 9790 4678 17846 4730
rect 17898 4678 17950 4730
rect 18002 4678 18054 4730
rect 18106 4678 26162 4730
rect 26214 4678 26266 4730
rect 26318 4678 26370 4730
rect 26422 4678 34478 4730
rect 34530 4678 34582 4730
rect 34634 4678 34686 4730
rect 34738 4678 34768 4730
rect 1344 4644 34768 4678
rect 6414 4562 6466 4574
rect 4722 4510 4734 4562
rect 4786 4510 4798 4562
rect 6066 4510 6078 4562
rect 6130 4510 6142 4562
rect 6414 4498 6466 4510
rect 7086 4562 7138 4574
rect 7086 4498 7138 4510
rect 7534 4562 7586 4574
rect 7534 4498 7586 4510
rect 7758 4562 7810 4574
rect 17502 4562 17554 4574
rect 11330 4510 11342 4562
rect 11394 4510 11406 4562
rect 11890 4510 11902 4562
rect 11954 4510 11966 4562
rect 7758 4498 7810 4510
rect 17502 4498 17554 4510
rect 18622 4562 18674 4574
rect 22754 4510 22766 4562
rect 22818 4510 22830 4562
rect 33058 4510 33070 4562
rect 33122 4510 33134 4562
rect 18622 4498 18674 4510
rect 5182 4450 5234 4462
rect 2482 4398 2494 4450
rect 2546 4398 2558 4450
rect 5182 4386 5234 4398
rect 5630 4450 5682 4462
rect 5630 4386 5682 4398
rect 6862 4450 6914 4462
rect 6862 4386 6914 4398
rect 7422 4450 7474 4462
rect 8654 4450 8706 4462
rect 16046 4450 16098 4462
rect 8306 4398 8318 4450
rect 8370 4398 8382 4450
rect 8978 4398 8990 4450
rect 9042 4398 9054 4450
rect 9538 4398 9550 4450
rect 9602 4398 9614 4450
rect 13346 4398 13358 4450
rect 13410 4398 13422 4450
rect 7422 4386 7474 4398
rect 8654 4386 8706 4398
rect 16046 4386 16098 4398
rect 18846 4450 18898 4462
rect 27906 4398 27918 4450
rect 27970 4398 27982 4450
rect 31154 4398 31166 4450
rect 31218 4398 31230 4450
rect 18846 4386 18898 4398
rect 5518 4338 5570 4350
rect 1810 4286 1822 4338
rect 1874 4286 1886 4338
rect 5518 4274 5570 4286
rect 5742 4338 5794 4350
rect 5742 4274 5794 4286
rect 6750 4338 6802 4350
rect 11006 4338 11058 4350
rect 16158 4338 16210 4350
rect 8082 4286 8094 4338
rect 8146 4286 8158 4338
rect 9762 4286 9774 4338
rect 9826 4286 9838 4338
rect 12114 4286 12126 4338
rect 12178 4286 12190 4338
rect 12562 4286 12574 4338
rect 12626 4286 12638 4338
rect 6750 4274 6802 4286
rect 11006 4274 11058 4286
rect 16158 4274 16210 4286
rect 16382 4338 16434 4350
rect 23102 4338 23154 4350
rect 16594 4286 16606 4338
rect 16658 4286 16670 4338
rect 19170 4286 19182 4338
rect 19234 4286 19246 4338
rect 19618 4286 19630 4338
rect 19682 4286 19694 4338
rect 16382 4274 16434 4286
rect 23102 4274 23154 4286
rect 23774 4338 23826 4350
rect 33406 4338 33458 4350
rect 24210 4286 24222 4338
rect 24274 4286 24286 4338
rect 28578 4286 28590 4338
rect 28642 4286 28654 4338
rect 31938 4286 31950 4338
rect 32002 4286 32014 4338
rect 23774 4274 23826 4286
rect 33406 4274 33458 4286
rect 33630 4338 33682 4350
rect 33630 4274 33682 4286
rect 10782 4226 10834 4238
rect 23326 4226 23378 4238
rect 15474 4174 15486 4226
rect 15538 4174 15550 4226
rect 19058 4174 19070 4226
rect 19122 4174 19134 4226
rect 20290 4174 20302 4226
rect 20354 4174 20366 4226
rect 22418 4174 22430 4226
rect 22482 4174 22494 4226
rect 10782 4162 10834 4174
rect 23326 4162 23378 4174
rect 23662 4226 23714 4238
rect 25778 4174 25790 4226
rect 25842 4174 25854 4226
rect 29026 4174 29038 4226
rect 29090 4174 29102 4226
rect 23662 4162 23714 4174
rect 23998 4114 24050 4126
rect 23998 4050 24050 4062
rect 1344 3946 34608 3980
rect 1344 3894 5372 3946
rect 5424 3894 5476 3946
rect 5528 3894 5580 3946
rect 5632 3894 13688 3946
rect 13740 3894 13792 3946
rect 13844 3894 13896 3946
rect 13948 3894 22004 3946
rect 22056 3894 22108 3946
rect 22160 3894 22212 3946
rect 22264 3894 30320 3946
rect 30372 3894 30424 3946
rect 30476 3894 30528 3946
rect 30580 3894 34608 3946
rect 1344 3860 34608 3894
rect 6638 3778 6690 3790
rect 6638 3714 6690 3726
rect 8206 3778 8258 3790
rect 8206 3714 8258 3726
rect 14926 3778 14978 3790
rect 14926 3714 14978 3726
rect 15262 3778 15314 3790
rect 15262 3714 15314 3726
rect 5742 3666 5794 3678
rect 5742 3602 5794 3614
rect 8318 3666 8370 3678
rect 15486 3666 15538 3678
rect 24558 3666 24610 3678
rect 10210 3614 10222 3666
rect 10274 3614 10286 3666
rect 12450 3614 12462 3666
rect 12514 3614 12526 3666
rect 16930 3614 16942 3666
rect 16994 3614 17006 3666
rect 19058 3614 19070 3666
rect 19122 3614 19134 3666
rect 21522 3614 21534 3666
rect 21586 3614 21598 3666
rect 23650 3614 23662 3666
rect 23714 3614 23726 3666
rect 8318 3602 8370 3614
rect 15486 3602 15538 3614
rect 24558 3602 24610 3614
rect 24670 3666 24722 3678
rect 24670 3602 24722 3614
rect 32958 3666 33010 3678
rect 32958 3602 33010 3614
rect 6526 3554 6578 3566
rect 9538 3502 9550 3554
rect 9602 3502 9614 3554
rect 19730 3502 19742 3554
rect 19794 3502 19806 3554
rect 20738 3502 20750 3554
rect 20802 3502 20814 3554
rect 24882 3502 24894 3554
rect 24946 3502 24958 3554
rect 25218 3502 25230 3554
rect 25282 3502 25294 3554
rect 31602 3502 31614 3554
rect 31666 3502 31678 3554
rect 32386 3502 32398 3554
rect 32450 3502 32462 3554
rect 6526 3490 6578 3502
rect 32174 3442 32226 3454
rect 26898 3390 26910 3442
rect 26962 3390 26974 3442
rect 30034 3390 30046 3442
rect 30098 3390 30110 3442
rect 32174 3378 32226 3390
rect 1344 3162 34768 3196
rect 1344 3110 9530 3162
rect 9582 3110 9634 3162
rect 9686 3110 9738 3162
rect 9790 3110 17846 3162
rect 17898 3110 17950 3162
rect 18002 3110 18054 3162
rect 18106 3110 26162 3162
rect 26214 3110 26266 3162
rect 26318 3110 26370 3162
rect 26422 3110 34478 3162
rect 34530 3110 34582 3162
rect 34634 3110 34686 3162
rect 34738 3110 34768 3162
rect 1344 3076 34768 3110
<< via1 >>
rect 5372 32118 5424 32170
rect 5476 32118 5528 32170
rect 5580 32118 5632 32170
rect 13688 32118 13740 32170
rect 13792 32118 13844 32170
rect 13896 32118 13948 32170
rect 22004 32118 22056 32170
rect 22108 32118 22160 32170
rect 22212 32118 22264 32170
rect 30320 32118 30372 32170
rect 30424 32118 30476 32170
rect 30528 32118 30580 32170
rect 9530 31334 9582 31386
rect 9634 31334 9686 31386
rect 9738 31334 9790 31386
rect 17846 31334 17898 31386
rect 17950 31334 18002 31386
rect 18054 31334 18106 31386
rect 26162 31334 26214 31386
rect 26266 31334 26318 31386
rect 26370 31334 26422 31386
rect 34478 31334 34530 31386
rect 34582 31334 34634 31386
rect 34686 31334 34738 31386
rect 5372 30550 5424 30602
rect 5476 30550 5528 30602
rect 5580 30550 5632 30602
rect 13688 30550 13740 30602
rect 13792 30550 13844 30602
rect 13896 30550 13948 30602
rect 22004 30550 22056 30602
rect 22108 30550 22160 30602
rect 22212 30550 22264 30602
rect 30320 30550 30372 30602
rect 30424 30550 30476 30602
rect 30528 30550 30580 30602
rect 9530 29766 9582 29818
rect 9634 29766 9686 29818
rect 9738 29766 9790 29818
rect 17846 29766 17898 29818
rect 17950 29766 18002 29818
rect 18054 29766 18106 29818
rect 26162 29766 26214 29818
rect 26266 29766 26318 29818
rect 26370 29766 26422 29818
rect 34478 29766 34530 29818
rect 34582 29766 34634 29818
rect 34686 29766 34738 29818
rect 5372 28982 5424 29034
rect 5476 28982 5528 29034
rect 5580 28982 5632 29034
rect 13688 28982 13740 29034
rect 13792 28982 13844 29034
rect 13896 28982 13948 29034
rect 22004 28982 22056 29034
rect 22108 28982 22160 29034
rect 22212 28982 22264 29034
rect 30320 28982 30372 29034
rect 30424 28982 30476 29034
rect 30528 28982 30580 29034
rect 11230 28702 11282 28754
rect 8430 28590 8482 28642
rect 9102 28478 9154 28530
rect 9530 28198 9582 28250
rect 9634 28198 9686 28250
rect 9738 28198 9790 28250
rect 17846 28198 17898 28250
rect 17950 28198 18002 28250
rect 18054 28198 18106 28250
rect 26162 28198 26214 28250
rect 26266 28198 26318 28250
rect 26370 28198 26422 28250
rect 34478 28198 34530 28250
rect 34582 28198 34634 28250
rect 34686 28198 34738 28250
rect 5070 27918 5122 27970
rect 4286 27806 4338 27858
rect 4510 27806 4562 27858
rect 4846 27806 4898 27858
rect 5182 27806 5234 27858
rect 10222 27806 10274 27858
rect 20078 27806 20130 27858
rect 20302 27806 20354 27858
rect 20638 27806 20690 27858
rect 3614 27694 3666 27746
rect 11006 27694 11058 27746
rect 13134 27694 13186 27746
rect 20526 27694 20578 27746
rect 5372 27414 5424 27466
rect 5476 27414 5528 27466
rect 5580 27414 5632 27466
rect 13688 27414 13740 27466
rect 13792 27414 13844 27466
rect 13896 27414 13948 27466
rect 22004 27414 22056 27466
rect 22108 27414 22160 27466
rect 22212 27414 22264 27466
rect 30320 27414 30372 27466
rect 30424 27414 30476 27466
rect 30528 27414 30580 27466
rect 5854 27246 5906 27298
rect 4622 27134 4674 27186
rect 4958 27134 5010 27186
rect 10222 27134 10274 27186
rect 12238 27134 12290 27186
rect 17054 27134 17106 27186
rect 20302 27134 20354 27186
rect 1822 27022 1874 27074
rect 5966 27022 6018 27074
rect 6190 27022 6242 27074
rect 6750 27022 6802 27074
rect 7422 27022 7474 27074
rect 12014 27022 12066 27074
rect 14254 27022 14306 27074
rect 17502 27022 17554 27074
rect 2494 26910 2546 26962
rect 5070 26910 5122 26962
rect 6302 26910 6354 26962
rect 6638 26910 6690 26962
rect 6862 26910 6914 26962
rect 8094 26910 8146 26962
rect 12462 26910 12514 26962
rect 12686 26910 12738 26962
rect 14926 26910 14978 26962
rect 18174 26910 18226 26962
rect 20638 26910 20690 26962
rect 20750 26910 20802 26962
rect 9530 26630 9582 26682
rect 9634 26630 9686 26682
rect 9738 26630 9790 26682
rect 17846 26630 17898 26682
rect 17950 26630 18002 26682
rect 18054 26630 18106 26682
rect 26162 26630 26214 26682
rect 26266 26630 26318 26682
rect 26370 26630 26422 26682
rect 34478 26630 34530 26682
rect 34582 26630 34634 26682
rect 34686 26630 34738 26682
rect 9886 26462 9938 26514
rect 16382 26462 16434 26514
rect 18174 26462 18226 26514
rect 18958 26462 19010 26514
rect 7310 26350 7362 26402
rect 18286 26350 18338 26402
rect 18510 26350 18562 26402
rect 19070 26350 19122 26402
rect 20526 26350 20578 26402
rect 25230 26350 25282 26402
rect 1822 26238 1874 26290
rect 7982 26238 8034 26290
rect 11790 26238 11842 26290
rect 12350 26238 12402 26290
rect 13134 26238 13186 26290
rect 16270 26238 16322 26290
rect 16494 26238 16546 26290
rect 16942 26238 16994 26290
rect 17838 26238 17890 26290
rect 18846 26238 18898 26290
rect 19518 26238 19570 26290
rect 19742 26238 19794 26290
rect 22990 26238 23042 26290
rect 23214 26238 23266 26290
rect 23326 26238 23378 26290
rect 25566 26238 25618 26290
rect 25678 26238 25730 26290
rect 2494 26126 2546 26178
rect 4622 26126 4674 26178
rect 5182 26126 5234 26178
rect 9998 26126 10050 26178
rect 12462 26126 12514 26178
rect 13806 26126 13858 26178
rect 15934 26126 15986 26178
rect 22654 26126 22706 26178
rect 25342 26126 25394 26178
rect 23774 26014 23826 26066
rect 5372 25846 5424 25898
rect 5476 25846 5528 25898
rect 5580 25846 5632 25898
rect 13688 25846 13740 25898
rect 13792 25846 13844 25898
rect 13896 25846 13948 25898
rect 22004 25846 22056 25898
rect 22108 25846 22160 25898
rect 22212 25846 22264 25898
rect 30320 25846 30372 25898
rect 30424 25846 30476 25898
rect 30528 25846 30580 25898
rect 2606 25678 2658 25730
rect 2942 25678 2994 25730
rect 3278 25678 3330 25730
rect 18958 25678 19010 25730
rect 4958 25566 5010 25618
rect 9886 25566 9938 25618
rect 12462 25566 12514 25618
rect 13582 25566 13634 25618
rect 14478 25566 14530 25618
rect 15374 25566 15426 25618
rect 19966 25566 20018 25618
rect 23102 25566 23154 25618
rect 25230 25566 25282 25618
rect 27358 25566 27410 25618
rect 2606 25454 2658 25506
rect 3278 25454 3330 25506
rect 4622 25454 4674 25506
rect 7086 25454 7138 25506
rect 12574 25454 12626 25506
rect 13694 25454 13746 25506
rect 14142 25454 14194 25506
rect 14254 25454 14306 25506
rect 14702 25454 14754 25506
rect 15150 25454 15202 25506
rect 15486 25454 15538 25506
rect 15822 25454 15874 25506
rect 16158 25454 16210 25506
rect 19294 25454 19346 25506
rect 19854 25454 19906 25506
rect 20078 25454 20130 25506
rect 20526 25454 20578 25506
rect 21646 25454 21698 25506
rect 22542 25454 22594 25506
rect 26014 25454 26066 25506
rect 26350 25454 26402 25506
rect 3614 25342 3666 25394
rect 4062 25342 4114 25394
rect 7758 25342 7810 25394
rect 14926 25342 14978 25394
rect 16270 25342 16322 25394
rect 19518 25342 19570 25394
rect 22766 25342 22818 25394
rect 26686 25342 26738 25394
rect 27022 25342 27074 25394
rect 12126 25230 12178 25282
rect 12350 25230 12402 25282
rect 13470 25230 13522 25282
rect 16382 25230 16434 25282
rect 16606 25230 16658 25282
rect 21870 25230 21922 25282
rect 27246 25230 27298 25282
rect 9530 25062 9582 25114
rect 9634 25062 9686 25114
rect 9738 25062 9790 25114
rect 17846 25062 17898 25114
rect 17950 25062 18002 25114
rect 18054 25062 18106 25114
rect 26162 25062 26214 25114
rect 26266 25062 26318 25114
rect 26370 25062 26422 25114
rect 34478 25062 34530 25114
rect 34582 25062 34634 25114
rect 34686 25062 34738 25114
rect 4734 24894 4786 24946
rect 6302 24894 6354 24946
rect 8878 24894 8930 24946
rect 11006 24894 11058 24946
rect 11118 24894 11170 24946
rect 11230 24894 11282 24946
rect 15150 24894 15202 24946
rect 18846 24894 18898 24946
rect 23662 24894 23714 24946
rect 25678 24894 25730 24946
rect 25790 24894 25842 24946
rect 4062 24782 4114 24834
rect 5854 24782 5906 24834
rect 6414 24782 6466 24834
rect 12350 24782 12402 24834
rect 13246 24782 13298 24834
rect 15710 24782 15762 24834
rect 18174 24782 18226 24834
rect 28478 24782 28530 24834
rect 4398 24670 4450 24722
rect 5070 24670 5122 24722
rect 5294 24670 5346 24722
rect 5630 24670 5682 24722
rect 11454 24670 11506 24722
rect 11678 24670 11730 24722
rect 12238 24670 12290 24722
rect 12574 24670 12626 24722
rect 12686 24670 12738 24722
rect 14590 24670 14642 24722
rect 15038 24670 15090 24722
rect 15262 24670 15314 24722
rect 18510 24670 18562 24722
rect 19070 24670 19122 24722
rect 20190 24670 20242 24722
rect 20862 24670 20914 24722
rect 22878 24670 22930 24722
rect 22990 24670 23042 24722
rect 23886 24670 23938 24722
rect 24334 24670 24386 24722
rect 24446 24670 24498 24722
rect 24558 24670 24610 24722
rect 25118 24670 25170 24722
rect 25566 24670 25618 24722
rect 29262 24670 29314 24722
rect 8990 24558 9042 24610
rect 12462 24558 12514 24610
rect 13358 24558 13410 24610
rect 13470 24558 13522 24610
rect 14142 24558 14194 24610
rect 20414 24558 20466 24610
rect 26350 24558 26402 24610
rect 15598 24446 15650 24498
rect 5372 24278 5424 24330
rect 5476 24278 5528 24330
rect 5580 24278 5632 24330
rect 13688 24278 13740 24330
rect 13792 24278 13844 24330
rect 13896 24278 13948 24330
rect 22004 24278 22056 24330
rect 22108 24278 22160 24330
rect 22212 24278 22264 24330
rect 30320 24278 30372 24330
rect 30424 24278 30476 24330
rect 30528 24278 30580 24330
rect 12126 24110 12178 24162
rect 13582 24110 13634 24162
rect 9998 23998 10050 24050
rect 11006 23998 11058 24050
rect 15038 23998 15090 24050
rect 20302 23998 20354 24050
rect 26238 23998 26290 24050
rect 27022 23998 27074 24050
rect 7086 23886 7138 23938
rect 10894 23886 10946 23938
rect 11678 23886 11730 23938
rect 13470 23886 13522 23938
rect 14142 23886 14194 23938
rect 17950 23886 18002 23938
rect 19182 23886 19234 23938
rect 26126 23886 26178 23938
rect 5070 23774 5122 23826
rect 7870 23774 7922 23826
rect 11118 23774 11170 23826
rect 11230 23774 11282 23826
rect 12014 23774 12066 23826
rect 14478 23774 14530 23826
rect 17166 23774 17218 23826
rect 18846 23774 18898 23826
rect 26686 23774 26738 23826
rect 4846 23662 4898 23714
rect 4958 23662 5010 23714
rect 12126 23662 12178 23714
rect 13022 23662 13074 23714
rect 13694 23662 13746 23714
rect 13918 23662 13970 23714
rect 14590 23662 14642 23714
rect 14814 23662 14866 23714
rect 18510 23662 18562 23714
rect 18958 23662 19010 23714
rect 19518 23662 19570 23714
rect 19854 23662 19906 23714
rect 25902 23662 25954 23714
rect 26350 23662 26402 23714
rect 26910 23662 26962 23714
rect 9530 23494 9582 23546
rect 9634 23494 9686 23546
rect 9738 23494 9790 23546
rect 17846 23494 17898 23546
rect 17950 23494 18002 23546
rect 18054 23494 18106 23546
rect 26162 23494 26214 23546
rect 26266 23494 26318 23546
rect 26370 23494 26422 23546
rect 34478 23494 34530 23546
rect 34582 23494 34634 23546
rect 34686 23494 34738 23546
rect 5854 23326 5906 23378
rect 8430 23326 8482 23378
rect 8878 23326 8930 23378
rect 9998 23326 10050 23378
rect 11006 23326 11058 23378
rect 12910 23326 12962 23378
rect 14142 23326 14194 23378
rect 15934 23326 15986 23378
rect 17390 23326 17442 23378
rect 18846 23326 18898 23378
rect 19070 23326 19122 23378
rect 25790 23326 25842 23378
rect 9886 23214 9938 23266
rect 10222 23214 10274 23266
rect 10894 23214 10946 23266
rect 11790 23214 11842 23266
rect 12686 23214 12738 23266
rect 13694 23214 13746 23266
rect 13806 23214 13858 23266
rect 14814 23214 14866 23266
rect 15822 23214 15874 23266
rect 18622 23214 18674 23266
rect 20302 23214 20354 23266
rect 22766 23214 22818 23266
rect 23102 23214 23154 23266
rect 24670 23214 24722 23266
rect 29150 23214 29202 23266
rect 2046 23102 2098 23154
rect 5518 23102 5570 23154
rect 6190 23102 6242 23154
rect 6414 23102 6466 23154
rect 6638 23102 6690 23154
rect 10334 23102 10386 23154
rect 10670 23102 10722 23154
rect 11342 23102 11394 23154
rect 11678 23102 11730 23154
rect 12126 23102 12178 23154
rect 12462 23102 12514 23154
rect 13470 23102 13522 23154
rect 14478 23102 14530 23154
rect 15038 23102 15090 23154
rect 15374 23102 15426 23154
rect 16046 23102 16098 23154
rect 18398 23102 18450 23154
rect 19182 23102 19234 23154
rect 19518 23102 19570 23154
rect 24446 23102 24498 23154
rect 25230 23102 25282 23154
rect 26126 23102 26178 23154
rect 26462 23102 26514 23154
rect 26686 23102 26738 23154
rect 29822 23102 29874 23154
rect 2830 22990 2882 23042
rect 4958 22990 5010 23042
rect 5294 22990 5346 23042
rect 6750 22990 6802 23042
rect 8542 22990 8594 23042
rect 8990 22990 9042 23042
rect 12574 22990 12626 23042
rect 17726 22990 17778 23042
rect 17950 22990 18002 23042
rect 22430 22990 22482 23042
rect 27022 22990 27074 23042
rect 11454 22878 11506 22930
rect 25454 22878 25506 22930
rect 5372 22710 5424 22762
rect 5476 22710 5528 22762
rect 5580 22710 5632 22762
rect 13688 22710 13740 22762
rect 13792 22710 13844 22762
rect 13896 22710 13948 22762
rect 22004 22710 22056 22762
rect 22108 22710 22160 22762
rect 22212 22710 22264 22762
rect 30320 22710 30372 22762
rect 30424 22710 30476 22762
rect 30528 22710 30580 22762
rect 5742 22542 5794 22594
rect 5966 22542 6018 22594
rect 19294 22542 19346 22594
rect 4622 22430 4674 22482
rect 7870 22430 7922 22482
rect 19406 22430 19458 22482
rect 24222 22430 24274 22482
rect 25342 22430 25394 22482
rect 1822 22318 1874 22370
rect 6078 22318 6130 22370
rect 12910 22318 12962 22370
rect 15038 22318 15090 22370
rect 19630 22318 19682 22370
rect 19966 22318 20018 22370
rect 20302 22318 20354 22370
rect 21310 22318 21362 22370
rect 25230 22318 25282 22370
rect 26126 22318 26178 22370
rect 26350 22318 26402 22370
rect 26910 22318 26962 22370
rect 2494 22206 2546 22258
rect 5630 22206 5682 22258
rect 18622 22206 18674 22258
rect 20526 22206 20578 22258
rect 20638 22206 20690 22258
rect 20750 22206 20802 22258
rect 22094 22206 22146 22258
rect 27022 22206 27074 22258
rect 27470 22206 27522 22258
rect 25454 22094 25506 22146
rect 25678 22094 25730 22146
rect 26574 22094 26626 22146
rect 26686 22094 26738 22146
rect 27246 22094 27298 22146
rect 27582 22094 27634 22146
rect 9530 21926 9582 21978
rect 9634 21926 9686 21978
rect 9738 21926 9790 21978
rect 17846 21926 17898 21978
rect 17950 21926 18002 21978
rect 18054 21926 18106 21978
rect 26162 21926 26214 21978
rect 26266 21926 26318 21978
rect 26370 21926 26422 21978
rect 34478 21926 34530 21978
rect 34582 21926 34634 21978
rect 34686 21926 34738 21978
rect 3614 21758 3666 21810
rect 5518 21758 5570 21810
rect 12686 21758 12738 21810
rect 13582 21758 13634 21810
rect 13694 21758 13746 21810
rect 13806 21758 13858 21810
rect 14702 21758 14754 21810
rect 14926 21758 14978 21810
rect 15710 21758 15762 21810
rect 16830 21758 16882 21810
rect 17950 21758 18002 21810
rect 19406 21758 19458 21810
rect 19966 21758 20018 21810
rect 21086 21758 21138 21810
rect 23662 21758 23714 21810
rect 3950 21646 4002 21698
rect 4622 21646 4674 21698
rect 5406 21646 5458 21698
rect 10782 21646 10834 21698
rect 11342 21646 11394 21698
rect 12350 21646 12402 21698
rect 13470 21646 13522 21698
rect 14814 21646 14866 21698
rect 16494 21646 16546 21698
rect 19294 21646 19346 21698
rect 20638 21646 20690 21698
rect 20862 21646 20914 21698
rect 21758 21646 21810 21698
rect 22542 21646 22594 21698
rect 24222 21646 24274 21698
rect 26126 21646 26178 21698
rect 26238 21646 26290 21698
rect 3390 21534 3442 21586
rect 3614 21534 3666 21586
rect 4398 21534 4450 21586
rect 4510 21534 4562 21586
rect 5742 21534 5794 21586
rect 10670 21534 10722 21586
rect 11566 21534 11618 21586
rect 11902 21534 11954 21586
rect 13022 21534 13074 21586
rect 14142 21534 14194 21586
rect 14478 21534 14530 21586
rect 15150 21534 15202 21586
rect 15486 21534 15538 21586
rect 18174 21534 18226 21586
rect 20302 21534 20354 21586
rect 21310 21534 21362 21586
rect 21870 21534 21922 21586
rect 22094 21534 22146 21586
rect 22430 21534 22482 21586
rect 24110 21534 24162 21586
rect 24446 21534 24498 21586
rect 29486 21534 29538 21586
rect 5070 21422 5122 21474
rect 11678 21422 11730 21474
rect 15374 21422 15426 21474
rect 17614 21422 17666 21474
rect 18958 21422 19010 21474
rect 20750 21422 20802 21474
rect 24670 21422 24722 21474
rect 26574 21422 26626 21474
rect 28702 21422 28754 21474
rect 10782 21310 10834 21362
rect 19406 21310 19458 21362
rect 26126 21310 26178 21362
rect 5372 21142 5424 21194
rect 5476 21142 5528 21194
rect 5580 21142 5632 21194
rect 13688 21142 13740 21194
rect 13792 21142 13844 21194
rect 13896 21142 13948 21194
rect 22004 21142 22056 21194
rect 22108 21142 22160 21194
rect 22212 21142 22264 21194
rect 30320 21142 30372 21194
rect 30424 21142 30476 21194
rect 30528 21142 30580 21194
rect 2606 20974 2658 21026
rect 11454 20974 11506 21026
rect 12686 20974 12738 21026
rect 11006 20862 11058 20914
rect 15822 20862 15874 20914
rect 25902 20862 25954 20914
rect 28030 20862 28082 20914
rect 3278 20750 3330 20802
rect 4958 20750 5010 20802
rect 5630 20750 5682 20802
rect 7646 20750 7698 20802
rect 12574 20750 12626 20802
rect 13806 20750 13858 20802
rect 14142 20750 14194 20802
rect 16046 20750 16098 20802
rect 16942 20750 16994 20802
rect 23102 20750 23154 20802
rect 26462 20750 26514 20802
rect 26686 20750 26738 20802
rect 27582 20750 27634 20802
rect 27806 20750 27858 20802
rect 3950 20638 4002 20690
rect 5742 20638 5794 20690
rect 8206 20638 8258 20690
rect 10558 20638 10610 20690
rect 10782 20638 10834 20690
rect 11342 20638 11394 20690
rect 11454 20638 11506 20690
rect 12686 20638 12738 20690
rect 13470 20638 13522 20690
rect 14366 20638 14418 20690
rect 16718 20638 16770 20690
rect 17390 20638 17442 20690
rect 17726 20638 17778 20690
rect 23774 20638 23826 20690
rect 26238 20638 26290 20690
rect 28142 20638 28194 20690
rect 2382 20526 2434 20578
rect 2494 20526 2546 20578
rect 2942 20526 2994 20578
rect 3614 20526 3666 20578
rect 4286 20526 4338 20578
rect 4398 20526 4450 20578
rect 4510 20526 4562 20578
rect 7758 20526 7810 20578
rect 10222 20526 10274 20578
rect 10446 20526 10498 20578
rect 13582 20526 13634 20578
rect 16382 20526 16434 20578
rect 18062 20526 18114 20578
rect 18398 20526 18450 20578
rect 9530 20358 9582 20410
rect 9634 20358 9686 20410
rect 9738 20358 9790 20410
rect 17846 20358 17898 20410
rect 17950 20358 18002 20410
rect 18054 20358 18106 20410
rect 26162 20358 26214 20410
rect 26266 20358 26318 20410
rect 26370 20358 26422 20410
rect 34478 20358 34530 20410
rect 34582 20358 34634 20410
rect 34686 20358 34738 20410
rect 5070 20078 5122 20130
rect 8206 20078 8258 20130
rect 8878 20078 8930 20130
rect 12014 20078 12066 20130
rect 12574 20078 12626 20130
rect 14254 20078 14306 20130
rect 14926 20078 14978 20130
rect 15262 20078 15314 20130
rect 16830 20078 16882 20130
rect 1822 19966 1874 20018
rect 5294 19966 5346 20018
rect 5518 19966 5570 20018
rect 7534 19966 7586 20018
rect 9998 19966 10050 20018
rect 10558 19966 10610 20018
rect 10782 19966 10834 20018
rect 11454 19966 11506 20018
rect 11902 19966 11954 20018
rect 12126 19966 12178 20018
rect 12686 19966 12738 20018
rect 14030 19966 14082 20018
rect 14702 19966 14754 20018
rect 15486 19966 15538 20018
rect 16606 19966 16658 20018
rect 17502 19966 17554 20018
rect 17950 19966 18002 20018
rect 18174 19966 18226 20018
rect 18510 19966 18562 20018
rect 18846 19966 18898 20018
rect 19070 19966 19122 20018
rect 20302 19966 20354 20018
rect 20750 19966 20802 20018
rect 21646 19966 21698 20018
rect 25678 19966 25730 20018
rect 2606 19854 2658 19906
rect 4734 19854 4786 19906
rect 5182 19854 5234 19906
rect 7422 19854 7474 19906
rect 9662 19854 9714 19906
rect 16046 19854 16098 19906
rect 18062 19854 18114 19906
rect 18958 19854 19010 19906
rect 21198 19854 21250 19906
rect 22318 19854 22370 19906
rect 24446 19854 24498 19906
rect 26462 19854 26514 19906
rect 28590 19854 28642 19906
rect 8654 19742 8706 19794
rect 8990 19742 9042 19794
rect 10222 19742 10274 19794
rect 12574 19742 12626 19794
rect 5372 19574 5424 19626
rect 5476 19574 5528 19626
rect 5580 19574 5632 19626
rect 13688 19574 13740 19626
rect 13792 19574 13844 19626
rect 13896 19574 13948 19626
rect 22004 19574 22056 19626
rect 22108 19574 22160 19626
rect 22212 19574 22264 19626
rect 30320 19574 30372 19626
rect 30424 19574 30476 19626
rect 30528 19574 30580 19626
rect 9774 19406 9826 19458
rect 12686 19406 12738 19458
rect 17614 19406 17666 19458
rect 21870 19406 21922 19458
rect 22206 19406 22258 19458
rect 2494 19294 2546 19346
rect 4622 19294 4674 19346
rect 7982 19294 8034 19346
rect 8990 19294 9042 19346
rect 9438 19294 9490 19346
rect 11342 19294 11394 19346
rect 12238 19294 12290 19346
rect 17390 19294 17442 19346
rect 18398 19294 18450 19346
rect 22878 19294 22930 19346
rect 26014 19294 26066 19346
rect 1822 19182 1874 19234
rect 7086 19182 7138 19234
rect 7310 19182 7362 19234
rect 8654 19182 8706 19234
rect 8878 19182 8930 19234
rect 9214 19182 9266 19234
rect 10782 19182 10834 19234
rect 27246 19182 27298 19234
rect 9998 19070 10050 19122
rect 10558 19070 10610 19122
rect 11230 19070 11282 19122
rect 12798 19070 12850 19122
rect 11006 18958 11058 19010
rect 11902 18958 11954 19010
rect 12126 18958 12178 19010
rect 12350 18958 12402 19010
rect 14926 18958 14978 19010
rect 17950 18958 18002 19010
rect 22094 18958 22146 19010
rect 9530 18790 9582 18842
rect 9634 18790 9686 18842
rect 9738 18790 9790 18842
rect 17846 18790 17898 18842
rect 17950 18790 18002 18842
rect 18054 18790 18106 18842
rect 26162 18790 26214 18842
rect 26266 18790 26318 18842
rect 26370 18790 26422 18842
rect 34478 18790 34530 18842
rect 34582 18790 34634 18842
rect 34686 18790 34738 18842
rect 7422 18622 7474 18674
rect 8206 18622 8258 18674
rect 10782 18622 10834 18674
rect 12686 18622 12738 18674
rect 22654 18622 22706 18674
rect 23326 18622 23378 18674
rect 5854 18510 5906 18562
rect 6526 18510 6578 18562
rect 7982 18510 8034 18562
rect 8766 18510 8818 18562
rect 8878 18510 8930 18562
rect 9550 18510 9602 18562
rect 9662 18510 9714 18562
rect 11454 18510 11506 18562
rect 19518 18510 19570 18562
rect 22990 18510 23042 18562
rect 26686 18510 26738 18562
rect 5630 18398 5682 18450
rect 6302 18398 6354 18450
rect 7870 18398 7922 18450
rect 8318 18398 8370 18450
rect 9886 18398 9938 18450
rect 10558 18398 10610 18450
rect 10670 18398 10722 18450
rect 11342 18398 11394 18450
rect 11678 18398 11730 18450
rect 11790 18398 11842 18450
rect 14030 18398 14082 18450
rect 17390 18398 17442 18450
rect 17614 18398 17666 18450
rect 18062 18398 18114 18450
rect 18734 18398 18786 18450
rect 23662 18398 23714 18450
rect 23886 18398 23938 18450
rect 23998 18398 24050 18450
rect 26238 18398 26290 18450
rect 27246 18398 27298 18450
rect 6862 18286 6914 18338
rect 7086 18286 7138 18338
rect 8094 18286 8146 18338
rect 10334 18286 10386 18338
rect 12126 18286 12178 18338
rect 12350 18286 12402 18338
rect 14702 18286 14754 18338
rect 16830 18286 16882 18338
rect 17502 18286 17554 18338
rect 21646 18286 21698 18338
rect 26574 18286 26626 18338
rect 29262 18286 29314 18338
rect 8878 18174 8930 18226
rect 10110 18174 10162 18226
rect 26910 18174 26962 18226
rect 5372 18006 5424 18058
rect 5476 18006 5528 18058
rect 5580 18006 5632 18058
rect 13688 18006 13740 18058
rect 13792 18006 13844 18058
rect 13896 18006 13948 18058
rect 22004 18006 22056 18058
rect 22108 18006 22160 18058
rect 22212 18006 22264 18058
rect 30320 18006 30372 18058
rect 30424 18006 30476 18058
rect 30528 18006 30580 18058
rect 6414 17838 6466 17890
rect 6750 17838 6802 17890
rect 9550 17838 9602 17890
rect 9886 17838 9938 17890
rect 26238 17838 26290 17890
rect 28478 17838 28530 17890
rect 4622 17726 4674 17778
rect 8430 17726 8482 17778
rect 10446 17726 10498 17778
rect 16046 17726 16098 17778
rect 25902 17726 25954 17778
rect 27918 17726 27970 17778
rect 29150 17726 29202 17778
rect 1822 17614 1874 17666
rect 6190 17614 6242 17666
rect 7086 17614 7138 17666
rect 7646 17614 7698 17666
rect 7870 17614 7922 17666
rect 9102 17614 9154 17666
rect 10222 17614 10274 17666
rect 10894 17614 10946 17666
rect 11230 17614 11282 17666
rect 15822 17614 15874 17666
rect 16158 17614 16210 17666
rect 16494 17614 16546 17666
rect 27246 17614 27298 17666
rect 27470 17614 27522 17666
rect 28142 17614 28194 17666
rect 31950 17614 32002 17666
rect 2494 17502 2546 17554
rect 10670 17502 10722 17554
rect 17390 17502 17442 17554
rect 18062 17502 18114 17554
rect 18958 17502 19010 17554
rect 26014 17502 26066 17554
rect 26574 17502 26626 17554
rect 31278 17502 31330 17554
rect 5070 17390 5122 17442
rect 7198 17390 7250 17442
rect 7422 17390 7474 17442
rect 8878 17390 8930 17442
rect 9774 17390 9826 17442
rect 10446 17390 10498 17442
rect 11118 17390 11170 17442
rect 17726 17390 17778 17442
rect 18398 17390 18450 17442
rect 19070 17390 19122 17442
rect 9530 17222 9582 17274
rect 9634 17222 9686 17274
rect 9738 17222 9790 17274
rect 17846 17222 17898 17274
rect 17950 17222 18002 17274
rect 18054 17222 18106 17274
rect 26162 17222 26214 17274
rect 26266 17222 26318 17274
rect 26370 17222 26422 17274
rect 34478 17222 34530 17274
rect 34582 17222 34634 17274
rect 34686 17222 34738 17274
rect 7086 17054 7138 17106
rect 7422 17054 7474 17106
rect 8206 17054 8258 17106
rect 8430 17054 8482 17106
rect 8654 17054 8706 17106
rect 9886 17054 9938 17106
rect 14366 17054 14418 17106
rect 15822 17054 15874 17106
rect 17390 17054 17442 17106
rect 28926 17054 28978 17106
rect 33070 17054 33122 17106
rect 8094 16942 8146 16994
rect 14142 16942 14194 16994
rect 15262 16942 15314 16994
rect 15934 16942 15986 16994
rect 16718 16942 16770 16994
rect 17614 16942 17666 16994
rect 17726 16942 17778 16994
rect 17950 16942 18002 16994
rect 20638 16942 20690 16994
rect 29038 16942 29090 16994
rect 3278 16830 3330 16882
rect 3950 16830 4002 16882
rect 6750 16830 6802 16882
rect 7534 16830 7586 16882
rect 8878 16830 8930 16882
rect 9550 16830 9602 16882
rect 12126 16830 12178 16882
rect 12238 16830 12290 16882
rect 13582 16830 13634 16882
rect 13918 16830 13970 16882
rect 15374 16830 15426 16882
rect 15710 16830 15762 16882
rect 16382 16830 16434 16882
rect 16830 16830 16882 16882
rect 21422 16830 21474 16882
rect 24558 16830 24610 16882
rect 25342 16830 25394 16882
rect 28590 16830 28642 16882
rect 29262 16830 29314 16882
rect 29598 16830 29650 16882
rect 33294 16830 33346 16882
rect 33630 16830 33682 16882
rect 6078 16718 6130 16770
rect 12798 16718 12850 16770
rect 14030 16718 14082 16770
rect 18174 16718 18226 16770
rect 18510 16718 18562 16770
rect 21758 16718 21810 16770
rect 23886 16718 23938 16770
rect 26014 16718 26066 16770
rect 28142 16718 28194 16770
rect 30382 16718 30434 16770
rect 32510 16718 32562 16770
rect 33182 16718 33234 16770
rect 12686 16606 12738 16658
rect 15262 16606 15314 16658
rect 16718 16606 16770 16658
rect 5372 16438 5424 16490
rect 5476 16438 5528 16490
rect 5580 16438 5632 16490
rect 13688 16438 13740 16490
rect 13792 16438 13844 16490
rect 13896 16438 13948 16490
rect 22004 16438 22056 16490
rect 22108 16438 22160 16490
rect 22212 16438 22264 16490
rect 30320 16438 30372 16490
rect 30424 16438 30476 16490
rect 30528 16438 30580 16490
rect 5742 16270 5794 16322
rect 6302 16270 6354 16322
rect 17950 16270 18002 16322
rect 5070 16158 5122 16210
rect 5742 16158 5794 16210
rect 6302 16158 6354 16210
rect 10782 16158 10834 16210
rect 12910 16158 12962 16210
rect 13694 16158 13746 16210
rect 17390 16158 17442 16210
rect 17726 16158 17778 16210
rect 23438 16158 23490 16210
rect 24446 16158 24498 16210
rect 28030 16158 28082 16210
rect 29262 16158 29314 16210
rect 34190 16158 34242 16210
rect 2270 16046 2322 16098
rect 10110 16046 10162 16098
rect 13806 16046 13858 16098
rect 14814 16046 14866 16098
rect 15486 16046 15538 16098
rect 15710 16046 15762 16098
rect 15934 16046 15986 16098
rect 16606 16046 16658 16098
rect 17278 16046 17330 16098
rect 19070 16046 19122 16098
rect 22430 16046 22482 16098
rect 23662 16046 23714 16098
rect 24670 16046 24722 16098
rect 27022 16046 27074 16098
rect 27918 16046 27970 16098
rect 28142 16046 28194 16098
rect 29150 16046 29202 16098
rect 29374 16046 29426 16098
rect 29822 16046 29874 16098
rect 30046 16046 30098 16098
rect 31390 16046 31442 16098
rect 2942 15934 2994 15986
rect 14142 15934 14194 15986
rect 14478 15934 14530 15986
rect 15038 15934 15090 15986
rect 15150 15934 15202 15986
rect 16046 15934 16098 15986
rect 16158 15934 16210 15986
rect 16942 15934 16994 15986
rect 18510 15934 18562 15986
rect 18622 15934 18674 15986
rect 21422 15934 21474 15986
rect 22206 15934 22258 15986
rect 22654 15934 22706 15986
rect 22766 15934 22818 15986
rect 24334 15934 24386 15986
rect 27582 15934 27634 15986
rect 28366 15934 28418 15986
rect 32062 15934 32114 15986
rect 9662 15822 9714 15874
rect 14254 15822 14306 15874
rect 16830 15822 16882 15874
rect 18286 15822 18338 15874
rect 18846 15822 18898 15874
rect 21534 15822 21586 15874
rect 21646 15822 21698 15874
rect 23998 15822 24050 15874
rect 27358 15822 27410 15874
rect 27694 15822 27746 15874
rect 30382 15822 30434 15874
rect 9530 15654 9582 15706
rect 9634 15654 9686 15706
rect 9738 15654 9790 15706
rect 17846 15654 17898 15706
rect 17950 15654 18002 15706
rect 18054 15654 18106 15706
rect 26162 15654 26214 15706
rect 26266 15654 26318 15706
rect 26370 15654 26422 15706
rect 34478 15654 34530 15706
rect 34582 15654 34634 15706
rect 34686 15654 34738 15706
rect 14814 15486 14866 15538
rect 15486 15486 15538 15538
rect 15598 15486 15650 15538
rect 27358 15486 27410 15538
rect 27582 15486 27634 15538
rect 29934 15486 29986 15538
rect 33070 15486 33122 15538
rect 11902 15374 11954 15426
rect 14702 15374 14754 15426
rect 16270 15374 16322 15426
rect 16718 15374 16770 15426
rect 16830 15374 16882 15426
rect 22878 15374 22930 15426
rect 26126 15374 26178 15426
rect 26350 15374 26402 15426
rect 27694 15374 27746 15426
rect 28814 15374 28866 15426
rect 29262 15374 29314 15426
rect 29486 15374 29538 15426
rect 30382 15374 30434 15426
rect 30942 15374 30994 15426
rect 32398 15374 32450 15426
rect 5742 15262 5794 15314
rect 8990 15262 9042 15314
rect 11230 15262 11282 15314
rect 15262 15262 15314 15314
rect 15374 15262 15426 15314
rect 15710 15262 15762 15314
rect 17950 15262 18002 15314
rect 18174 15262 18226 15314
rect 28590 15262 28642 15314
rect 31054 15262 31106 15314
rect 31502 15262 31554 15314
rect 31726 15262 31778 15314
rect 32062 15262 32114 15314
rect 33630 15262 33682 15314
rect 6414 15150 6466 15202
rect 8542 15150 8594 15202
rect 14030 15150 14082 15202
rect 16382 15150 16434 15202
rect 26014 15150 26066 15202
rect 29262 15150 29314 15202
rect 29822 15150 29874 15202
rect 30494 15150 30546 15202
rect 30606 15150 30658 15202
rect 33406 15150 33458 15202
rect 31278 15038 31330 15090
rect 32062 15038 32114 15090
rect 5372 14870 5424 14922
rect 5476 14870 5528 14922
rect 5580 14870 5632 14922
rect 13688 14870 13740 14922
rect 13792 14870 13844 14922
rect 13896 14870 13948 14922
rect 22004 14870 22056 14922
rect 22108 14870 22160 14922
rect 22212 14870 22264 14922
rect 30320 14870 30372 14922
rect 30424 14870 30476 14922
rect 30528 14870 30580 14922
rect 17950 14702 18002 14754
rect 18174 14702 18226 14754
rect 28254 14702 28306 14754
rect 29262 14702 29314 14754
rect 30830 14702 30882 14754
rect 32174 14702 32226 14754
rect 32622 14702 32674 14754
rect 4622 14590 4674 14642
rect 16494 14590 16546 14642
rect 20638 14590 20690 14642
rect 21310 14590 21362 14642
rect 23438 14590 23490 14642
rect 29598 14590 29650 14642
rect 31166 14590 31218 14642
rect 1822 14478 1874 14530
rect 5630 14478 5682 14530
rect 12686 14478 12738 14530
rect 16158 14478 16210 14530
rect 17054 14478 17106 14530
rect 17390 14478 17442 14530
rect 17502 14478 17554 14530
rect 19630 14478 19682 14530
rect 20750 14478 20802 14530
rect 24222 14478 24274 14530
rect 27246 14478 27298 14530
rect 28030 14478 28082 14530
rect 29374 14478 29426 14530
rect 31838 14478 31890 14530
rect 32398 14478 32450 14530
rect 32846 14478 32898 14530
rect 2494 14366 2546 14418
rect 8430 14366 8482 14418
rect 15822 14366 15874 14418
rect 17726 14366 17778 14418
rect 19406 14366 19458 14418
rect 20078 14366 20130 14418
rect 27470 14366 27522 14418
rect 27582 14366 27634 14418
rect 29710 14366 29762 14418
rect 30718 14366 30770 14418
rect 31278 14366 31330 14418
rect 31614 14366 31666 14418
rect 5070 14254 5122 14306
rect 5966 14254 6018 14306
rect 13582 14254 13634 14306
rect 15934 14254 15986 14306
rect 20302 14254 20354 14306
rect 20526 14254 20578 14306
rect 32510 14254 32562 14306
rect 9530 14086 9582 14138
rect 9634 14086 9686 14138
rect 9738 14086 9790 14138
rect 17846 14086 17898 14138
rect 17950 14086 18002 14138
rect 18054 14086 18106 14138
rect 26162 14086 26214 14138
rect 26266 14086 26318 14138
rect 26370 14086 26422 14138
rect 34478 14086 34530 14138
rect 34582 14086 34634 14138
rect 34686 14086 34738 14138
rect 6526 13918 6578 13970
rect 10670 13918 10722 13970
rect 11118 13918 11170 13970
rect 17390 13918 17442 13970
rect 18398 13918 18450 13970
rect 18846 13918 18898 13970
rect 22878 13918 22930 13970
rect 23662 13918 23714 13970
rect 24222 13918 24274 13970
rect 25678 13918 25730 13970
rect 31278 13918 31330 13970
rect 32286 13918 32338 13970
rect 10558 13806 10610 13858
rect 10894 13806 10946 13858
rect 11790 13806 11842 13858
rect 15934 13806 15986 13858
rect 19406 13806 19458 13858
rect 20414 13806 20466 13858
rect 29934 13806 29986 13858
rect 5406 13694 5458 13746
rect 5630 13694 5682 13746
rect 6302 13694 6354 13746
rect 6414 13694 6466 13746
rect 6750 13694 6802 13746
rect 10110 13694 10162 13746
rect 10334 13694 10386 13746
rect 11342 13694 11394 13746
rect 15262 13694 15314 13746
rect 15822 13694 15874 13746
rect 17726 13694 17778 13746
rect 18174 13694 18226 13746
rect 18734 13694 18786 13746
rect 19070 13694 19122 13746
rect 20078 13694 20130 13746
rect 22206 13694 22258 13746
rect 22654 13694 22706 13746
rect 23550 13694 23602 13746
rect 23886 13694 23938 13746
rect 25454 13694 25506 13746
rect 26126 13694 26178 13746
rect 26350 13694 26402 13746
rect 26686 13694 26738 13746
rect 27022 13694 27074 13746
rect 30718 13694 30770 13746
rect 31726 13694 31778 13746
rect 33182 13694 33234 13746
rect 33630 13694 33682 13746
rect 5854 13582 5906 13634
rect 7758 13582 7810 13634
rect 10894 13582 10946 13634
rect 26462 13582 26514 13634
rect 27246 13582 27298 13634
rect 27806 13582 27858 13634
rect 7870 13470 7922 13522
rect 11678 13470 11730 13522
rect 21310 13470 21362 13522
rect 21758 13470 21810 13522
rect 21982 13470 22034 13522
rect 26910 13470 26962 13522
rect 27358 13470 27410 13522
rect 31054 13470 31106 13522
rect 31390 13470 31442 13522
rect 31950 13470 32002 13522
rect 33294 13470 33346 13522
rect 33518 13470 33570 13522
rect 5372 13302 5424 13354
rect 5476 13302 5528 13354
rect 5580 13302 5632 13354
rect 13688 13302 13740 13354
rect 13792 13302 13844 13354
rect 13896 13302 13948 13354
rect 22004 13302 22056 13354
rect 22108 13302 22160 13354
rect 22212 13302 22264 13354
rect 30320 13302 30372 13354
rect 30424 13302 30476 13354
rect 30528 13302 30580 13354
rect 6526 13134 6578 13186
rect 18622 13134 18674 13186
rect 20302 13134 20354 13186
rect 22094 13134 22146 13186
rect 29150 13134 29202 13186
rect 29486 13134 29538 13186
rect 4622 13022 4674 13074
rect 7422 13022 7474 13074
rect 10782 13022 10834 13074
rect 11230 13022 11282 13074
rect 12126 13022 12178 13074
rect 15374 13022 15426 13074
rect 17054 13022 17106 13074
rect 17950 13022 18002 13074
rect 20078 13022 20130 13074
rect 22318 13022 22370 13074
rect 22990 13022 23042 13074
rect 24782 13022 24834 13074
rect 26910 13022 26962 13074
rect 29710 13022 29762 13074
rect 31278 13022 31330 13074
rect 33406 13022 33458 13074
rect 3614 12910 3666 12962
rect 4286 12910 4338 12962
rect 5070 12910 5122 12962
rect 5630 12910 5682 12962
rect 5854 12910 5906 12962
rect 6078 12910 6130 12962
rect 6750 12910 6802 12962
rect 7086 12910 7138 12962
rect 7982 12910 8034 12962
rect 11678 12910 11730 12962
rect 12574 12910 12626 12962
rect 18846 12910 18898 12962
rect 19518 12910 19570 12962
rect 20526 12910 20578 12962
rect 20862 12910 20914 12962
rect 21870 12910 21922 12962
rect 24110 12910 24162 12962
rect 27470 12910 27522 12962
rect 34078 12910 34130 12962
rect 7534 12798 7586 12850
rect 8654 12798 8706 12850
rect 13806 12798 13858 12850
rect 14142 12798 14194 12850
rect 19294 12798 19346 12850
rect 19854 12798 19906 12850
rect 21646 12798 21698 12850
rect 22542 12798 22594 12850
rect 22878 12798 22930 12850
rect 27358 12798 27410 12850
rect 3726 12686 3778 12738
rect 3838 12686 3890 12738
rect 4510 12686 4562 12738
rect 4734 12686 4786 12738
rect 6862 12686 6914 12738
rect 11118 12686 11170 12738
rect 11342 12686 11394 12738
rect 12014 12686 12066 12738
rect 18398 12686 18450 12738
rect 18510 12686 18562 12738
rect 19406 12686 19458 12738
rect 19742 12686 19794 12738
rect 22430 12686 22482 12738
rect 27134 12686 27186 12738
rect 9530 12518 9582 12570
rect 9634 12518 9686 12570
rect 9738 12518 9790 12570
rect 17846 12518 17898 12570
rect 17950 12518 18002 12570
rect 18054 12518 18106 12570
rect 26162 12518 26214 12570
rect 26266 12518 26318 12570
rect 26370 12518 26422 12570
rect 34478 12518 34530 12570
rect 34582 12518 34634 12570
rect 34686 12518 34738 12570
rect 4174 12350 4226 12402
rect 5294 12350 5346 12402
rect 5630 12350 5682 12402
rect 6414 12350 6466 12402
rect 7086 12350 7138 12402
rect 9886 12350 9938 12402
rect 20638 12350 20690 12402
rect 20974 12350 21026 12402
rect 3166 12238 3218 12290
rect 3614 12238 3666 12290
rect 6750 12238 6802 12290
rect 7982 12238 8034 12290
rect 8654 12238 8706 12290
rect 8990 12238 9042 12290
rect 9550 12238 9602 12290
rect 10558 12238 10610 12290
rect 18174 12238 18226 12290
rect 23662 12238 23714 12290
rect 2830 12126 2882 12178
rect 3502 12126 3554 12178
rect 3838 12126 3890 12178
rect 4398 12126 4450 12178
rect 4510 12126 4562 12178
rect 4734 12126 4786 12178
rect 4958 12126 5010 12178
rect 7422 12126 7474 12178
rect 8318 12126 8370 12178
rect 10334 12126 10386 12178
rect 11006 12126 11058 12178
rect 12686 12126 12738 12178
rect 17502 12126 17554 12178
rect 24334 12126 24386 12178
rect 26014 12126 26066 12178
rect 26574 12126 26626 12178
rect 31502 12126 31554 12178
rect 6078 12014 6130 12066
rect 10782 12014 10834 12066
rect 13582 12014 13634 12066
rect 20302 12014 20354 12066
rect 21534 12014 21586 12066
rect 26686 12014 26738 12066
rect 5854 11902 5906 11954
rect 6190 11902 6242 11954
rect 31390 11902 31442 11954
rect 31726 11902 31778 11954
rect 31838 11902 31890 11954
rect 5372 11734 5424 11786
rect 5476 11734 5528 11786
rect 5580 11734 5632 11786
rect 13688 11734 13740 11786
rect 13792 11734 13844 11786
rect 13896 11734 13948 11786
rect 22004 11734 22056 11786
rect 22108 11734 22160 11786
rect 22212 11734 22264 11786
rect 30320 11734 30372 11786
rect 30424 11734 30476 11786
rect 30528 11734 30580 11786
rect 6862 11566 6914 11618
rect 8654 11566 8706 11618
rect 8878 11566 8930 11618
rect 17614 11566 17666 11618
rect 20414 11566 20466 11618
rect 22766 11566 22818 11618
rect 2382 11454 2434 11506
rect 3054 11454 3106 11506
rect 4286 11454 4338 11506
rect 6414 11454 6466 11506
rect 9886 11454 9938 11506
rect 10670 11454 10722 11506
rect 14254 11454 14306 11506
rect 16382 11454 16434 11506
rect 17838 11454 17890 11506
rect 18734 11454 18786 11506
rect 19518 11454 19570 11506
rect 20526 11454 20578 11506
rect 21422 11454 21474 11506
rect 22878 11454 22930 11506
rect 27358 11454 27410 11506
rect 32062 11454 32114 11506
rect 34190 11454 34242 11506
rect 2158 11342 2210 11394
rect 3278 11342 3330 11394
rect 3502 11342 3554 11394
rect 3614 11342 3666 11394
rect 4174 11342 4226 11394
rect 5518 11342 5570 11394
rect 6078 11342 6130 11394
rect 6302 11342 6354 11394
rect 6526 11342 6578 11394
rect 7086 11342 7138 11394
rect 7534 11342 7586 11394
rect 8990 11342 9042 11394
rect 9550 11342 9602 11394
rect 10446 11342 10498 11394
rect 13470 11342 13522 11394
rect 19406 11342 19458 11394
rect 19630 11342 19682 11394
rect 19854 11342 19906 11394
rect 20078 11342 20130 11394
rect 21534 11342 21586 11394
rect 21870 11342 21922 11394
rect 24446 11342 24498 11394
rect 29150 11342 29202 11394
rect 29486 11342 29538 11394
rect 30270 11342 30322 11394
rect 31278 11342 31330 11394
rect 4510 11230 4562 11282
rect 4622 11230 4674 11282
rect 5854 11230 5906 11282
rect 7422 11230 7474 11282
rect 7870 11230 7922 11282
rect 8206 11230 8258 11282
rect 8542 11230 8594 11282
rect 9662 11230 9714 11282
rect 9998 11230 10050 11282
rect 16718 11230 16770 11282
rect 25230 11230 25282 11282
rect 2270 11118 2322 11170
rect 2494 11118 2546 11170
rect 2606 11118 2658 11170
rect 3726 11118 3778 11170
rect 4398 11118 4450 11170
rect 7310 11118 7362 11170
rect 8094 11118 8146 11170
rect 10670 11118 10722 11170
rect 16830 11118 16882 11170
rect 17278 11118 17330 11170
rect 18286 11118 18338 11170
rect 29598 11118 29650 11170
rect 29710 11118 29762 11170
rect 30046 11118 30098 11170
rect 9530 10950 9582 11002
rect 9634 10950 9686 11002
rect 9738 10950 9790 11002
rect 17846 10950 17898 11002
rect 17950 10950 18002 11002
rect 18054 10950 18106 11002
rect 26162 10950 26214 11002
rect 26266 10950 26318 11002
rect 26370 10950 26422 11002
rect 34478 10950 34530 11002
rect 34582 10950 34634 11002
rect 34686 10950 34738 11002
rect 3278 10782 3330 10834
rect 3726 10782 3778 10834
rect 4734 10782 4786 10834
rect 4958 10782 5010 10834
rect 10334 10782 10386 10834
rect 10894 10782 10946 10834
rect 17390 10782 17442 10834
rect 25790 10782 25842 10834
rect 3838 10670 3890 10722
rect 7982 10670 8034 10722
rect 8990 10670 9042 10722
rect 10446 10670 10498 10722
rect 11118 10670 11170 10722
rect 13022 10670 13074 10722
rect 26014 10670 26066 10722
rect 30718 10670 30770 10722
rect 33294 10670 33346 10722
rect 2718 10558 2770 10610
rect 3054 10558 3106 10610
rect 5070 10558 5122 10610
rect 7870 10558 7922 10610
rect 8206 10558 8258 10610
rect 8542 10558 8594 10610
rect 8878 10558 8930 10610
rect 9550 10558 9602 10610
rect 9886 10558 9938 10610
rect 9998 10558 10050 10610
rect 10670 10558 10722 10610
rect 11342 10558 11394 10610
rect 12350 10558 12402 10610
rect 16270 10558 16322 10610
rect 16494 10558 16546 10610
rect 16606 10558 16658 10610
rect 16830 10558 16882 10610
rect 18510 10558 18562 10610
rect 22318 10558 22370 10610
rect 26910 10558 26962 10610
rect 27246 10558 27298 10610
rect 2942 10446 2994 10498
rect 10222 10446 10274 10498
rect 15150 10446 15202 10498
rect 17838 10446 17890 10498
rect 19182 10446 19234 10498
rect 21310 10446 21362 10498
rect 25678 10446 25730 10498
rect 3614 10334 3666 10386
rect 8654 10334 8706 10386
rect 15822 10334 15874 10386
rect 33070 10334 33122 10386
rect 33406 10334 33458 10386
rect 5372 10166 5424 10218
rect 5476 10166 5528 10218
rect 5580 10166 5632 10218
rect 13688 10166 13740 10218
rect 13792 10166 13844 10218
rect 13896 10166 13948 10218
rect 22004 10166 22056 10218
rect 22108 10166 22160 10218
rect 22212 10166 22264 10218
rect 30320 10166 30372 10218
rect 30424 10166 30476 10218
rect 30528 10166 30580 10218
rect 2270 9998 2322 10050
rect 2718 9998 2770 10050
rect 9214 9998 9266 10050
rect 19630 9998 19682 10050
rect 31054 9998 31106 10050
rect 6078 9886 6130 9938
rect 8878 9886 8930 9938
rect 10558 9886 10610 9938
rect 12462 9886 12514 9938
rect 14478 9886 14530 9938
rect 20414 9886 20466 9938
rect 21758 9886 21810 9938
rect 30046 9886 30098 9938
rect 34190 9886 34242 9938
rect 2942 9774 2994 9826
rect 3166 9774 3218 9826
rect 5630 9774 5682 9826
rect 9102 9774 9154 9826
rect 9550 9774 9602 9826
rect 11454 9774 11506 9826
rect 11566 9774 11618 9826
rect 12910 9774 12962 9826
rect 14030 9774 14082 9826
rect 17838 9774 17890 9826
rect 19294 9774 19346 9826
rect 19742 9774 19794 9826
rect 26910 9774 26962 9826
rect 29262 9774 29314 9826
rect 29486 9774 29538 9826
rect 29710 9774 29762 9826
rect 30382 9774 30434 9826
rect 30830 9774 30882 9826
rect 31278 9774 31330 9826
rect 3502 9662 3554 9714
rect 3950 9662 4002 9714
rect 5854 9662 5906 9714
rect 6190 9662 6242 9714
rect 8766 9662 8818 9714
rect 9998 9662 10050 9714
rect 10110 9662 10162 9714
rect 10670 9662 10722 9714
rect 10894 9662 10946 9714
rect 11230 9662 11282 9714
rect 13694 9662 13746 9714
rect 14142 9662 14194 9714
rect 17278 9662 17330 9714
rect 18622 9662 18674 9714
rect 18958 9662 19010 9714
rect 19854 9662 19906 9714
rect 21422 9662 21474 9714
rect 22094 9662 22146 9714
rect 22878 9662 22930 9714
rect 30270 9662 30322 9714
rect 32062 9662 32114 9714
rect 3614 9550 3666 9602
rect 3726 9550 3778 9602
rect 10334 9550 10386 9602
rect 12014 9550 12066 9602
rect 13582 9550 13634 9602
rect 18286 9550 18338 9602
rect 21870 9550 21922 9602
rect 28254 9550 28306 9602
rect 28590 9550 28642 9602
rect 29486 9550 29538 9602
rect 9530 9382 9582 9434
rect 9634 9382 9686 9434
rect 9738 9382 9790 9434
rect 17846 9382 17898 9434
rect 17950 9382 18002 9434
rect 18054 9382 18106 9434
rect 26162 9382 26214 9434
rect 26266 9382 26318 9434
rect 26370 9382 26422 9434
rect 34478 9382 34530 9434
rect 34582 9382 34634 9434
rect 34686 9382 34738 9434
rect 3390 9214 3442 9266
rect 5294 9214 5346 9266
rect 5406 9214 5458 9266
rect 6862 9214 6914 9266
rect 7870 9214 7922 9266
rect 26238 9214 26290 9266
rect 26574 9214 26626 9266
rect 33182 9214 33234 9266
rect 2494 9102 2546 9154
rect 2830 9102 2882 9154
rect 7758 9102 7810 9154
rect 3166 8990 3218 9042
rect 3502 8990 3554 9042
rect 3726 8990 3778 9042
rect 4846 8990 4898 9042
rect 5182 8990 5234 9042
rect 5518 8990 5570 9042
rect 6414 8990 6466 9042
rect 6638 8990 6690 9042
rect 7646 8990 7698 9042
rect 8318 8990 8370 9042
rect 9550 8990 9602 9042
rect 9774 9046 9826 9098
rect 10110 9102 10162 9154
rect 16270 9102 16322 9154
rect 9886 9046 9938 9098
rect 17278 9102 17330 9154
rect 18846 9102 18898 9154
rect 19742 9102 19794 9154
rect 21758 9102 21810 9154
rect 27806 9102 27858 9154
rect 30382 9102 30434 9154
rect 31838 9102 31890 9154
rect 33630 9102 33682 9154
rect 11902 8990 11954 9042
rect 13246 8990 13298 9042
rect 15038 8990 15090 9042
rect 15374 8990 15426 9042
rect 18958 8990 19010 9042
rect 19294 8990 19346 9042
rect 20974 8990 21026 9042
rect 24334 8990 24386 9042
rect 24558 8990 24610 9042
rect 27022 8990 27074 9042
rect 30270 8990 30322 9042
rect 31278 8990 31330 9042
rect 33070 8990 33122 9042
rect 33294 8990 33346 9042
rect 6526 8878 6578 8930
rect 10334 8878 10386 8930
rect 12238 8878 12290 8930
rect 13134 8878 13186 8930
rect 14478 8878 14530 8930
rect 23886 8878 23938 8930
rect 29934 8878 29986 8930
rect 30606 8878 30658 8930
rect 3726 8766 3778 8818
rect 11342 8766 11394 8818
rect 11678 8766 11730 8818
rect 24222 8766 24274 8818
rect 5372 8598 5424 8650
rect 5476 8598 5528 8650
rect 5580 8598 5632 8650
rect 13688 8598 13740 8650
rect 13792 8598 13844 8650
rect 13896 8598 13948 8650
rect 22004 8598 22056 8650
rect 22108 8598 22160 8650
rect 22212 8598 22264 8650
rect 30320 8598 30372 8650
rect 30424 8598 30476 8650
rect 30528 8598 30580 8650
rect 12574 8430 12626 8482
rect 19070 8430 19122 8482
rect 2718 8318 2770 8370
rect 3838 8318 3890 8370
rect 7198 8318 7250 8370
rect 9214 8318 9266 8370
rect 9662 8318 9714 8370
rect 12238 8318 12290 8370
rect 12798 8318 12850 8370
rect 13358 8318 13410 8370
rect 18286 8318 18338 8370
rect 22318 8318 22370 8370
rect 23774 8318 23826 8370
rect 25902 8318 25954 8370
rect 28142 8318 28194 8370
rect 29934 8318 29986 8370
rect 30046 8318 30098 8370
rect 30382 8318 30434 8370
rect 34190 8318 34242 8370
rect 3166 8206 3218 8258
rect 3390 8206 3442 8258
rect 3614 8206 3666 8258
rect 4958 8206 5010 8258
rect 5630 8206 5682 8258
rect 5854 8206 5906 8258
rect 6078 8206 6130 8258
rect 6862 8206 6914 8258
rect 9438 8206 9490 8258
rect 9886 8206 9938 8258
rect 11678 8206 11730 8258
rect 15150 8206 15202 8258
rect 16718 8206 16770 8258
rect 18062 8206 18114 8258
rect 18958 8206 19010 8258
rect 22094 8206 22146 8258
rect 22990 8206 23042 8258
rect 26238 8206 26290 8258
rect 27134 8206 27186 8258
rect 27694 8206 27746 8258
rect 28030 8206 28082 8258
rect 30606 8206 30658 8258
rect 31278 8206 31330 8258
rect 2830 8094 2882 8146
rect 3838 8094 3890 8146
rect 4622 8094 4674 8146
rect 6302 8094 6354 8146
rect 6526 8094 6578 8146
rect 7534 8094 7586 8146
rect 8766 8094 8818 8146
rect 8990 8094 9042 8146
rect 10110 8094 10162 8146
rect 10446 8094 10498 8146
rect 11118 8094 11170 8146
rect 11454 8094 11506 8146
rect 12014 8094 12066 8146
rect 12238 8094 12290 8146
rect 14926 8094 14978 8146
rect 15822 8094 15874 8146
rect 32062 8094 32114 8146
rect 2606 7982 2658 8034
rect 4062 7982 4114 8034
rect 4734 7982 4786 8034
rect 5518 7982 5570 8034
rect 7086 7982 7138 8034
rect 7310 7982 7362 8034
rect 8430 7982 8482 8034
rect 8654 7982 8706 8034
rect 17166 7982 17218 8034
rect 21534 7982 21586 8034
rect 21758 7982 21810 8034
rect 26574 7982 26626 8034
rect 26910 7982 26962 8034
rect 28254 7982 28306 8034
rect 30942 7982 30994 8034
rect 9530 7814 9582 7866
rect 9634 7814 9686 7866
rect 9738 7814 9790 7866
rect 17846 7814 17898 7866
rect 17950 7814 18002 7866
rect 18054 7814 18106 7866
rect 26162 7814 26214 7866
rect 26266 7814 26318 7866
rect 26370 7814 26422 7866
rect 34478 7814 34530 7866
rect 34582 7814 34634 7866
rect 34686 7814 34738 7866
rect 2942 7646 2994 7698
rect 5182 7646 5234 7698
rect 6750 7646 6802 7698
rect 6862 7646 6914 7698
rect 8094 7646 8146 7698
rect 8878 7646 8930 7698
rect 9662 7646 9714 7698
rect 10558 7646 10610 7698
rect 11566 7646 11618 7698
rect 12574 7646 12626 7698
rect 12910 7646 12962 7698
rect 27470 7646 27522 7698
rect 28142 7646 28194 7698
rect 30270 7646 30322 7698
rect 31726 7646 31778 7698
rect 2158 7534 2210 7586
rect 2494 7534 2546 7586
rect 4510 7534 4562 7586
rect 4846 7534 4898 7586
rect 14366 7534 14418 7586
rect 22430 7534 22482 7586
rect 23326 7534 23378 7586
rect 23550 7534 23602 7586
rect 25902 7534 25954 7586
rect 27918 7534 27970 7586
rect 29486 7534 29538 7586
rect 33070 7534 33122 7586
rect 2830 7422 2882 7474
rect 3054 7422 3106 7474
rect 3502 7422 3554 7474
rect 4398 7422 4450 7474
rect 5182 7422 5234 7474
rect 5294 7422 5346 7474
rect 5518 7422 5570 7474
rect 5742 7422 5794 7474
rect 6638 7422 6690 7474
rect 7198 7422 7250 7474
rect 7870 7422 7922 7474
rect 7982 7422 8034 7474
rect 8206 7422 8258 7474
rect 8430 7422 8482 7474
rect 8990 7422 9042 7474
rect 9550 7422 9602 7474
rect 9774 7422 9826 7474
rect 10222 7422 10274 7474
rect 10894 7422 10946 7474
rect 11454 7422 11506 7474
rect 11678 7422 11730 7474
rect 12014 7422 12066 7474
rect 13134 7422 13186 7474
rect 13358 7422 13410 7474
rect 14142 7422 14194 7474
rect 15262 7422 15314 7474
rect 15486 7422 15538 7474
rect 16270 7422 16322 7474
rect 16494 7422 16546 7474
rect 17838 7422 17890 7474
rect 18286 7422 18338 7474
rect 18734 7422 18786 7474
rect 21982 7422 22034 7474
rect 22206 7422 22258 7474
rect 22766 7422 22818 7474
rect 22990 7422 23042 7474
rect 26014 7422 26066 7474
rect 26238 7422 26290 7474
rect 27582 7422 27634 7474
rect 29262 7422 29314 7474
rect 29598 7422 29650 7474
rect 29822 7422 29874 7474
rect 31614 7422 31666 7474
rect 31838 7422 31890 7474
rect 32286 7422 32338 7474
rect 32510 7422 32562 7474
rect 33406 7422 33458 7474
rect 33518 7422 33570 7474
rect 4174 7310 4226 7362
rect 13918 7310 13970 7362
rect 14254 7310 14306 7362
rect 16606 7310 16658 7362
rect 17390 7310 17442 7362
rect 19518 7310 19570 7362
rect 21646 7310 21698 7362
rect 23438 7310 23490 7362
rect 25678 7310 25730 7362
rect 28030 7310 28082 7362
rect 3838 7198 3890 7250
rect 3950 7198 4002 7250
rect 8878 7198 8930 7250
rect 12798 7198 12850 7250
rect 26686 7198 26738 7250
rect 27134 7198 27186 7250
rect 27358 7198 27410 7250
rect 31390 7198 31442 7250
rect 32174 7198 32226 7250
rect 33182 7198 33234 7250
rect 5372 7030 5424 7082
rect 5476 7030 5528 7082
rect 5580 7030 5632 7082
rect 13688 7030 13740 7082
rect 13792 7030 13844 7082
rect 13896 7030 13948 7082
rect 22004 7030 22056 7082
rect 22108 7030 22160 7082
rect 22212 7030 22264 7082
rect 30320 7030 30372 7082
rect 30424 7030 30476 7082
rect 30528 7030 30580 7082
rect 9998 6862 10050 6914
rect 27134 6862 27186 6914
rect 29374 6862 29426 6914
rect 5742 6750 5794 6802
rect 7758 6750 7810 6802
rect 18174 6750 18226 6802
rect 23774 6750 23826 6802
rect 29150 6750 29202 6802
rect 29710 6750 29762 6802
rect 30382 6750 30434 6802
rect 33966 6750 34018 6802
rect 4958 6638 5010 6690
rect 5630 6638 5682 6690
rect 6414 6638 6466 6690
rect 7646 6638 7698 6690
rect 8654 6638 8706 6690
rect 10222 6638 10274 6690
rect 10894 6638 10946 6690
rect 12910 6638 12962 6690
rect 13358 6638 13410 6690
rect 14590 6638 14642 6690
rect 15262 6638 15314 6690
rect 21758 6638 21810 6690
rect 22094 6638 22146 6690
rect 22318 6638 22370 6690
rect 23214 6638 23266 6690
rect 26462 6638 26514 6690
rect 27246 6638 27298 6690
rect 27470 6638 27522 6690
rect 28142 6638 28194 6690
rect 30158 6638 30210 6690
rect 30718 6638 30770 6690
rect 31054 6638 31106 6690
rect 5070 6526 5122 6578
rect 6078 6526 6130 6578
rect 6638 6526 6690 6578
rect 6750 6526 6802 6578
rect 7982 6526 8034 6578
rect 10558 6526 10610 6578
rect 11230 6526 11282 6578
rect 12574 6526 12626 6578
rect 13806 6526 13858 6578
rect 14254 6526 14306 6578
rect 16046 6526 16098 6578
rect 19070 6526 19122 6578
rect 22990 6526 23042 6578
rect 24110 6526 24162 6578
rect 24782 6526 24834 6578
rect 27582 6526 27634 6578
rect 31838 6526 31890 6578
rect 5854 6414 5906 6466
rect 8878 6414 8930 6466
rect 9662 6414 9714 6466
rect 11566 6414 11618 6466
rect 18734 6414 18786 6466
rect 27918 6414 27970 6466
rect 9530 6246 9582 6298
rect 9634 6246 9686 6298
rect 9738 6246 9790 6298
rect 17846 6246 17898 6298
rect 17950 6246 18002 6298
rect 18054 6246 18106 6298
rect 26162 6246 26214 6298
rect 26266 6246 26318 6298
rect 26370 6246 26422 6298
rect 34478 6246 34530 6298
rect 34582 6246 34634 6298
rect 34686 6246 34738 6298
rect 3054 6078 3106 6130
rect 4622 6078 4674 6130
rect 5518 6078 5570 6130
rect 6190 6078 6242 6130
rect 7198 6078 7250 6130
rect 7646 6078 7698 6130
rect 3502 5966 3554 6018
rect 5854 5966 5906 6018
rect 6750 5966 6802 6018
rect 6862 5966 6914 6018
rect 2830 5854 2882 5906
rect 4398 5854 4450 5906
rect 5182 5854 5234 5906
rect 6526 5854 6578 5906
rect 7982 6078 8034 6130
rect 8206 6078 8258 6130
rect 13694 6078 13746 6130
rect 20974 6078 21026 6130
rect 33294 6078 33346 6130
rect 7870 5966 7922 6018
rect 8430 5966 8482 6018
rect 12014 5966 12066 6018
rect 12686 5966 12738 6018
rect 13022 5966 13074 6018
rect 16606 5966 16658 6018
rect 21310 5966 21362 6018
rect 22990 5966 23042 6018
rect 25678 5966 25730 6018
rect 26686 5966 26738 6018
rect 28702 5966 28754 6018
rect 29822 5966 29874 6018
rect 30942 5966 30994 6018
rect 7422 5854 7474 5906
rect 8654 5854 8706 5906
rect 8878 5854 8930 5906
rect 13246 5854 13298 5906
rect 14142 5854 14194 5906
rect 14366 5854 14418 5906
rect 15710 5854 15762 5906
rect 15934 5854 15986 5906
rect 17390 5854 17442 5906
rect 17838 5854 17890 5906
rect 18846 5854 18898 5906
rect 19294 5854 19346 5906
rect 21646 5854 21698 5906
rect 21758 5854 21810 5906
rect 22654 5854 22706 5906
rect 24446 5854 24498 5906
rect 25342 5854 25394 5906
rect 25566 5854 25618 5906
rect 26126 5854 26178 5906
rect 26462 5854 26514 5906
rect 27022 5854 27074 5906
rect 27694 5854 27746 5906
rect 29038 5854 29090 5906
rect 30046 5854 30098 5906
rect 30606 5854 30658 5906
rect 31166 5854 31218 5906
rect 31502 5854 31554 5906
rect 31950 5854 32002 5906
rect 33070 5854 33122 5906
rect 33630 5854 33682 5906
rect 8990 5742 9042 5794
rect 14590 5742 14642 5794
rect 18398 5742 18450 5794
rect 21422 5742 21474 5794
rect 22542 5742 22594 5794
rect 24334 5742 24386 5794
rect 26910 5742 26962 5794
rect 27806 5742 27858 5794
rect 30718 5742 30770 5794
rect 31726 5742 31778 5794
rect 33182 5742 33234 5794
rect 3390 5630 3442 5682
rect 7198 5630 7250 5682
rect 24110 5630 24162 5682
rect 27358 5630 27410 5682
rect 27470 5630 27522 5682
rect 29038 5630 29090 5682
rect 32062 5630 32114 5682
rect 5372 5462 5424 5514
rect 5476 5462 5528 5514
rect 5580 5462 5632 5514
rect 13688 5462 13740 5514
rect 13792 5462 13844 5514
rect 13896 5462 13948 5514
rect 22004 5462 22056 5514
rect 22108 5462 22160 5514
rect 22212 5462 22264 5514
rect 30320 5462 30372 5514
rect 30424 5462 30476 5514
rect 30528 5462 30580 5514
rect 3950 5294 4002 5346
rect 4510 5294 4562 5346
rect 13582 5294 13634 5346
rect 21982 5294 22034 5346
rect 27358 5294 27410 5346
rect 27694 5294 27746 5346
rect 29262 5294 29314 5346
rect 3390 5182 3442 5234
rect 10782 5182 10834 5234
rect 10894 5182 10946 5234
rect 12126 5182 12178 5234
rect 19182 5182 19234 5234
rect 21646 5182 21698 5234
rect 24110 5182 24162 5234
rect 26238 5182 26290 5234
rect 30494 5182 30546 5234
rect 32062 5182 32114 5234
rect 34190 5182 34242 5234
rect 2158 5070 2210 5122
rect 2718 5070 2770 5122
rect 3614 5070 3666 5122
rect 4286 5070 4338 5122
rect 4846 5070 4898 5122
rect 5966 5070 6018 5122
rect 7422 5070 7474 5122
rect 8094 5070 8146 5122
rect 8878 5070 8930 5122
rect 9102 5070 9154 5122
rect 10110 5070 10162 5122
rect 11230 5070 11282 5122
rect 11790 5070 11842 5122
rect 12798 5070 12850 5122
rect 13470 5070 13522 5122
rect 13918 5070 13970 5122
rect 15934 5070 15986 5122
rect 18174 5070 18226 5122
rect 21870 5070 21922 5122
rect 22766 5070 22818 5122
rect 23326 5070 23378 5122
rect 27022 5070 27074 5122
rect 27358 5070 27410 5122
rect 29486 5070 29538 5122
rect 29710 5070 29762 5122
rect 30270 5070 30322 5122
rect 30718 5070 30770 5122
rect 30942 5070 30994 5122
rect 31278 5070 31330 5122
rect 2382 4958 2434 5010
rect 3054 4958 3106 5010
rect 5070 4958 5122 5010
rect 7198 4958 7250 5010
rect 7870 4958 7922 5010
rect 9438 4958 9490 5010
rect 9662 4958 9714 5010
rect 12686 4958 12738 5010
rect 14030 4958 14082 5010
rect 17726 4958 17778 5010
rect 21534 4958 21586 5010
rect 4286 4846 4338 4898
rect 6190 4846 6242 4898
rect 6302 4846 6354 4898
rect 14142 4846 14194 4898
rect 29598 4846 29650 4898
rect 9530 4678 9582 4730
rect 9634 4678 9686 4730
rect 9738 4678 9790 4730
rect 17846 4678 17898 4730
rect 17950 4678 18002 4730
rect 18054 4678 18106 4730
rect 26162 4678 26214 4730
rect 26266 4678 26318 4730
rect 26370 4678 26422 4730
rect 34478 4678 34530 4730
rect 34582 4678 34634 4730
rect 34686 4678 34738 4730
rect 4734 4510 4786 4562
rect 6078 4510 6130 4562
rect 6414 4510 6466 4562
rect 7086 4510 7138 4562
rect 7534 4510 7586 4562
rect 7758 4510 7810 4562
rect 11342 4510 11394 4562
rect 11902 4510 11954 4562
rect 17502 4510 17554 4562
rect 18622 4510 18674 4562
rect 22766 4510 22818 4562
rect 33070 4510 33122 4562
rect 2494 4398 2546 4450
rect 5182 4398 5234 4450
rect 5630 4398 5682 4450
rect 6862 4398 6914 4450
rect 7422 4398 7474 4450
rect 8318 4398 8370 4450
rect 8654 4398 8706 4450
rect 8990 4398 9042 4450
rect 9550 4398 9602 4450
rect 13358 4398 13410 4450
rect 16046 4398 16098 4450
rect 18846 4398 18898 4450
rect 27918 4398 27970 4450
rect 31166 4398 31218 4450
rect 1822 4286 1874 4338
rect 5518 4286 5570 4338
rect 5742 4286 5794 4338
rect 6750 4286 6802 4338
rect 8094 4286 8146 4338
rect 9774 4286 9826 4338
rect 11006 4286 11058 4338
rect 12126 4286 12178 4338
rect 12574 4286 12626 4338
rect 16158 4286 16210 4338
rect 16382 4286 16434 4338
rect 16606 4286 16658 4338
rect 19182 4286 19234 4338
rect 19630 4286 19682 4338
rect 23102 4286 23154 4338
rect 23774 4286 23826 4338
rect 24222 4286 24274 4338
rect 28590 4286 28642 4338
rect 31950 4286 32002 4338
rect 33406 4286 33458 4338
rect 33630 4286 33682 4338
rect 10782 4174 10834 4226
rect 15486 4174 15538 4226
rect 19070 4174 19122 4226
rect 20302 4174 20354 4226
rect 22430 4174 22482 4226
rect 23326 4174 23378 4226
rect 23662 4174 23714 4226
rect 25790 4174 25842 4226
rect 29038 4174 29090 4226
rect 23998 4062 24050 4114
rect 5372 3894 5424 3946
rect 5476 3894 5528 3946
rect 5580 3894 5632 3946
rect 13688 3894 13740 3946
rect 13792 3894 13844 3946
rect 13896 3894 13948 3946
rect 22004 3894 22056 3946
rect 22108 3894 22160 3946
rect 22212 3894 22264 3946
rect 30320 3894 30372 3946
rect 30424 3894 30476 3946
rect 30528 3894 30580 3946
rect 6638 3726 6690 3778
rect 8206 3726 8258 3778
rect 14926 3726 14978 3778
rect 15262 3726 15314 3778
rect 5742 3614 5794 3666
rect 8318 3614 8370 3666
rect 10222 3614 10274 3666
rect 12462 3614 12514 3666
rect 15486 3614 15538 3666
rect 16942 3614 16994 3666
rect 19070 3614 19122 3666
rect 21534 3614 21586 3666
rect 23662 3614 23714 3666
rect 24558 3614 24610 3666
rect 24670 3614 24722 3666
rect 32958 3614 33010 3666
rect 6526 3502 6578 3554
rect 9550 3502 9602 3554
rect 19742 3502 19794 3554
rect 20750 3502 20802 3554
rect 24894 3502 24946 3554
rect 25230 3502 25282 3554
rect 31614 3502 31666 3554
rect 32398 3502 32450 3554
rect 26910 3390 26962 3442
rect 30046 3390 30098 3442
rect 32174 3390 32226 3442
rect 9530 3110 9582 3162
rect 9634 3110 9686 3162
rect 9738 3110 9790 3162
rect 17846 3110 17898 3162
rect 17950 3110 18002 3162
rect 18054 3110 18106 3162
rect 26162 3110 26214 3162
rect 26266 3110 26318 3162
rect 26370 3110 26422 3162
rect 34478 3110 34530 3162
rect 34582 3110 34634 3162
rect 34686 3110 34738 3162
<< metal2 >>
rect 5370 32172 5634 32182
rect 5426 32116 5474 32172
rect 5530 32116 5578 32172
rect 5370 32106 5634 32116
rect 13686 32172 13950 32182
rect 13742 32116 13790 32172
rect 13846 32116 13894 32172
rect 13686 32106 13950 32116
rect 22002 32172 22266 32182
rect 22058 32116 22106 32172
rect 22162 32116 22210 32172
rect 22002 32106 22266 32116
rect 30318 32172 30582 32182
rect 30374 32116 30422 32172
rect 30478 32116 30526 32172
rect 30318 32106 30582 32116
rect 9528 31388 9792 31398
rect 9584 31332 9632 31388
rect 9688 31332 9736 31388
rect 9528 31322 9792 31332
rect 17844 31388 18108 31398
rect 17900 31332 17948 31388
rect 18004 31332 18052 31388
rect 17844 31322 18108 31332
rect 26160 31388 26424 31398
rect 26216 31332 26264 31388
rect 26320 31332 26368 31388
rect 26160 31322 26424 31332
rect 34476 31388 34740 31398
rect 34532 31332 34580 31388
rect 34636 31332 34684 31388
rect 34476 31322 34740 31332
rect 5370 30604 5634 30614
rect 5426 30548 5474 30604
rect 5530 30548 5578 30604
rect 5370 30538 5634 30548
rect 13686 30604 13950 30614
rect 13742 30548 13790 30604
rect 13846 30548 13894 30604
rect 13686 30538 13950 30548
rect 22002 30604 22266 30614
rect 22058 30548 22106 30604
rect 22162 30548 22210 30604
rect 22002 30538 22266 30548
rect 30318 30604 30582 30614
rect 30374 30548 30422 30604
rect 30478 30548 30526 30604
rect 30318 30538 30582 30548
rect 9528 29820 9792 29830
rect 9584 29764 9632 29820
rect 9688 29764 9736 29820
rect 9528 29754 9792 29764
rect 17844 29820 18108 29830
rect 17900 29764 17948 29820
rect 18004 29764 18052 29820
rect 17844 29754 18108 29764
rect 26160 29820 26424 29830
rect 26216 29764 26264 29820
rect 26320 29764 26368 29820
rect 26160 29754 26424 29764
rect 34476 29820 34740 29830
rect 34532 29764 34580 29820
rect 34636 29764 34684 29820
rect 34476 29754 34740 29764
rect 5370 29036 5634 29046
rect 5426 28980 5474 29036
rect 5530 28980 5578 29036
rect 5370 28970 5634 28980
rect 13686 29036 13950 29046
rect 13742 28980 13790 29036
rect 13846 28980 13894 29036
rect 13686 28970 13950 28980
rect 22002 29036 22266 29046
rect 22058 28980 22106 29036
rect 22162 28980 22210 29036
rect 22002 28970 22266 28980
rect 30318 29036 30582 29046
rect 30374 28980 30422 29036
rect 30478 28980 30526 29036
rect 30318 28970 30582 28980
rect 11228 28756 11284 28766
rect 11228 28754 11732 28756
rect 11228 28702 11230 28754
rect 11282 28702 11732 28754
rect 11228 28700 11732 28702
rect 11228 28690 11284 28700
rect 8428 28642 8484 28654
rect 8428 28590 8430 28642
rect 8482 28590 8484 28642
rect 5068 27970 5124 27982
rect 5068 27918 5070 27970
rect 5122 27918 5124 27970
rect 4284 27858 4340 27870
rect 4284 27806 4286 27858
rect 4338 27806 4340 27858
rect 3612 27748 3668 27758
rect 2940 27746 3668 27748
rect 2940 27694 3614 27746
rect 3666 27694 3668 27746
rect 2940 27692 3668 27694
rect 1820 27074 1876 27086
rect 1820 27022 1822 27074
rect 1874 27022 1876 27074
rect 1820 26290 1876 27022
rect 2492 26962 2548 26974
rect 2492 26910 2494 26962
rect 2546 26910 2548 26962
rect 2492 26404 2548 26910
rect 2492 26338 2548 26348
rect 1820 26238 1822 26290
rect 1874 26238 1876 26290
rect 1820 25508 1876 26238
rect 2492 26180 2548 26190
rect 2492 26178 2660 26180
rect 2492 26126 2494 26178
rect 2546 26126 2660 26178
rect 2492 26124 2660 26126
rect 2492 26114 2548 26124
rect 2604 25730 2660 26124
rect 2604 25678 2606 25730
rect 2658 25678 2660 25730
rect 2604 25666 2660 25678
rect 2940 25730 2996 27692
rect 3612 27682 3668 27692
rect 4284 26908 4340 27806
rect 4508 27860 4564 27870
rect 4844 27860 4900 27870
rect 4508 27858 4900 27860
rect 4508 27806 4510 27858
rect 4562 27806 4846 27858
rect 4898 27806 4900 27858
rect 4508 27804 4900 27806
rect 4508 27794 4564 27804
rect 4844 27794 4900 27804
rect 4620 27188 4676 27198
rect 4956 27188 5012 27198
rect 5068 27188 5124 27918
rect 5180 27858 5236 27870
rect 5180 27806 5182 27858
rect 5234 27806 5236 27858
rect 5180 27300 5236 27806
rect 8428 27860 8484 28590
rect 9100 28532 9156 28542
rect 9100 28530 9940 28532
rect 9100 28478 9102 28530
rect 9154 28478 9940 28530
rect 9100 28476 9940 28478
rect 9100 28466 9156 28476
rect 9528 28252 9792 28262
rect 9584 28196 9632 28252
rect 9688 28196 9736 28252
rect 9528 28186 9792 28196
rect 5370 27468 5634 27478
rect 5426 27412 5474 27468
rect 5530 27412 5578 27468
rect 5370 27402 5634 27412
rect 5180 27234 5236 27244
rect 5852 27300 5908 27310
rect 5852 27206 5908 27244
rect 4620 27186 5124 27188
rect 4620 27134 4622 27186
rect 4674 27134 4958 27186
rect 5010 27134 5124 27186
rect 4620 27132 5124 27134
rect 4620 27122 4676 27132
rect 4956 27122 5012 27132
rect 5964 27076 6020 27086
rect 5964 26982 6020 27020
rect 6188 27074 6244 27086
rect 6188 27022 6190 27074
rect 6242 27022 6244 27074
rect 4956 26964 5012 26974
rect 4284 26852 4564 26908
rect 2940 25678 2942 25730
rect 2994 25678 2996 25730
rect 2940 25666 2996 25678
rect 3276 26404 3332 26414
rect 3276 25730 3332 26348
rect 3276 25678 3278 25730
rect 3330 25678 3332 25730
rect 3276 25666 3332 25678
rect 4508 26180 4564 26852
rect 4620 26180 4676 26190
rect 4508 26178 4676 26180
rect 4508 26126 4622 26178
rect 4674 26126 4676 26178
rect 4508 26124 4676 26126
rect 1820 23156 1876 25452
rect 2604 25508 2660 25518
rect 3276 25508 3332 25518
rect 2604 25506 3332 25508
rect 2604 25454 2606 25506
rect 2658 25454 3278 25506
rect 3330 25454 3332 25506
rect 2604 25452 3332 25454
rect 2044 23156 2100 23166
rect 1820 23154 2100 23156
rect 1820 23102 2046 23154
rect 2098 23102 2100 23154
rect 1820 23100 2100 23102
rect 1820 22372 1876 22382
rect 2044 22372 2100 23100
rect 1820 22370 2100 22372
rect 1820 22318 1822 22370
rect 1874 22318 2100 22370
rect 1820 22316 2100 22318
rect 1820 20018 1876 22316
rect 2492 22260 2548 22270
rect 2492 22166 2548 22204
rect 2604 21026 2660 25452
rect 3276 24948 3332 25452
rect 3612 25396 3668 25406
rect 4060 25396 4116 25406
rect 3612 25394 4116 25396
rect 3612 25342 3614 25394
rect 3666 25342 4062 25394
rect 4114 25342 4116 25394
rect 3612 25340 4116 25342
rect 3612 25330 3668 25340
rect 4060 25330 4116 25340
rect 3276 24882 3332 24892
rect 4060 24836 4116 24846
rect 4060 23604 4116 24780
rect 4396 24722 4452 24734
rect 4396 24670 4398 24722
rect 4450 24670 4452 24722
rect 4396 24500 4452 24670
rect 4508 24724 4564 26124
rect 4620 26114 4676 26124
rect 4956 25620 5012 26908
rect 4732 25618 5012 25620
rect 4732 25566 4958 25618
rect 5010 25566 5012 25618
rect 4732 25564 5012 25566
rect 4620 25506 4676 25518
rect 4620 25454 4622 25506
rect 4674 25454 4676 25506
rect 4620 25396 4676 25454
rect 4620 25330 4676 25340
rect 4732 24946 4788 25564
rect 4956 25554 5012 25564
rect 5068 26962 5124 26974
rect 5068 26910 5070 26962
rect 5122 26910 5124 26962
rect 5068 25396 5124 26910
rect 5068 25330 5124 25340
rect 5180 26964 5236 26974
rect 5180 26178 5236 26908
rect 5180 26126 5182 26178
rect 5234 26126 5236 26178
rect 4732 24894 4734 24946
rect 4786 24894 4788 24946
rect 4732 24882 4788 24894
rect 5068 24836 5124 24846
rect 4620 24724 4676 24734
rect 4508 24668 4620 24724
rect 4620 24658 4676 24668
rect 5068 24722 5124 24780
rect 5068 24670 5070 24722
rect 5122 24670 5124 24722
rect 5068 24658 5124 24670
rect 5180 24724 5236 26126
rect 5370 25900 5634 25910
rect 5426 25844 5474 25900
rect 5530 25844 5578 25900
rect 5370 25834 5634 25844
rect 5852 25396 5908 25406
rect 5852 24834 5908 25340
rect 5852 24782 5854 24834
rect 5906 24782 5908 24834
rect 5852 24770 5908 24782
rect 5964 24836 6020 24846
rect 5292 24724 5348 24734
rect 5180 24722 5348 24724
rect 5180 24670 5294 24722
rect 5346 24670 5348 24722
rect 5180 24668 5348 24670
rect 5292 24658 5348 24668
rect 5628 24724 5684 24734
rect 5628 24630 5684 24668
rect 4396 24434 4452 24444
rect 5370 24332 5634 24342
rect 5426 24276 5474 24332
rect 5530 24276 5578 24332
rect 5370 24266 5634 24276
rect 5068 23828 5124 23838
rect 5068 23826 5572 23828
rect 5068 23774 5070 23826
rect 5122 23774 5572 23826
rect 5068 23772 5572 23774
rect 5068 23762 5124 23772
rect 4060 23538 4116 23548
rect 4844 23714 4900 23726
rect 4844 23662 4846 23714
rect 4898 23662 4900 23714
rect 2828 23044 2884 23054
rect 4844 23044 4900 23662
rect 4956 23714 5012 23726
rect 4956 23662 4958 23714
rect 5010 23662 5012 23714
rect 4956 23268 5012 23662
rect 4956 23202 5012 23212
rect 5404 23604 5460 23614
rect 4956 23044 5012 23054
rect 4844 23042 5012 23044
rect 4844 22990 4958 23042
rect 5010 22990 5012 23042
rect 4844 22988 5012 22990
rect 2828 22950 2884 22988
rect 4956 22932 5012 22988
rect 5292 23042 5348 23054
rect 5292 22990 5294 23042
rect 5346 22990 5348 23042
rect 5292 22932 5348 22990
rect 4956 22876 5348 22932
rect 5404 22932 5460 23548
rect 5516 23156 5572 23772
rect 5852 23380 5908 23390
rect 5964 23380 6020 24780
rect 6188 24500 6244 27022
rect 6748 27076 6804 27086
rect 6748 26982 6804 27020
rect 7420 27074 7476 27086
rect 7420 27022 7422 27074
rect 7474 27022 7476 27074
rect 6300 26962 6356 26974
rect 6300 26910 6302 26962
rect 6354 26910 6356 26962
rect 6300 26404 6356 26910
rect 6300 26338 6356 26348
rect 6412 26964 6468 26974
rect 6188 24434 6244 24444
rect 6300 24946 6356 24958
rect 6300 24894 6302 24946
rect 6354 24894 6356 24946
rect 5852 23378 6020 23380
rect 5852 23326 5854 23378
rect 5906 23326 6020 23378
rect 5852 23324 6020 23326
rect 5852 23314 5908 23324
rect 6188 23268 6244 23278
rect 5516 23154 6020 23156
rect 5516 23102 5518 23154
rect 5570 23102 6020 23154
rect 5516 23100 6020 23102
rect 5516 23090 5572 23100
rect 5404 22876 5796 22932
rect 5180 22596 5236 22876
rect 5370 22764 5634 22774
rect 5426 22708 5474 22764
rect 5530 22708 5578 22764
rect 5370 22698 5634 22708
rect 5180 22540 5572 22596
rect 4620 22482 4676 22494
rect 4620 22430 4622 22482
rect 4674 22430 4676 22482
rect 3612 22372 3668 22382
rect 3612 21810 3668 22316
rect 3612 21758 3614 21810
rect 3666 21758 3668 21810
rect 3612 21746 3668 21758
rect 3948 21700 4004 21710
rect 3948 21606 4004 21644
rect 4620 21700 4676 22430
rect 5516 21810 5572 22540
rect 5740 22594 5796 22876
rect 5964 22596 6020 23100
rect 6188 23154 6244 23212
rect 6188 23102 6190 23154
rect 6242 23102 6244 23154
rect 6188 23090 6244 23102
rect 5740 22542 5742 22594
rect 5794 22542 5796 22594
rect 5740 22530 5796 22542
rect 5852 22594 6020 22596
rect 5852 22542 5966 22594
rect 6018 22542 6020 22594
rect 5852 22540 6020 22542
rect 5628 22260 5684 22270
rect 5628 22166 5684 22204
rect 5852 21924 5908 22540
rect 5964 22530 6020 22540
rect 6076 22372 6132 22382
rect 6076 22278 6132 22316
rect 5516 21758 5518 21810
rect 5570 21758 5572 21810
rect 5516 21746 5572 21758
rect 5628 21868 5908 21924
rect 4620 21606 4676 21644
rect 5404 21700 5460 21710
rect 5404 21606 5460 21644
rect 2604 20974 2606 21026
rect 2658 20974 2660 21026
rect 2604 20962 2660 20974
rect 3388 21586 3444 21598
rect 3388 21534 3390 21586
rect 3442 21534 3444 21586
rect 3276 20804 3332 20814
rect 3276 20710 3332 20748
rect 2380 20580 2436 20590
rect 2380 20486 2436 20524
rect 2492 20578 2548 20590
rect 2492 20526 2494 20578
rect 2546 20526 2548 20578
rect 1820 19966 1822 20018
rect 1874 19966 1876 20018
rect 1820 19234 1876 19966
rect 2492 19346 2548 20526
rect 2940 20580 2996 20590
rect 2940 20486 2996 20524
rect 3388 20580 3444 21534
rect 3388 20514 3444 20524
rect 3612 21586 3668 21598
rect 3612 21534 3614 21586
rect 3666 21534 3668 21586
rect 3612 20578 3668 21534
rect 4396 21586 4452 21598
rect 4396 21534 4398 21586
rect 4450 21534 4452 21586
rect 4396 20916 4452 21534
rect 4508 21586 4564 21598
rect 5628 21588 5684 21868
rect 4508 21534 4510 21586
rect 4562 21534 4564 21586
rect 4508 21028 4564 21534
rect 5516 21532 5684 21588
rect 5740 21586 5796 21598
rect 5740 21534 5742 21586
rect 5794 21534 5796 21586
rect 5068 21476 5124 21486
rect 5516 21476 5572 21532
rect 5068 21474 5572 21476
rect 5068 21422 5070 21474
rect 5122 21422 5572 21474
rect 5068 21420 5572 21422
rect 5068 21410 5124 21420
rect 5370 21196 5634 21206
rect 5426 21140 5474 21196
rect 5530 21140 5578 21196
rect 5370 21130 5634 21140
rect 4508 20972 4676 21028
rect 4396 20860 4564 20916
rect 3948 20692 4004 20702
rect 3948 20598 4004 20636
rect 3612 20526 3614 20578
rect 3666 20526 3668 20578
rect 3612 20020 3668 20526
rect 4284 20580 4340 20590
rect 4284 20486 4340 20524
rect 4396 20578 4452 20590
rect 4396 20526 4398 20578
rect 4450 20526 4452 20578
rect 4396 20132 4452 20526
rect 4396 20066 4452 20076
rect 4508 20578 4564 20860
rect 4508 20526 4510 20578
rect 4562 20526 4564 20578
rect 3612 19954 3668 19964
rect 4508 20020 4564 20526
rect 4508 19954 4564 19964
rect 4620 20804 4676 20972
rect 4732 20804 4788 20814
rect 4620 20748 4732 20804
rect 2604 19908 2660 19918
rect 2604 19814 2660 19852
rect 2492 19294 2494 19346
rect 2546 19294 2548 19346
rect 2492 19282 2548 19294
rect 4620 19346 4676 20748
rect 4732 20738 4788 20748
rect 4956 20802 5012 20814
rect 4956 20750 4958 20802
rect 5010 20750 5012 20802
rect 4844 20692 4900 20702
rect 4732 19908 4788 19918
rect 4844 19908 4900 20636
rect 4732 19906 4900 19908
rect 4732 19854 4734 19906
rect 4786 19854 4900 19906
rect 4732 19852 4900 19854
rect 4732 19842 4788 19852
rect 4956 19460 5012 20750
rect 5628 20802 5684 20814
rect 5628 20750 5630 20802
rect 5682 20750 5684 20802
rect 5068 20580 5124 20590
rect 5068 20130 5124 20524
rect 5628 20468 5684 20750
rect 5740 20690 5796 21534
rect 5740 20638 5742 20690
rect 5794 20638 5796 20690
rect 5740 20626 5796 20638
rect 6300 20468 6356 24894
rect 6412 24834 6468 26908
rect 6636 26962 6692 26974
rect 6636 26910 6638 26962
rect 6690 26910 6692 26962
rect 6636 24836 6692 26910
rect 6860 26964 6916 26974
rect 6860 26870 6916 26908
rect 7308 26404 7364 26414
rect 7308 26310 7364 26348
rect 6412 24782 6414 24834
rect 6466 24782 6468 24834
rect 6412 24770 6468 24782
rect 6524 24780 6636 24836
rect 6412 23156 6468 23166
rect 6524 23156 6580 24780
rect 6636 24770 6692 24780
rect 7084 25508 7140 25518
rect 6412 23154 6580 23156
rect 6412 23102 6414 23154
rect 6466 23102 6580 23154
rect 6412 23100 6580 23102
rect 6636 24500 6692 24510
rect 6636 23156 6692 24444
rect 6412 23090 6468 23100
rect 6636 23062 6692 23100
rect 7084 23938 7140 25452
rect 7420 25508 7476 27022
rect 8092 26962 8148 26974
rect 8428 26964 8484 27804
rect 8092 26910 8094 26962
rect 8146 26910 8148 26962
rect 8092 26516 8148 26910
rect 8092 26450 8148 26460
rect 8316 26908 8484 26964
rect 7420 25442 7476 25452
rect 7980 26292 8036 26302
rect 8316 26292 8372 26908
rect 9528 26684 9792 26694
rect 9584 26628 9632 26684
rect 9688 26628 9736 26684
rect 9528 26618 9792 26628
rect 7980 26290 8372 26292
rect 7980 26238 7982 26290
rect 8034 26238 8372 26290
rect 7980 26236 8372 26238
rect 8876 26516 8932 26526
rect 7980 25508 8036 26236
rect 7980 25442 8036 25452
rect 7756 25394 7812 25406
rect 7756 25342 7758 25394
rect 7810 25342 7812 25394
rect 7756 24164 7812 25342
rect 8876 24946 8932 26460
rect 9884 26514 9940 28476
rect 10220 27860 10276 27870
rect 10220 27766 10276 27804
rect 11004 27748 11060 27758
rect 11004 27654 11060 27692
rect 9884 26462 9886 26514
rect 9938 26462 9940 26514
rect 9884 26450 9940 26462
rect 10220 27186 10276 27198
rect 10220 27134 10222 27186
rect 10274 27134 10276 27186
rect 9996 26178 10052 26190
rect 9996 26126 9998 26178
rect 10050 26126 10052 26178
rect 9884 25618 9940 25630
rect 9884 25566 9886 25618
rect 9938 25566 9940 25618
rect 9528 25116 9792 25126
rect 9584 25060 9632 25116
rect 9688 25060 9736 25116
rect 9528 25050 9792 25060
rect 8876 24894 8878 24946
rect 8930 24894 8932 24946
rect 8876 24882 8932 24894
rect 8988 24610 9044 24622
rect 8988 24558 8990 24610
rect 9042 24558 9044 24610
rect 7756 24098 7812 24108
rect 8876 24164 8932 24174
rect 7084 23886 7086 23938
rect 7138 23886 7140 23938
rect 6748 23044 6804 23054
rect 6748 22950 6804 22988
rect 7084 22484 7140 23886
rect 7868 23828 7924 23838
rect 7868 23826 8372 23828
rect 7868 23774 7870 23826
rect 7922 23774 8372 23826
rect 7868 23772 8372 23774
rect 7868 23762 7924 23772
rect 8316 23380 8372 23772
rect 8428 23380 8484 23390
rect 8316 23378 8484 23380
rect 8316 23326 8430 23378
rect 8482 23326 8484 23378
rect 8316 23324 8484 23326
rect 8428 23314 8484 23324
rect 8876 23378 8932 24108
rect 8988 24052 9044 24558
rect 8988 23986 9044 23996
rect 9528 23548 9792 23558
rect 9584 23492 9632 23548
rect 9688 23492 9736 23548
rect 9528 23482 9792 23492
rect 8876 23326 8878 23378
rect 8930 23326 8932 23378
rect 8876 23314 8932 23326
rect 9884 23266 9940 25566
rect 9996 24948 10052 26126
rect 9996 24882 10052 24892
rect 10220 24388 10276 27134
rect 11676 26964 11732 28700
rect 17844 28252 18108 28262
rect 17900 28196 17948 28252
rect 18004 28196 18052 28252
rect 17844 28186 18108 28196
rect 26160 28252 26424 28262
rect 26216 28196 26264 28252
rect 26320 28196 26368 28252
rect 26160 28186 26424 28196
rect 34476 28252 34740 28262
rect 34532 28196 34580 28252
rect 34636 28196 34684 28252
rect 34476 28186 34740 28196
rect 19292 27860 19348 27870
rect 19180 27804 19292 27860
rect 12236 27748 12292 27758
rect 13132 27748 13188 27758
rect 12236 27186 12292 27692
rect 12236 27134 12238 27186
rect 12290 27134 12292 27186
rect 12236 27122 12292 27134
rect 13020 27746 13188 27748
rect 13020 27694 13134 27746
rect 13186 27694 13188 27746
rect 13020 27692 13188 27694
rect 12012 27074 12068 27086
rect 12012 27022 12014 27074
rect 12066 27022 12068 27074
rect 11676 26908 11844 26964
rect 11788 26290 11844 26908
rect 11788 26238 11790 26290
rect 11842 26238 11844 26290
rect 11004 25396 11060 25406
rect 11004 24948 11060 25340
rect 11788 25172 11844 26238
rect 11228 25116 11844 25172
rect 10220 24322 10276 24332
rect 10892 24946 11060 24948
rect 10892 24894 11006 24946
rect 11058 24894 11060 24946
rect 10892 24892 11060 24894
rect 9996 24050 10052 24062
rect 9996 23998 9998 24050
rect 10050 23998 10052 24050
rect 9996 23604 10052 23998
rect 10892 23938 10948 24892
rect 11004 24882 11060 24892
rect 11116 24948 11172 24958
rect 11116 24854 11172 24892
rect 11228 24946 11284 25116
rect 11228 24894 11230 24946
rect 11282 24894 11284 24946
rect 11228 24882 11284 24894
rect 11788 24836 11844 25116
rect 11788 24770 11844 24780
rect 11452 24724 11508 24734
rect 11452 24722 11620 24724
rect 11452 24670 11454 24722
rect 11506 24670 11620 24722
rect 11452 24668 11620 24670
rect 11452 24658 11508 24668
rect 11116 24388 11172 24398
rect 11004 24052 11060 24062
rect 11004 23958 11060 23996
rect 11116 24052 11172 24332
rect 11116 23996 11396 24052
rect 10892 23886 10894 23938
rect 10946 23886 10948 23938
rect 10892 23874 10948 23886
rect 11116 23826 11172 23996
rect 11116 23774 11118 23826
rect 11170 23774 11172 23826
rect 11116 23762 11172 23774
rect 11228 23826 11284 23838
rect 11228 23774 11230 23826
rect 11282 23774 11284 23826
rect 9996 23538 10052 23548
rect 11228 23492 11284 23774
rect 11004 23436 11284 23492
rect 11340 23828 11396 23996
rect 9996 23380 10052 23390
rect 9996 23286 10052 23324
rect 11004 23378 11060 23436
rect 11004 23326 11006 23378
rect 11058 23326 11060 23378
rect 11004 23314 11060 23326
rect 9884 23214 9886 23266
rect 9938 23214 9940 23266
rect 8540 23042 8596 23054
rect 8540 22990 8542 23042
rect 8594 22990 8596 23042
rect 7084 22418 7140 22428
rect 7868 22484 7924 22494
rect 7868 22390 7924 22428
rect 8540 22260 8596 22990
rect 8988 23044 9044 23054
rect 8988 22950 9044 22988
rect 9884 22932 9940 23214
rect 10220 23266 10276 23278
rect 10220 23214 10222 23266
rect 10274 23214 10276 23266
rect 10220 23156 10276 23214
rect 10892 23266 10948 23278
rect 10892 23214 10894 23266
rect 10946 23214 10948 23266
rect 10332 23156 10388 23166
rect 10220 23154 10388 23156
rect 10220 23102 10334 23154
rect 10386 23102 10388 23154
rect 10220 23100 10388 23102
rect 10332 23090 10388 23100
rect 10668 23154 10724 23166
rect 10668 23102 10670 23154
rect 10722 23102 10724 23154
rect 9884 22866 9940 22876
rect 8540 22194 8596 22204
rect 9528 21980 9792 21990
rect 9584 21924 9632 21980
rect 9688 21924 9736 21980
rect 9528 21914 9792 21924
rect 10668 21812 10724 23102
rect 10892 22148 10948 23214
rect 11340 23154 11396 23772
rect 11340 23102 11342 23154
rect 11394 23102 11396 23154
rect 11340 23090 11396 23102
rect 11452 22932 11508 22942
rect 11564 22932 11620 24668
rect 11676 24722 11732 24734
rect 11676 24670 11678 24722
rect 11730 24670 11732 24722
rect 11676 24052 11732 24670
rect 12012 24612 12068 27022
rect 12460 26964 12516 26974
rect 12460 26870 12516 26908
rect 12684 26962 12740 26974
rect 12684 26910 12686 26962
rect 12738 26910 12740 26962
rect 12348 26292 12404 26302
rect 12348 26198 12404 26236
rect 12460 26180 12516 26190
rect 12460 26178 12628 26180
rect 12460 26126 12462 26178
rect 12514 26126 12628 26178
rect 12460 26124 12628 26126
rect 12460 26114 12516 26124
rect 12348 25732 12404 25742
rect 12348 25620 12404 25676
rect 12460 25620 12516 25630
rect 12348 25618 12516 25620
rect 12348 25566 12462 25618
rect 12514 25566 12516 25618
rect 12348 25564 12516 25566
rect 12460 25554 12516 25564
rect 12572 25506 12628 26124
rect 12684 25620 12740 26910
rect 12684 25554 12740 25564
rect 13020 26292 13076 27692
rect 13132 27682 13188 27692
rect 13686 27468 13950 27478
rect 13742 27412 13790 27468
rect 13846 27412 13894 27468
rect 13686 27402 13950 27412
rect 17052 27188 17108 27198
rect 16716 27186 17108 27188
rect 16716 27134 17054 27186
rect 17106 27134 17108 27186
rect 16716 27132 17108 27134
rect 12572 25454 12574 25506
rect 12626 25454 12628 25506
rect 12572 25442 12628 25454
rect 13020 25508 13076 26236
rect 13132 27076 13188 27086
rect 13132 26290 13188 27020
rect 14252 27076 14308 27086
rect 14252 26982 14308 27020
rect 14924 26964 14980 26974
rect 14924 26962 15092 26964
rect 14924 26910 14926 26962
rect 14978 26910 15092 26962
rect 14924 26908 15092 26910
rect 16716 26908 16772 27132
rect 17052 27122 17108 27132
rect 14924 26898 14980 26908
rect 13132 26238 13134 26290
rect 13186 26238 13188 26290
rect 13132 26226 13188 26238
rect 13804 26180 13860 26190
rect 13804 26178 14532 26180
rect 13804 26126 13806 26178
rect 13858 26126 14532 26178
rect 13804 26124 14532 26126
rect 13804 26114 13860 26124
rect 13686 25900 13950 25910
rect 13742 25844 13790 25900
rect 13846 25844 13894 25900
rect 13686 25834 13950 25844
rect 14252 25732 14308 25742
rect 13580 25620 13636 25630
rect 13580 25526 13636 25564
rect 14140 25620 14196 25630
rect 13020 25442 13076 25452
rect 13692 25508 13748 25518
rect 12012 24546 12068 24556
rect 12124 25282 12180 25294
rect 12124 25230 12126 25282
rect 12178 25230 12180 25282
rect 12124 24500 12180 25230
rect 12348 25282 12404 25294
rect 12348 25230 12350 25282
rect 12402 25230 12404 25282
rect 12348 24948 12404 25230
rect 12348 24834 12404 24892
rect 13468 25282 13524 25294
rect 13468 25230 13470 25282
rect 13522 25230 13524 25282
rect 12348 24782 12350 24834
rect 12402 24782 12404 24834
rect 12348 24770 12404 24782
rect 13244 24834 13300 24846
rect 13244 24782 13246 24834
rect 13298 24782 13300 24834
rect 12236 24724 12292 24734
rect 12236 24630 12292 24668
rect 12572 24722 12628 24734
rect 12572 24670 12574 24722
rect 12626 24670 12628 24722
rect 12460 24612 12516 24650
rect 12460 24546 12516 24556
rect 12124 24434 12180 24444
rect 12124 24164 12180 24174
rect 11676 23938 11732 23996
rect 11676 23886 11678 23938
rect 11730 23886 11732 23938
rect 11676 23874 11732 23886
rect 11900 24162 12180 24164
rect 11900 24110 12126 24162
rect 12178 24110 12180 24162
rect 11900 24108 12180 24110
rect 12572 24164 12628 24670
rect 12684 24724 12740 24734
rect 12684 24630 12740 24668
rect 13244 24724 13300 24782
rect 13468 24836 13524 25230
rect 13468 24770 13524 24780
rect 13244 24658 13300 24668
rect 13356 24610 13412 24622
rect 13356 24558 13358 24610
rect 13410 24558 13412 24610
rect 12572 24108 13188 24164
rect 11788 23716 11844 23726
rect 11676 23604 11732 23614
rect 11676 23154 11732 23548
rect 11788 23266 11844 23660
rect 11788 23214 11790 23266
rect 11842 23214 11844 23266
rect 11788 23202 11844 23214
rect 11676 23102 11678 23154
rect 11730 23102 11732 23154
rect 11676 23090 11732 23102
rect 11564 22876 11732 22932
rect 11452 22838 11508 22876
rect 10892 22092 11172 22148
rect 10668 21746 10724 21756
rect 10780 21700 10836 21710
rect 11004 21700 11060 21710
rect 10780 21698 10948 21700
rect 10780 21646 10782 21698
rect 10834 21646 10948 21698
rect 10780 21644 10948 21646
rect 10780 21634 10836 21644
rect 10668 21586 10724 21598
rect 10668 21534 10670 21586
rect 10722 21534 10724 21586
rect 10668 20916 10724 21534
rect 10780 21364 10836 21374
rect 10780 21270 10836 21308
rect 10220 20860 10724 20916
rect 7644 20804 7700 20814
rect 7644 20710 7700 20748
rect 8204 20692 8260 20702
rect 8204 20598 8260 20636
rect 7756 20580 7812 20590
rect 5628 20412 6356 20468
rect 7644 20578 7812 20580
rect 7644 20526 7758 20578
rect 7810 20526 7812 20578
rect 7644 20524 7812 20526
rect 5068 20078 5070 20130
rect 5122 20078 5124 20130
rect 5068 20066 5124 20078
rect 5516 20132 5572 20142
rect 5292 20020 5348 20030
rect 5292 19926 5348 19964
rect 5516 20018 5572 20076
rect 5516 19966 5518 20018
rect 5570 19966 5572 20018
rect 5516 19954 5572 19966
rect 7532 20018 7588 20030
rect 7532 19966 7534 20018
rect 7586 19966 7588 20018
rect 5180 19908 5236 19918
rect 5180 19814 5236 19852
rect 6748 19908 6804 19918
rect 5370 19628 5634 19638
rect 5426 19572 5474 19628
rect 5530 19572 5578 19628
rect 5370 19562 5634 19572
rect 4956 19394 5012 19404
rect 4620 19294 4622 19346
rect 4674 19294 4676 19346
rect 4620 19282 4676 19294
rect 1820 19182 1822 19234
rect 1874 19182 1876 19234
rect 1820 19170 1876 19182
rect 5852 18562 5908 18574
rect 5852 18510 5854 18562
rect 5906 18510 5908 18562
rect 4620 18452 4676 18462
rect 4620 17778 4676 18396
rect 5628 18452 5684 18462
rect 5628 18358 5684 18396
rect 5852 18340 5908 18510
rect 6524 18562 6580 18574
rect 6524 18510 6526 18562
rect 6578 18510 6580 18562
rect 5852 18274 5908 18284
rect 6300 18450 6356 18462
rect 6300 18398 6302 18450
rect 6354 18398 6356 18450
rect 6300 18228 6356 18398
rect 6300 18162 6356 18172
rect 6412 18452 6468 18462
rect 6524 18452 6580 18510
rect 6636 18452 6692 18462
rect 6524 18396 6636 18452
rect 5370 18060 5634 18070
rect 5426 18004 5474 18060
rect 5530 18004 5578 18060
rect 5370 17994 5634 18004
rect 6412 17890 6468 18396
rect 6636 18386 6692 18396
rect 6412 17838 6414 17890
rect 6466 17838 6468 17890
rect 6412 17826 6468 17838
rect 6748 17890 6804 19852
rect 7420 19908 7476 19918
rect 7420 19814 7476 19852
rect 7084 19234 7140 19246
rect 7084 19182 7086 19234
rect 7138 19182 7140 19234
rect 6972 18788 7028 18798
rect 6748 17838 6750 17890
rect 6802 17838 6804 17890
rect 6748 17826 6804 17838
rect 6860 18338 6916 18350
rect 6860 18286 6862 18338
rect 6914 18286 6916 18338
rect 6860 18228 6916 18286
rect 4620 17726 4622 17778
rect 4674 17726 4676 17778
rect 4620 17714 4676 17726
rect 1820 17666 1876 17678
rect 1820 17614 1822 17666
rect 1874 17614 1876 17666
rect 1596 15204 1652 15214
rect 1596 4228 1652 15148
rect 1820 15092 1876 17614
rect 6188 17668 6244 17678
rect 2492 17556 2548 17566
rect 2380 17554 2548 17556
rect 2380 17502 2494 17554
rect 2546 17502 2548 17554
rect 2380 17500 2548 17502
rect 1820 14530 1876 15036
rect 2268 16098 2324 16110
rect 2268 16046 2270 16098
rect 2322 16046 2324 16098
rect 2268 15092 2324 16046
rect 2268 15026 2324 15036
rect 1820 14478 1822 14530
rect 1874 14478 1876 14530
rect 1820 14466 1876 14478
rect 2044 12180 2100 12190
rect 2044 9156 2100 12124
rect 2380 11506 2436 17500
rect 2492 17490 2548 17500
rect 5068 17444 5124 17454
rect 5068 17442 5796 17444
rect 5068 17390 5070 17442
rect 5122 17390 5796 17442
rect 5068 17388 5796 17390
rect 5068 17378 5124 17388
rect 3276 16882 3332 16894
rect 3276 16830 3278 16882
rect 3330 16830 3332 16882
rect 2940 15986 2996 15998
rect 2940 15934 2942 15986
rect 2994 15934 2996 15986
rect 2492 14418 2548 14430
rect 2492 14366 2494 14418
rect 2546 14366 2548 14418
rect 2492 13524 2548 14366
rect 2940 14308 2996 15934
rect 2940 14242 2996 14252
rect 3276 15092 3332 16830
rect 3948 16884 4004 16894
rect 3948 16790 4004 16828
rect 5068 16884 5124 16894
rect 5124 16828 5236 16884
rect 5068 16818 5124 16828
rect 5068 16660 5124 16670
rect 5068 16210 5124 16604
rect 5068 16158 5070 16210
rect 5122 16158 5124 16210
rect 5068 16146 5124 16158
rect 3276 14084 3332 15036
rect 5180 14756 5236 16828
rect 5370 16492 5634 16502
rect 5426 16436 5474 16492
rect 5530 16436 5578 16492
rect 5370 16426 5634 16436
rect 5740 16322 5796 17388
rect 6076 16772 6132 16782
rect 6188 16772 6244 17612
rect 6748 16884 6804 16894
rect 6860 16884 6916 18172
rect 6972 17108 7028 18732
rect 7084 18340 7140 19182
rect 7084 18246 7140 18284
rect 7308 19236 7364 19246
rect 7532 19236 7588 19966
rect 7308 19234 7588 19236
rect 7308 19182 7310 19234
rect 7362 19182 7588 19234
rect 7308 19180 7588 19182
rect 7308 18452 7364 19180
rect 7420 18676 7476 18686
rect 7420 18582 7476 18620
rect 7644 18564 7700 20524
rect 7756 20514 7812 20524
rect 10220 20578 10276 20860
rect 10780 20804 10836 20814
rect 10556 20690 10612 20702
rect 10556 20638 10558 20690
rect 10610 20638 10612 20690
rect 10220 20526 10222 20578
rect 10274 20526 10276 20578
rect 9528 20412 9792 20422
rect 9584 20356 9632 20412
rect 9688 20356 9736 20412
rect 9528 20346 9792 20356
rect 8204 20244 8260 20254
rect 8204 20130 8260 20188
rect 10220 20244 10276 20526
rect 10220 20178 10276 20188
rect 10444 20578 10500 20590
rect 10444 20526 10446 20578
rect 10498 20526 10500 20578
rect 8204 20078 8206 20130
rect 8258 20078 8260 20130
rect 8204 20066 8260 20078
rect 8876 20130 8932 20142
rect 8876 20078 8878 20130
rect 8930 20078 8932 20130
rect 8876 20020 8932 20078
rect 8876 19954 8932 19964
rect 9436 20020 9492 20030
rect 9996 20020 10052 20030
rect 9492 19964 9604 20020
rect 9436 19954 9492 19964
rect 7980 19908 8036 19918
rect 7980 19346 8036 19852
rect 7980 19294 7982 19346
rect 8034 19294 8036 19346
rect 7980 19282 8036 19294
rect 8652 19794 8708 19806
rect 8652 19742 8654 19794
rect 8706 19742 8708 19794
rect 8652 19236 8708 19742
rect 8428 19234 8708 19236
rect 8428 19182 8654 19234
rect 8706 19182 8708 19234
rect 8428 19180 8708 19182
rect 8204 18788 8260 18798
rect 8204 18674 8260 18732
rect 8204 18622 8206 18674
rect 8258 18622 8260 18674
rect 7308 17780 7364 18396
rect 7532 18508 7700 18564
rect 7980 18564 8036 18574
rect 7420 17780 7476 17790
rect 7308 17724 7420 17780
rect 7420 17714 7476 17724
rect 7084 17668 7140 17678
rect 7084 17574 7140 17612
rect 7196 17444 7252 17454
rect 7196 17442 7364 17444
rect 7196 17390 7198 17442
rect 7250 17390 7364 17442
rect 7196 17388 7364 17390
rect 7196 17378 7252 17388
rect 7084 17108 7140 17118
rect 6972 17106 7140 17108
rect 6972 17054 7086 17106
rect 7138 17054 7140 17106
rect 6972 17052 7140 17054
rect 7308 17108 7364 17388
rect 7420 17442 7476 17454
rect 7420 17390 7422 17442
rect 7474 17390 7476 17442
rect 7420 17332 7476 17390
rect 7420 17266 7476 17276
rect 7532 17220 7588 18508
rect 7980 18470 8036 18508
rect 7868 18450 7924 18462
rect 7868 18398 7870 18450
rect 7922 18398 7924 18450
rect 7644 18340 7700 18350
rect 7644 17666 7700 18284
rect 7644 17614 7646 17666
rect 7698 17614 7700 17666
rect 7644 17602 7700 17614
rect 7868 17668 7924 18398
rect 8092 18338 8148 18350
rect 8092 18286 8094 18338
rect 8146 18286 8148 18338
rect 8092 18116 8148 18286
rect 8092 18050 8148 18060
rect 8204 18004 8260 18622
rect 8316 18450 8372 18462
rect 8316 18398 8318 18450
rect 8370 18398 8372 18450
rect 8316 18340 8372 18398
rect 8316 18274 8372 18284
rect 8204 17938 8260 17948
rect 8428 17892 8484 19180
rect 8652 19170 8708 19180
rect 8876 19796 8932 19806
rect 8876 19234 8932 19740
rect 8988 19796 9044 19806
rect 8988 19794 9156 19796
rect 8988 19742 8990 19794
rect 9042 19742 9156 19794
rect 8988 19740 9156 19742
rect 8988 19730 9044 19740
rect 8988 19348 9044 19358
rect 8988 19254 9044 19292
rect 8876 19182 8878 19234
rect 8930 19182 8932 19234
rect 8876 18788 8932 19182
rect 9100 19124 9156 19740
rect 9548 19572 9604 19964
rect 9996 19926 10052 19964
rect 10444 20020 10500 20526
rect 10556 20356 10612 20638
rect 10780 20690 10836 20748
rect 10780 20638 10782 20690
rect 10834 20638 10836 20690
rect 10556 20300 10724 20356
rect 10444 19954 10500 19964
rect 10556 20018 10612 20030
rect 10556 19966 10558 20018
rect 10610 19966 10612 20018
rect 9660 19908 9716 19918
rect 9660 19814 9716 19852
rect 10220 19794 10276 19806
rect 10220 19742 10222 19794
rect 10274 19742 10276 19794
rect 10220 19572 10276 19742
rect 9548 19516 9828 19572
rect 9772 19458 9828 19516
rect 10220 19506 10276 19516
rect 9772 19406 9774 19458
rect 9826 19406 9828 19458
rect 9436 19348 9492 19358
rect 9212 19346 9492 19348
rect 9212 19294 9438 19346
rect 9490 19294 9492 19346
rect 9212 19292 9492 19294
rect 9212 19234 9268 19292
rect 9436 19282 9492 19292
rect 9212 19182 9214 19234
rect 9266 19182 9268 19234
rect 9212 19170 9268 19182
rect 9100 18788 9156 19068
rect 9772 19012 9828 19406
rect 10556 19348 10612 19966
rect 10668 19684 10724 20300
rect 10780 20018 10836 20638
rect 10780 19966 10782 20018
rect 10834 19966 10836 20018
rect 10780 19954 10836 19966
rect 10668 19618 10724 19628
rect 10892 19572 10948 21644
rect 11004 20914 11060 21644
rect 11116 21588 11172 22092
rect 11340 21698 11396 21710
rect 11340 21646 11342 21698
rect 11394 21646 11396 21698
rect 11340 21588 11396 21646
rect 11564 21588 11620 21598
rect 11116 21532 11396 21588
rect 11340 21252 11396 21532
rect 11340 21186 11396 21196
rect 11452 21586 11620 21588
rect 11452 21534 11566 21586
rect 11618 21534 11620 21586
rect 11452 21532 11620 21534
rect 11452 21026 11508 21532
rect 11564 21522 11620 21532
rect 11676 21474 11732 22876
rect 11900 21586 11956 24108
rect 12124 24098 12180 24108
rect 12572 23940 12628 23950
rect 12012 23828 12068 23866
rect 12572 23828 12628 23884
rect 12796 23940 12852 23950
rect 12012 23762 12068 23772
rect 12236 23772 12628 23828
rect 12684 23828 12740 23838
rect 12124 23714 12180 23726
rect 12124 23662 12126 23714
rect 12178 23662 12180 23714
rect 12124 23380 12180 23662
rect 12124 23314 12180 23324
rect 12124 23154 12180 23166
rect 12124 23102 12126 23154
rect 12178 23102 12180 23154
rect 12124 22036 12180 23102
rect 12124 21970 12180 21980
rect 11900 21534 11902 21586
rect 11954 21534 11956 21586
rect 11900 21522 11956 21534
rect 12012 21812 12068 21822
rect 11676 21422 11678 21474
rect 11730 21422 11732 21474
rect 11676 21410 11732 21422
rect 11452 20974 11454 21026
rect 11506 20974 11508 21026
rect 11452 20962 11508 20974
rect 11004 20862 11006 20914
rect 11058 20862 11060 20914
rect 11004 20850 11060 20862
rect 11340 20692 11396 20702
rect 10556 19282 10612 19292
rect 10780 19516 10948 19572
rect 11116 20690 11396 20692
rect 11116 20638 11342 20690
rect 11394 20638 11396 20690
rect 11116 20636 11396 20638
rect 10668 19236 10724 19246
rect 9772 18946 9828 18956
rect 9996 19122 10052 19134
rect 9996 19070 9998 19122
rect 10050 19070 10052 19122
rect 9528 18844 9792 18854
rect 9584 18788 9632 18844
rect 9688 18788 9736 18844
rect 8876 18732 9044 18788
rect 9100 18732 9380 18788
rect 9528 18778 9792 18788
rect 8988 18676 9044 18732
rect 8988 18620 9268 18676
rect 8764 18564 8820 18574
rect 8428 17780 8484 17836
rect 7868 17574 7924 17612
rect 8092 17778 8484 17780
rect 8092 17726 8430 17778
rect 8482 17726 8484 17778
rect 8092 17724 8484 17726
rect 7532 17164 7812 17220
rect 7420 17108 7476 17118
rect 7308 17106 7476 17108
rect 7308 17054 7422 17106
rect 7474 17054 7476 17106
rect 7308 17052 7476 17054
rect 7084 17042 7140 17052
rect 7420 17042 7476 17052
rect 6804 16828 6916 16884
rect 7532 16884 7588 16894
rect 6748 16790 6804 16828
rect 7532 16790 7588 16828
rect 6076 16770 6244 16772
rect 6076 16718 6078 16770
rect 6130 16718 6244 16770
rect 6076 16716 6244 16718
rect 6076 16706 6132 16716
rect 5740 16270 5742 16322
rect 5794 16270 5796 16322
rect 5740 16210 5796 16270
rect 5740 16158 5742 16210
rect 5794 16158 5796 16210
rect 5740 15314 5796 16158
rect 6300 16322 6356 16334
rect 6300 16270 6302 16322
rect 6354 16270 6356 16322
rect 6300 16210 6356 16270
rect 6300 16158 6302 16210
rect 6354 16158 6356 16210
rect 6300 16146 6356 16158
rect 5740 15262 5742 15314
rect 5794 15262 5796 15314
rect 5370 14924 5634 14934
rect 5426 14868 5474 14924
rect 5530 14868 5578 14924
rect 5370 14858 5634 14868
rect 5180 14700 5348 14756
rect 4620 14644 4676 14654
rect 4620 14550 4676 14588
rect 3276 14018 3332 14028
rect 3500 14308 3556 14318
rect 2492 13458 2548 13468
rect 2828 13076 2884 13086
rect 2828 12180 2884 13020
rect 3388 12740 3444 12750
rect 3500 12740 3556 14252
rect 5068 14306 5124 14318
rect 5068 14254 5070 14306
rect 5122 14254 5124 14306
rect 5068 14084 5124 14254
rect 5068 14018 5124 14028
rect 5292 13524 5348 14700
rect 5628 14644 5684 14654
rect 5628 14532 5684 14588
rect 5404 14530 5684 14532
rect 5404 14478 5630 14530
rect 5682 14478 5684 14530
rect 5404 14476 5684 14478
rect 5404 13746 5460 14476
rect 5628 14466 5684 14476
rect 5740 14084 5796 15262
rect 6412 15202 6468 15214
rect 6412 15150 6414 15202
rect 6466 15150 6468 15202
rect 5964 14308 6020 14346
rect 5964 14242 6020 14252
rect 5964 14084 6020 14094
rect 5740 14028 5964 14084
rect 5404 13694 5406 13746
rect 5458 13694 5460 13746
rect 5404 13682 5460 13694
rect 5628 13746 5684 13758
rect 5628 13694 5630 13746
rect 5682 13694 5684 13746
rect 5628 13636 5684 13694
rect 5852 13636 5908 13646
rect 5628 13570 5684 13580
rect 5740 13634 5908 13636
rect 5740 13582 5854 13634
rect 5906 13582 5908 13634
rect 5740 13580 5908 13582
rect 5180 13468 5348 13524
rect 5068 13188 5124 13198
rect 3612 13132 4452 13188
rect 3612 12962 3668 13132
rect 4396 13076 4452 13132
rect 4620 13076 4676 13086
rect 4396 13074 4676 13076
rect 4396 13022 4622 13074
rect 4674 13022 4676 13074
rect 4396 13020 4676 13022
rect 4620 13010 4676 13020
rect 3612 12910 3614 12962
rect 3666 12910 3668 12962
rect 3612 12898 3668 12910
rect 4284 12962 4340 12974
rect 4284 12910 4286 12962
rect 4338 12910 4340 12962
rect 3724 12740 3780 12750
rect 3500 12738 3780 12740
rect 3500 12686 3726 12738
rect 3778 12686 3780 12738
rect 3500 12684 3780 12686
rect 2828 12086 2884 12124
rect 3164 12290 3220 12302
rect 3164 12238 3166 12290
rect 3218 12238 3220 12290
rect 3164 11620 3220 12238
rect 3388 11732 3444 12684
rect 3724 12674 3780 12684
rect 3836 12738 3892 12750
rect 3836 12686 3838 12738
rect 3890 12686 3892 12738
rect 3836 12404 3892 12686
rect 4172 12404 4228 12414
rect 3836 12402 4228 12404
rect 3836 12350 4174 12402
rect 4226 12350 4228 12402
rect 3836 12348 4228 12350
rect 4172 12338 4228 12348
rect 3612 12292 3668 12302
rect 3612 12198 3668 12236
rect 3500 12180 3556 12190
rect 3500 12086 3556 12124
rect 3836 12180 3892 12190
rect 3836 12178 4004 12180
rect 3836 12126 3838 12178
rect 3890 12126 4004 12178
rect 3836 12124 4004 12126
rect 3836 12114 3892 12124
rect 3948 11956 4004 12124
rect 3388 11676 3556 11732
rect 3164 11564 3444 11620
rect 2380 11454 2382 11506
rect 2434 11454 2436 11506
rect 2380 11442 2436 11454
rect 3052 11508 3108 11518
rect 3052 11414 3108 11452
rect 2156 11396 2212 11406
rect 3276 11396 3332 11406
rect 2156 11302 2212 11340
rect 3164 11394 3332 11396
rect 3164 11342 3278 11394
rect 3330 11342 3332 11394
rect 3164 11340 3332 11342
rect 2268 11172 2324 11182
rect 2044 9090 2100 9100
rect 2156 11170 2324 11172
rect 2156 11118 2270 11170
rect 2322 11118 2324 11170
rect 2156 11116 2324 11118
rect 2156 8708 2212 11116
rect 2268 11106 2324 11116
rect 2492 11170 2548 11182
rect 2492 11118 2494 11170
rect 2546 11118 2548 11170
rect 2492 10836 2548 11118
rect 2604 11172 2660 11182
rect 2604 11078 2660 11116
rect 2492 10780 2884 10836
rect 2716 10612 2772 10622
rect 2268 10610 2772 10612
rect 2268 10558 2718 10610
rect 2770 10558 2772 10610
rect 2268 10556 2772 10558
rect 2268 10050 2324 10556
rect 2716 10546 2772 10556
rect 2828 10500 2884 10780
rect 3052 10610 3108 10622
rect 3052 10558 3054 10610
rect 3106 10558 3108 10610
rect 2940 10500 2996 10510
rect 2828 10498 2996 10500
rect 2828 10446 2942 10498
rect 2994 10446 2996 10498
rect 2828 10444 2996 10446
rect 2940 10434 2996 10444
rect 2716 10052 2772 10062
rect 2268 9998 2270 10050
rect 2322 9998 2324 10050
rect 2268 9986 2324 9998
rect 2380 9996 2716 10052
rect 2156 8642 2212 8652
rect 2156 7586 2212 7598
rect 2156 7534 2158 7586
rect 2210 7534 2212 7586
rect 2156 7364 2212 7534
rect 2156 7298 2212 7308
rect 2380 7140 2436 9996
rect 2716 9958 2772 9996
rect 2604 9828 2660 9838
rect 2492 9156 2548 9166
rect 2492 9062 2548 9100
rect 2604 8034 2660 9772
rect 2940 9826 2996 9838
rect 2940 9774 2942 9826
rect 2994 9774 2996 9826
rect 2940 9268 2996 9774
rect 3052 9604 3108 10558
rect 3164 10052 3220 11340
rect 3276 11330 3332 11340
rect 3388 11172 3444 11564
rect 3276 11116 3444 11172
rect 3500 11396 3556 11676
rect 3948 11620 4004 11900
rect 4284 11788 4340 12910
rect 5068 12962 5124 13132
rect 5068 12910 5070 12962
rect 5122 12910 5124 12962
rect 5068 12898 5124 12910
rect 4508 12740 4564 12750
rect 4732 12740 4788 12750
rect 4508 12738 4676 12740
rect 4508 12686 4510 12738
rect 4562 12686 4676 12738
rect 4508 12684 4676 12686
rect 4508 12674 4564 12684
rect 4508 12292 4564 12302
rect 4172 11732 4340 11788
rect 4396 12178 4452 12190
rect 4396 12126 4398 12178
rect 4450 12126 4452 12178
rect 4396 12068 4452 12126
rect 4508 12178 4564 12236
rect 4508 12126 4510 12178
rect 4562 12126 4564 12178
rect 4508 12114 4564 12126
rect 4396 11788 4452 12012
rect 4620 11844 4676 12684
rect 4732 12646 4788 12684
rect 4396 11732 4564 11788
rect 4620 11778 4676 11788
rect 4732 12180 4788 12190
rect 4732 11788 4788 12124
rect 4956 12180 5012 12190
rect 4956 12086 5012 12124
rect 4732 11732 4900 11788
rect 4172 11620 4228 11732
rect 4508 11666 4564 11676
rect 4172 11564 4340 11620
rect 3948 11554 4004 11564
rect 4284 11506 4340 11564
rect 4284 11454 4286 11506
rect 4338 11454 4340 11506
rect 4284 11442 4340 11454
rect 3276 11060 3332 11116
rect 3276 10834 3332 11004
rect 3276 10782 3278 10834
rect 3330 10782 3332 10834
rect 3276 10770 3332 10782
rect 3500 10724 3556 11340
rect 3612 11396 3668 11406
rect 4172 11396 4228 11406
rect 3612 11394 4228 11396
rect 3612 11342 3614 11394
rect 3666 11342 4174 11394
rect 4226 11342 4228 11394
rect 3612 11340 4228 11342
rect 3612 11330 3668 11340
rect 4172 11330 4228 11340
rect 4284 11284 4340 11294
rect 3612 11172 3668 11182
rect 3612 10836 3668 11116
rect 3724 11172 3780 11182
rect 3724 11170 4004 11172
rect 3724 11118 3726 11170
rect 3778 11118 4004 11170
rect 3724 11116 4004 11118
rect 3724 11106 3780 11116
rect 3724 10836 3780 10846
rect 3612 10834 3780 10836
rect 3612 10782 3726 10834
rect 3778 10782 3780 10834
rect 3612 10780 3780 10782
rect 3724 10770 3780 10780
rect 3500 10668 3668 10724
rect 3612 10612 3668 10668
rect 3836 10722 3892 10734
rect 3836 10670 3838 10722
rect 3890 10670 3892 10722
rect 3836 10612 3892 10670
rect 3612 10556 3892 10612
rect 3612 10388 3668 10398
rect 3388 10386 3668 10388
rect 3388 10334 3614 10386
rect 3666 10334 3668 10386
rect 3388 10332 3668 10334
rect 3276 10052 3332 10062
rect 3164 9996 3276 10052
rect 3276 9986 3332 9996
rect 3164 9828 3220 9838
rect 3164 9734 3220 9772
rect 3052 9538 3108 9548
rect 2940 9202 2996 9212
rect 3388 9266 3444 10332
rect 3612 10322 3668 10332
rect 3948 10276 4004 11116
rect 4284 10724 4340 11228
rect 4508 11282 4564 11294
rect 4508 11230 4510 11282
rect 4562 11230 4564 11282
rect 4284 10388 4340 10668
rect 4396 11170 4452 11182
rect 4396 11118 4398 11170
rect 4450 11118 4452 11170
rect 4396 10612 4452 11118
rect 4508 11060 4564 11230
rect 4620 11284 4676 11294
rect 4620 11190 4676 11228
rect 4508 11004 4788 11060
rect 4732 10834 4788 11004
rect 4732 10782 4734 10834
rect 4786 10782 4788 10834
rect 4732 10770 4788 10782
rect 4396 10546 4452 10556
rect 4284 10332 4452 10388
rect 3948 10220 4340 10276
rect 3948 10052 4004 10062
rect 3500 9716 3556 9726
rect 3500 9622 3556 9660
rect 3948 9714 4004 9996
rect 3948 9662 3950 9714
rect 4002 9662 4004 9714
rect 3948 9650 4004 9662
rect 3612 9604 3668 9614
rect 3612 9510 3668 9548
rect 3724 9604 3780 9614
rect 3724 9602 3892 9604
rect 3724 9550 3726 9602
rect 3778 9550 3892 9602
rect 3724 9548 3892 9550
rect 3724 9538 3780 9548
rect 3388 9214 3390 9266
rect 3442 9214 3444 9266
rect 3388 9202 3444 9214
rect 3500 9492 3556 9502
rect 2828 9156 2884 9166
rect 2828 9062 2884 9100
rect 3164 9042 3220 9054
rect 3164 8990 3166 9042
rect 3218 8990 3220 9042
rect 3164 8428 3220 8990
rect 3500 9042 3556 9436
rect 3836 9268 3892 9548
rect 3836 9212 4116 9268
rect 3500 8990 3502 9042
rect 3554 8990 3556 9042
rect 3500 8978 3556 8990
rect 3612 9044 3668 9054
rect 3724 9044 3780 9054
rect 3668 9042 3780 9044
rect 3668 8990 3726 9042
rect 3778 8990 3780 9042
rect 3668 8988 3780 8990
rect 2716 8372 3220 8428
rect 2716 8370 2772 8372
rect 2716 8318 2718 8370
rect 2770 8318 2772 8370
rect 2716 8306 2772 8318
rect 3164 8260 3220 8270
rect 2940 8258 3220 8260
rect 2940 8206 3166 8258
rect 3218 8206 3220 8258
rect 2940 8204 3220 8206
rect 2828 8148 2884 8158
rect 2828 8054 2884 8092
rect 2604 7982 2606 8034
rect 2658 7982 2660 8034
rect 2492 7812 2548 7822
rect 2492 7586 2548 7756
rect 2492 7534 2494 7586
rect 2546 7534 2548 7586
rect 2492 7522 2548 7534
rect 2604 7364 2660 7982
rect 2940 7698 2996 8204
rect 3164 8194 3220 8204
rect 3388 8258 3444 8270
rect 3388 8206 3390 8258
rect 3442 8206 3444 8258
rect 3388 8148 3444 8206
rect 3612 8260 3668 8988
rect 3724 8978 3780 8988
rect 3948 9044 4004 9054
rect 3612 8166 3668 8204
rect 3724 8818 3780 8830
rect 3724 8766 3726 8818
rect 3778 8766 3780 8818
rect 3388 8082 3444 8092
rect 2940 7646 2942 7698
rect 2994 7646 2996 7698
rect 2940 7634 2996 7646
rect 3276 7812 3332 7822
rect 2828 7476 2884 7486
rect 2604 7298 2660 7308
rect 2716 7474 2996 7476
rect 2716 7422 2830 7474
rect 2882 7422 2996 7474
rect 2716 7420 2996 7422
rect 2716 7140 2772 7420
rect 2828 7410 2884 7420
rect 2380 7084 2772 7140
rect 2828 5906 2884 5918
rect 2828 5854 2830 5906
rect 2882 5854 2884 5906
rect 2716 5236 2772 5246
rect 2156 5124 2212 5134
rect 2716 5124 2772 5180
rect 2156 5030 2212 5068
rect 2380 5122 2772 5124
rect 2380 5070 2718 5122
rect 2770 5070 2772 5122
rect 2380 5068 2772 5070
rect 2380 5010 2436 5068
rect 2716 5058 2772 5068
rect 2828 5124 2884 5854
rect 2940 5684 2996 7420
rect 3052 7474 3108 7486
rect 3052 7422 3054 7474
rect 3106 7422 3108 7474
rect 3052 6244 3108 7422
rect 3276 7028 3332 7756
rect 3500 7474 3556 7486
rect 3500 7422 3502 7474
rect 3554 7422 3556 7474
rect 3500 7252 3556 7422
rect 3500 7186 3556 7196
rect 3276 6972 3556 7028
rect 3052 6130 3108 6188
rect 3052 6078 3054 6130
rect 3106 6078 3108 6130
rect 3052 6066 3108 6078
rect 3164 6916 3220 6926
rect 3052 5684 3108 5694
rect 2940 5628 3052 5684
rect 3052 5618 3108 5628
rect 2828 5058 2884 5068
rect 3052 5012 3108 5022
rect 3164 5012 3220 6860
rect 3500 6018 3556 6972
rect 3500 5966 3502 6018
rect 3554 5966 3556 6018
rect 3500 5954 3556 5966
rect 3388 5682 3444 5694
rect 3388 5630 3390 5682
rect 3442 5630 3444 5682
rect 3388 5234 3444 5630
rect 3388 5182 3390 5234
rect 3442 5182 3444 5234
rect 3388 5124 3444 5182
rect 3388 5058 3444 5068
rect 3612 5122 3668 5134
rect 3612 5070 3614 5122
rect 3666 5070 3668 5122
rect 2380 4958 2382 5010
rect 2434 4958 2436 5010
rect 2380 4946 2436 4958
rect 2940 5010 3220 5012
rect 2940 4958 3054 5010
rect 3106 4958 3220 5010
rect 2940 4956 3220 4958
rect 2940 4900 2996 4956
rect 3052 4946 3108 4956
rect 2492 4844 2996 4900
rect 2492 4450 2548 4844
rect 3612 4788 3668 5070
rect 3724 4900 3780 8766
rect 3836 8708 3892 8718
rect 3836 8370 3892 8652
rect 3836 8318 3838 8370
rect 3890 8318 3892 8370
rect 3836 8306 3892 8318
rect 3836 8148 3892 8158
rect 3948 8148 4004 8988
rect 4060 8372 4116 9212
rect 4060 8306 4116 8316
rect 3836 8146 4004 8148
rect 3836 8094 3838 8146
rect 3890 8094 4004 8146
rect 3836 8092 4004 8094
rect 3836 8082 3892 8092
rect 4060 8034 4116 8046
rect 4060 7982 4062 8034
rect 4114 7982 4116 8034
rect 3948 7924 4004 7934
rect 3836 7250 3892 7262
rect 3836 7198 3838 7250
rect 3890 7198 3892 7250
rect 3836 6692 3892 7198
rect 3948 7250 4004 7868
rect 3948 7198 3950 7250
rect 4002 7198 4004 7250
rect 3948 7028 4004 7198
rect 3948 6962 4004 6972
rect 3836 6626 3892 6636
rect 4060 6692 4116 7982
rect 4284 7924 4340 10220
rect 4172 7364 4228 7374
rect 4172 7270 4228 7308
rect 4060 6626 4116 6636
rect 4284 6468 4340 7868
rect 4396 8148 4452 10332
rect 4396 7474 4452 8092
rect 4620 9716 4676 9726
rect 4620 9268 4676 9660
rect 4844 9492 4900 11732
rect 4956 11732 5012 11742
rect 4956 10834 5012 11676
rect 4956 10782 4958 10834
rect 5010 10782 5012 10834
rect 4956 10770 5012 10782
rect 5068 10612 5124 10650
rect 5068 10546 5124 10556
rect 5068 10388 5124 10398
rect 5068 9492 5124 10332
rect 5180 10052 5236 13468
rect 5370 13356 5634 13366
rect 5426 13300 5474 13356
rect 5530 13300 5578 13356
rect 5370 13290 5634 13300
rect 5628 12964 5684 12974
rect 5740 12964 5796 13580
rect 5852 13570 5908 13580
rect 5684 12908 5796 12964
rect 5852 12962 5908 12974
rect 5852 12910 5854 12962
rect 5906 12910 5908 12962
rect 5628 12870 5684 12908
rect 5292 12740 5348 12750
rect 5292 12402 5348 12684
rect 5292 12350 5294 12402
rect 5346 12350 5348 12402
rect 5292 12338 5348 12350
rect 5628 12404 5684 12414
rect 5628 12310 5684 12348
rect 5852 12180 5908 12910
rect 5852 11954 5908 12124
rect 5852 11902 5854 11954
rect 5906 11902 5908 11954
rect 5852 11890 5908 11902
rect 5370 11788 5634 11798
rect 5426 11732 5474 11788
rect 5530 11732 5578 11788
rect 5370 11722 5634 11732
rect 5516 11396 5572 11406
rect 5516 10388 5572 11340
rect 5852 11284 5908 11294
rect 5852 11190 5908 11228
rect 5516 10322 5572 10332
rect 5370 10220 5634 10230
rect 5426 10164 5474 10220
rect 5530 10164 5578 10220
rect 5370 10154 5634 10164
rect 5180 9996 5460 10052
rect 4844 9426 4900 9436
rect 4956 9436 5124 9492
rect 4620 8146 4676 9212
rect 4844 9268 4900 9278
rect 4844 9042 4900 9212
rect 4844 8990 4846 9042
rect 4898 8990 4900 9042
rect 4844 8978 4900 8990
rect 4956 8428 5012 9436
rect 5292 9268 5348 9278
rect 4844 8372 5012 8428
rect 5068 9266 5348 9268
rect 5068 9214 5294 9266
rect 5346 9214 5348 9266
rect 5068 9212 5348 9214
rect 4620 8094 4622 8146
rect 4674 8094 4676 8146
rect 4508 7700 4564 7710
rect 4508 7586 4564 7644
rect 4508 7534 4510 7586
rect 4562 7534 4564 7586
rect 4508 7522 4564 7534
rect 4396 7422 4398 7474
rect 4450 7422 4452 7474
rect 4396 7410 4452 7422
rect 4620 6804 4676 8094
rect 4732 8260 4788 8270
rect 4732 8034 4788 8204
rect 4732 7982 4734 8034
rect 4786 7982 4788 8034
rect 4732 7476 4788 7982
rect 4732 7410 4788 7420
rect 4844 7586 4900 8372
rect 4956 8260 5012 8270
rect 4956 8166 5012 8204
rect 5068 7700 5124 9212
rect 5292 9202 5348 9212
rect 5404 9266 5460 9996
rect 5628 9828 5684 9838
rect 5628 9734 5684 9772
rect 5852 9714 5908 9726
rect 5852 9662 5854 9714
rect 5906 9662 5908 9714
rect 5404 9214 5406 9266
rect 5458 9214 5460 9266
rect 5404 9202 5460 9214
rect 5740 9492 5796 9502
rect 5180 9042 5236 9054
rect 5180 8990 5182 9042
rect 5234 8990 5236 9042
rect 5180 8036 5236 8990
rect 5516 9042 5572 9054
rect 5516 8990 5518 9042
rect 5570 8990 5572 9042
rect 5516 8932 5572 8990
rect 5516 8866 5572 8876
rect 5370 8652 5634 8662
rect 5426 8596 5474 8652
rect 5530 8596 5578 8652
rect 5370 8586 5634 8596
rect 5628 8372 5684 8382
rect 5628 8258 5684 8316
rect 5628 8206 5630 8258
rect 5682 8206 5684 8258
rect 5628 8194 5684 8206
rect 5516 8036 5572 8046
rect 5180 8034 5572 8036
rect 5180 7982 5518 8034
rect 5570 7982 5572 8034
rect 5180 7980 5572 7982
rect 5516 7970 5572 7980
rect 5628 8036 5684 8046
rect 5180 7700 5236 7710
rect 5068 7698 5236 7700
rect 5068 7646 5182 7698
rect 5234 7646 5236 7698
rect 5068 7644 5236 7646
rect 5180 7634 5236 7644
rect 4844 7534 4846 7586
rect 4898 7534 4900 7586
rect 4844 6916 4900 7534
rect 5180 7474 5236 7486
rect 5180 7422 5182 7474
rect 5234 7422 5236 7474
rect 5180 6916 5236 7422
rect 5292 7476 5348 7486
rect 5292 7382 5348 7420
rect 5516 7476 5572 7486
rect 5628 7476 5684 7980
rect 5740 7700 5796 9436
rect 5852 8484 5908 9662
rect 5852 8418 5908 8428
rect 5852 8260 5908 8270
rect 5852 8166 5908 8204
rect 5740 7644 5908 7700
rect 5516 7474 5684 7476
rect 5516 7422 5518 7474
rect 5570 7422 5684 7474
rect 5516 7420 5684 7422
rect 5740 7476 5796 7486
rect 5516 7410 5572 7420
rect 5740 7382 5796 7420
rect 5370 7084 5634 7094
rect 5426 7028 5474 7084
rect 5530 7028 5578 7084
rect 5370 7018 5634 7028
rect 5180 6860 5796 6916
rect 4844 6850 4900 6860
rect 4732 6804 4788 6814
rect 4620 6748 4732 6804
rect 4732 6738 4788 6748
rect 5740 6802 5796 6860
rect 5740 6750 5742 6802
rect 5794 6750 5796 6802
rect 5740 6738 5796 6750
rect 4956 6692 5012 6702
rect 4956 6598 5012 6636
rect 5628 6692 5684 6702
rect 5628 6598 5684 6636
rect 5852 6692 5908 7644
rect 5852 6626 5908 6636
rect 5068 6580 5124 6590
rect 5068 6486 5124 6524
rect 3948 6412 4340 6468
rect 5852 6466 5908 6478
rect 5852 6414 5854 6466
rect 5906 6414 5908 6466
rect 3948 5346 4004 6412
rect 5852 6356 5908 6414
rect 5852 6290 5908 6300
rect 4620 6244 4676 6254
rect 4620 6130 4676 6188
rect 4620 6078 4622 6130
rect 4674 6078 4676 6130
rect 4620 6066 4676 6078
rect 5516 6132 5572 6142
rect 5516 6038 5572 6076
rect 4508 6020 4564 6030
rect 3948 5294 3950 5346
rect 4002 5294 4004 5346
rect 3948 5282 4004 5294
rect 4396 5906 4452 5918
rect 4396 5854 4398 5906
rect 4450 5854 4452 5906
rect 4284 5236 4340 5246
rect 4284 5122 4340 5180
rect 4284 5070 4286 5122
rect 4338 5070 4340 5122
rect 4284 5058 4340 5070
rect 4284 4900 4340 4910
rect 3724 4898 4340 4900
rect 3724 4846 4286 4898
rect 4338 4846 4340 4898
rect 3724 4844 4340 4846
rect 4284 4834 4340 4844
rect 3612 4722 3668 4732
rect 4396 4788 4452 5854
rect 4508 5346 4564 5964
rect 5852 6020 5908 6030
rect 5852 5926 5908 5964
rect 5180 5908 5236 5918
rect 4508 5294 4510 5346
rect 4562 5294 4564 5346
rect 4508 5282 4564 5294
rect 4844 5906 5236 5908
rect 4844 5854 5182 5906
rect 5234 5854 5236 5906
rect 4844 5852 5236 5854
rect 4844 5124 4900 5852
rect 5180 5842 5236 5852
rect 5370 5516 5634 5526
rect 5426 5460 5474 5516
rect 5530 5460 5578 5516
rect 5370 5450 5634 5460
rect 5964 5348 6020 14028
rect 6412 13972 6468 15150
rect 6860 14308 6916 14318
rect 6916 14252 7028 14308
rect 6860 14242 6916 14252
rect 6524 13972 6580 13982
rect 6412 13970 6580 13972
rect 6412 13918 6526 13970
rect 6578 13918 6580 13970
rect 6412 13916 6580 13918
rect 6524 13906 6580 13916
rect 6300 13746 6356 13758
rect 6300 13694 6302 13746
rect 6354 13694 6356 13746
rect 6076 12962 6132 12974
rect 6076 12910 6078 12962
rect 6130 12910 6132 12962
rect 6076 12292 6132 12910
rect 6076 12226 6132 12236
rect 6076 12066 6132 12078
rect 6076 12014 6078 12066
rect 6130 12014 6132 12066
rect 6076 11956 6132 12014
rect 6076 11890 6132 11900
rect 6188 11954 6244 11966
rect 6188 11902 6190 11954
rect 6242 11902 6244 11954
rect 6076 11394 6132 11406
rect 6076 11342 6078 11394
rect 6130 11342 6132 11394
rect 6076 11060 6132 11342
rect 6076 10994 6132 11004
rect 6076 9940 6132 9950
rect 6188 9940 6244 11902
rect 6300 11956 6356 13694
rect 6412 13746 6468 13758
rect 6748 13748 6804 13758
rect 6412 13694 6414 13746
rect 6466 13694 6468 13746
rect 6412 13412 6468 13694
rect 6412 13346 6468 13356
rect 6524 13746 6804 13748
rect 6524 13694 6750 13746
rect 6802 13694 6804 13746
rect 6524 13692 6804 13694
rect 6412 13188 6468 13198
rect 6412 12404 6468 13132
rect 6524 13186 6580 13692
rect 6748 13682 6804 13692
rect 6972 13748 7028 14252
rect 7756 13972 7812 17164
rect 8092 16994 8148 17724
rect 8428 17714 8484 17724
rect 8540 18562 8820 18564
rect 8540 18510 8766 18562
rect 8818 18510 8820 18562
rect 8540 18508 8820 18510
rect 8540 17668 8596 18508
rect 8764 18498 8820 18508
rect 8876 18564 8932 18574
rect 8932 18508 9156 18564
rect 8876 18470 8932 18508
rect 8876 18228 8932 18238
rect 8876 18134 8932 18172
rect 9100 17668 9156 18508
rect 8204 17556 8260 17566
rect 8204 17106 8260 17500
rect 8204 17054 8206 17106
rect 8258 17054 8260 17106
rect 8204 17042 8260 17054
rect 8428 17108 8484 17118
rect 8540 17108 8596 17612
rect 8428 17106 8596 17108
rect 8428 17054 8430 17106
rect 8482 17054 8596 17106
rect 8428 17052 8596 17054
rect 8652 17666 9156 17668
rect 8652 17614 9102 17666
rect 9154 17614 9156 17666
rect 8652 17612 9156 17614
rect 8652 17106 8708 17612
rect 9100 17556 9156 17612
rect 9100 17490 9156 17500
rect 8876 17442 8932 17454
rect 8876 17390 8878 17442
rect 8930 17390 8932 17442
rect 8876 17332 8932 17390
rect 9212 17332 9268 18620
rect 9324 18564 9380 18732
rect 9548 18564 9604 18574
rect 9324 18562 9604 18564
rect 9324 18510 9550 18562
rect 9602 18510 9604 18562
rect 9324 18508 9604 18510
rect 9548 18498 9604 18508
rect 9660 18564 9716 18574
rect 9660 18470 9716 18508
rect 9884 18450 9940 18462
rect 9884 18398 9886 18450
rect 9938 18398 9940 18450
rect 9884 18340 9940 18398
rect 9884 18274 9940 18284
rect 9996 18116 10052 19070
rect 10556 19124 10612 19134
rect 10556 19030 10612 19068
rect 10556 18676 10612 18686
rect 10444 18620 10556 18676
rect 10332 18340 10388 18350
rect 10220 18338 10388 18340
rect 10220 18286 10334 18338
rect 10386 18286 10388 18338
rect 10220 18284 10388 18286
rect 10108 18228 10164 18238
rect 10108 18134 10164 18172
rect 9660 18060 10052 18116
rect 9660 18004 9716 18060
rect 10220 18004 10276 18284
rect 10332 18274 10388 18284
rect 9548 17892 9604 17902
rect 9548 17798 9604 17836
rect 9660 17444 9716 17948
rect 9884 17948 10276 18004
rect 9884 17890 9940 17948
rect 9884 17838 9886 17890
rect 9938 17838 9940 17890
rect 9884 17826 9940 17838
rect 10444 17778 10500 18620
rect 10556 18610 10612 18620
rect 10556 18452 10612 18462
rect 10556 18358 10612 18396
rect 10668 18450 10724 19180
rect 10780 19236 10836 19516
rect 11116 19236 11172 20636
rect 11340 20626 11396 20636
rect 11452 20692 11508 20702
rect 11340 20132 11396 20142
rect 11340 19346 11396 20076
rect 11452 20018 11508 20636
rect 12012 20130 12068 21756
rect 12124 20244 12180 20254
rect 12236 20244 12292 23772
rect 12684 23716 12740 23772
rect 12348 23660 12740 23716
rect 12348 21924 12404 23660
rect 12796 23548 12852 23884
rect 12460 23436 12852 23548
rect 13020 23714 13076 23726
rect 13020 23662 13022 23714
rect 13074 23662 13076 23714
rect 12684 23266 12740 23278
rect 12684 23214 12686 23266
rect 12738 23214 12740 23266
rect 12348 21858 12404 21868
rect 12460 23154 12516 23166
rect 12460 23102 12462 23154
rect 12514 23102 12516 23154
rect 12348 21698 12404 21710
rect 12348 21646 12350 21698
rect 12402 21646 12404 21698
rect 12348 21588 12404 21646
rect 12348 20804 12404 21532
rect 12460 21476 12516 23102
rect 12572 23044 12628 23054
rect 12572 22950 12628 22988
rect 12684 22932 12740 23214
rect 12684 22866 12740 22876
rect 12460 21410 12516 21420
rect 12684 22372 12740 22382
rect 12684 21810 12740 22316
rect 12684 21758 12686 21810
rect 12738 21758 12740 21810
rect 12348 20738 12404 20748
rect 12572 21364 12628 21374
rect 12572 20802 12628 21308
rect 12684 21252 12740 21758
rect 12796 21588 12852 23436
rect 12908 23492 12964 23502
rect 12908 23378 12964 23436
rect 12908 23326 12910 23378
rect 12962 23326 12964 23378
rect 12908 23314 12964 23326
rect 12908 22372 12964 22382
rect 13020 22372 13076 23662
rect 13132 23268 13188 24108
rect 13356 23940 13412 24558
rect 13468 24612 13524 24622
rect 13692 24612 13748 25452
rect 14140 25506 14196 25564
rect 14140 25454 14142 25506
rect 14194 25454 14196 25506
rect 14140 25442 14196 25454
rect 14252 25506 14308 25676
rect 14476 25618 14532 26124
rect 15036 25844 15092 26908
rect 16492 26852 16772 26908
rect 17500 27076 17556 27086
rect 16380 26516 16436 26526
rect 16044 26514 16436 26516
rect 16044 26462 16382 26514
rect 16434 26462 16436 26514
rect 16044 26460 16436 26462
rect 15932 26180 15988 26190
rect 15708 26178 15988 26180
rect 15708 26126 15934 26178
rect 15986 26126 15988 26178
rect 15708 26124 15988 26126
rect 15036 25788 15316 25844
rect 14476 25566 14478 25618
rect 14530 25566 14532 25618
rect 14476 25554 14532 25566
rect 15260 25620 15316 25788
rect 15372 25620 15428 25630
rect 15260 25618 15428 25620
rect 15260 25566 15374 25618
rect 15426 25566 15428 25618
rect 15260 25564 15428 25566
rect 15372 25554 15428 25564
rect 14252 25454 14254 25506
rect 14306 25454 14308 25506
rect 14252 25442 14308 25454
rect 14700 25508 14756 25518
rect 14588 24724 14644 24734
rect 14140 24612 14196 24650
rect 14588 24630 14644 24668
rect 13468 24610 13748 24612
rect 13468 24558 13470 24610
rect 13522 24558 13748 24610
rect 13468 24556 13748 24558
rect 14028 24556 14140 24612
rect 13468 24546 13524 24556
rect 13686 24332 13950 24342
rect 13742 24276 13790 24332
rect 13846 24276 13894 24332
rect 13686 24266 13950 24276
rect 13580 24164 13636 24174
rect 13580 24162 13860 24164
rect 13580 24110 13582 24162
rect 13634 24110 13860 24162
rect 13580 24108 13860 24110
rect 13580 24098 13636 24108
rect 13468 23940 13524 23950
rect 13356 23938 13524 23940
rect 13356 23886 13470 23938
rect 13522 23886 13524 23938
rect 13356 23884 13524 23886
rect 13468 23874 13524 23884
rect 13580 23828 13636 23838
rect 13468 23604 13524 23614
rect 13468 23380 13524 23548
rect 13132 23202 13188 23212
rect 13356 23324 13524 23380
rect 12908 22370 13076 22372
rect 12908 22318 12910 22370
rect 12962 22318 13076 22370
rect 12908 22316 13076 22318
rect 12908 22148 12964 22316
rect 12908 22082 12964 22092
rect 12796 21522 12852 21532
rect 13020 22036 13076 22046
rect 13356 22036 13412 23324
rect 13580 23268 13636 23772
rect 13692 23716 13748 23726
rect 13692 23622 13748 23660
rect 13692 23268 13748 23278
rect 13580 23266 13748 23268
rect 13580 23214 13694 23266
rect 13746 23214 13748 23266
rect 13580 23212 13748 23214
rect 13468 23154 13524 23166
rect 13468 23102 13470 23154
rect 13522 23102 13524 23154
rect 13468 22372 13524 23102
rect 13692 22932 13748 23212
rect 13804 23266 13860 24108
rect 14028 23828 14084 24556
rect 14140 24546 14196 24556
rect 14140 24388 14196 24398
rect 14140 23938 14196 24332
rect 14700 24052 14756 25452
rect 15148 25506 15204 25518
rect 15148 25454 15150 25506
rect 15202 25454 15204 25506
rect 14924 25396 14980 25406
rect 14924 25302 14980 25340
rect 15148 24946 15204 25454
rect 15484 25508 15540 25518
rect 15484 25414 15540 25452
rect 15148 24894 15150 24946
rect 15202 24894 15204 24946
rect 15148 24882 15204 24894
rect 15260 25172 15316 25182
rect 14140 23886 14142 23938
rect 14194 23886 14196 23938
rect 14140 23874 14196 23886
rect 14252 23996 14756 24052
rect 15036 24722 15092 24734
rect 15036 24670 15038 24722
rect 15090 24670 15092 24722
rect 15036 24052 15092 24670
rect 15260 24722 15316 25116
rect 15708 25172 15764 26124
rect 15932 26114 15988 26124
rect 15820 25508 15876 25518
rect 16044 25508 16100 26460
rect 16380 26450 16436 26460
rect 16268 26290 16324 26302
rect 16268 26238 16270 26290
rect 16322 26238 16324 26290
rect 16268 26180 16324 26238
rect 16268 25620 16324 26124
rect 15820 25506 16100 25508
rect 15820 25454 15822 25506
rect 15874 25454 16100 25506
rect 15820 25452 16100 25454
rect 16156 25564 16324 25620
rect 16492 26290 16548 26852
rect 16492 26238 16494 26290
rect 16546 26238 16548 26290
rect 16156 25506 16212 25564
rect 16156 25454 16158 25506
rect 16210 25454 16212 25506
rect 15820 25442 15876 25452
rect 16156 25442 16212 25454
rect 16268 25396 16324 25406
rect 16268 25302 16324 25340
rect 15708 25106 15764 25116
rect 16380 25282 16436 25294
rect 16380 25230 16382 25282
rect 16434 25230 16436 25282
rect 16380 25172 16436 25230
rect 16380 25106 16436 25116
rect 15708 24836 15764 24846
rect 16492 24836 16548 26238
rect 16940 26290 16996 26302
rect 16940 26238 16942 26290
rect 16994 26238 16996 26290
rect 16604 25284 16660 25294
rect 16604 25190 16660 25228
rect 16940 25284 16996 26238
rect 17500 26292 17556 27020
rect 17612 26964 17668 26974
rect 17668 26908 17780 26964
rect 17612 26898 17668 26908
rect 17724 26292 17780 26908
rect 18172 26962 18228 26974
rect 18172 26910 18174 26962
rect 18226 26910 18228 26962
rect 17844 26684 18108 26694
rect 17900 26628 17948 26684
rect 18004 26628 18052 26684
rect 17844 26618 18108 26628
rect 18172 26514 18228 26910
rect 18172 26462 18174 26514
rect 18226 26462 18228 26514
rect 18172 26450 18228 26462
rect 18284 26964 18340 26974
rect 18284 26402 18340 26908
rect 18956 26516 19012 26526
rect 18284 26350 18286 26402
rect 18338 26350 18340 26402
rect 18284 26338 18340 26350
rect 18508 26514 19012 26516
rect 18508 26462 18958 26514
rect 19010 26462 19012 26514
rect 18508 26460 19012 26462
rect 18508 26402 18564 26460
rect 18956 26450 19012 26460
rect 18508 26350 18510 26402
rect 18562 26350 18564 26402
rect 18508 26338 18564 26350
rect 19068 26404 19124 26414
rect 19068 26310 19124 26348
rect 17836 26292 17892 26302
rect 17724 26290 17892 26292
rect 17724 26238 17838 26290
rect 17890 26238 17892 26290
rect 17724 26236 17892 26238
rect 17500 26226 17556 26236
rect 17836 26226 17892 26236
rect 18844 26290 18900 26302
rect 18844 26238 18846 26290
rect 18898 26238 18900 26290
rect 18844 26180 18900 26238
rect 18844 25508 18900 26124
rect 19180 26068 19236 27804
rect 19292 27794 19348 27804
rect 20076 27858 20132 27870
rect 20076 27806 20078 27858
rect 20130 27806 20132 27858
rect 19516 27188 19572 27198
rect 19572 27132 19684 27188
rect 19516 27122 19572 27132
rect 18956 26012 19236 26068
rect 19516 26290 19572 26302
rect 19516 26238 19518 26290
rect 19570 26238 19572 26290
rect 18956 25730 19012 26012
rect 18956 25678 18958 25730
rect 19010 25678 19012 25730
rect 18956 25666 19012 25678
rect 19516 25620 19572 26238
rect 19516 25554 19572 25564
rect 16940 25218 16996 25228
rect 17500 25284 17556 25294
rect 15708 24834 16548 24836
rect 15708 24782 15710 24834
rect 15762 24782 16548 24834
rect 15708 24780 16548 24782
rect 15708 24770 15764 24780
rect 15260 24670 15262 24722
rect 15314 24670 15316 24722
rect 15260 24388 15316 24670
rect 15260 24322 15316 24332
rect 15596 24498 15652 24510
rect 15596 24446 15598 24498
rect 15650 24446 15652 24498
rect 15372 24052 15428 24062
rect 15036 24050 15316 24052
rect 15036 23998 15038 24050
rect 15090 23998 15316 24050
rect 15036 23996 15316 23998
rect 14028 23762 14084 23772
rect 13916 23716 13972 23754
rect 13916 23650 13972 23660
rect 13916 23492 13972 23502
rect 13972 23436 14084 23492
rect 13916 23426 13972 23436
rect 13804 23214 13806 23266
rect 13858 23214 13860 23266
rect 13804 23202 13860 23214
rect 13916 22932 13972 22942
rect 13692 22876 13916 22932
rect 13916 22866 13972 22876
rect 13686 22764 13950 22774
rect 13742 22708 13790 22764
rect 13846 22708 13894 22764
rect 13686 22698 13950 22708
rect 14028 22596 14084 23436
rect 14140 23380 14196 23390
rect 14252 23380 14308 23996
rect 15036 23958 15092 23996
rect 14476 23826 14532 23838
rect 14476 23774 14478 23826
rect 14530 23774 14532 23826
rect 14476 23604 14532 23774
rect 14476 23538 14532 23548
rect 14588 23714 14644 23726
rect 14588 23662 14590 23714
rect 14642 23662 14644 23714
rect 14140 23378 14308 23380
rect 14140 23326 14142 23378
rect 14194 23326 14308 23378
rect 14140 23324 14308 23326
rect 14140 23314 14196 23324
rect 14476 23154 14532 23166
rect 14476 23102 14478 23154
rect 14530 23102 14532 23154
rect 13468 22306 13524 22316
rect 13804 22540 14084 22596
rect 14364 22932 14420 22942
rect 13580 22260 13636 22270
rect 13636 22204 13748 22260
rect 13580 22194 13636 22204
rect 13356 21980 13636 22036
rect 13020 21586 13076 21980
rect 13580 21810 13636 21980
rect 13580 21758 13582 21810
rect 13634 21758 13636 21810
rect 13580 21746 13636 21758
rect 13692 21810 13748 22204
rect 13692 21758 13694 21810
rect 13746 21758 13748 21810
rect 13692 21746 13748 21758
rect 13804 21810 13860 22540
rect 13804 21758 13806 21810
rect 13858 21758 13860 21810
rect 13804 21746 13860 21758
rect 13468 21700 13524 21738
rect 13468 21634 13524 21644
rect 14140 21588 14196 21598
rect 13020 21534 13022 21586
rect 13074 21534 13076 21586
rect 12684 21196 12852 21252
rect 12684 21028 12740 21038
rect 12684 20934 12740 20972
rect 12572 20750 12574 20802
rect 12626 20750 12628 20802
rect 12572 20738 12628 20750
rect 12684 20692 12740 20702
rect 12684 20598 12740 20636
rect 12796 20580 12852 21196
rect 12796 20514 12852 20524
rect 12180 20188 12292 20244
rect 12124 20178 12180 20188
rect 12012 20078 12014 20130
rect 12066 20078 12068 20130
rect 12012 20066 12068 20078
rect 12572 20130 12628 20142
rect 12572 20078 12574 20130
rect 12626 20078 12628 20130
rect 11900 20020 11956 20030
rect 11452 19966 11454 20018
rect 11506 19966 11508 20018
rect 11452 19954 11508 19966
rect 11676 20018 11956 20020
rect 11676 19966 11902 20018
rect 11954 19966 11956 20018
rect 11676 19964 11956 19966
rect 11340 19294 11342 19346
rect 11394 19294 11396 19346
rect 11340 19282 11396 19294
rect 10780 19234 10948 19236
rect 10780 19182 10782 19234
rect 10834 19182 10948 19234
rect 10780 19180 10948 19182
rect 10780 19170 10836 19180
rect 10780 19012 10836 19022
rect 10780 18674 10836 18956
rect 10780 18622 10782 18674
rect 10834 18622 10836 18674
rect 10780 18610 10836 18622
rect 10668 18398 10670 18450
rect 10722 18398 10724 18450
rect 10668 18386 10724 18398
rect 10444 17726 10446 17778
rect 10498 17726 10500 17778
rect 10444 17714 10500 17726
rect 10220 17668 10276 17678
rect 10220 17574 10276 17612
rect 10892 17666 10948 19180
rect 11116 19170 11172 19180
rect 11228 19122 11284 19134
rect 11228 19070 11230 19122
rect 11282 19070 11284 19122
rect 10892 17614 10894 17666
rect 10946 17614 10948 17666
rect 10892 17602 10948 17614
rect 11004 19010 11060 19022
rect 11004 18958 11006 19010
rect 11058 18958 11060 19010
rect 11004 18228 11060 18958
rect 11228 18788 11284 19070
rect 11452 18788 11508 18798
rect 11228 18732 11452 18788
rect 11340 18564 11396 18574
rect 11340 18452 11396 18508
rect 10668 17556 10724 17566
rect 9772 17444 9828 17482
rect 10668 17462 10724 17500
rect 9660 17388 9772 17444
rect 9772 17378 9828 17388
rect 10444 17442 10500 17454
rect 10444 17390 10446 17442
rect 10498 17390 10500 17442
rect 8876 17276 9268 17332
rect 9884 17332 9940 17342
rect 9528 17276 9792 17286
rect 9584 17220 9632 17276
rect 9688 17220 9736 17276
rect 9528 17210 9792 17220
rect 8652 17054 8654 17106
rect 8706 17054 8708 17106
rect 8428 17042 8484 17052
rect 8652 17042 8708 17054
rect 9884 17106 9940 17276
rect 9884 17054 9886 17106
rect 9938 17054 9940 17106
rect 9884 17042 9940 17054
rect 10444 17332 10500 17390
rect 11004 17332 11060 18172
rect 11228 18450 11396 18452
rect 11228 18398 11342 18450
rect 11394 18398 11396 18450
rect 11228 18396 11396 18398
rect 11228 17666 11284 18396
rect 11340 18386 11396 18396
rect 11452 18562 11508 18732
rect 11452 18510 11454 18562
rect 11506 18510 11508 18562
rect 11452 18452 11508 18510
rect 11452 18386 11508 18396
rect 11676 18450 11732 19964
rect 11900 19954 11956 19964
rect 12124 20020 12180 20030
rect 12572 20020 12628 20078
rect 13020 20132 13076 21534
rect 14028 21586 14196 21588
rect 14028 21534 14142 21586
rect 14194 21534 14196 21586
rect 14028 21532 14196 21534
rect 13686 21196 13950 21206
rect 13742 21140 13790 21196
rect 13846 21140 13894 21196
rect 13686 21130 13950 21140
rect 14028 20916 14084 21532
rect 14140 21522 14196 21532
rect 14364 21364 14420 22876
rect 14476 21812 14532 23102
rect 14476 21586 14532 21756
rect 14476 21534 14478 21586
rect 14530 21534 14532 21586
rect 14476 21522 14532 21534
rect 14588 23044 14644 23662
rect 14364 21308 14532 21364
rect 13804 20860 14084 20916
rect 13804 20802 13860 20860
rect 13804 20750 13806 20802
rect 13858 20750 13860 20802
rect 13804 20738 13860 20750
rect 14140 20802 14196 20814
rect 14140 20750 14142 20802
rect 14194 20750 14196 20802
rect 13468 20692 13524 20702
rect 13020 20066 13076 20076
rect 13356 20690 13524 20692
rect 13356 20638 13470 20690
rect 13522 20638 13524 20690
rect 13356 20636 13524 20638
rect 12124 20018 12516 20020
rect 12124 19966 12126 20018
rect 12178 19966 12516 20018
rect 12124 19964 12516 19966
rect 12124 19954 12180 19964
rect 12460 19460 12516 19964
rect 12572 19954 12628 19964
rect 12684 20020 12740 20030
rect 12684 20018 12964 20020
rect 12684 19966 12686 20018
rect 12738 19966 12964 20018
rect 12684 19964 12964 19966
rect 12684 19954 12740 19964
rect 12572 19794 12628 19806
rect 12572 19742 12574 19794
rect 12626 19742 12628 19794
rect 12572 19684 12628 19742
rect 12572 19618 12628 19628
rect 12684 19460 12740 19470
rect 12460 19458 12740 19460
rect 12460 19406 12686 19458
rect 12738 19406 12740 19458
rect 12460 19404 12740 19406
rect 12684 19394 12740 19404
rect 12236 19348 12292 19358
rect 12236 19254 12292 19292
rect 12796 19122 12852 19134
rect 12796 19070 12798 19122
rect 12850 19070 12852 19122
rect 11900 19010 11956 19022
rect 11900 18958 11902 19010
rect 11954 18958 11956 19010
rect 11900 18676 11956 18958
rect 11900 18610 11956 18620
rect 12124 19010 12180 19022
rect 12124 18958 12126 19010
rect 12178 18958 12180 19010
rect 12124 18564 12180 18958
rect 12348 19012 12404 19022
rect 12348 19010 12628 19012
rect 12348 18958 12350 19010
rect 12402 18958 12628 19010
rect 12348 18956 12628 18958
rect 12348 18946 12404 18956
rect 12572 18676 12628 18956
rect 12684 18676 12740 18686
rect 12572 18674 12740 18676
rect 12572 18622 12686 18674
rect 12738 18622 12740 18674
rect 12572 18620 12740 18622
rect 12684 18610 12740 18620
rect 12124 18498 12180 18508
rect 11676 18398 11678 18450
rect 11730 18398 11732 18450
rect 11676 18386 11732 18398
rect 11788 18450 11844 18462
rect 11788 18398 11790 18450
rect 11842 18398 11844 18450
rect 11788 18228 11844 18398
rect 11900 18452 11956 18462
rect 11956 18396 12068 18452
rect 11900 18386 11956 18396
rect 12012 18340 12068 18396
rect 12124 18340 12180 18350
rect 12012 18338 12180 18340
rect 12012 18286 12126 18338
rect 12178 18286 12180 18338
rect 12012 18284 12180 18286
rect 12124 18274 12180 18284
rect 12348 18340 12404 18350
rect 12348 18246 12404 18284
rect 11788 18162 11844 18172
rect 12796 18116 12852 19070
rect 12908 18228 12964 19964
rect 13356 19348 13412 20636
rect 13468 20626 13524 20636
rect 13580 20580 13636 20590
rect 13580 20486 13636 20524
rect 14140 20580 14196 20750
rect 14364 20804 14420 20814
rect 14364 20690 14420 20748
rect 14364 20638 14366 20690
rect 14418 20638 14420 20690
rect 14364 20626 14420 20638
rect 14140 20514 14196 20524
rect 13580 20132 13636 20142
rect 13580 19796 13636 20076
rect 14252 20132 14308 20142
rect 14252 20038 14308 20076
rect 13356 19282 13412 19292
rect 13468 19740 13636 19796
rect 14028 20018 14084 20030
rect 14028 19966 14030 20018
rect 14082 19966 14084 20018
rect 14028 19908 14084 19966
rect 14476 20020 14532 21308
rect 14588 21028 14644 22988
rect 14700 23716 14756 23726
rect 14700 22820 14756 23660
rect 14812 23716 14868 23726
rect 14812 23714 15092 23716
rect 14812 23662 14814 23714
rect 14866 23662 15092 23714
rect 14812 23660 15092 23662
rect 14812 23650 14868 23660
rect 15036 23380 15092 23660
rect 15036 23324 15204 23380
rect 14812 23268 14868 23278
rect 14812 23174 14868 23212
rect 15036 23154 15092 23166
rect 15036 23102 15038 23154
rect 15090 23102 15092 23154
rect 14924 23044 14980 23054
rect 15036 23044 15092 23102
rect 14980 22988 15092 23044
rect 14924 22978 14980 22988
rect 14700 22764 14980 22820
rect 14700 21924 14756 21934
rect 14700 21810 14756 21868
rect 14700 21758 14702 21810
rect 14754 21758 14756 21810
rect 14700 21746 14756 21758
rect 14924 21810 14980 22764
rect 15036 22370 15092 22382
rect 15036 22318 15038 22370
rect 15090 22318 15092 22370
rect 15036 22148 15092 22318
rect 15036 22082 15092 22092
rect 14924 21758 14926 21810
rect 14978 21758 14980 21810
rect 14924 21746 14980 21758
rect 14812 21700 14868 21710
rect 14812 21606 14868 21644
rect 15148 21586 15204 23324
rect 15260 21924 15316 23996
rect 15372 23492 15428 23996
rect 15596 23940 15652 24446
rect 15596 23874 15652 23884
rect 15372 23154 15428 23436
rect 15932 23828 15988 23838
rect 15932 23378 15988 23772
rect 17164 23828 17220 23838
rect 17164 23734 17220 23772
rect 15932 23326 15934 23378
rect 15986 23326 15988 23378
rect 15932 23314 15988 23326
rect 17388 23380 17444 23390
rect 17388 23286 17444 23324
rect 15820 23268 15876 23278
rect 15820 23174 15876 23212
rect 15372 23102 15374 23154
rect 15426 23102 15428 23154
rect 15372 23090 15428 23102
rect 16044 23154 16100 23166
rect 16044 23102 16046 23154
rect 16098 23102 16100 23154
rect 16044 22932 16100 23102
rect 16044 22866 16100 22876
rect 15260 21858 15316 21868
rect 15708 21812 15764 21822
rect 16828 21812 16884 21822
rect 15764 21756 15876 21812
rect 15708 21718 15764 21756
rect 15148 21534 15150 21586
rect 15202 21534 15204 21586
rect 15148 21522 15204 21534
rect 15484 21586 15540 21598
rect 15484 21534 15486 21586
rect 15538 21534 15540 21586
rect 15372 21476 15428 21486
rect 15372 21382 15428 21420
rect 15484 21028 15540 21534
rect 14588 20972 14868 21028
rect 14812 20132 14868 20972
rect 15484 20962 15540 20972
rect 15596 21476 15652 21486
rect 14924 20132 14980 20142
rect 14812 20130 14980 20132
rect 14812 20078 14926 20130
rect 14978 20078 14980 20130
rect 14812 20076 14980 20078
rect 14700 20020 14756 20030
rect 14476 20018 14756 20020
rect 14476 19966 14702 20018
rect 14754 19966 14756 20018
rect 14476 19964 14756 19966
rect 12908 18162 12964 18172
rect 12796 18050 12852 18060
rect 11228 17614 11230 17666
rect 11282 17614 11284 17666
rect 11116 17444 11172 17454
rect 11116 17350 11172 17388
rect 10444 17276 11060 17332
rect 11228 17332 11284 17614
rect 10444 17108 10500 17276
rect 11228 17266 11284 17276
rect 10444 17042 10500 17052
rect 8092 16942 8094 16994
rect 8146 16942 8148 16994
rect 8092 16930 8148 16942
rect 8876 16884 8932 16894
rect 9548 16884 9604 16894
rect 8876 16882 9604 16884
rect 8876 16830 8878 16882
rect 8930 16830 9550 16882
rect 9602 16830 9604 16882
rect 8876 16828 9604 16830
rect 8540 15204 8596 15214
rect 8876 15204 8932 16828
rect 9548 16818 9604 16828
rect 10780 16884 10836 16894
rect 10780 16210 10836 16828
rect 12124 16884 12180 16894
rect 12124 16790 12180 16828
rect 12236 16882 12292 16894
rect 12236 16830 12238 16882
rect 12290 16830 12292 16882
rect 12236 16772 12292 16830
rect 12908 16884 12964 16894
rect 12236 16706 12292 16716
rect 12796 16770 12852 16782
rect 12796 16718 12798 16770
rect 12850 16718 12852 16770
rect 12684 16660 12740 16670
rect 10780 16158 10782 16210
rect 10834 16158 10836 16210
rect 10780 16146 10836 16158
rect 12348 16658 12740 16660
rect 12348 16606 12686 16658
rect 12738 16606 12740 16658
rect 12348 16604 12740 16606
rect 10108 16098 10164 16110
rect 10108 16046 10110 16098
rect 10162 16046 10164 16098
rect 9660 15876 9716 15886
rect 10108 15876 10164 16046
rect 12348 15876 12404 16604
rect 12684 16594 12740 16604
rect 12796 16212 12852 16718
rect 12796 16146 12852 16156
rect 12908 16210 12964 16828
rect 12908 16158 12910 16210
rect 12962 16158 12964 16210
rect 12908 16146 12964 16158
rect 13468 16884 13524 19740
rect 13686 19628 13950 19638
rect 13742 19572 13790 19628
rect 13846 19572 13894 19628
rect 13686 19562 13950 19572
rect 13916 19460 13972 19470
rect 14028 19460 14084 19852
rect 14700 19796 14756 19964
rect 14700 19730 14756 19740
rect 13972 19404 14084 19460
rect 13916 19394 13972 19404
rect 14028 18452 14084 18462
rect 14028 18358 14084 18396
rect 14700 18340 14756 18350
rect 14700 18246 14756 18284
rect 13686 18060 13950 18070
rect 13742 18004 13790 18060
rect 13846 18004 13894 18060
rect 13686 17994 13950 18004
rect 14364 17556 14420 17566
rect 14364 17106 14420 17500
rect 14364 17054 14366 17106
rect 14418 17054 14420 17106
rect 14140 16994 14196 17006
rect 14140 16942 14142 16994
rect 14194 16942 14196 16994
rect 13580 16884 13636 16894
rect 13468 16882 13636 16884
rect 13468 16830 13582 16882
rect 13634 16830 13636 16882
rect 13468 16828 13636 16830
rect 13468 15988 13524 16828
rect 13580 16818 13636 16828
rect 13916 16882 13972 16894
rect 13916 16830 13918 16882
rect 13970 16830 13972 16882
rect 13916 16660 13972 16830
rect 14140 16884 14196 16942
rect 14140 16818 14196 16828
rect 14028 16772 14084 16782
rect 14028 16678 14084 16716
rect 13916 16594 13972 16604
rect 13686 16492 13950 16502
rect 13742 16436 13790 16492
rect 13846 16436 13894 16492
rect 13686 16426 13950 16436
rect 13692 16212 13748 16222
rect 13692 16118 13748 16156
rect 13804 16098 13860 16110
rect 13804 16046 13806 16098
rect 13858 16046 13860 16098
rect 13804 15988 13860 16046
rect 13468 15932 13860 15988
rect 14140 15988 14196 15998
rect 14364 15988 14420 17054
rect 14812 16324 14868 20076
rect 14924 20066 14980 20076
rect 15260 20130 15316 20142
rect 15260 20078 15262 20130
rect 15314 20078 15316 20130
rect 15260 19908 15316 20078
rect 15260 19842 15316 19852
rect 15484 20020 15540 20030
rect 15596 20020 15652 21420
rect 15820 20916 15876 21756
rect 16492 21698 16548 21710
rect 16492 21646 16494 21698
rect 16546 21646 16548 21698
rect 16492 21364 16548 21646
rect 16492 21298 16548 21308
rect 15820 20822 15876 20860
rect 16716 20916 16772 20926
rect 16044 20804 16100 20814
rect 16044 20710 16100 20748
rect 16716 20690 16772 20860
rect 16828 20804 16884 21756
rect 17500 21252 17556 25228
rect 17844 25116 18108 25126
rect 17900 25060 17948 25116
rect 18004 25060 18052 25116
rect 17844 25050 18108 25060
rect 18844 24946 18900 25452
rect 19292 25506 19348 25518
rect 19292 25454 19294 25506
rect 19346 25454 19348 25506
rect 19292 25284 19348 25454
rect 19516 25396 19572 25406
rect 19516 25302 19572 25340
rect 19292 25218 19348 25228
rect 18844 24894 18846 24946
rect 18898 24894 18900 24946
rect 18844 24882 18900 24894
rect 18172 24836 18228 24846
rect 18228 24780 18340 24836
rect 18172 24742 18228 24780
rect 17948 23940 18004 23950
rect 17948 23938 18228 23940
rect 17948 23886 17950 23938
rect 18002 23886 18228 23938
rect 17948 23884 18228 23886
rect 17948 23874 18004 23884
rect 17844 23548 18108 23558
rect 17900 23492 17948 23548
rect 18004 23492 18052 23548
rect 17844 23482 18108 23492
rect 17836 23380 17892 23390
rect 17724 23044 17780 23054
rect 17724 22950 17780 22988
rect 17836 22148 17892 23324
rect 18172 23156 18228 23884
rect 18284 23716 18340 24780
rect 18508 24724 18564 24734
rect 18508 24722 18676 24724
rect 18508 24670 18510 24722
rect 18562 24670 18676 24722
rect 18508 24668 18676 24670
rect 18508 24658 18564 24668
rect 18620 24612 18676 24668
rect 19068 24722 19124 24734
rect 19068 24670 19070 24722
rect 19122 24670 19124 24722
rect 19068 24612 19124 24670
rect 18620 24556 19124 24612
rect 18284 23650 18340 23660
rect 18508 23714 18564 23726
rect 18508 23662 18510 23714
rect 18562 23662 18564 23714
rect 18508 23380 18564 23662
rect 18172 23090 18228 23100
rect 18284 23324 18564 23380
rect 17724 22092 17892 22148
rect 17948 23042 18004 23054
rect 17948 22990 17950 23042
rect 18002 22990 18004 23042
rect 17948 22148 18004 22990
rect 18284 22148 18340 23324
rect 18620 23268 18676 24556
rect 19180 23940 19236 23950
rect 19180 23938 19460 23940
rect 19180 23886 19182 23938
rect 19234 23886 19460 23938
rect 19180 23884 19460 23886
rect 19180 23874 19236 23884
rect 18844 23826 18900 23838
rect 18844 23774 18846 23826
rect 18898 23774 18900 23826
rect 18844 23378 18900 23774
rect 18844 23326 18846 23378
rect 18898 23326 18900 23378
rect 18844 23314 18900 23326
rect 18956 23714 19012 23726
rect 18956 23662 18958 23714
rect 19010 23662 19012 23714
rect 18956 23268 19012 23662
rect 19292 23716 19348 23726
rect 19068 23380 19124 23390
rect 19068 23286 19124 23324
rect 18620 23266 18788 23268
rect 18620 23214 18622 23266
rect 18674 23214 18788 23266
rect 18620 23212 18788 23214
rect 18620 23202 18676 23212
rect 17948 22092 18340 22148
rect 17724 21812 17780 22092
rect 17844 21980 18108 21990
rect 17900 21924 17948 21980
rect 18004 21924 18052 21980
rect 17844 21914 18108 21924
rect 17948 21812 18004 21822
rect 17724 21810 18004 21812
rect 17724 21758 17950 21810
rect 18002 21758 18004 21810
rect 17724 21756 18004 21758
rect 17948 21746 18004 21756
rect 18172 21586 18228 21598
rect 18172 21534 18174 21586
rect 18226 21534 18228 21586
rect 17612 21476 17668 21486
rect 17612 21382 17668 21420
rect 18172 21476 18228 21534
rect 18172 21410 18228 21420
rect 17500 21196 17892 21252
rect 16940 20804 16996 20814
rect 16828 20802 17444 20804
rect 16828 20750 16942 20802
rect 16994 20750 17444 20802
rect 16828 20748 17444 20750
rect 16940 20738 16996 20748
rect 16716 20638 16718 20690
rect 16770 20638 16772 20690
rect 16716 20626 16772 20638
rect 17388 20692 17444 20748
rect 17724 20692 17780 20702
rect 17388 20690 17668 20692
rect 17388 20638 17390 20690
rect 17442 20638 17668 20690
rect 17388 20636 17668 20638
rect 17388 20626 17444 20636
rect 15484 20018 15652 20020
rect 15484 19966 15486 20018
rect 15538 19966 15652 20018
rect 15484 19964 15652 19966
rect 16380 20578 16436 20590
rect 16380 20526 16382 20578
rect 16434 20526 16436 20578
rect 16380 20020 16436 20526
rect 17500 20468 17556 20478
rect 16828 20132 16884 20142
rect 16940 20132 16996 20142
rect 16828 20130 16940 20132
rect 16828 20078 16830 20130
rect 16882 20078 16940 20130
rect 16828 20076 16940 20078
rect 16828 20066 16884 20076
rect 14812 16258 14868 16268
rect 14924 19012 14980 19022
rect 15484 19012 15540 19964
rect 16380 19954 16436 19964
rect 16604 20018 16660 20030
rect 16604 19966 16606 20018
rect 16658 19966 16660 20018
rect 16044 19908 16100 19918
rect 14924 19010 15540 19012
rect 14924 18958 14926 19010
rect 14978 18958 15540 19010
rect 14924 18956 15540 18958
rect 15932 19906 16100 19908
rect 15932 19854 16046 19906
rect 16098 19854 16100 19906
rect 15932 19852 16100 19854
rect 15932 19796 15988 19852
rect 16044 19842 16100 19852
rect 16604 19908 16660 19966
rect 16604 19842 16660 19852
rect 14812 16100 14868 16110
rect 14700 16098 14868 16100
rect 14700 16046 14814 16098
rect 14866 16046 14868 16098
rect 14700 16044 14868 16046
rect 14476 15988 14532 15998
rect 14364 15986 14532 15988
rect 14364 15934 14478 15986
rect 14530 15934 14532 15986
rect 14364 15932 14532 15934
rect 14140 15894 14196 15932
rect 14476 15922 14532 15932
rect 14700 15988 14756 16044
rect 14812 16034 14868 16044
rect 14700 15922 14756 15932
rect 9660 15874 10164 15876
rect 9660 15822 9662 15874
rect 9714 15822 10164 15874
rect 9660 15820 10164 15822
rect 9660 15810 9716 15820
rect 9528 15708 9792 15718
rect 9584 15652 9632 15708
rect 9688 15652 9736 15708
rect 9528 15642 9792 15652
rect 8540 15202 8932 15204
rect 8540 15150 8542 15202
rect 8594 15150 8932 15202
rect 8540 15148 8932 15150
rect 8988 15314 9044 15326
rect 8988 15262 8990 15314
rect 9042 15262 9044 15314
rect 8540 15138 8596 15148
rect 8988 15092 9044 15262
rect 10108 15148 10164 15820
rect 11900 15820 12404 15876
rect 14252 15874 14308 15886
rect 14252 15822 14254 15874
rect 14306 15822 14308 15874
rect 11900 15426 11956 15820
rect 11900 15374 11902 15426
rect 11954 15374 11956 15426
rect 11900 15362 11956 15374
rect 11228 15316 11284 15326
rect 11228 15222 11284 15260
rect 13468 15316 13524 15326
rect 7756 13906 7812 13916
rect 8428 14420 8484 14430
rect 8988 14420 9044 15036
rect 9996 15092 10164 15148
rect 9996 15026 10052 15036
rect 8428 14418 9044 14420
rect 8428 14366 8430 14418
rect 8482 14366 9044 14418
rect 8428 14364 9044 14366
rect 12684 14530 12740 14542
rect 12684 14478 12686 14530
rect 12738 14478 12740 14530
rect 8428 14084 8484 14364
rect 12684 14308 12740 14478
rect 9528 14140 9792 14150
rect 9584 14084 9632 14140
rect 9688 14084 9736 14140
rect 9528 14074 9792 14084
rect 6524 13134 6526 13186
rect 6578 13134 6580 13186
rect 6524 13122 6580 13134
rect 6636 13524 6692 13534
rect 6636 12404 6692 13468
rect 6748 12964 6804 12974
rect 6748 12870 6804 12908
rect 6860 12740 6916 12750
rect 6860 12646 6916 12684
rect 6412 12310 6468 12348
rect 6524 12348 6636 12404
rect 6300 11900 6468 11956
rect 6412 11506 6468 11900
rect 6412 11454 6414 11506
rect 6466 11454 6468 11506
rect 6412 11442 6468 11454
rect 6076 9938 6244 9940
rect 6076 9886 6078 9938
rect 6130 9886 6244 9938
rect 6076 9884 6244 9886
rect 6300 11396 6356 11406
rect 6300 10612 6356 11340
rect 6524 11396 6580 12348
rect 6636 12338 6692 12348
rect 6748 12292 6804 12302
rect 6748 12198 6804 12236
rect 6860 11620 6916 11630
rect 6972 11620 7028 13692
rect 7756 13634 7812 13646
rect 7756 13582 7758 13634
rect 7810 13582 7812 13634
rect 7084 13188 7140 13198
rect 7084 12962 7140 13132
rect 7756 13188 7812 13582
rect 7756 13122 7812 13132
rect 7868 13522 7924 13534
rect 7868 13470 7870 13522
rect 7922 13470 7924 13522
rect 7420 13076 7476 13086
rect 7420 12982 7476 13020
rect 7084 12910 7086 12962
rect 7138 12910 7140 12962
rect 7084 12898 7140 12910
rect 7532 12850 7588 12862
rect 7532 12798 7534 12850
rect 7586 12798 7588 12850
rect 7196 12740 7252 12750
rect 7084 12404 7140 12414
rect 7084 12310 7140 12348
rect 6860 11618 6972 11620
rect 6860 11566 6862 11618
rect 6914 11566 6972 11618
rect 6860 11564 6972 11566
rect 6860 11554 6916 11564
rect 6972 11526 7028 11564
rect 7084 11396 7140 11406
rect 6524 11394 6692 11396
rect 6524 11342 6526 11394
rect 6578 11342 6692 11394
rect 6524 11340 6692 11342
rect 6524 11330 6580 11340
rect 6636 10948 6692 11340
rect 7084 11302 7140 11340
rect 7196 11172 7252 12684
rect 7532 12404 7588 12798
rect 7532 12338 7588 12348
rect 7308 12292 7364 12302
rect 7308 11508 7364 12236
rect 7420 12178 7476 12190
rect 7420 12126 7422 12178
rect 7474 12126 7476 12178
rect 7420 11732 7476 12126
rect 7420 11666 7476 11676
rect 7868 11732 7924 13470
rect 7980 12964 8036 12974
rect 8428 12964 8484 14028
rect 10668 14028 11060 14084
rect 10668 13970 10724 14028
rect 10668 13918 10670 13970
rect 10722 13918 10724 13970
rect 10668 13906 10724 13918
rect 11004 13972 11060 14028
rect 11116 13972 11172 13982
rect 11004 13970 11172 13972
rect 11004 13918 11118 13970
rect 11170 13918 11172 13970
rect 11004 13916 11172 13918
rect 11116 13906 11172 13916
rect 11900 13972 11956 13982
rect 10556 13860 10612 13870
rect 10108 13746 10164 13758
rect 10108 13694 10110 13746
rect 10162 13694 10164 13746
rect 10108 13524 10164 13694
rect 10332 13748 10388 13758
rect 10332 13654 10388 13692
rect 10108 13458 10164 13468
rect 8652 13412 8708 13422
rect 7980 12962 8428 12964
rect 7980 12910 7982 12962
rect 8034 12910 8428 12962
rect 7980 12908 8428 12910
rect 7980 12898 8036 12908
rect 8428 12870 8484 12908
rect 8540 13076 8596 13086
rect 7980 12290 8036 12302
rect 8540 12292 8596 13020
rect 8652 12852 8708 13356
rect 10556 13300 10612 13804
rect 10892 13860 10948 13870
rect 11788 13860 11844 13870
rect 10892 13858 11060 13860
rect 10892 13806 10894 13858
rect 10946 13806 11060 13858
rect 10892 13804 11060 13806
rect 10892 13794 10948 13804
rect 10892 13634 10948 13646
rect 10892 13582 10894 13634
rect 10946 13582 10948 13634
rect 10556 13244 10836 13300
rect 10780 13074 10836 13244
rect 10780 13022 10782 13074
rect 10834 13022 10836 13074
rect 10780 13010 10836 13022
rect 8652 12850 8820 12852
rect 8652 12798 8654 12850
rect 8706 12798 8820 12850
rect 8652 12796 8820 12798
rect 8652 12786 8708 12796
rect 8652 12292 8708 12302
rect 7980 12238 7982 12290
rect 8034 12238 8036 12290
rect 7980 12068 8036 12238
rect 8428 12290 8708 12292
rect 8428 12238 8654 12290
rect 8706 12238 8708 12290
rect 8428 12236 8708 12238
rect 8764 12292 8820 12796
rect 9528 12572 9792 12582
rect 9584 12516 9632 12572
rect 9688 12516 9736 12572
rect 9528 12506 9792 12516
rect 9884 12404 9940 12414
rect 9884 12310 9940 12348
rect 10892 12404 10948 13582
rect 11004 12740 11060 13804
rect 11788 13766 11844 13804
rect 11340 13748 11396 13758
rect 11228 13746 11396 13748
rect 11228 13694 11342 13746
rect 11394 13694 11396 13746
rect 11228 13692 11396 13694
rect 11228 13074 11284 13692
rect 11340 13682 11396 13692
rect 11228 13022 11230 13074
rect 11282 13022 11284 13074
rect 11228 13010 11284 13022
rect 11676 13522 11732 13534
rect 11676 13470 11678 13522
rect 11730 13470 11732 13522
rect 11676 12962 11732 13470
rect 11900 13076 11956 13916
rect 11900 13010 11956 13020
rect 12124 13748 12180 13758
rect 12124 13074 12180 13692
rect 12124 13022 12126 13074
rect 12178 13022 12180 13074
rect 12124 13010 12180 13022
rect 12236 13524 12292 13534
rect 11676 12910 11678 12962
rect 11730 12910 11732 12962
rect 11676 12898 11732 12910
rect 11004 12674 11060 12684
rect 11116 12740 11172 12750
rect 11340 12740 11396 12750
rect 11116 12738 11284 12740
rect 11116 12686 11118 12738
rect 11170 12686 11284 12738
rect 11116 12684 11284 12686
rect 11116 12674 11172 12684
rect 10892 12338 10948 12348
rect 8988 12292 9044 12302
rect 8764 12236 8988 12292
rect 8316 12178 8372 12190
rect 8316 12126 8318 12178
rect 8370 12126 8372 12178
rect 8036 12012 8148 12068
rect 7980 12002 8036 12012
rect 7868 11666 7924 11676
rect 7308 11452 7588 11508
rect 7532 11394 7588 11452
rect 7532 11342 7534 11394
rect 7586 11342 7588 11394
rect 7420 11284 7476 11294
rect 7420 11190 7476 11228
rect 6972 11116 7252 11172
rect 7308 11170 7364 11182
rect 7308 11118 7310 11170
rect 7362 11118 7364 11170
rect 6636 10892 6916 10948
rect 6300 9940 6356 10556
rect 6076 9874 6132 9884
rect 6300 9874 6356 9884
rect 6188 9716 6244 9726
rect 6188 9622 6244 9660
rect 6860 9268 6916 10892
rect 6860 9174 6916 9212
rect 6412 9044 6468 9054
rect 6412 8950 6468 8988
rect 6636 9044 6692 9054
rect 6636 8950 6692 8988
rect 6524 8932 6580 8942
rect 6524 8838 6580 8876
rect 6076 8258 6132 8270
rect 6076 8206 6078 8258
rect 6130 8206 6132 8258
rect 6076 7700 6132 8206
rect 6860 8258 6916 8270
rect 6860 8206 6862 8258
rect 6914 8206 6916 8258
rect 6300 8148 6356 8158
rect 6524 8148 6580 8158
rect 6300 8146 6468 8148
rect 6300 8094 6302 8146
rect 6354 8094 6468 8146
rect 6300 8092 6468 8094
rect 6300 8082 6356 8092
rect 6412 7812 6468 8092
rect 6524 8054 6580 8092
rect 6860 7924 6916 8206
rect 6972 8260 7028 11116
rect 7196 10052 7252 10062
rect 6972 8194 7028 8204
rect 7084 8484 7140 8494
rect 7084 8036 7140 8428
rect 7196 8370 7252 9996
rect 7308 8708 7364 11118
rect 7532 10052 7588 11342
rect 7868 11284 7924 11294
rect 7868 11190 7924 11228
rect 8092 11170 8148 12012
rect 8316 11732 8372 12126
rect 8316 11666 8372 11676
rect 8204 11284 8260 11294
rect 8204 11282 8372 11284
rect 8204 11230 8206 11282
rect 8258 11230 8372 11282
rect 8204 11228 8372 11230
rect 8204 11218 8260 11228
rect 8092 11118 8094 11170
rect 8146 11118 8148 11170
rect 7868 10948 7924 10958
rect 7868 10610 7924 10892
rect 7868 10558 7870 10610
rect 7922 10558 7924 10610
rect 7868 10052 7924 10558
rect 7532 9986 7588 9996
rect 7644 9996 7924 10052
rect 7980 10722 8036 10734
rect 7980 10670 7982 10722
rect 8034 10670 8036 10722
rect 7644 9042 7700 9996
rect 7868 9828 7924 9838
rect 7980 9828 8036 10670
rect 8092 10612 8148 11118
rect 8092 10546 8148 10556
rect 8204 10610 8260 10622
rect 8204 10558 8206 10610
rect 8258 10558 8260 10610
rect 8204 10500 8260 10558
rect 8204 10434 8260 10444
rect 8316 10276 8372 11228
rect 7924 9772 8036 9828
rect 8204 10220 8372 10276
rect 7868 9266 7924 9772
rect 8204 9492 8260 10220
rect 8428 9940 8484 12236
rect 8652 12226 8708 12236
rect 8988 12198 9044 12236
rect 9548 12290 9604 12302
rect 9548 12238 9550 12290
rect 9602 12238 9604 12290
rect 9548 11788 9604 12238
rect 10556 12292 10612 12302
rect 10556 12198 10612 12236
rect 10332 12180 10388 12190
rect 9324 11732 9604 11788
rect 9996 12178 10388 12180
rect 9996 12126 10334 12178
rect 10386 12126 10388 12178
rect 9996 12124 10388 12126
rect 8652 11620 8708 11630
rect 8652 11526 8708 11564
rect 8876 11620 8932 11630
rect 8876 11526 8932 11564
rect 8988 11394 9044 11406
rect 8988 11342 8990 11394
rect 9042 11342 9044 11394
rect 8540 11282 8596 11294
rect 8540 11230 8542 11282
rect 8594 11230 8596 11282
rect 8540 10610 8596 11230
rect 8540 10558 8542 10610
rect 8594 10558 8596 10610
rect 8540 10546 8596 10558
rect 8876 11060 8932 11070
rect 8876 10610 8932 11004
rect 8988 10948 9044 11342
rect 8988 10882 9044 10892
rect 9100 11396 9156 11406
rect 8988 10724 9044 10734
rect 9100 10724 9156 11340
rect 8988 10722 9156 10724
rect 8988 10670 8990 10722
rect 9042 10670 9156 10722
rect 8988 10668 9156 10670
rect 9324 10724 9380 11732
rect 9884 11508 9940 11518
rect 9996 11508 10052 12124
rect 10332 12114 10388 12124
rect 11004 12178 11060 12190
rect 11004 12126 11006 12178
rect 11058 12126 11060 12178
rect 10780 12066 10836 12078
rect 10780 12014 10782 12066
rect 10834 12014 10836 12066
rect 9884 11506 10052 11508
rect 9884 11454 9886 11506
rect 9938 11454 10052 11506
rect 9884 11452 10052 11454
rect 10668 11508 10724 11518
rect 9884 11442 9940 11452
rect 10668 11414 10724 11452
rect 9548 11394 9604 11406
rect 9548 11342 9550 11394
rect 9602 11342 9604 11394
rect 9548 11172 9604 11342
rect 10444 11396 10500 11406
rect 10444 11302 10500 11340
rect 9660 11284 9716 11294
rect 9996 11284 10052 11294
rect 9660 11190 9716 11228
rect 9884 11282 10052 11284
rect 9884 11230 9998 11282
rect 10050 11230 10052 11282
rect 9884 11228 10052 11230
rect 9548 11106 9604 11116
rect 9528 11004 9792 11014
rect 9584 10948 9632 11004
rect 9688 10948 9736 11004
rect 9528 10938 9792 10948
rect 9884 10836 9940 11228
rect 9996 11218 10052 11228
rect 10780 11284 10836 12014
rect 10780 11218 10836 11228
rect 10668 11172 10724 11182
rect 10556 11170 10724 11172
rect 10556 11118 10670 11170
rect 10722 11118 10724 11170
rect 10556 11116 10724 11118
rect 10556 11060 10612 11116
rect 10668 11106 10724 11116
rect 8988 10658 9044 10668
rect 9324 10658 9380 10668
rect 9436 10780 9940 10836
rect 10332 11004 10612 11060
rect 10332 10834 10388 11004
rect 10892 10836 10948 10846
rect 10332 10782 10334 10834
rect 10386 10782 10388 10834
rect 8876 10558 8878 10610
rect 8930 10558 8932 10610
rect 8876 10546 8932 10558
rect 8204 9426 8260 9436
rect 8316 9884 8484 9940
rect 8652 10386 8708 10398
rect 8652 10334 8654 10386
rect 8706 10334 8708 10386
rect 8652 9940 8708 10334
rect 9212 10052 9268 10062
rect 8988 9996 9212 10052
rect 8876 9940 8932 9950
rect 8652 9938 8932 9940
rect 8652 9886 8878 9938
rect 8930 9886 8932 9938
rect 8652 9884 8932 9886
rect 7868 9214 7870 9266
rect 7922 9214 7924 9266
rect 7868 9202 7924 9214
rect 7756 9156 7812 9166
rect 7756 9062 7812 9100
rect 7644 8990 7646 9042
rect 7698 8990 7700 9042
rect 7644 8820 7700 8990
rect 8316 9042 8372 9884
rect 8876 9874 8932 9884
rect 8316 8990 8318 9042
rect 8370 8990 8372 9042
rect 8316 8978 8372 8990
rect 8540 9716 8596 9726
rect 8764 9716 8820 9726
rect 8596 9714 8820 9716
rect 8596 9662 8766 9714
rect 8818 9662 8820 9714
rect 8596 9660 8820 9662
rect 7644 8754 7700 8764
rect 7308 8484 7364 8652
rect 7308 8418 7364 8428
rect 7196 8318 7198 8370
rect 7250 8318 7252 8370
rect 7196 8306 7252 8318
rect 7532 8146 7588 8158
rect 7532 8094 7534 8146
rect 7586 8094 7588 8146
rect 6860 7858 6916 7868
rect 6972 8034 7140 8036
rect 6972 7982 7086 8034
rect 7138 7982 7140 8034
rect 6972 7980 7140 7982
rect 6412 7756 6804 7812
rect 6076 7634 6132 7644
rect 6748 7698 6804 7756
rect 6748 7646 6750 7698
rect 6802 7646 6804 7698
rect 6748 7634 6804 7646
rect 6860 7700 6916 7710
rect 6860 7606 6916 7644
rect 6188 7476 6244 7486
rect 6636 7476 6692 7486
rect 6188 7028 6244 7420
rect 6188 6962 6244 6972
rect 6524 7474 6692 7476
rect 6524 7422 6638 7474
rect 6690 7422 6692 7474
rect 6524 7420 6692 7422
rect 6076 6692 6132 6702
rect 6076 6578 6132 6636
rect 6412 6692 6468 6702
rect 6412 6598 6468 6636
rect 6076 6526 6078 6578
rect 6130 6526 6132 6578
rect 6076 6514 6132 6526
rect 6188 6468 6244 6478
rect 6188 6130 6244 6412
rect 6524 6356 6580 7420
rect 6636 7410 6692 7420
rect 6972 7364 7028 7980
rect 7084 7970 7140 7980
rect 7308 8034 7364 8046
rect 7308 7982 7310 8034
rect 7362 7982 7364 8034
rect 7308 7700 7364 7982
rect 6972 7298 7028 7308
rect 7084 7644 7364 7700
rect 6636 6692 6692 6702
rect 6636 6578 6692 6636
rect 6636 6526 6638 6578
rect 6690 6526 6692 6578
rect 6636 6514 6692 6526
rect 6748 6580 6804 6590
rect 6748 6578 7028 6580
rect 6748 6526 6750 6578
rect 6802 6526 7028 6578
rect 6748 6524 7028 6526
rect 6748 6514 6804 6524
rect 6860 6356 6916 6366
rect 6580 6300 6692 6356
rect 6524 6262 6580 6300
rect 6188 6078 6190 6130
rect 6242 6078 6244 6130
rect 6188 6066 6244 6078
rect 6524 5906 6580 5918
rect 6524 5854 6526 5906
rect 6578 5854 6580 5906
rect 5852 5292 6020 5348
rect 6300 5796 6356 5806
rect 4844 5030 4900 5068
rect 4956 5236 5012 5246
rect 4396 4722 4452 4732
rect 4732 4564 4788 4574
rect 4732 4470 4788 4508
rect 2492 4398 2494 4450
rect 2546 4398 2548 4450
rect 2492 4386 2548 4398
rect 4956 4452 5012 5180
rect 5516 5124 5572 5134
rect 5068 5010 5124 5022
rect 5068 4958 5070 5010
rect 5122 4958 5124 5010
rect 5068 4900 5124 4958
rect 5068 4834 5124 4844
rect 5180 4452 5236 4462
rect 4956 4396 5180 4452
rect 5180 4358 5236 4396
rect 1820 4340 1876 4350
rect 1820 4246 1876 4284
rect 5516 4338 5572 5068
rect 5740 4564 5796 4574
rect 5628 4508 5740 4564
rect 5628 4450 5684 4508
rect 5740 4498 5796 4508
rect 5628 4398 5630 4450
rect 5682 4398 5684 4450
rect 5628 4386 5684 4398
rect 5516 4286 5518 4338
rect 5570 4286 5572 4338
rect 5516 4274 5572 4286
rect 5740 4338 5796 4350
rect 5740 4286 5742 4338
rect 5794 4286 5796 4338
rect 1596 4162 1652 4172
rect 3612 4228 3668 4238
rect 3612 800 3668 4172
rect 5740 4228 5796 4286
rect 5740 4162 5796 4172
rect 5852 4340 5908 5292
rect 5964 5124 6020 5134
rect 5964 4564 6020 5068
rect 6188 4900 6244 4910
rect 6188 4806 6244 4844
rect 6300 4898 6356 5740
rect 6300 4846 6302 4898
rect 6354 4846 6356 4898
rect 6300 4834 6356 4846
rect 6076 4564 6132 4574
rect 5964 4562 6132 4564
rect 5964 4510 6078 4562
rect 6130 4510 6132 4562
rect 5964 4508 6132 4510
rect 6076 4498 6132 4508
rect 6412 4564 6468 4574
rect 6524 4564 6580 5854
rect 6636 5012 6692 6300
rect 6748 6018 6804 6030
rect 6748 5966 6750 6018
rect 6802 5966 6804 6018
rect 6748 5796 6804 5966
rect 6860 6018 6916 6300
rect 6860 5966 6862 6018
rect 6914 5966 6916 6018
rect 6860 5954 6916 5966
rect 6972 6020 7028 6524
rect 7084 6468 7140 7644
rect 7084 6402 7140 6412
rect 7196 7476 7252 7486
rect 7196 6130 7252 7420
rect 7196 6078 7198 6130
rect 7250 6078 7252 6130
rect 7196 6066 7252 6078
rect 7532 6132 7588 8094
rect 8428 8036 8484 8046
rect 8092 8034 8484 8036
rect 8092 7982 8430 8034
rect 8482 7982 8484 8034
rect 8092 7980 8484 7982
rect 7868 7700 7924 7710
rect 7868 7474 7924 7644
rect 8092 7698 8148 7980
rect 8428 7970 8484 7980
rect 8092 7646 8094 7698
rect 8146 7646 8148 7698
rect 8092 7634 8148 7646
rect 7868 7422 7870 7474
rect 7922 7422 7924 7474
rect 7756 6804 7812 6842
rect 7756 6738 7812 6748
rect 7644 6692 7700 6702
rect 7644 6598 7700 6636
rect 7868 6244 7924 7422
rect 7980 7476 8036 7486
rect 7980 7474 8148 7476
rect 7980 7422 7982 7474
rect 8034 7422 8148 7474
rect 7980 7420 8148 7422
rect 7980 7410 8036 7420
rect 7980 6692 8036 6702
rect 7980 6578 8036 6636
rect 7980 6526 7982 6578
rect 8034 6526 8036 6578
rect 7980 6356 8036 6526
rect 7980 6290 8036 6300
rect 8092 6468 8148 7420
rect 8204 7474 8260 7486
rect 8204 7422 8206 7474
rect 8258 7422 8260 7474
rect 8204 7364 8260 7422
rect 8204 7298 8260 7308
rect 8428 7476 8484 7486
rect 8540 7476 8596 9660
rect 8764 9650 8820 9660
rect 8988 9044 9044 9996
rect 9212 9958 9268 9996
rect 9324 9940 9380 9950
rect 9100 9828 9156 9838
rect 9324 9828 9380 9884
rect 9100 9826 9380 9828
rect 9100 9774 9102 9826
rect 9154 9774 9380 9826
rect 9100 9772 9380 9774
rect 9100 9762 9156 9772
rect 9436 9604 9492 10780
rect 10332 10770 10388 10782
rect 10444 10834 10948 10836
rect 10444 10782 10894 10834
rect 10946 10782 10948 10834
rect 10444 10780 10948 10782
rect 9996 10724 10052 10734
rect 9548 10612 9604 10622
rect 9548 10518 9604 10556
rect 9884 10610 9940 10622
rect 9884 10558 9886 10610
rect 9938 10558 9940 10610
rect 9548 10052 9604 10062
rect 9548 9828 9604 9996
rect 9548 9734 9604 9772
rect 9212 9548 9492 9604
rect 8764 8146 8820 8158
rect 8764 8094 8766 8146
rect 8818 8094 8820 8146
rect 8428 7474 8596 7476
rect 8428 7422 8430 7474
rect 8482 7422 8596 7474
rect 8428 7420 8596 7422
rect 8652 8034 8708 8046
rect 8652 7982 8654 8034
rect 8706 7982 8708 8034
rect 8428 6804 8484 7420
rect 8652 6916 8708 7982
rect 7756 6188 7924 6244
rect 7644 6132 7700 6170
rect 7532 6076 7644 6132
rect 7644 6066 7700 6076
rect 6860 5796 6916 5806
rect 6748 5740 6860 5796
rect 6860 5730 6916 5740
rect 6636 4946 6692 4956
rect 6412 4562 6580 4564
rect 6412 4510 6414 4562
rect 6466 4510 6580 4562
rect 6412 4508 6580 4510
rect 6412 4498 6468 4508
rect 5370 3948 5634 3958
rect 5426 3892 5474 3948
rect 5530 3892 5578 3948
rect 5370 3882 5634 3892
rect 5740 3668 5796 3678
rect 5852 3668 5908 4284
rect 5740 3666 5908 3668
rect 5740 3614 5742 3666
rect 5794 3614 5908 3666
rect 5740 3612 5908 3614
rect 5740 3602 5796 3612
rect 6524 3554 6580 4508
rect 6748 4788 6804 4798
rect 6636 4340 6692 4350
rect 6636 3778 6692 4284
rect 6636 3726 6638 3778
rect 6690 3726 6692 3778
rect 6636 3714 6692 3726
rect 6748 4338 6804 4732
rect 6860 4452 6916 4462
rect 6860 4358 6916 4396
rect 6748 4286 6750 4338
rect 6802 4286 6804 4338
rect 6748 3780 6804 4286
rect 6860 4228 6916 4238
rect 6972 4228 7028 5964
rect 7420 5906 7476 5918
rect 7420 5854 7422 5906
rect 7474 5854 7476 5906
rect 7196 5682 7252 5694
rect 7196 5630 7198 5682
rect 7250 5630 7252 5682
rect 7196 5010 7252 5630
rect 7196 4958 7198 5010
rect 7250 4958 7252 5010
rect 7196 4676 7252 4958
rect 7196 4610 7252 4620
rect 7308 5572 7364 5582
rect 7084 4564 7140 4574
rect 7084 4470 7140 4508
rect 7308 4452 7364 5516
rect 7420 5122 7476 5854
rect 7420 5070 7422 5122
rect 7474 5070 7476 5122
rect 7420 5012 7476 5070
rect 7756 5012 7812 6188
rect 7980 6132 8036 6142
rect 7980 6038 8036 6076
rect 7868 6018 7924 6030
rect 7868 5966 7870 6018
rect 7922 5966 7924 6018
rect 7868 5908 7924 5966
rect 7868 5842 7924 5852
rect 8092 5122 8148 6412
rect 8316 6748 8484 6804
rect 8540 6860 8708 6916
rect 8204 6244 8260 6254
rect 8316 6244 8372 6748
rect 8540 6580 8596 6860
rect 8260 6188 8372 6244
rect 8428 6524 8596 6580
rect 8652 6690 8708 6702
rect 8652 6638 8654 6690
rect 8706 6638 8708 6690
rect 8204 6130 8260 6188
rect 8204 6078 8206 6130
rect 8258 6078 8260 6130
rect 8204 6066 8260 6078
rect 8428 6018 8484 6524
rect 8652 6356 8708 6638
rect 8652 6290 8708 6300
rect 8428 5966 8430 6018
rect 8482 5966 8484 6018
rect 8428 5908 8484 5966
rect 8428 5842 8484 5852
rect 8540 6244 8596 6254
rect 8092 5070 8094 5122
rect 8146 5070 8148 5122
rect 8092 5058 8148 5070
rect 7868 5012 7924 5022
rect 7420 4956 7700 5012
rect 7756 5010 7924 5012
rect 7756 4958 7870 5010
rect 7922 4958 7924 5010
rect 7756 4956 7924 4958
rect 7532 4788 7588 4798
rect 7532 4562 7588 4732
rect 7532 4510 7534 4562
rect 7586 4510 7588 4562
rect 7532 4498 7588 4510
rect 7420 4452 7476 4462
rect 7308 4396 7420 4452
rect 7420 4358 7476 4396
rect 7644 4340 7700 4956
rect 7868 4788 7924 4956
rect 7868 4722 7924 4732
rect 8204 5012 8260 5022
rect 7756 4564 7812 4574
rect 7756 4470 7812 4508
rect 8204 4452 8260 4956
rect 8316 4452 8372 4462
rect 8204 4450 8372 4452
rect 8204 4398 8318 4450
rect 8370 4398 8372 4450
rect 8204 4396 8372 4398
rect 8092 4340 8148 4350
rect 8316 4340 8372 4396
rect 7644 4338 8260 4340
rect 7644 4286 8094 4338
rect 8146 4286 8260 4338
rect 7644 4284 8260 4286
rect 8092 4274 8148 4284
rect 6916 4172 7028 4228
rect 6860 4162 6916 4172
rect 6748 3714 6804 3724
rect 8204 3778 8260 4284
rect 8316 4274 8372 4284
rect 8204 3726 8206 3778
rect 8258 3726 8260 3778
rect 8204 3714 8260 3726
rect 8316 3668 8372 3678
rect 8540 3668 8596 6188
rect 8764 6132 8820 8094
rect 8988 8146 9044 8988
rect 8988 8094 8990 8146
rect 9042 8094 9044 8146
rect 8988 8082 9044 8094
rect 9100 9492 9156 9502
rect 8876 7700 8932 7710
rect 8876 7606 8932 7644
rect 8988 7474 9044 7486
rect 8988 7422 8990 7474
rect 9042 7422 9044 7474
rect 8876 7252 8932 7262
rect 8876 7158 8932 7196
rect 8876 6466 8932 6478
rect 8876 6414 8878 6466
rect 8930 6414 8932 6466
rect 8876 6244 8932 6414
rect 8988 6468 9044 7422
rect 8988 6402 9044 6412
rect 8876 6178 8932 6188
rect 8764 6066 8820 6076
rect 8876 6020 8932 6030
rect 8652 5906 8708 5918
rect 8652 5854 8654 5906
rect 8706 5854 8708 5906
rect 8652 5348 8708 5854
rect 8876 5906 8932 5964
rect 8876 5854 8878 5906
rect 8930 5854 8932 5906
rect 8876 5842 8932 5854
rect 8988 5796 9044 5806
rect 9100 5796 9156 9436
rect 9212 8370 9268 9548
rect 9528 9436 9792 9446
rect 9584 9380 9632 9436
rect 9688 9380 9736 9436
rect 9528 9370 9792 9380
rect 9884 9380 9940 10558
rect 9996 10610 10052 10668
rect 10444 10722 10500 10780
rect 10892 10770 10948 10780
rect 10444 10670 10446 10722
rect 10498 10670 10500 10722
rect 10444 10658 10500 10670
rect 9996 10558 9998 10610
rect 10050 10558 10052 10610
rect 9996 10546 10052 10558
rect 10668 10610 10724 10622
rect 10668 10558 10670 10610
rect 10722 10558 10724 10610
rect 10220 10500 10276 10510
rect 10220 10406 10276 10444
rect 10668 10388 10724 10558
rect 10668 10322 10724 10332
rect 10556 9940 10612 9950
rect 10108 9938 10612 9940
rect 10108 9886 10558 9938
rect 10610 9886 10612 9938
rect 10108 9884 10612 9886
rect 9996 9714 10052 9726
rect 9996 9662 9998 9714
rect 10050 9662 10052 9714
rect 9996 9380 10052 9662
rect 10108 9714 10164 9884
rect 10556 9874 10612 9884
rect 10668 9940 10724 9950
rect 11004 9940 11060 12126
rect 11116 11620 11172 11630
rect 11116 10722 11172 11564
rect 11116 10670 11118 10722
rect 11170 10670 11172 10722
rect 11116 10164 11172 10670
rect 11116 10098 11172 10108
rect 10444 9716 10500 9726
rect 10668 9716 10724 9884
rect 10108 9662 10110 9714
rect 10162 9662 10164 9714
rect 10108 9650 10164 9662
rect 10332 9660 10444 9716
rect 10332 9602 10388 9660
rect 10444 9650 10500 9660
rect 10556 9714 10724 9716
rect 10556 9662 10670 9714
rect 10722 9662 10724 9714
rect 10556 9660 10724 9662
rect 10332 9550 10334 9602
rect 10386 9550 10388 9602
rect 10332 9538 10388 9550
rect 9996 9324 10388 9380
rect 9884 9314 9940 9324
rect 9660 9268 9716 9278
rect 9548 9042 9604 9054
rect 9548 8990 9550 9042
rect 9602 8990 9604 9042
rect 9548 8820 9604 8990
rect 9548 8754 9604 8764
rect 9212 8318 9214 8370
rect 9266 8318 9268 8370
rect 9212 8306 9268 8318
rect 9660 8370 9716 9212
rect 10108 9154 10164 9166
rect 9660 8318 9662 8370
rect 9714 8318 9716 8370
rect 9660 8306 9716 8318
rect 9772 9098 9828 9110
rect 9772 9046 9774 9098
rect 9826 9046 9828 9098
rect 9436 8260 9492 8270
rect 9324 8258 9492 8260
rect 9324 8206 9438 8258
rect 9490 8206 9492 8258
rect 9324 8204 9492 8206
rect 9212 7252 9268 7262
rect 9324 7252 9380 8204
rect 9436 8194 9492 8204
rect 9772 8148 9828 9046
rect 9884 9098 9940 9110
rect 9884 9046 9886 9098
rect 9938 9046 9940 9098
rect 9884 8596 9940 9046
rect 10108 9102 10110 9154
rect 10162 9102 10164 9154
rect 10108 9044 10164 9102
rect 10108 8978 10164 8988
rect 10332 8930 10388 9324
rect 10332 8878 10334 8930
rect 10386 8878 10388 8930
rect 10332 8866 10388 8878
rect 9884 8540 10052 8596
rect 9884 8372 9940 8382
rect 9884 8258 9940 8316
rect 9884 8206 9886 8258
rect 9938 8206 9940 8258
rect 9884 8194 9940 8206
rect 9772 8082 9828 8092
rect 9996 7924 10052 8540
rect 10556 8484 10612 9660
rect 10668 9650 10724 9660
rect 10780 9884 11060 9940
rect 11228 9940 11284 12684
rect 11340 12646 11396 12684
rect 12012 12740 12068 12750
rect 12012 12646 12068 12684
rect 10780 9716 10836 9884
rect 11228 9874 11284 9884
rect 11340 11732 11396 11742
rect 11340 10610 11396 11676
rect 11340 10558 11342 10610
rect 11394 10558 11396 10610
rect 10780 9650 10836 9660
rect 10892 9716 10948 9726
rect 11228 9716 11284 9726
rect 11340 9716 11396 10558
rect 10892 9714 11060 9716
rect 10892 9662 10894 9714
rect 10946 9662 11060 9714
rect 10892 9660 11060 9662
rect 10892 9650 10948 9660
rect 10108 8146 10164 8158
rect 10444 8148 10500 8158
rect 10108 8094 10110 8146
rect 10162 8094 10164 8146
rect 10108 8036 10164 8094
rect 10108 7970 10164 7980
rect 10332 8146 10500 8148
rect 10332 8094 10446 8146
rect 10498 8094 10500 8146
rect 10332 8092 10500 8094
rect 9528 7868 9792 7878
rect 9584 7812 9632 7868
rect 9688 7812 9736 7868
rect 9528 7802 9792 7812
rect 9884 7868 10052 7924
rect 9660 7700 9716 7710
rect 9884 7700 9940 7868
rect 9660 7698 9940 7700
rect 9660 7646 9662 7698
rect 9714 7646 9940 7698
rect 9660 7644 9940 7646
rect 9996 7700 10052 7710
rect 9660 7634 9716 7644
rect 9268 7196 9380 7252
rect 9548 7474 9604 7486
rect 9548 7422 9550 7474
rect 9602 7422 9604 7474
rect 9212 7186 9268 7196
rect 9548 6692 9604 7422
rect 9772 7476 9828 7486
rect 9996 7476 10052 7644
rect 10332 7588 10388 8092
rect 10444 8082 10500 8092
rect 10556 7698 10612 8428
rect 10556 7646 10558 7698
rect 10610 7646 10612 7698
rect 10556 7634 10612 7646
rect 10668 9268 10724 9278
rect 10332 7522 10388 7532
rect 9772 7474 10052 7476
rect 9772 7422 9774 7474
rect 9826 7422 10052 7474
rect 9772 7420 10052 7422
rect 10220 7474 10276 7486
rect 10220 7422 10222 7474
rect 10274 7422 10276 7474
rect 9660 6804 9716 6814
rect 9772 6804 9828 7420
rect 10220 7252 10276 7422
rect 10668 7364 10724 9212
rect 11004 9044 11060 9660
rect 11228 9714 11396 9716
rect 11228 9662 11230 9714
rect 11282 9662 11396 9714
rect 11228 9660 11396 9662
rect 11452 10052 11508 10062
rect 11452 9826 11508 9996
rect 11900 9940 11956 9950
rect 11452 9774 11454 9826
rect 11506 9774 11508 9826
rect 11228 9650 11284 9660
rect 11452 9268 11508 9774
rect 11564 9828 11620 9838
rect 11564 9826 11844 9828
rect 11564 9774 11566 9826
rect 11618 9774 11844 9826
rect 11564 9772 11844 9774
rect 11564 9762 11620 9772
rect 11452 9202 11508 9212
rect 11788 9716 11844 9772
rect 11004 8988 11620 9044
rect 11340 8818 11396 8830
rect 11340 8766 11342 8818
rect 11394 8766 11396 8818
rect 11340 8372 11396 8766
rect 11340 8306 11396 8316
rect 11452 8820 11508 8830
rect 11116 8146 11172 8158
rect 11116 8094 11118 8146
rect 11170 8094 11172 8146
rect 11004 7588 11060 7598
rect 10892 7532 11004 7588
rect 10892 7474 10948 7532
rect 11004 7522 11060 7532
rect 10892 7422 10894 7474
rect 10946 7422 10948 7474
rect 10892 7410 10948 7422
rect 9996 7196 10220 7252
rect 9716 6748 9828 6804
rect 9884 7028 9940 7038
rect 9660 6738 9716 6748
rect 9212 6636 9604 6692
rect 9212 6020 9268 6636
rect 9660 6468 9716 6478
rect 9212 5954 9268 5964
rect 9324 6466 9716 6468
rect 9324 6414 9662 6466
rect 9714 6414 9716 6466
rect 9324 6412 9716 6414
rect 8988 5794 9156 5796
rect 8988 5742 8990 5794
rect 9042 5742 9156 5794
rect 8988 5740 9156 5742
rect 8988 5730 9044 5740
rect 9324 5684 9380 6412
rect 9660 6402 9716 6412
rect 9528 6300 9792 6310
rect 9584 6244 9632 6300
rect 9688 6244 9736 6300
rect 9528 6234 9792 6244
rect 9436 5908 9492 5918
rect 9492 5852 9716 5908
rect 9436 5842 9492 5852
rect 9324 5618 9380 5628
rect 8652 4900 8708 5292
rect 8876 5236 8932 5246
rect 8876 5122 8932 5180
rect 8876 5070 8878 5122
rect 8930 5070 8932 5122
rect 8876 5058 8932 5070
rect 9100 5122 9156 5134
rect 9100 5070 9102 5122
rect 9154 5070 9156 5122
rect 8652 4834 8708 4844
rect 8988 4788 9044 4798
rect 8652 4452 8708 4462
rect 8652 4358 8708 4396
rect 8988 4450 9044 4732
rect 9100 4564 9156 5070
rect 9436 5012 9492 5022
rect 9436 4918 9492 4956
rect 9660 5010 9716 5852
rect 9660 4958 9662 5010
rect 9714 4958 9716 5010
rect 9660 4946 9716 4958
rect 9884 5124 9940 6972
rect 9996 6914 10052 7196
rect 10220 7186 10276 7196
rect 10556 7308 10724 7364
rect 9996 6862 9998 6914
rect 10050 6862 10052 6914
rect 9996 6850 10052 6862
rect 10220 6690 10276 6702
rect 10220 6638 10222 6690
rect 10274 6638 10276 6690
rect 10220 6132 10276 6638
rect 10556 6578 10612 7308
rect 10892 7252 10948 7262
rect 10892 6690 10948 7196
rect 10892 6638 10894 6690
rect 10946 6638 10948 6690
rect 10892 6626 10948 6638
rect 10556 6526 10558 6578
rect 10610 6526 10612 6578
rect 10556 6514 10612 6526
rect 10220 6066 10276 6076
rect 10780 5348 10836 5358
rect 10780 5234 10836 5292
rect 10780 5182 10782 5234
rect 10834 5182 10836 5234
rect 10780 5170 10836 5182
rect 10892 5236 10948 5246
rect 10892 5142 10948 5180
rect 10108 5124 10164 5134
rect 9884 5122 10164 5124
rect 9884 5070 10110 5122
rect 10162 5070 10164 5122
rect 9884 5068 10164 5070
rect 11116 5124 11172 8094
rect 11452 8146 11508 8764
rect 11452 8094 11454 8146
rect 11506 8094 11508 8146
rect 11452 8082 11508 8094
rect 11564 7698 11620 8988
rect 11676 8818 11732 8830
rect 11676 8766 11678 8818
rect 11730 8766 11732 8818
rect 11676 8372 11732 8766
rect 11788 8596 11844 9660
rect 11900 9042 11956 9884
rect 12236 9940 12292 13468
rect 12572 12964 12628 12974
rect 12572 12870 12628 12908
rect 12684 12178 12740 14252
rect 12684 12126 12686 12178
rect 12738 12126 12740 12178
rect 12684 12114 12740 12126
rect 13468 12068 13524 15260
rect 14028 15316 14084 15326
rect 14252 15316 14308 15822
rect 14812 15876 14868 15886
rect 14812 15538 14868 15820
rect 14812 15486 14814 15538
rect 14866 15486 14868 15538
rect 14812 15474 14868 15486
rect 14700 15428 14756 15438
rect 14700 15334 14756 15372
rect 14084 15260 14308 15316
rect 14028 15202 14084 15260
rect 14028 15150 14030 15202
rect 14082 15150 14084 15202
rect 14028 15138 14084 15150
rect 13686 14924 13950 14934
rect 13742 14868 13790 14924
rect 13846 14868 13894 14924
rect 13686 14858 13950 14868
rect 13580 14308 13636 14318
rect 13580 14214 13636 14252
rect 13686 13356 13950 13366
rect 13742 13300 13790 13356
rect 13846 13300 13894 13356
rect 13686 13290 13950 13300
rect 13804 12852 13860 12862
rect 13804 12758 13860 12796
rect 14140 12852 14196 12862
rect 14140 12758 14196 12796
rect 14924 12852 14980 18956
rect 15820 17666 15876 17678
rect 15820 17614 15822 17666
rect 15874 17614 15876 17666
rect 15820 17106 15876 17614
rect 15932 17556 15988 19740
rect 16828 18564 16884 18574
rect 16044 18340 16100 18350
rect 16044 17778 16100 18284
rect 16044 17726 16046 17778
rect 16098 17726 16100 17778
rect 16044 17714 16100 17726
rect 16492 18340 16548 18350
rect 16156 17666 16212 17678
rect 16156 17614 16158 17666
rect 16210 17614 16212 17666
rect 16156 17556 16212 17614
rect 16492 17666 16548 18284
rect 16492 17614 16494 17666
rect 16546 17614 16548 17666
rect 16492 17602 16548 17614
rect 16828 18338 16884 18508
rect 16828 18286 16830 18338
rect 16882 18286 16884 18338
rect 15932 17500 16100 17556
rect 15820 17054 15822 17106
rect 15874 17054 15876 17106
rect 15820 17042 15876 17054
rect 15260 16996 15316 17006
rect 15036 16994 15316 16996
rect 15036 16942 15262 16994
rect 15314 16942 15316 16994
rect 15036 16940 15316 16942
rect 15036 15986 15092 16940
rect 15260 16884 15316 16940
rect 15932 16996 15988 17006
rect 15932 16902 15988 16940
rect 15260 16818 15316 16828
rect 15372 16882 15428 16894
rect 15372 16830 15374 16882
rect 15426 16830 15428 16882
rect 15260 16660 15316 16670
rect 15260 16566 15316 16604
rect 15260 16100 15316 16110
rect 15036 15934 15038 15986
rect 15090 15934 15092 15986
rect 15036 15922 15092 15934
rect 15148 15988 15204 16026
rect 15148 15922 15204 15932
rect 15148 15764 15204 15774
rect 15148 15148 15204 15708
rect 15260 15540 15316 16044
rect 15372 15652 15428 16830
rect 15708 16882 15764 16894
rect 15708 16830 15710 16882
rect 15762 16830 15764 16882
rect 15708 16436 15764 16830
rect 16044 16772 16100 17500
rect 16156 17490 16212 17500
rect 16716 16996 16772 17006
rect 16716 16902 16772 16940
rect 16380 16884 16436 16894
rect 16380 16882 16660 16884
rect 16380 16830 16382 16882
rect 16434 16830 16660 16882
rect 16380 16828 16660 16830
rect 16380 16818 16436 16828
rect 15596 16380 15764 16436
rect 15820 16716 16100 16772
rect 15484 16098 15540 16110
rect 15484 16046 15486 16098
rect 15538 16046 15540 16098
rect 15484 15876 15540 16046
rect 15484 15810 15540 15820
rect 15372 15596 15540 15652
rect 15260 15484 15428 15540
rect 15260 15316 15316 15326
rect 15260 15222 15316 15260
rect 15372 15314 15428 15484
rect 15484 15538 15540 15596
rect 15484 15486 15486 15538
rect 15538 15486 15540 15538
rect 15484 15474 15540 15486
rect 15596 15538 15652 16380
rect 15708 16098 15764 16110
rect 15708 16046 15710 16098
rect 15762 16046 15764 16098
rect 15708 15764 15764 16046
rect 15708 15698 15764 15708
rect 15596 15486 15598 15538
rect 15650 15486 15652 15538
rect 15372 15262 15374 15314
rect 15426 15262 15428 15314
rect 15372 15250 15428 15262
rect 15596 15428 15652 15486
rect 15148 15092 15316 15148
rect 14924 12786 14980 12796
rect 15260 13746 15316 15092
rect 15596 14196 15652 15372
rect 15596 14130 15652 14140
rect 15708 15314 15764 15326
rect 15708 15262 15710 15314
rect 15762 15262 15764 15314
rect 15708 13972 15764 15262
rect 15820 14644 15876 16716
rect 16492 16660 16548 16670
rect 16380 16604 16492 16660
rect 15932 16436 15988 16446
rect 15932 16098 15988 16380
rect 15932 16046 15934 16098
rect 15986 16046 15988 16098
rect 15932 15764 15988 16046
rect 16044 15988 16100 15998
rect 16044 15894 16100 15932
rect 16156 15988 16212 15998
rect 16380 15988 16436 16604
rect 16492 16594 16548 16604
rect 16156 15986 16380 15988
rect 16156 15934 16158 15986
rect 16210 15934 16380 15986
rect 16156 15932 16380 15934
rect 16156 15922 16212 15932
rect 16380 15894 16436 15932
rect 16604 16098 16660 16828
rect 16828 16882 16884 18286
rect 16940 17108 16996 20076
rect 17500 20018 17556 20412
rect 17500 19966 17502 20018
rect 17554 19966 17556 20018
rect 17500 19954 17556 19966
rect 17612 19458 17668 20636
rect 17612 19406 17614 19458
rect 17666 19406 17668 19458
rect 17612 19394 17668 19406
rect 17388 19348 17444 19358
rect 17388 19254 17444 19292
rect 17500 18564 17556 18574
rect 17556 18508 17668 18564
rect 17500 18498 17556 18508
rect 17388 18450 17444 18462
rect 17388 18398 17390 18450
rect 17442 18398 17444 18450
rect 17164 17556 17220 17566
rect 17388 17556 17444 18398
rect 17612 18450 17668 18508
rect 17612 18398 17614 18450
rect 17666 18398 17668 18450
rect 17612 18386 17668 18398
rect 17500 18340 17556 18350
rect 17500 18246 17556 18284
rect 17724 18004 17780 20636
rect 17836 20580 17892 21196
rect 18060 20580 18116 20590
rect 17892 20578 18116 20580
rect 17892 20526 18062 20578
rect 18114 20526 18116 20578
rect 17892 20524 18116 20526
rect 17836 20514 17892 20524
rect 18060 20514 18116 20524
rect 17844 20412 18108 20422
rect 17900 20356 17948 20412
rect 18004 20356 18052 20412
rect 17844 20346 18108 20356
rect 17948 20018 18004 20030
rect 17948 19966 17950 20018
rect 18002 19966 18004 20018
rect 17948 19796 18004 19966
rect 18172 20020 18228 20030
rect 18172 19926 18228 19964
rect 17948 19730 18004 19740
rect 18060 19906 18116 19918
rect 18060 19854 18062 19906
rect 18114 19854 18116 19906
rect 18060 19684 18116 19854
rect 18060 19618 18116 19628
rect 17948 19012 18004 19022
rect 17948 19010 18228 19012
rect 17948 18958 17950 19010
rect 18002 18958 18228 19010
rect 17948 18956 18228 18958
rect 17948 18946 18004 18956
rect 17844 18844 18108 18854
rect 17900 18788 17948 18844
rect 18004 18788 18052 18844
rect 17844 18778 18108 18788
rect 18060 18450 18116 18462
rect 18060 18398 18062 18450
rect 18114 18398 18116 18450
rect 18060 18228 18116 18398
rect 18060 18162 18116 18172
rect 17612 17948 17780 18004
rect 17220 17500 17332 17556
rect 17164 17490 17220 17500
rect 17164 17332 17220 17342
rect 17052 17108 17108 17118
rect 16940 17052 17052 17108
rect 17052 17042 17108 17052
rect 16828 16830 16830 16882
rect 16882 16830 16884 16882
rect 16716 16660 16772 16670
rect 16716 16566 16772 16604
rect 16828 16324 16884 16830
rect 17052 16324 17108 16334
rect 16828 16268 17052 16324
rect 17052 16258 17108 16268
rect 16604 16046 16606 16098
rect 16658 16046 16660 16098
rect 15932 15708 16324 15764
rect 16268 15426 16324 15708
rect 16268 15374 16270 15426
rect 16322 15374 16324 15426
rect 16268 15362 16324 15374
rect 16380 15202 16436 15214
rect 16380 15150 16382 15202
rect 16434 15150 16436 15202
rect 15820 14578 15876 14588
rect 16156 14756 16212 14766
rect 16156 14530 16212 14700
rect 16156 14478 16158 14530
rect 16210 14478 16212 14530
rect 16156 14466 16212 14478
rect 16380 14532 16436 15150
rect 16604 14756 16660 16046
rect 16716 15988 16772 15998
rect 16716 15426 16772 15932
rect 16940 15988 16996 15998
rect 16940 15894 16996 15932
rect 16828 15874 16884 15886
rect 16828 15822 16830 15874
rect 16882 15822 16884 15874
rect 16828 15764 16884 15822
rect 17164 15876 17220 17276
rect 17276 17108 17332 17500
rect 17388 17554 17556 17556
rect 17388 17502 17390 17554
rect 17442 17502 17556 17554
rect 17388 17500 17556 17502
rect 17388 17490 17444 17500
rect 17388 17108 17444 17118
rect 17276 17106 17444 17108
rect 17276 17054 17390 17106
rect 17442 17054 17444 17106
rect 17276 17052 17444 17054
rect 17388 17042 17444 17052
rect 17276 16884 17332 16894
rect 17500 16884 17556 17500
rect 17612 17332 17668 17948
rect 18172 17780 18228 18956
rect 17724 17724 18228 17780
rect 17724 17444 17780 17724
rect 17836 17556 17892 17566
rect 18060 17556 18116 17566
rect 17892 17554 18116 17556
rect 17892 17502 18062 17554
rect 18114 17502 18116 17554
rect 17892 17500 18116 17502
rect 17836 17490 17892 17500
rect 18060 17490 18116 17500
rect 18172 17556 18228 17566
rect 17724 17350 17780 17388
rect 17612 17266 17668 17276
rect 17844 17276 18108 17286
rect 17900 17220 17948 17276
rect 18004 17220 18052 17276
rect 17844 17210 18108 17220
rect 17948 17108 18004 17118
rect 17332 16828 17556 16884
rect 17612 16994 17668 17006
rect 17612 16942 17614 16994
rect 17666 16942 17668 16994
rect 17276 16098 17332 16828
rect 17612 16772 17668 16942
rect 17612 16706 17668 16716
rect 17724 16994 17780 17006
rect 17724 16942 17726 16994
rect 17778 16942 17780 16994
rect 17724 16436 17780 16942
rect 17388 16380 17780 16436
rect 17836 16996 17892 17006
rect 17388 16210 17444 16380
rect 17388 16158 17390 16210
rect 17442 16158 17444 16210
rect 17388 16146 17444 16158
rect 17724 16212 17780 16222
rect 17836 16212 17892 16940
rect 17948 16994 18004 17052
rect 17948 16942 17950 16994
rect 18002 16942 18004 16994
rect 17948 16930 18004 16942
rect 18172 16770 18228 17500
rect 18172 16718 18174 16770
rect 18226 16718 18228 16770
rect 18172 16706 18228 16718
rect 18284 16436 18340 22092
rect 18396 23154 18452 23166
rect 18396 23102 18398 23154
rect 18450 23102 18452 23154
rect 18396 21812 18452 23102
rect 18732 23044 18788 23212
rect 18956 23202 19012 23212
rect 18620 22258 18676 22270
rect 18620 22206 18622 22258
rect 18674 22206 18676 22258
rect 18620 21812 18676 22206
rect 18732 22036 18788 22988
rect 18732 21970 18788 21980
rect 18844 23156 18900 23166
rect 18844 21812 18900 23100
rect 18620 21756 18900 21812
rect 18396 21746 18452 21756
rect 18396 20578 18452 20590
rect 18396 20526 18398 20578
rect 18450 20526 18452 20578
rect 18396 19908 18452 20526
rect 18844 20244 18900 21756
rect 19180 23154 19236 23166
rect 19180 23102 19182 23154
rect 19234 23102 19236 23154
rect 18620 20188 18900 20244
rect 18956 21474 19012 21486
rect 18956 21422 18958 21474
rect 19010 21422 19012 21474
rect 18956 20244 19012 21422
rect 19180 21364 19236 23102
rect 19292 22594 19348 23660
rect 19292 22542 19294 22594
rect 19346 22542 19348 22594
rect 19292 22530 19348 22542
rect 19404 22482 19460 23884
rect 19516 23716 19572 23726
rect 19628 23716 19684 27132
rect 20076 26908 20132 27806
rect 20300 27860 20356 27870
rect 20300 27766 20356 27804
rect 20636 27858 20692 27870
rect 20636 27806 20638 27858
rect 20690 27806 20692 27858
rect 20524 27746 20580 27758
rect 20524 27694 20526 27746
rect 20578 27694 20580 27746
rect 19964 26852 20132 26908
rect 20300 27186 20356 27198
rect 20300 27134 20302 27186
rect 20354 27134 20356 27186
rect 19516 23714 19684 23716
rect 19516 23662 19518 23714
rect 19570 23662 19684 23714
rect 19516 23660 19684 23662
rect 19516 23650 19572 23660
rect 19516 23156 19572 23194
rect 19516 23090 19572 23100
rect 19516 22932 19572 22942
rect 19628 22932 19684 23660
rect 19740 26292 19796 26302
rect 19740 23156 19796 26236
rect 19964 25618 20020 26852
rect 20300 26404 20356 27134
rect 20300 25732 20356 26348
rect 20524 26402 20580 27694
rect 20636 27188 20692 27806
rect 22002 27468 22266 27478
rect 22058 27412 22106 27468
rect 22162 27412 22210 27468
rect 22002 27402 22266 27412
rect 30318 27468 30582 27478
rect 30374 27412 30422 27468
rect 30478 27412 30526 27468
rect 30318 27402 30582 27412
rect 20636 27122 20692 27132
rect 20636 26964 20692 26974
rect 20636 26870 20692 26908
rect 20748 26962 20804 26974
rect 20748 26910 20750 26962
rect 20802 26910 20804 26962
rect 20524 26350 20526 26402
rect 20578 26350 20580 26402
rect 20524 26338 20580 26350
rect 20300 25666 20356 25676
rect 19964 25566 19966 25618
rect 20018 25566 20020 25618
rect 19964 25554 20020 25566
rect 20524 25620 20580 25630
rect 19852 25508 19908 25518
rect 19852 25414 19908 25452
rect 20076 25508 20132 25518
rect 20076 25414 20132 25452
rect 20524 25506 20580 25564
rect 20524 25454 20526 25506
rect 20578 25454 20580 25506
rect 20524 25442 20580 25454
rect 20748 25508 20804 26910
rect 26160 26684 26424 26694
rect 26216 26628 26264 26684
rect 26320 26628 26368 26684
rect 26160 26618 26424 26628
rect 34476 26684 34740 26694
rect 34532 26628 34580 26684
rect 34636 26628 34684 26684
rect 34476 26618 34740 26628
rect 25228 26404 25284 26414
rect 25228 26402 25508 26404
rect 25228 26350 25230 26402
rect 25282 26350 25508 26402
rect 25228 26348 25508 26350
rect 25228 26338 25284 26348
rect 22988 26290 23044 26302
rect 22988 26238 22990 26290
rect 23042 26238 23044 26290
rect 22652 26180 22708 26190
rect 22988 26180 23044 26238
rect 22652 26178 23044 26180
rect 22652 26126 22654 26178
rect 22706 26126 23044 26178
rect 22652 26124 23044 26126
rect 23212 26290 23268 26302
rect 23212 26238 23214 26290
rect 23266 26238 23268 26290
rect 22002 25900 22266 25910
rect 22058 25844 22106 25900
rect 22162 25844 22210 25900
rect 22002 25834 22266 25844
rect 21980 25620 22036 25630
rect 20748 25442 20804 25452
rect 21644 25508 21700 25518
rect 21644 25414 21700 25452
rect 20860 25396 20916 25406
rect 20188 24722 20244 24734
rect 20188 24670 20190 24722
rect 20242 24670 20244 24722
rect 20188 24612 20244 24670
rect 20860 24722 20916 25340
rect 21756 25396 21812 25406
rect 21756 25284 21812 25340
rect 21868 25284 21924 25294
rect 21756 25282 21924 25284
rect 21756 25230 21870 25282
rect 21922 25230 21924 25282
rect 21756 25228 21924 25230
rect 21868 25218 21924 25228
rect 20860 24670 20862 24722
rect 20914 24670 20916 24722
rect 20860 24658 20916 24670
rect 20244 24556 20356 24612
rect 20188 24546 20244 24556
rect 20300 24050 20356 24556
rect 20300 23998 20302 24050
rect 20354 23998 20356 24050
rect 20300 23986 20356 23998
rect 20412 24610 20468 24622
rect 20412 24558 20414 24610
rect 20466 24558 20468 24610
rect 19740 23090 19796 23100
rect 19852 23714 19908 23726
rect 19852 23662 19854 23714
rect 19906 23662 19908 23714
rect 19572 22876 19684 22932
rect 19516 22866 19572 22876
rect 19852 22484 19908 23662
rect 20300 23268 20356 23278
rect 20300 23174 20356 23212
rect 19404 22430 19406 22482
rect 19458 22430 19460 22482
rect 19404 22418 19460 22430
rect 19740 22428 19908 22484
rect 19628 22370 19684 22382
rect 19628 22318 19630 22370
rect 19682 22318 19684 22370
rect 19292 22036 19348 22046
rect 19292 21698 19348 21980
rect 19404 21812 19460 21822
rect 19628 21812 19684 22318
rect 19404 21810 19684 21812
rect 19404 21758 19406 21810
rect 19458 21758 19684 21810
rect 19404 21756 19684 21758
rect 19404 21746 19460 21756
rect 19292 21646 19294 21698
rect 19346 21646 19348 21698
rect 19292 21634 19348 21646
rect 19628 21700 19684 21756
rect 19628 21634 19684 21644
rect 19404 21364 19460 21374
rect 19180 21362 19460 21364
rect 19180 21310 19406 21362
rect 19458 21310 19460 21362
rect 19180 21308 19460 21310
rect 18956 20188 19236 20244
rect 18396 19842 18452 19852
rect 18508 20018 18564 20030
rect 18508 19966 18510 20018
rect 18562 19966 18564 20018
rect 18508 19684 18564 19966
rect 18508 19618 18564 19628
rect 18396 19348 18452 19358
rect 18396 19254 18452 19292
rect 18620 18452 18676 20188
rect 18844 20018 18900 20030
rect 18844 19966 18846 20018
rect 18898 19966 18900 20018
rect 18844 19796 18900 19966
rect 19068 20020 19124 20030
rect 19068 19926 19124 19964
rect 18844 18676 18900 19740
rect 18956 19906 19012 19918
rect 18956 19854 18958 19906
rect 19010 19854 19012 19906
rect 18956 19124 19012 19854
rect 19180 19572 19236 20188
rect 19404 20020 19460 21308
rect 19740 21364 19796 22428
rect 19964 22372 20020 22382
rect 19740 21298 19796 21308
rect 19852 22370 20020 22372
rect 19852 22318 19966 22370
rect 20018 22318 20020 22370
rect 19852 22316 20020 22318
rect 19516 20020 19572 20030
rect 19404 19964 19516 20020
rect 19516 19954 19572 19964
rect 19852 19572 19908 22316
rect 19964 22306 20020 22316
rect 20300 22372 20356 22382
rect 20300 22278 20356 22316
rect 19964 22148 20020 22158
rect 19964 21812 20020 22092
rect 19964 21718 20020 21756
rect 20300 21586 20356 21598
rect 20300 21534 20302 21586
rect 20354 21534 20356 21586
rect 20300 21364 20356 21534
rect 20300 21298 20356 21308
rect 20300 20020 20356 20030
rect 20300 19926 20356 19964
rect 19180 19516 19908 19572
rect 18956 19068 19572 19124
rect 18844 18610 18900 18620
rect 19516 18562 19572 19068
rect 19516 18510 19518 18562
rect 19570 18510 19572 18562
rect 19516 18498 19572 18510
rect 18732 18452 18788 18462
rect 18620 18396 18732 18452
rect 18732 18358 18788 18396
rect 18956 17556 19012 17566
rect 18956 17462 19012 17500
rect 18396 17444 18452 17454
rect 18396 16548 18452 17388
rect 19068 17444 19124 17454
rect 19068 17350 19124 17388
rect 18508 16772 18564 16782
rect 18508 16678 18564 16716
rect 19068 16660 19124 16670
rect 18396 16492 18788 16548
rect 18284 16380 18452 16436
rect 17948 16324 18004 16334
rect 17948 16230 18004 16268
rect 17724 16210 17892 16212
rect 17724 16158 17726 16210
rect 17778 16158 17892 16210
rect 17724 16156 17892 16158
rect 17724 16146 17780 16156
rect 17276 16046 17278 16098
rect 17330 16046 17332 16098
rect 17276 16034 17332 16046
rect 18284 15876 18340 15886
rect 17164 15820 17668 15876
rect 16828 15698 16884 15708
rect 16716 15374 16718 15426
rect 16770 15374 16772 15426
rect 16716 15362 16772 15374
rect 16828 15428 16884 15438
rect 16828 15426 17556 15428
rect 16828 15374 16830 15426
rect 16882 15374 17556 15426
rect 16828 15372 17556 15374
rect 16828 15362 16884 15372
rect 16604 14690 16660 14700
rect 17276 15092 17332 15102
rect 16380 14466 16436 14476
rect 16492 14644 16548 14654
rect 15820 14418 15876 14430
rect 15820 14366 15822 14418
rect 15874 14366 15876 14418
rect 15820 14196 15876 14366
rect 15932 14308 15988 14318
rect 15932 14306 16100 14308
rect 15932 14254 15934 14306
rect 15986 14254 16100 14306
rect 15932 14252 16100 14254
rect 15932 14242 15988 14252
rect 15820 14130 15876 14140
rect 15708 13916 15988 13972
rect 15932 13858 15988 13916
rect 15932 13806 15934 13858
rect 15986 13806 15988 13858
rect 15932 13794 15988 13806
rect 15260 13694 15262 13746
rect 15314 13694 15316 13746
rect 13580 12068 13636 12078
rect 13468 12066 13636 12068
rect 13468 12014 13582 12066
rect 13634 12014 13636 12066
rect 13468 12012 13636 12014
rect 13468 11394 13524 12012
rect 13580 12002 13636 12012
rect 13686 11788 13950 11798
rect 13742 11732 13790 11788
rect 13846 11732 13894 11788
rect 13686 11722 13950 11732
rect 14252 11508 14308 11518
rect 14252 11414 14308 11452
rect 13468 11342 13470 11394
rect 13522 11342 13524 11394
rect 13020 11284 13076 11294
rect 13020 10722 13076 11228
rect 13020 10670 13022 10722
rect 13074 10670 13076 10722
rect 13020 10658 13076 10670
rect 12348 10610 12404 10622
rect 12348 10558 12350 10610
rect 12402 10558 12404 10610
rect 12348 10388 12404 10558
rect 12348 10322 12404 10332
rect 13468 10388 13524 11342
rect 15148 10500 15204 10510
rect 15260 10500 15316 13694
rect 15820 13746 15876 13758
rect 15820 13694 15822 13746
rect 15874 13694 15876 13746
rect 15820 13636 15876 13694
rect 16044 13636 16100 14252
rect 16492 13860 16548 14588
rect 17052 14532 17108 14542
rect 17052 14438 17108 14476
rect 17276 14308 17332 15036
rect 17388 14532 17444 14542
rect 17388 14438 17444 14476
rect 17500 14530 17556 15372
rect 17500 14478 17502 14530
rect 17554 14478 17556 14530
rect 17500 14466 17556 14478
rect 16492 13794 16548 13804
rect 17164 14252 17276 14308
rect 15820 13580 16100 13636
rect 15372 13076 15428 13086
rect 15372 12982 15428 13020
rect 15820 11508 15876 13580
rect 16380 13076 16436 13086
rect 17052 13076 17108 13086
rect 17164 13076 17220 14252
rect 17276 14242 17332 14252
rect 17388 14196 17444 14206
rect 17388 13970 17444 14140
rect 17388 13918 17390 13970
rect 17442 13918 17444 13970
rect 17388 13906 17444 13918
rect 16436 13020 16548 13076
rect 16380 13010 16436 13020
rect 16380 11508 16436 11518
rect 15820 11506 16436 11508
rect 15820 11454 16382 11506
rect 16434 11454 16436 11506
rect 15820 11452 16436 11454
rect 16380 11442 16436 11452
rect 16492 10836 16548 13020
rect 17052 13074 17220 13076
rect 17052 13022 17054 13074
rect 17106 13022 17220 13074
rect 17052 13020 17220 13022
rect 17052 13010 17108 13020
rect 17612 12516 17668 15820
rect 17844 15708 18108 15718
rect 17900 15652 17948 15708
rect 18004 15652 18052 15708
rect 17844 15642 18108 15652
rect 17836 15316 17892 15326
rect 17836 14756 17892 15260
rect 17948 15316 18004 15326
rect 18172 15316 18228 15326
rect 17948 15314 18228 15316
rect 17948 15262 17950 15314
rect 18002 15262 18174 15314
rect 18226 15262 18228 15314
rect 17948 15260 18228 15262
rect 17948 15204 18004 15260
rect 18172 15250 18228 15260
rect 17948 15138 18004 15148
rect 17948 14756 18004 14766
rect 17836 14754 18004 14756
rect 17836 14702 17950 14754
rect 18002 14702 18004 14754
rect 17836 14700 18004 14702
rect 17948 14690 18004 14700
rect 18172 14756 18228 14766
rect 18284 14756 18340 15820
rect 18172 14754 18340 14756
rect 18172 14702 18174 14754
rect 18226 14702 18340 14754
rect 18172 14700 18340 14702
rect 18172 14690 18228 14700
rect 17388 12460 17668 12516
rect 17724 14418 17780 14430
rect 17724 14366 17726 14418
rect 17778 14366 17780 14418
rect 17724 13748 17780 14366
rect 18396 14196 18452 16380
rect 18620 16100 18676 16110
rect 18508 15988 18564 15998
rect 18508 15894 18564 15932
rect 18620 15986 18676 16044
rect 18620 15934 18622 15986
rect 18674 15934 18676 15986
rect 18620 15922 18676 15934
rect 17844 14140 18108 14150
rect 17900 14084 17948 14140
rect 18004 14084 18052 14140
rect 17844 14074 18108 14084
rect 18172 14140 18564 14196
rect 15148 10498 15316 10500
rect 15148 10446 15150 10498
rect 15202 10446 15316 10498
rect 15148 10444 15316 10446
rect 16268 10610 16324 10622
rect 16268 10558 16270 10610
rect 16322 10558 16324 10610
rect 15148 10434 15204 10444
rect 13468 10322 13524 10332
rect 14924 10388 14980 10398
rect 13686 10220 13950 10230
rect 13742 10164 13790 10220
rect 13846 10164 13894 10220
rect 13686 10154 13950 10164
rect 12236 9874 12292 9884
rect 12460 9938 12516 9950
rect 12460 9886 12462 9938
rect 12514 9886 12516 9938
rect 12012 9604 12068 9614
rect 12012 9510 12068 9548
rect 12348 9604 12404 9614
rect 11900 8990 11902 9042
rect 11954 8990 11956 9042
rect 11900 8820 11956 8990
rect 11900 8754 11956 8764
rect 12236 8930 12292 8942
rect 12236 8878 12238 8930
rect 12290 8878 12292 8930
rect 12236 8708 12292 8878
rect 12236 8642 12292 8652
rect 11788 8530 11844 8540
rect 12236 8372 12292 8382
rect 11676 8370 12292 8372
rect 11676 8318 12238 8370
rect 12290 8318 12292 8370
rect 11676 8316 12292 8318
rect 11676 8258 11732 8316
rect 12236 8306 12292 8316
rect 11676 8206 11678 8258
rect 11730 8206 11732 8258
rect 11676 8194 11732 8206
rect 12012 8148 12068 8158
rect 12236 8148 12292 8158
rect 12012 8146 12180 8148
rect 12012 8094 12014 8146
rect 12066 8094 12180 8146
rect 12012 8092 12180 8094
rect 12012 8082 12068 8092
rect 12124 7924 12180 8092
rect 12236 8054 12292 8092
rect 12348 7924 12404 9548
rect 12460 8484 12516 9886
rect 14476 9940 14532 9950
rect 14476 9846 14532 9884
rect 12908 9828 12964 9838
rect 14028 9828 14084 9838
rect 12908 9734 12964 9772
rect 13916 9826 14084 9828
rect 13916 9774 14030 9826
rect 14082 9774 14084 9826
rect 13916 9772 14084 9774
rect 13692 9714 13748 9726
rect 13692 9662 13694 9714
rect 13746 9662 13748 9714
rect 13580 9604 13636 9614
rect 13580 9510 13636 9548
rect 12572 9492 12628 9502
rect 13692 9492 13748 9662
rect 13804 9716 13860 9726
rect 13916 9716 13972 9772
rect 14028 9762 14084 9772
rect 13860 9660 13972 9716
rect 14140 9714 14196 9726
rect 14140 9662 14142 9714
rect 14194 9662 14196 9714
rect 13804 9650 13860 9660
rect 14028 9604 14084 9614
rect 14140 9604 14196 9662
rect 14084 9548 14196 9604
rect 14028 9538 14084 9548
rect 12628 9436 12740 9492
rect 12572 9426 12628 9436
rect 12572 8484 12628 8494
rect 12460 8428 12572 8484
rect 12572 8390 12628 8428
rect 12124 7868 12404 7924
rect 12684 8148 12740 9436
rect 13692 9426 13748 9436
rect 13244 9042 13300 9054
rect 13244 8990 13246 9042
rect 13298 8990 13300 9042
rect 13132 8930 13188 8942
rect 13132 8878 13134 8930
rect 13186 8878 13188 8930
rect 12908 8708 12964 8718
rect 12964 8652 13076 8708
rect 12908 8642 12964 8652
rect 12908 8484 12964 8494
rect 12796 8372 12852 8382
rect 12796 8278 12852 8316
rect 11564 7646 11566 7698
rect 11618 7646 11620 7698
rect 11564 7634 11620 7646
rect 12572 7700 12628 7710
rect 12684 7700 12740 8092
rect 12572 7698 12740 7700
rect 12572 7646 12574 7698
rect 12626 7646 12740 7698
rect 12572 7644 12740 7646
rect 12908 7698 12964 8428
rect 12908 7646 12910 7698
rect 12962 7646 12964 7698
rect 12572 7634 12628 7644
rect 12908 7634 12964 7646
rect 11452 7474 11508 7486
rect 11452 7422 11454 7474
rect 11506 7422 11508 7474
rect 11228 7364 11284 7374
rect 11228 6578 11284 7308
rect 11228 6526 11230 6578
rect 11282 6526 11284 6578
rect 11228 6514 11284 6526
rect 11228 5124 11284 5134
rect 11116 5122 11396 5124
rect 11116 5070 11230 5122
rect 11282 5070 11396 5122
rect 11116 5068 11396 5070
rect 9528 4732 9792 4742
rect 9584 4676 9632 4732
rect 9688 4676 9736 4732
rect 9528 4666 9792 4676
rect 9100 4498 9156 4508
rect 9772 4564 9828 4574
rect 8988 4398 8990 4450
rect 9042 4398 9044 4450
rect 8316 3666 8596 3668
rect 8316 3614 8318 3666
rect 8370 3614 8596 3666
rect 8316 3612 8596 3614
rect 8988 3668 9044 4398
rect 9548 4450 9604 4462
rect 9548 4398 9550 4450
rect 9602 4398 9604 4450
rect 9548 4116 9604 4398
rect 9772 4338 9828 4508
rect 9772 4286 9774 4338
rect 9826 4286 9828 4338
rect 9772 4274 9828 4286
rect 9884 4116 9940 5068
rect 10108 5058 10164 5068
rect 11228 5058 11284 5068
rect 11340 4564 11396 5068
rect 11340 4470 11396 4508
rect 11452 4452 11508 7422
rect 11676 7476 11732 7486
rect 11564 6468 11620 6478
rect 11564 4900 11620 6412
rect 11676 6244 11732 7420
rect 12012 7476 12068 7486
rect 12012 6916 12068 7420
rect 12796 7252 12852 7262
rect 12796 7158 12852 7196
rect 12012 6850 12068 6860
rect 12572 6916 12628 6926
rect 12460 6804 12516 6814
rect 11676 6188 12068 6244
rect 12012 6018 12068 6188
rect 12012 5966 12014 6018
rect 12066 5966 12068 6018
rect 12012 5954 12068 5966
rect 11900 5796 11956 5806
rect 11788 5124 11844 5134
rect 11788 5030 11844 5068
rect 11564 4834 11620 4844
rect 11900 4562 11956 5740
rect 12124 5348 12180 5358
rect 12124 5234 12180 5292
rect 12124 5182 12126 5234
rect 12178 5182 12180 5234
rect 12124 5170 12180 5182
rect 11900 4510 11902 4562
rect 11954 4510 11956 4562
rect 11900 4498 11956 4510
rect 12124 4564 12180 4574
rect 11452 4386 11508 4396
rect 11004 4338 11060 4350
rect 11004 4286 11006 4338
rect 11058 4286 11060 4338
rect 9548 4060 9940 4116
rect 10780 4228 10836 4238
rect 11004 4228 11060 4286
rect 12124 4338 12180 4508
rect 12124 4286 12126 4338
rect 12178 4286 12180 4338
rect 12124 4274 12180 4286
rect 10780 4226 11060 4228
rect 10780 4174 10782 4226
rect 10834 4174 11060 4226
rect 10780 4172 11060 4174
rect 8316 3602 8372 3612
rect 8988 3602 9044 3612
rect 10220 3668 10276 3678
rect 10220 3574 10276 3612
rect 6524 3502 6526 3554
rect 6578 3502 6580 3554
rect 6524 3490 6580 3502
rect 9548 3556 9604 3566
rect 9548 3462 9604 3500
rect 9528 3164 9792 3174
rect 9584 3108 9632 3164
rect 9688 3108 9736 3164
rect 9528 3098 9792 3108
rect 10780 800 10836 4172
rect 12460 3666 12516 6748
rect 12572 6578 12628 6860
rect 12908 6916 12964 6926
rect 12908 6690 12964 6860
rect 12908 6638 12910 6690
rect 12962 6638 12964 6690
rect 12908 6626 12964 6638
rect 12572 6526 12574 6578
rect 12626 6526 12628 6578
rect 12572 6514 12628 6526
rect 12684 6580 12740 6590
rect 12684 6018 12740 6524
rect 12684 5966 12686 6018
rect 12738 5966 12740 6018
rect 12684 5124 12740 5966
rect 13020 6244 13076 8652
rect 13132 8036 13188 8878
rect 13132 7970 13188 7980
rect 13244 7700 13300 8990
rect 14476 8930 14532 8942
rect 14476 8878 14478 8930
rect 14530 8878 14532 8930
rect 13356 8820 13412 8830
rect 13356 8370 13412 8764
rect 13686 8652 13950 8662
rect 13742 8596 13790 8652
rect 13846 8596 13894 8652
rect 13686 8586 13950 8596
rect 13356 8318 13358 8370
rect 13410 8318 13412 8370
rect 13356 8306 13412 8318
rect 13244 7634 13300 7644
rect 14140 8036 14196 8046
rect 14140 7588 14196 7980
rect 13132 7474 13188 7486
rect 13356 7476 13412 7486
rect 13132 7422 13134 7474
rect 13186 7422 13188 7474
rect 13132 6580 13188 7422
rect 13132 6514 13188 6524
rect 13244 7474 13412 7476
rect 13244 7422 13358 7474
rect 13410 7422 13412 7474
rect 13244 7420 13412 7422
rect 13020 6018 13076 6188
rect 13020 5966 13022 6018
rect 13074 5966 13076 6018
rect 13020 5954 13076 5966
rect 13244 6468 13300 7420
rect 13356 7410 13412 7420
rect 14140 7474 14196 7532
rect 14140 7422 14142 7474
rect 14194 7422 14196 7474
rect 14140 7410 14196 7422
rect 14364 7700 14420 7710
rect 14364 7586 14420 7644
rect 14364 7534 14366 7586
rect 14418 7534 14420 7586
rect 13916 7364 13972 7374
rect 13916 7270 13972 7308
rect 14252 7362 14308 7374
rect 14252 7310 14254 7362
rect 14306 7310 14308 7362
rect 13686 7084 13950 7094
rect 13742 7028 13790 7084
rect 13846 7028 13894 7084
rect 13686 7018 13950 7028
rect 14252 6804 14308 7310
rect 14140 6748 14308 6804
rect 14364 6804 14420 7534
rect 13356 6692 13412 6702
rect 13356 6598 13412 6636
rect 13804 6580 13860 6590
rect 13804 6486 13860 6524
rect 13244 5906 13300 6412
rect 13692 6132 13748 6142
rect 13692 6038 13748 6076
rect 14140 5908 14196 6748
rect 14364 6738 14420 6748
rect 14252 6578 14308 6590
rect 14252 6526 14254 6578
rect 14306 6526 14308 6578
rect 14252 6244 14308 6526
rect 14252 6178 14308 6188
rect 13244 5854 13246 5906
rect 13298 5854 13300 5906
rect 12684 5010 12740 5068
rect 12796 5124 12852 5134
rect 13244 5124 13300 5854
rect 14028 5906 14196 5908
rect 14028 5854 14142 5906
rect 14194 5854 14196 5906
rect 14028 5852 14196 5854
rect 13686 5516 13950 5526
rect 13742 5460 13790 5516
rect 13846 5460 13894 5516
rect 13686 5450 13950 5460
rect 13580 5348 13636 5358
rect 13580 5254 13636 5292
rect 12796 5122 13244 5124
rect 12796 5070 12798 5122
rect 12850 5070 13244 5122
rect 12796 5068 13244 5070
rect 12796 5058 12852 5068
rect 13244 5058 13300 5068
rect 13468 5122 13524 5134
rect 13468 5070 13470 5122
rect 13522 5070 13524 5122
rect 12684 4958 12686 5010
rect 12738 4958 12740 5010
rect 12684 4946 12740 4958
rect 13468 4564 13524 5070
rect 13916 5124 13972 5134
rect 13916 5030 13972 5068
rect 14028 5012 14084 5852
rect 14140 5842 14196 5852
rect 14364 5908 14420 5918
rect 14476 5908 14532 8878
rect 14924 8708 14980 10332
rect 15820 10386 15876 10398
rect 15820 10334 15822 10386
rect 15874 10334 15876 10386
rect 15036 9716 15092 9726
rect 15036 9044 15092 9660
rect 15036 8950 15092 8988
rect 15372 9042 15428 9054
rect 15372 8990 15374 9042
rect 15426 8990 15428 9042
rect 14924 8652 15092 8708
rect 14924 8148 14980 8158
rect 14924 8054 14980 8092
rect 14588 6692 14644 6702
rect 14588 6598 14644 6636
rect 15036 6692 15092 8652
rect 15372 8484 15428 8990
rect 15148 8260 15204 8270
rect 15148 8258 15316 8260
rect 15148 8206 15150 8258
rect 15202 8206 15316 8258
rect 15148 8204 15316 8206
rect 15148 8194 15204 8204
rect 15260 7474 15316 8204
rect 15372 7812 15428 8428
rect 15820 8148 15876 10334
rect 16268 10164 16324 10558
rect 16492 10610 16548 10780
rect 16716 11282 16772 11294
rect 16716 11230 16718 11282
rect 16770 11230 16772 11282
rect 16492 10558 16494 10610
rect 16546 10558 16548 10610
rect 16492 10546 16548 10558
rect 16604 10612 16660 10622
rect 16604 10518 16660 10556
rect 16268 10098 16324 10108
rect 16268 9156 16324 9166
rect 16268 8372 16324 9100
rect 16268 8306 16324 8316
rect 16492 8260 16548 8270
rect 15820 8146 16100 8148
rect 15820 8094 15822 8146
rect 15874 8094 16100 8146
rect 15820 8092 16100 8094
rect 15820 8082 15876 8092
rect 15372 7756 15876 7812
rect 15708 7588 15764 7598
rect 15260 7422 15262 7474
rect 15314 7422 15316 7474
rect 15260 7140 15316 7422
rect 15484 7476 15540 7486
rect 15484 7382 15540 7420
rect 15260 7074 15316 7084
rect 15260 6692 15316 6702
rect 15036 6690 15316 6692
rect 15036 6638 15262 6690
rect 15314 6638 15316 6690
rect 15036 6636 15316 6638
rect 14364 5906 14476 5908
rect 14364 5854 14366 5906
rect 14418 5854 14476 5906
rect 14364 5852 14476 5854
rect 14364 5842 14420 5852
rect 14476 5814 14532 5852
rect 14588 5796 14644 5806
rect 14588 5348 14644 5740
rect 14588 5282 14644 5292
rect 14028 4918 14084 4956
rect 13468 4498 13524 4508
rect 14140 4898 14196 4910
rect 14140 4846 14142 4898
rect 14194 4846 14196 4898
rect 13356 4452 13412 4462
rect 13356 4358 13412 4396
rect 12460 3614 12462 3666
rect 12514 3614 12516 3666
rect 12460 3602 12516 3614
rect 12572 4340 12628 4350
rect 12572 3556 12628 4284
rect 14140 4228 14196 4846
rect 15036 4340 15092 6636
rect 15260 6626 15316 6636
rect 15596 5908 15652 5918
rect 15484 5572 15540 5582
rect 15036 4274 15092 4284
rect 15260 5012 15316 5022
rect 14140 4162 14196 4172
rect 13686 3948 13950 3958
rect 13742 3892 13790 3948
rect 13846 3892 13894 3948
rect 13686 3882 13950 3892
rect 14924 3780 14980 3790
rect 14924 3686 14980 3724
rect 15260 3778 15316 4956
rect 15484 4226 15540 5516
rect 15484 4174 15486 4226
rect 15538 4174 15540 4226
rect 15484 4162 15540 4174
rect 15596 5124 15652 5852
rect 15708 5906 15764 7532
rect 15708 5854 15710 5906
rect 15762 5854 15764 5906
rect 15708 5842 15764 5854
rect 15820 5908 15876 7756
rect 16044 7588 16100 8092
rect 16044 7522 16100 7532
rect 16268 7474 16324 7486
rect 16268 7422 16270 7474
rect 16322 7422 16324 7474
rect 16156 7364 16212 7374
rect 16044 6578 16100 6590
rect 16044 6526 16046 6578
rect 16098 6526 16100 6578
rect 15932 5908 15988 5918
rect 15820 5906 15988 5908
rect 15820 5854 15934 5906
rect 15986 5854 15988 5906
rect 15820 5852 15988 5854
rect 15932 5842 15988 5852
rect 16044 5348 16100 6526
rect 16044 5282 16100 5292
rect 15932 5124 15988 5134
rect 15596 5122 15988 5124
rect 15596 5070 15934 5122
rect 15986 5070 15988 5122
rect 15596 5068 15988 5070
rect 15260 3726 15262 3778
rect 15314 3726 15316 3778
rect 15260 3714 15316 3726
rect 15484 3668 15540 3678
rect 15596 3668 15652 5068
rect 15932 5058 15988 5068
rect 16044 4900 16100 4910
rect 16044 4450 16100 4844
rect 16044 4398 16046 4450
rect 16098 4398 16100 4450
rect 16044 4386 16100 4398
rect 16156 4564 16212 7308
rect 16268 7140 16324 7422
rect 16492 7476 16548 8204
rect 16716 8258 16772 11230
rect 16828 11172 16884 11182
rect 16828 11170 16996 11172
rect 16828 11118 16830 11170
rect 16882 11118 16996 11170
rect 16828 11116 16996 11118
rect 16828 11106 16884 11116
rect 16716 8206 16718 8258
rect 16770 8206 16772 8258
rect 16716 7700 16772 8206
rect 16828 10610 16884 10622
rect 16828 10558 16830 10610
rect 16882 10558 16884 10610
rect 16828 8260 16884 10558
rect 16940 9828 16996 11116
rect 17276 11170 17332 11182
rect 17276 11118 17278 11170
rect 17330 11118 17332 11170
rect 17276 10164 17332 11118
rect 17388 11172 17444 12460
rect 17612 12292 17668 12302
rect 17388 11106 17444 11116
rect 17500 12178 17556 12190
rect 17500 12126 17502 12178
rect 17554 12126 17556 12178
rect 17388 10836 17444 10846
rect 17388 10742 17444 10780
rect 17500 10724 17556 12126
rect 17612 11618 17668 12236
rect 17612 11566 17614 11618
rect 17666 11566 17668 11618
rect 17612 11554 17668 11566
rect 17724 11508 17780 13692
rect 17948 13860 18004 13870
rect 17948 13074 18004 13804
rect 18172 13860 18228 14140
rect 18396 13972 18452 13982
rect 18396 13878 18452 13916
rect 18172 13746 18228 13804
rect 18172 13694 18174 13746
rect 18226 13694 18228 13746
rect 18172 13682 18228 13694
rect 17948 13022 17950 13074
rect 18002 13022 18004 13074
rect 17948 12964 18004 13022
rect 18508 12964 18564 14140
rect 18732 13972 18788 16492
rect 19068 16098 19124 16604
rect 19068 16046 19070 16098
rect 19122 16046 19124 16098
rect 19068 16034 19124 16046
rect 18844 15876 18900 15886
rect 18844 15782 18900 15820
rect 19628 15148 19684 19516
rect 19964 19348 20020 19358
rect 19964 15148 20020 19292
rect 20412 19348 20468 24558
rect 21980 24500 22036 25564
rect 22540 25506 22596 25518
rect 22540 25454 22542 25506
rect 22594 25454 22596 25506
rect 22540 25396 22596 25454
rect 22652 25508 22708 26124
rect 22652 25442 22708 25452
rect 22876 25732 22932 25742
rect 22540 25330 22596 25340
rect 22764 25394 22820 25406
rect 22764 25342 22766 25394
rect 22818 25342 22820 25394
rect 22764 24948 22820 25342
rect 22764 24882 22820 24892
rect 22876 24722 22932 25676
rect 23100 25620 23156 25630
rect 23100 25526 23156 25564
rect 22876 24670 22878 24722
rect 22930 24670 22932 24722
rect 22876 24658 22932 24670
rect 22988 25284 23044 25294
rect 22988 24722 23044 25228
rect 23212 24948 23268 26238
rect 23324 26290 23380 26302
rect 23324 26238 23326 26290
rect 23378 26238 23380 26290
rect 23324 25396 23380 26238
rect 25340 26178 25396 26190
rect 25340 26126 25342 26178
rect 25394 26126 25396 26178
rect 23772 26066 23828 26078
rect 23772 26014 23774 26066
rect 23826 26014 23828 26066
rect 23548 25396 23604 25406
rect 23324 25340 23548 25396
rect 23212 24882 23268 24892
rect 22988 24670 22990 24722
rect 23042 24670 23044 24722
rect 22988 24658 23044 24670
rect 23100 24724 23156 24734
rect 21980 24434 22036 24444
rect 22002 24332 22266 24342
rect 22058 24276 22106 24332
rect 22162 24276 22210 24332
rect 22002 24266 22266 24276
rect 22764 23268 22820 23278
rect 23100 23268 23156 24668
rect 21868 23266 22820 23268
rect 21868 23214 22766 23266
rect 22818 23214 22820 23266
rect 21868 23212 22820 23214
rect 21084 22372 21140 22382
rect 20524 22258 20580 22270
rect 20524 22206 20526 22258
rect 20578 22206 20580 22258
rect 20524 21588 20580 22206
rect 20636 22260 20692 22270
rect 20636 22166 20692 22204
rect 20748 22258 20804 22270
rect 20748 22206 20750 22258
rect 20802 22206 20804 22258
rect 20636 21700 20692 21710
rect 20636 21606 20692 21644
rect 20524 21522 20580 21532
rect 20748 21474 20804 22206
rect 21084 21810 21140 22316
rect 21308 22370 21364 22382
rect 21308 22318 21310 22370
rect 21362 22318 21364 22370
rect 21308 21924 21364 22318
rect 21308 21858 21364 21868
rect 21868 21812 21924 23212
rect 22764 23202 22820 23212
rect 22876 23266 23156 23268
rect 22876 23214 23102 23266
rect 23154 23214 23156 23266
rect 22876 23212 23156 23214
rect 22428 23044 22484 23054
rect 22876 23044 22932 23212
rect 23100 23202 23156 23212
rect 23212 24500 23268 24510
rect 22428 23042 22932 23044
rect 22428 22990 22430 23042
rect 22482 22990 22932 23042
rect 22428 22988 22932 22990
rect 22428 22978 22484 22988
rect 22002 22764 22266 22774
rect 22058 22708 22106 22764
rect 22162 22708 22210 22764
rect 22002 22698 22266 22708
rect 22092 22260 22148 22270
rect 22092 22166 22148 22204
rect 21084 21758 21086 21810
rect 21138 21758 21140 21810
rect 21084 21746 21140 21758
rect 21756 21756 21924 21812
rect 21980 21924 22036 21934
rect 20748 21422 20750 21474
rect 20802 21422 20804 21474
rect 20748 21410 20804 21422
rect 20860 21698 20916 21710
rect 20860 21646 20862 21698
rect 20914 21646 20916 21698
rect 20860 21476 20916 21646
rect 21756 21700 21812 21756
rect 21756 21606 21812 21644
rect 20748 20020 20804 20030
rect 20860 20020 20916 21420
rect 21308 21586 21364 21598
rect 21308 21534 21310 21586
rect 21362 21534 21364 21586
rect 21308 20692 21364 21534
rect 21868 21586 21924 21598
rect 21868 21534 21870 21586
rect 21922 21534 21924 21586
rect 21756 21476 21812 21486
rect 21868 21476 21924 21534
rect 21812 21420 21924 21476
rect 21756 21410 21812 21420
rect 21980 21364 22036 21868
rect 22876 21812 22932 21822
rect 22092 21700 22148 21710
rect 22092 21586 22148 21644
rect 22540 21700 22596 21710
rect 22540 21606 22596 21644
rect 22092 21534 22094 21586
rect 22146 21534 22148 21586
rect 22092 21522 22148 21534
rect 22428 21588 22484 21598
rect 22428 21494 22484 21532
rect 21308 20626 21364 20636
rect 21868 21308 22036 21364
rect 22652 21364 22708 21374
rect 21868 20804 21924 21308
rect 22002 21196 22266 21206
rect 22058 21140 22106 21196
rect 22162 21140 22210 21196
rect 22002 21130 22266 21140
rect 21868 20132 21924 20748
rect 21644 20076 21924 20132
rect 21644 20020 21700 20076
rect 20748 20018 20916 20020
rect 20748 19966 20750 20018
rect 20802 19966 20916 20018
rect 20748 19964 20916 19966
rect 21420 20018 21700 20020
rect 21420 19966 21646 20018
rect 21698 19966 21700 20018
rect 21420 19964 21700 19966
rect 20748 19954 20804 19964
rect 21196 19908 21252 19918
rect 21196 19814 21252 19852
rect 20412 19282 20468 19292
rect 20636 17444 20692 17454
rect 20636 16994 20692 17388
rect 20636 16942 20638 16994
rect 20690 16942 20692 16994
rect 20636 16930 20692 16942
rect 21420 16882 21476 19964
rect 21644 19954 21700 19964
rect 21868 19908 21924 19918
rect 21868 19458 21924 19852
rect 22316 19908 22372 19918
rect 22316 19906 22484 19908
rect 22316 19854 22318 19906
rect 22370 19854 22484 19906
rect 22316 19852 22484 19854
rect 22316 19842 22372 19852
rect 22002 19628 22266 19638
rect 22058 19572 22106 19628
rect 22162 19572 22210 19628
rect 22002 19562 22266 19572
rect 21868 19406 21870 19458
rect 21922 19406 21924 19458
rect 21868 19394 21924 19406
rect 22204 19460 22260 19470
rect 22428 19460 22484 19852
rect 22204 19458 22484 19460
rect 22204 19406 22206 19458
rect 22258 19406 22484 19458
rect 22204 19404 22484 19406
rect 22204 19394 22260 19404
rect 22092 19010 22148 19022
rect 22092 18958 22094 19010
rect 22146 18958 22148 19010
rect 21420 16830 21422 16882
rect 21474 16830 21476 16882
rect 21420 16818 21476 16830
rect 21644 18676 21700 18686
rect 21644 18338 21700 18620
rect 22092 18340 22148 18958
rect 22652 18676 22708 21308
rect 22652 18582 22708 18620
rect 22876 19346 22932 21756
rect 23100 20804 23156 20814
rect 23100 20710 23156 20748
rect 22876 19294 22878 19346
rect 22930 19294 22932 19346
rect 21644 18286 21646 18338
rect 21698 18286 21700 18338
rect 21644 16212 21700 18286
rect 21868 18284 22092 18340
rect 21644 16146 21700 16156
rect 21756 16770 21812 16782
rect 21756 16718 21758 16770
rect 21810 16718 21812 16770
rect 21756 16100 21812 16718
rect 21756 16034 21812 16044
rect 21420 15986 21476 15998
rect 21420 15934 21422 15986
rect 21474 15934 21476 15986
rect 21420 15148 21476 15934
rect 19404 15092 19684 15148
rect 19852 15092 20020 15148
rect 20636 15092 21476 15148
rect 21532 15874 21588 15886
rect 21532 15822 21534 15874
rect 21586 15822 21588 15874
rect 19404 14420 19460 15092
rect 19628 14530 19684 14542
rect 19628 14478 19630 14530
rect 19682 14478 19684 14530
rect 19404 14418 19572 14420
rect 19404 14366 19406 14418
rect 19458 14366 19572 14418
rect 19404 14364 19572 14366
rect 19404 14354 19460 14364
rect 18844 13972 18900 13982
rect 18732 13970 18900 13972
rect 18732 13918 18846 13970
rect 18898 13918 18900 13970
rect 18732 13916 18900 13918
rect 18844 13906 18900 13916
rect 19404 13860 19460 13870
rect 19404 13766 19460 13804
rect 18732 13748 18788 13758
rect 19068 13748 19124 13758
rect 18732 13654 18788 13692
rect 18844 13692 19068 13748
rect 19516 13748 19572 14364
rect 19628 13972 19684 14478
rect 19628 13906 19684 13916
rect 19516 13692 19684 13748
rect 18844 13300 18900 13692
rect 19068 13654 19124 13692
rect 18620 13244 18900 13300
rect 19516 13524 19572 13534
rect 18620 13186 18676 13244
rect 18620 13134 18622 13186
rect 18674 13134 18676 13186
rect 18620 13122 18676 13134
rect 18508 12908 18676 12964
rect 17948 12898 18004 12908
rect 18172 12740 18228 12750
rect 17844 12572 18108 12582
rect 17900 12516 17948 12572
rect 18004 12516 18052 12572
rect 17844 12506 18108 12516
rect 18172 12290 18228 12684
rect 18172 12238 18174 12290
rect 18226 12238 18228 12290
rect 18172 12226 18228 12238
rect 18396 12738 18452 12750
rect 18396 12686 18398 12738
rect 18450 12686 18452 12738
rect 18396 12292 18452 12686
rect 18508 12738 18564 12750
rect 18508 12686 18510 12738
rect 18562 12686 18564 12738
rect 18508 12404 18564 12686
rect 18508 12338 18564 12348
rect 18396 12226 18452 12236
rect 17836 11508 17892 11518
rect 17724 11506 17892 11508
rect 17724 11454 17838 11506
rect 17890 11454 17892 11506
rect 17724 11452 17892 11454
rect 17836 11442 17892 11452
rect 17500 10658 17556 10668
rect 17724 11172 17780 11182
rect 17724 10500 17780 11116
rect 18284 11170 18340 11182
rect 18284 11118 18286 11170
rect 18338 11118 18340 11170
rect 17844 11004 18108 11014
rect 17900 10948 17948 11004
rect 18004 10948 18052 11004
rect 17844 10938 18108 10948
rect 18284 10836 18340 11118
rect 18284 10770 18340 10780
rect 18396 10724 18452 10734
rect 18396 10612 18452 10668
rect 18508 10612 18564 10622
rect 18396 10610 18564 10612
rect 18396 10558 18510 10610
rect 18562 10558 18564 10610
rect 18396 10556 18564 10558
rect 18508 10546 18564 10556
rect 17836 10500 17892 10510
rect 17724 10444 17836 10500
rect 17836 10406 17892 10444
rect 17276 10098 17332 10108
rect 18620 9940 18676 12908
rect 18732 12068 18788 13244
rect 19068 13188 19124 13198
rect 18956 13132 19068 13188
rect 18844 12964 18900 12974
rect 18844 12870 18900 12908
rect 18732 12002 18788 12012
rect 18956 11620 19012 13132
rect 19068 13122 19124 13132
rect 19516 12962 19572 13468
rect 19516 12910 19518 12962
rect 19570 12910 19572 12962
rect 19516 12898 19572 12910
rect 19292 12850 19348 12862
rect 19292 12798 19294 12850
rect 19346 12798 19348 12850
rect 19292 12628 19348 12798
rect 19292 12562 19348 12572
rect 19404 12738 19460 12750
rect 19404 12686 19406 12738
rect 19458 12686 19460 12738
rect 19404 12292 19460 12686
rect 19404 12226 19460 12236
rect 18732 11564 19012 11620
rect 19404 12068 19460 12078
rect 18732 11506 18788 11564
rect 18732 11454 18734 11506
rect 18786 11454 18788 11506
rect 18732 11442 18788 11454
rect 18508 9884 18676 9940
rect 18732 10724 18788 10734
rect 16940 9762 16996 9772
rect 17836 9828 17892 9838
rect 17836 9734 17892 9772
rect 17276 9714 17332 9726
rect 17276 9662 17278 9714
rect 17330 9662 17332 9714
rect 17276 9156 17332 9662
rect 18284 9602 18340 9614
rect 18284 9550 18286 9602
rect 18338 9550 18340 9602
rect 17844 9436 18108 9446
rect 17900 9380 17948 9436
rect 18004 9380 18052 9436
rect 17844 9370 18108 9380
rect 17276 9062 17332 9100
rect 18060 9156 18116 9166
rect 18060 8260 18116 9100
rect 16828 8258 18116 8260
rect 16828 8206 18062 8258
rect 18114 8206 18116 8258
rect 16828 8204 18116 8206
rect 16716 7634 16772 7644
rect 17164 8034 17220 8046
rect 17164 7982 17166 8034
rect 17218 7982 17220 8034
rect 16492 7382 16548 7420
rect 16268 7074 16324 7084
rect 16604 7362 16660 7374
rect 16604 7310 16606 7362
rect 16658 7310 16660 7362
rect 16604 6020 16660 7310
rect 17164 6468 17220 7982
rect 17724 7476 17780 8204
rect 18060 8194 18116 8204
rect 18284 8370 18340 9550
rect 18284 8318 18286 8370
rect 18338 8318 18340 8370
rect 17844 7868 18108 7878
rect 17900 7812 17948 7868
rect 18004 7812 18052 7868
rect 17844 7802 18108 7812
rect 17836 7476 17892 7486
rect 17724 7474 18228 7476
rect 17724 7422 17838 7474
rect 17890 7422 18228 7474
rect 17724 7420 18228 7422
rect 17836 7410 17892 7420
rect 17388 7364 17444 7374
rect 17164 6402 17220 6412
rect 17276 7362 17444 7364
rect 17276 7310 17390 7362
rect 17442 7310 17444 7362
rect 17276 7308 17444 7310
rect 17276 6692 17332 7308
rect 17388 7298 17444 7308
rect 16156 4338 16212 4508
rect 16156 4286 16158 4338
rect 16210 4286 16212 4338
rect 16156 4274 16212 4286
rect 16380 6018 16660 6020
rect 16380 5966 16606 6018
rect 16658 5966 16660 6018
rect 16380 5964 16660 5966
rect 16380 4338 16436 5964
rect 16604 5954 16660 5964
rect 16380 4286 16382 4338
rect 16434 4286 16436 4338
rect 16380 4274 16436 4286
rect 16604 5684 16660 5694
rect 16604 4338 16660 5628
rect 17276 5684 17332 6636
rect 17388 7140 17444 7150
rect 17388 5906 17444 7084
rect 18172 6802 18228 7420
rect 18284 7474 18340 8318
rect 18508 8260 18564 9884
rect 18620 9716 18676 9726
rect 18620 9622 18676 9660
rect 18508 8194 18564 8204
rect 18732 8372 18788 10668
rect 18844 10612 18900 11564
rect 19404 11394 19460 12012
rect 19628 11956 19684 13692
rect 19852 13188 19908 15092
rect 20636 14642 20692 15092
rect 20636 14590 20638 14642
rect 20690 14590 20692 14642
rect 20636 14578 20692 14590
rect 21308 14644 21364 14654
rect 21532 14644 21588 15822
rect 21644 15876 21700 15886
rect 21868 15876 21924 18284
rect 22092 18274 22148 18284
rect 22876 18452 22932 19294
rect 22002 18060 22266 18070
rect 22058 18004 22106 18060
rect 22162 18004 22210 18060
rect 22002 17994 22266 18004
rect 22002 16492 22266 16502
rect 22058 16436 22106 16492
rect 22162 16436 22210 16492
rect 22002 16426 22266 16436
rect 22428 16100 22484 16110
rect 22428 16006 22484 16044
rect 21644 15874 21924 15876
rect 21644 15822 21646 15874
rect 21698 15822 21924 15874
rect 21644 15820 21924 15822
rect 22204 15986 22260 15998
rect 22204 15934 22206 15986
rect 22258 15934 22260 15986
rect 21644 15810 21700 15820
rect 21756 15204 21812 15820
rect 22204 15148 22260 15934
rect 22652 15988 22708 15998
rect 22652 15894 22708 15932
rect 22764 15986 22820 15998
rect 22764 15934 22766 15986
rect 22818 15934 22820 15986
rect 22764 15148 22820 15934
rect 22876 15428 22932 18396
rect 22988 18564 23044 18574
rect 23212 18564 23268 24444
rect 23548 21812 23604 25340
rect 23772 25284 23828 26014
rect 23772 25218 23828 25228
rect 24556 25620 24612 25630
rect 23660 24948 23716 24958
rect 23660 24854 23716 24892
rect 23884 24724 23940 24734
rect 23884 24630 23940 24668
rect 24332 24722 24388 24734
rect 24332 24670 24334 24722
rect 24386 24670 24388 24722
rect 24332 23268 24388 24670
rect 24444 24724 24500 24734
rect 24444 24630 24500 24668
rect 24556 24722 24612 25564
rect 25228 25620 25284 25630
rect 25340 25620 25396 26126
rect 25228 25618 25396 25620
rect 25228 25566 25230 25618
rect 25282 25566 25396 25618
rect 25228 25564 25396 25566
rect 25228 25554 25284 25564
rect 25452 25284 25508 26348
rect 25452 25218 25508 25228
rect 25564 26290 25620 26302
rect 25564 26238 25566 26290
rect 25618 26238 25620 26290
rect 25564 25396 25620 26238
rect 24556 24670 24558 24722
rect 24610 24670 24612 24722
rect 24556 24658 24612 24670
rect 25116 24722 25172 24734
rect 25564 24724 25620 25340
rect 25676 26290 25732 26302
rect 25676 26238 25678 26290
rect 25730 26238 25732 26290
rect 25676 24946 25732 26238
rect 30318 25900 30582 25910
rect 30374 25844 30422 25900
rect 30478 25844 30526 25900
rect 30318 25834 30582 25844
rect 26348 25620 26404 25630
rect 26012 25506 26068 25518
rect 26012 25454 26014 25506
rect 26066 25454 26068 25506
rect 25676 24894 25678 24946
rect 25730 24894 25732 24946
rect 25676 24882 25732 24894
rect 25788 25284 25844 25294
rect 25788 24946 25844 25228
rect 25788 24894 25790 24946
rect 25842 24894 25844 24946
rect 25788 24882 25844 24894
rect 25116 24670 25118 24722
rect 25170 24670 25172 24722
rect 25116 24500 25172 24670
rect 25116 24434 25172 24444
rect 25228 24722 25620 24724
rect 25228 24670 25566 24722
rect 25618 24670 25620 24722
rect 25228 24668 25620 24670
rect 25228 23380 25284 24668
rect 25564 24658 25620 24668
rect 25676 23828 25732 23838
rect 25228 23314 25284 23324
rect 25564 23772 25676 23828
rect 24332 23202 24388 23212
rect 24668 23266 24724 23278
rect 24668 23214 24670 23266
rect 24722 23214 24724 23266
rect 24444 23156 24500 23166
rect 24444 23062 24500 23100
rect 24668 22820 24724 23214
rect 24668 22754 24724 22764
rect 25116 23268 25172 23278
rect 25116 23156 25172 23212
rect 25228 23156 25284 23166
rect 25116 23154 25284 23156
rect 25116 23102 25230 23154
rect 25282 23102 25284 23154
rect 25116 23100 25284 23102
rect 24220 22482 24276 22494
rect 24220 22430 24222 22482
rect 24274 22430 24276 22482
rect 23660 21812 23716 21822
rect 23548 21810 23716 21812
rect 23548 21758 23662 21810
rect 23714 21758 23716 21810
rect 23548 21756 23716 21758
rect 23660 21746 23716 21756
rect 24220 21700 24276 22430
rect 25116 22148 25172 23100
rect 25228 23090 25284 23100
rect 25452 22932 25508 22942
rect 25228 22930 25508 22932
rect 25228 22878 25454 22930
rect 25506 22878 25508 22930
rect 25228 22876 25508 22878
rect 25228 22372 25284 22876
rect 25452 22866 25508 22876
rect 25340 22484 25396 22494
rect 25564 22484 25620 23772
rect 25676 23762 25732 23772
rect 25788 23716 25844 23726
rect 25788 23378 25844 23660
rect 25788 23326 25790 23378
rect 25842 23326 25844 23378
rect 25788 23314 25844 23326
rect 25900 23714 25956 23726
rect 25900 23662 25902 23714
rect 25954 23662 25956 23714
rect 25340 22482 25620 22484
rect 25340 22430 25342 22482
rect 25394 22430 25620 22482
rect 25340 22428 25620 22430
rect 25340 22418 25396 22428
rect 25228 22278 25284 22316
rect 25452 22148 25508 22158
rect 25116 22146 25508 22148
rect 25116 22094 25454 22146
rect 25506 22094 25508 22146
rect 25116 22092 25508 22094
rect 25452 22082 25508 22092
rect 25676 22148 25732 22158
rect 25900 22148 25956 23662
rect 25676 22146 25956 22148
rect 25676 22094 25678 22146
rect 25730 22094 25956 22146
rect 25676 22092 25956 22094
rect 24220 21606 24276 21644
rect 25676 21700 25732 22092
rect 24108 21586 24164 21598
rect 24108 21534 24110 21586
rect 24162 21534 24164 21586
rect 24108 21476 24164 21534
rect 24444 21588 24500 21598
rect 24444 21494 24500 21532
rect 23772 20692 23828 20702
rect 23772 20690 23940 20692
rect 23772 20638 23774 20690
rect 23826 20638 23940 20690
rect 23772 20636 23940 20638
rect 23772 20626 23828 20636
rect 22988 18562 23268 18564
rect 22988 18510 22990 18562
rect 23042 18510 23268 18562
rect 22988 18508 23268 18510
rect 23324 18676 23380 18686
rect 22988 18228 23044 18508
rect 23324 18340 23380 18620
rect 23660 18450 23716 18462
rect 23660 18398 23662 18450
rect 23714 18398 23716 18450
rect 23660 18340 23716 18398
rect 23884 18450 23940 20636
rect 23884 18398 23886 18450
rect 23938 18398 23940 18450
rect 23884 18386 23940 18398
rect 23996 20132 24052 20142
rect 23996 18450 24052 20076
rect 24108 19908 24164 21420
rect 24668 21476 24724 21486
rect 24668 21382 24724 21420
rect 24556 20804 24612 20814
rect 24444 19908 24500 19918
rect 24108 19906 24500 19908
rect 24108 19854 24446 19906
rect 24498 19854 24500 19906
rect 24108 19852 24500 19854
rect 24444 19842 24500 19852
rect 23996 18398 23998 18450
rect 24050 18398 24052 18450
rect 23996 18386 24052 18398
rect 23324 18284 23604 18340
rect 22988 18162 23044 18172
rect 23436 16212 23492 16222
rect 23436 16118 23492 16156
rect 22932 15372 23268 15428
rect 22876 15334 22932 15372
rect 21756 15138 21812 15148
rect 21308 14642 21476 14644
rect 21308 14590 21310 14642
rect 21362 14590 21476 14642
rect 21308 14588 21476 14590
rect 21308 14578 21364 14588
rect 20748 14530 20804 14542
rect 20748 14478 20750 14530
rect 20802 14478 20804 14530
rect 20076 14420 20132 14430
rect 19852 13122 19908 13132
rect 19964 14364 20076 14420
rect 19852 12850 19908 12862
rect 19852 12798 19854 12850
rect 19906 12798 19908 12850
rect 19740 12740 19796 12750
rect 19740 12646 19796 12684
rect 19852 12628 19908 12798
rect 19964 12628 20020 14364
rect 20076 14326 20132 14364
rect 20300 14306 20356 14318
rect 20300 14254 20302 14306
rect 20354 14254 20356 14306
rect 20188 13972 20244 13982
rect 20076 13748 20132 13758
rect 20076 13654 20132 13692
rect 20188 13188 20244 13916
rect 20300 13524 20356 14254
rect 20524 14308 20580 14318
rect 20524 14214 20580 14252
rect 20412 13860 20468 13870
rect 20748 13860 20804 14478
rect 20412 13858 20804 13860
rect 20412 13806 20414 13858
rect 20466 13806 20804 13858
rect 20412 13804 20804 13806
rect 20412 13794 20468 13804
rect 20300 13468 20468 13524
rect 20300 13188 20356 13198
rect 20188 13132 20300 13188
rect 20300 13094 20356 13132
rect 20076 13076 20132 13086
rect 20076 12982 20132 13020
rect 20412 12964 20468 13468
rect 20748 13076 20804 13804
rect 21420 14308 21476 14588
rect 21532 14578 21588 14588
rect 21868 15092 22260 15148
rect 22428 15092 22820 15148
rect 22876 15204 22932 15214
rect 21420 13636 21476 14252
rect 21420 13570 21476 13580
rect 21308 13524 21364 13534
rect 21756 13524 21812 13534
rect 21308 13430 21364 13468
rect 21532 13522 21812 13524
rect 21532 13470 21758 13522
rect 21810 13470 21812 13522
rect 21532 13468 21812 13470
rect 20748 13010 20804 13020
rect 20524 12964 20580 12974
rect 20412 12908 20524 12964
rect 20524 12870 20580 12908
rect 20860 12964 20916 12974
rect 20860 12962 21476 12964
rect 20860 12910 20862 12962
rect 20914 12910 21476 12962
rect 20860 12908 21476 12910
rect 20860 12898 20916 12908
rect 20972 12740 21028 12750
rect 19964 12572 20132 12628
rect 19628 11900 19796 11956
rect 19628 11732 19684 11742
rect 19404 11342 19406 11394
rect 19458 11342 19460 11394
rect 19404 11330 19460 11342
rect 19516 11506 19572 11518
rect 19516 11454 19518 11506
rect 19570 11454 19572 11506
rect 19516 10612 19572 11454
rect 19628 11394 19684 11676
rect 19628 11342 19630 11394
rect 19682 11342 19684 11394
rect 19628 11330 19684 11342
rect 19740 11172 19796 11900
rect 19852 11620 19908 12572
rect 19852 11554 19908 11564
rect 19964 12404 20020 12414
rect 19852 11396 19908 11406
rect 19964 11396 20020 12348
rect 20076 11732 20132 12572
rect 20636 12404 20692 12414
rect 20636 12310 20692 12348
rect 20972 12402 21028 12684
rect 20972 12350 20974 12402
rect 21026 12350 21028 12402
rect 20972 12338 21028 12350
rect 20300 12068 20356 12078
rect 20076 11666 20132 11676
rect 20188 12066 20580 12068
rect 20188 12014 20302 12066
rect 20354 12014 20580 12066
rect 20188 12012 20580 12014
rect 19852 11394 20020 11396
rect 19852 11342 19854 11394
rect 19906 11342 20020 11394
rect 19852 11340 20020 11342
rect 20076 11396 20132 11406
rect 20188 11396 20244 12012
rect 20300 12002 20356 12012
rect 20412 11620 20468 11630
rect 20412 11526 20468 11564
rect 20524 11506 20580 12012
rect 20524 11454 20526 11506
rect 20578 11454 20580 11506
rect 20524 11442 20580 11454
rect 21308 11732 21364 11742
rect 20076 11394 20244 11396
rect 20076 11342 20078 11394
rect 20130 11342 20244 11394
rect 20076 11340 20244 11342
rect 19852 11330 19908 11340
rect 20076 11330 20132 11340
rect 19740 11116 19908 11172
rect 19516 10556 19684 10612
rect 18844 9716 18900 10556
rect 18844 9492 18900 9660
rect 18956 10500 19012 10510
rect 18956 9716 19012 10444
rect 19180 10500 19236 10510
rect 19180 10498 19572 10500
rect 19180 10446 19182 10498
rect 19234 10446 19572 10498
rect 19180 10444 19572 10446
rect 19180 10434 19236 10444
rect 19292 10164 19348 10174
rect 19292 9828 19348 10108
rect 19516 9828 19572 10444
rect 19628 10050 19684 10556
rect 19628 9998 19630 10050
rect 19682 9998 19684 10050
rect 19628 9986 19684 9998
rect 19852 9940 19908 11116
rect 21308 10498 21364 11676
rect 21420 11506 21476 12908
rect 21420 11454 21422 11506
rect 21474 11454 21476 11506
rect 21420 11442 21476 11454
rect 21532 12066 21588 13468
rect 21756 13458 21812 13468
rect 21868 12964 21924 15092
rect 22002 14924 22266 14934
rect 22058 14868 22106 14924
rect 22162 14868 22210 14924
rect 22002 14858 22266 14868
rect 22204 14420 22260 14430
rect 22204 13746 22260 14364
rect 22204 13694 22206 13746
rect 22258 13694 22260 13746
rect 22204 13682 22260 13694
rect 21980 13524 22036 13562
rect 21980 13458 22036 13468
rect 22002 13356 22266 13366
rect 22058 13300 22106 13356
rect 22162 13300 22210 13356
rect 22002 13290 22266 13300
rect 22092 13188 22148 13198
rect 22092 13094 22148 13132
rect 22316 13076 22372 13086
rect 22428 13076 22484 15092
rect 22876 13970 22932 15148
rect 22876 13918 22878 13970
rect 22930 13918 22932 13970
rect 22876 13906 22932 13918
rect 22652 13746 22708 13758
rect 22652 13694 22654 13746
rect 22706 13694 22708 13746
rect 22652 13188 22708 13694
rect 22652 13122 22708 13132
rect 22988 13524 23044 13534
rect 22372 13020 22484 13076
rect 22988 13074 23044 13468
rect 22988 13022 22990 13074
rect 23042 13022 23044 13074
rect 22316 12982 22372 13020
rect 22988 13010 23044 13022
rect 21868 12870 21924 12908
rect 21644 12852 21700 12862
rect 22540 12852 22596 12862
rect 22876 12852 22932 12862
rect 21700 12796 21812 12852
rect 21644 12758 21700 12796
rect 21756 12292 21812 12796
rect 22540 12850 22820 12852
rect 22540 12798 22542 12850
rect 22594 12798 22820 12850
rect 22540 12796 22820 12798
rect 22540 12786 22596 12796
rect 22428 12740 22484 12750
rect 22428 12646 22484 12684
rect 21756 12236 21924 12292
rect 21532 12014 21534 12066
rect 21586 12014 21588 12066
rect 21532 11508 21588 12014
rect 21532 11394 21588 11452
rect 21532 11342 21534 11394
rect 21586 11342 21588 11394
rect 21532 11330 21588 11342
rect 21868 11394 21924 12236
rect 22002 11788 22266 11798
rect 22058 11732 22106 11788
rect 22162 11732 22210 11788
rect 22002 11722 22266 11732
rect 22764 11618 22820 12796
rect 22876 12758 22932 12796
rect 22764 11566 22766 11618
rect 22818 11566 22820 11618
rect 22764 11554 22820 11566
rect 22876 11508 22932 11518
rect 22876 11414 22932 11452
rect 21868 11342 21870 11394
rect 21922 11342 21924 11394
rect 21868 11330 21924 11342
rect 21308 10446 21310 10498
rect 21362 10446 21364 10498
rect 21308 10434 21364 10446
rect 21532 10836 21588 10846
rect 19740 9828 19796 9838
rect 19292 9826 19460 9828
rect 19292 9774 19294 9826
rect 19346 9774 19460 9826
rect 19292 9772 19460 9774
rect 19516 9826 19796 9828
rect 19516 9774 19742 9826
rect 19794 9774 19796 9826
rect 19516 9772 19796 9774
rect 19292 9762 19348 9772
rect 18956 9714 19236 9716
rect 18956 9662 18958 9714
rect 19010 9662 19236 9714
rect 18956 9660 19236 9662
rect 18956 9650 19012 9660
rect 18844 9436 19012 9492
rect 18844 9156 18900 9166
rect 18844 9062 18900 9100
rect 18956 9042 19012 9436
rect 18956 8990 18958 9042
rect 19010 8990 19012 9042
rect 18956 8978 19012 8990
rect 19180 9044 19236 9660
rect 19404 9156 19460 9772
rect 19740 9762 19796 9772
rect 19852 9714 19908 9884
rect 20412 9940 20468 9950
rect 20468 9884 20916 9940
rect 20412 9846 20468 9884
rect 19852 9662 19854 9714
rect 19906 9662 19908 9714
rect 19852 9650 19908 9662
rect 19740 9156 19796 9166
rect 19404 9154 19796 9156
rect 19404 9102 19742 9154
rect 19794 9102 19796 9154
rect 19404 9100 19796 9102
rect 19740 9090 19796 9100
rect 19292 9044 19348 9054
rect 19180 9042 19348 9044
rect 19180 8990 19294 9042
rect 19346 8990 19348 9042
rect 19180 8988 19348 8990
rect 19292 8978 19348 8988
rect 19068 8932 19124 8942
rect 19068 8482 19124 8876
rect 19068 8430 19070 8482
rect 19122 8430 19124 8482
rect 19068 8418 19124 8430
rect 18284 7422 18286 7474
rect 18338 7422 18340 7474
rect 18284 7410 18340 7422
rect 18732 7474 18788 8316
rect 19628 8372 19684 8382
rect 18732 7422 18734 7474
rect 18786 7422 18788 7474
rect 18732 7410 18788 7422
rect 18956 8258 19012 8270
rect 18956 8206 18958 8258
rect 19010 8206 19012 8258
rect 18172 6750 18174 6802
rect 18226 6750 18228 6802
rect 18172 6738 18228 6750
rect 17388 5854 17390 5906
rect 17442 5854 17444 5906
rect 17388 5842 17444 5854
rect 17724 6468 17780 6478
rect 17276 5618 17332 5628
rect 17724 5796 17780 6412
rect 18732 6468 18788 6478
rect 18732 6374 18788 6412
rect 17844 6300 18108 6310
rect 17900 6244 17948 6300
rect 18004 6244 18052 6300
rect 17844 6234 18108 6244
rect 16604 4286 16606 4338
rect 16658 4286 16660 4338
rect 16604 4274 16660 4286
rect 16940 5124 16996 5134
rect 15484 3666 15652 3668
rect 15484 3614 15486 3666
rect 15538 3614 15652 3666
rect 15484 3612 15652 3614
rect 16940 3666 16996 5068
rect 17724 5010 17780 5740
rect 17836 5906 17892 5918
rect 17836 5854 17838 5906
rect 17890 5854 17892 5906
rect 17836 5572 17892 5854
rect 18844 5906 18900 5918
rect 18844 5854 18846 5906
rect 18898 5854 18900 5906
rect 18396 5796 18452 5806
rect 18396 5794 18788 5796
rect 18396 5742 18398 5794
rect 18450 5742 18788 5794
rect 18396 5740 18788 5742
rect 18396 5730 18452 5740
rect 17836 5506 17892 5516
rect 18284 5236 18340 5246
rect 18172 5124 18228 5134
rect 18172 5030 18228 5068
rect 17724 4958 17726 5010
rect 17778 4958 17780 5010
rect 17724 4946 17780 4958
rect 17844 4732 18108 4742
rect 17900 4676 17948 4732
rect 18004 4676 18052 4732
rect 17844 4666 18108 4676
rect 17500 4564 17556 4574
rect 17500 4470 17556 4508
rect 16940 3614 16942 3666
rect 16994 3614 16996 3666
rect 15484 3602 15540 3612
rect 16940 3602 16996 3614
rect 12572 3490 12628 3500
rect 17844 3164 18108 3174
rect 17900 3108 17948 3164
rect 18004 3108 18052 3164
rect 17844 3098 18108 3108
rect 18284 2436 18340 5180
rect 18620 4564 18676 4574
rect 18620 4470 18676 4508
rect 18732 4452 18788 5740
rect 18844 5124 18900 5854
rect 18956 5572 19012 8206
rect 19068 8260 19124 8270
rect 19068 6578 19124 8204
rect 19068 6526 19070 6578
rect 19122 6526 19124 6578
rect 19068 6514 19124 6526
rect 19516 7362 19572 7374
rect 19516 7310 19518 7362
rect 19570 7310 19572 7362
rect 19516 6132 19572 7310
rect 19516 6066 19572 6076
rect 19292 5908 19348 5918
rect 19292 5814 19348 5852
rect 18956 5506 19012 5516
rect 19180 5236 19236 5246
rect 19180 5142 19236 5180
rect 18844 5058 18900 5068
rect 19180 4564 19236 4574
rect 18844 4452 18900 4462
rect 18732 4450 18900 4452
rect 18732 4398 18846 4450
rect 18898 4398 18900 4450
rect 18732 4396 18900 4398
rect 18844 4386 18900 4396
rect 19180 4338 19236 4508
rect 19180 4286 19182 4338
rect 19234 4286 19236 4338
rect 19180 4274 19236 4286
rect 19628 4338 19684 8316
rect 20860 6132 20916 9884
rect 21420 9716 21476 9726
rect 21420 9622 21476 9660
rect 20972 9044 21028 9054
rect 20972 8484 21028 8988
rect 20972 8418 21028 8428
rect 21532 8260 21588 10780
rect 22316 10612 22372 10622
rect 22316 10518 22372 10556
rect 23212 10612 23268 15372
rect 23436 14644 23492 14654
rect 23436 14550 23492 14588
rect 23548 13972 23604 18284
rect 23660 18274 23716 18284
rect 24556 16882 24612 20748
rect 25676 20244 25732 21644
rect 25900 21476 25956 21486
rect 25900 20916 25956 21420
rect 25900 20822 25956 20860
rect 25676 20178 25732 20188
rect 26012 20804 26068 25454
rect 26348 25506 26404 25564
rect 27356 25620 27412 25630
rect 27356 25618 28532 25620
rect 27356 25566 27358 25618
rect 27410 25566 28532 25618
rect 27356 25564 28532 25566
rect 27356 25554 27412 25564
rect 26348 25454 26350 25506
rect 26402 25454 26404 25506
rect 26348 25442 26404 25454
rect 26460 25396 26516 25406
rect 26684 25396 26740 25406
rect 27020 25396 27076 25406
rect 26516 25394 26740 25396
rect 26516 25342 26686 25394
rect 26738 25342 26740 25394
rect 26516 25340 26740 25342
rect 26460 25330 26516 25340
rect 26684 25330 26740 25340
rect 26796 25394 27076 25396
rect 26796 25342 27022 25394
rect 27074 25342 27076 25394
rect 26796 25340 27076 25342
rect 26160 25116 26424 25126
rect 26216 25060 26264 25116
rect 26320 25060 26368 25116
rect 26160 25050 26424 25060
rect 26348 24724 26404 24734
rect 26348 24612 26404 24668
rect 26124 24610 26404 24612
rect 26124 24558 26350 24610
rect 26402 24558 26404 24610
rect 26124 24556 26404 24558
rect 26124 24052 26180 24556
rect 26348 24546 26404 24556
rect 26796 24388 26852 25340
rect 27020 25330 27076 25340
rect 27244 25284 27300 25294
rect 27244 25190 27300 25228
rect 28476 24834 28532 25564
rect 34476 25116 34740 25126
rect 34532 25060 34580 25116
rect 34636 25060 34684 25116
rect 34476 25050 34740 25060
rect 28476 24782 28478 24834
rect 28530 24782 28532 24834
rect 28476 24770 28532 24782
rect 29260 24724 29316 24734
rect 29260 24722 29876 24724
rect 29260 24670 29262 24722
rect 29314 24670 29876 24722
rect 29260 24668 29876 24670
rect 29260 24658 29316 24668
rect 26124 23938 26180 23996
rect 26236 24332 26852 24388
rect 26236 24050 26292 24332
rect 26236 23998 26238 24050
rect 26290 23998 26292 24050
rect 26236 23986 26292 23998
rect 26684 24052 26740 24062
rect 26740 23996 26852 24052
rect 26684 23986 26740 23996
rect 26124 23886 26126 23938
rect 26178 23886 26180 23938
rect 26124 23874 26180 23886
rect 26684 23828 26740 23838
rect 26348 23716 26404 23754
rect 26684 23734 26740 23772
rect 26404 23660 26628 23716
rect 26348 23650 26404 23660
rect 26160 23548 26424 23558
rect 26216 23492 26264 23548
rect 26320 23492 26368 23548
rect 26160 23482 26424 23492
rect 26348 23380 26404 23390
rect 26124 23156 26180 23166
rect 26124 22370 26180 23100
rect 26124 22318 26126 22370
rect 26178 22318 26180 22370
rect 26124 22306 26180 22318
rect 26348 22372 26404 23324
rect 26460 23156 26516 23166
rect 26572 23156 26628 23660
rect 26460 23154 26628 23156
rect 26460 23102 26462 23154
rect 26514 23102 26628 23154
rect 26460 23100 26628 23102
rect 26684 23156 26740 23166
rect 26796 23156 26852 23996
rect 27020 24050 27076 24062
rect 27020 23998 27022 24050
rect 27074 23998 27076 24050
rect 26908 23716 26964 23726
rect 26908 23622 26964 23660
rect 27020 23268 27076 23998
rect 27020 23202 27076 23212
rect 29148 23268 29204 23278
rect 29148 23174 29204 23212
rect 26684 23154 26852 23156
rect 26684 23102 26686 23154
rect 26738 23102 26852 23154
rect 26684 23100 26852 23102
rect 26908 23156 26964 23166
rect 29820 23156 29876 24668
rect 30318 24332 30582 24342
rect 30374 24276 30422 24332
rect 30478 24276 30526 24332
rect 30318 24266 30582 24276
rect 34476 23548 34740 23558
rect 34532 23492 34580 23548
rect 34636 23492 34684 23548
rect 34476 23482 34740 23492
rect 26460 23090 26516 23100
rect 26684 23090 26740 23100
rect 26908 23044 26964 23100
rect 29484 23154 29876 23156
rect 29484 23102 29822 23154
rect 29874 23102 29876 23154
rect 29484 23100 29876 23102
rect 27020 23044 27076 23054
rect 26908 23042 27076 23044
rect 26908 22990 27022 23042
rect 27074 22990 27076 23042
rect 26908 22988 27076 22990
rect 27020 22978 27076 22988
rect 26348 22278 26404 22316
rect 26908 22820 26964 22830
rect 26908 22370 26964 22764
rect 26908 22318 26910 22370
rect 26962 22318 26964 22370
rect 26908 22306 26964 22318
rect 27020 22372 27076 22382
rect 27020 22258 27076 22316
rect 27020 22206 27022 22258
rect 27074 22206 27076 22258
rect 27020 22194 27076 22206
rect 27468 22258 27524 22270
rect 27468 22206 27470 22258
rect 27522 22206 27524 22258
rect 26572 22148 26628 22158
rect 26572 22054 26628 22092
rect 26684 22146 26740 22158
rect 26684 22094 26686 22146
rect 26738 22094 26740 22146
rect 26160 21980 26424 21990
rect 26216 21924 26264 21980
rect 26320 21924 26368 21980
rect 26160 21914 26424 21924
rect 26684 21812 26740 22094
rect 26236 21756 26740 21812
rect 26796 22148 26852 22158
rect 26124 21700 26180 21710
rect 26124 21606 26180 21644
rect 26236 21698 26292 21756
rect 26236 21646 26238 21698
rect 26290 21646 26292 21698
rect 26236 21634 26292 21646
rect 26124 21364 26180 21374
rect 26124 21270 26180 21308
rect 25676 20018 25732 20030
rect 25676 19966 25678 20018
rect 25730 19966 25732 20018
rect 25676 18340 25732 19966
rect 26012 19346 26068 20748
rect 26460 20802 26516 21756
rect 26572 21588 26628 21598
rect 26796 21588 26852 22092
rect 26628 21532 26852 21588
rect 27244 22146 27300 22158
rect 27244 22094 27246 22146
rect 27298 22094 27300 22146
rect 26572 21474 26628 21532
rect 26572 21422 26574 21474
rect 26626 21422 26628 21474
rect 26572 21410 26628 21422
rect 26460 20750 26462 20802
rect 26514 20750 26516 20802
rect 26460 20738 26516 20750
rect 26684 20916 26740 20926
rect 26684 20802 26740 20860
rect 26684 20750 26686 20802
rect 26738 20750 26740 20802
rect 26684 20738 26740 20750
rect 26236 20690 26292 20702
rect 26236 20638 26238 20690
rect 26290 20638 26292 20690
rect 26236 20580 26292 20638
rect 27244 20580 27300 22094
rect 27468 22148 27524 22206
rect 27468 22082 27524 22092
rect 27580 22148 27636 22158
rect 27580 22146 27860 22148
rect 27580 22094 27582 22146
rect 27634 22094 27860 22146
rect 27580 22092 27860 22094
rect 27580 22082 27636 22092
rect 27580 21364 27636 21374
rect 27580 20802 27636 21308
rect 27580 20750 27582 20802
rect 27634 20750 27636 20802
rect 27580 20738 27636 20750
rect 27804 20802 27860 22092
rect 29484 21586 29540 23100
rect 29820 23090 29876 23100
rect 30318 22764 30582 22774
rect 30374 22708 30422 22764
rect 30478 22708 30526 22764
rect 30318 22698 30582 22708
rect 34476 21980 34740 21990
rect 34532 21924 34580 21980
rect 34636 21924 34684 21980
rect 34476 21914 34740 21924
rect 29484 21534 29486 21586
rect 29538 21534 29540 21586
rect 28700 21474 28756 21486
rect 28700 21422 28702 21474
rect 28754 21422 28756 21474
rect 28028 20916 28084 20926
rect 28028 20822 28084 20860
rect 28700 20916 28756 21422
rect 28700 20850 28756 20860
rect 27804 20750 27806 20802
rect 27858 20750 27860 20802
rect 27804 20738 27860 20750
rect 28140 20690 28196 20702
rect 28140 20638 28142 20690
rect 28194 20638 28196 20690
rect 28140 20580 28196 20638
rect 26236 20524 26628 20580
rect 27244 20524 28196 20580
rect 26160 20412 26424 20422
rect 26216 20356 26264 20412
rect 26320 20356 26368 20412
rect 26160 20346 26424 20356
rect 26572 20132 26628 20524
rect 26572 20066 26628 20076
rect 26460 19908 26516 19918
rect 26460 19906 26628 19908
rect 26460 19854 26462 19906
rect 26514 19854 26628 19906
rect 26460 19852 26628 19854
rect 26460 19842 26516 19852
rect 26012 19294 26014 19346
rect 26066 19294 26068 19346
rect 26012 19282 26068 19294
rect 26160 18844 26424 18854
rect 26216 18788 26264 18844
rect 26320 18788 26368 18844
rect 26160 18778 26424 18788
rect 26236 18452 26292 18462
rect 26236 18358 26292 18396
rect 24556 16830 24558 16882
rect 24610 16830 24612 16882
rect 23884 16772 23940 16782
rect 23884 16770 24500 16772
rect 23884 16718 23886 16770
rect 23938 16718 24500 16770
rect 23884 16716 24500 16718
rect 23884 16706 23940 16716
rect 24444 16210 24500 16716
rect 24444 16158 24446 16210
rect 24498 16158 24500 16210
rect 24444 16146 24500 16158
rect 23660 16100 23716 16110
rect 23660 16006 23716 16044
rect 24332 15988 24388 15998
rect 24556 15988 24612 16830
rect 25340 16884 25396 16894
rect 25676 16884 25732 18284
rect 26572 18338 26628 19852
rect 28588 19906 28644 19918
rect 28588 19854 28590 19906
rect 28642 19854 28644 19906
rect 27244 19234 27300 19246
rect 27244 19182 27246 19234
rect 27298 19182 27300 19234
rect 26572 18286 26574 18338
rect 26626 18286 26628 18338
rect 26572 18274 26628 18286
rect 26684 18562 26740 18574
rect 26684 18510 26686 18562
rect 26738 18510 26740 18562
rect 26684 18004 26740 18510
rect 27244 18452 27300 19182
rect 27244 18358 27300 18396
rect 26684 17938 26740 17948
rect 26908 18226 26964 18238
rect 26908 18174 26910 18226
rect 26962 18174 26964 18226
rect 26236 17892 26292 17902
rect 26236 17798 26292 17836
rect 25340 16882 25732 16884
rect 25340 16830 25342 16882
rect 25394 16830 25732 16882
rect 25340 16828 25732 16830
rect 25900 17778 25956 17790
rect 25900 17726 25902 17778
rect 25954 17726 25956 17778
rect 25340 16818 25396 16828
rect 24332 15894 24388 15932
rect 24444 15932 24612 15988
rect 24668 16098 24724 16110
rect 24668 16046 24670 16098
rect 24722 16046 24724 16098
rect 23996 15874 24052 15886
rect 23996 15822 23998 15874
rect 24050 15822 24052 15874
rect 23996 14196 24052 15822
rect 24444 15148 24500 15932
rect 24220 15092 24500 15148
rect 24556 15204 24612 15214
rect 24668 15204 24724 16046
rect 25900 16100 25956 17726
rect 26012 17556 26068 17566
rect 26012 17462 26068 17500
rect 26572 17554 26628 17566
rect 26572 17502 26574 17554
rect 26626 17502 26628 17554
rect 26160 17276 26424 17286
rect 26216 17220 26264 17276
rect 26320 17220 26368 17276
rect 26160 17210 26424 17220
rect 25900 16034 25956 16044
rect 26012 16770 26068 16782
rect 26012 16718 26014 16770
rect 26066 16718 26068 16770
rect 24612 15148 24724 15204
rect 26012 15202 26068 16718
rect 26160 15708 26424 15718
rect 26216 15652 26264 15708
rect 26320 15652 26368 15708
rect 26160 15642 26424 15652
rect 26012 15150 26014 15202
rect 26066 15150 26068 15202
rect 24556 15138 24612 15148
rect 26012 15138 26068 15150
rect 26124 15426 26180 15438
rect 26124 15374 26126 15426
rect 26178 15374 26180 15426
rect 24220 14530 24276 15092
rect 24220 14478 24222 14530
rect 24274 14478 24276 14530
rect 24220 14466 24276 14478
rect 26124 14308 26180 15374
rect 26348 15428 26404 15438
rect 26572 15428 26628 17502
rect 26908 16212 26964 18174
rect 28476 18004 28532 18014
rect 27916 17892 27972 17902
rect 27916 17778 27972 17836
rect 28140 17892 28196 17902
rect 28196 17836 28308 17892
rect 28140 17826 28196 17836
rect 27916 17726 27918 17778
rect 27970 17726 27972 17778
rect 27916 17714 27972 17726
rect 27244 17666 27300 17678
rect 27244 17614 27246 17666
rect 27298 17614 27300 17666
rect 27244 16772 27300 17614
rect 27244 16706 27300 16716
rect 27468 17666 27524 17678
rect 28140 17668 28196 17678
rect 27468 17614 27470 17666
rect 27522 17614 27524 17666
rect 26908 16146 26964 16156
rect 27020 16100 27076 16110
rect 27020 16006 27076 16044
rect 27356 15876 27412 15886
rect 27356 15782 27412 15820
rect 27356 15540 27412 15550
rect 27468 15540 27524 17614
rect 28028 17666 28196 17668
rect 28028 17614 28142 17666
rect 28194 17614 28196 17666
rect 28028 17612 28196 17614
rect 27580 16772 27636 16782
rect 27580 15986 27636 16716
rect 28028 16436 28084 17612
rect 28140 17602 28196 17612
rect 28140 16772 28196 16782
rect 28140 16678 28196 16716
rect 27580 15934 27582 15986
rect 27634 15934 27636 15986
rect 27580 15922 27636 15934
rect 27916 16380 28084 16436
rect 27916 16098 27972 16380
rect 28028 16212 28084 16222
rect 28028 16118 28084 16156
rect 27916 16046 27918 16098
rect 27970 16046 27972 16098
rect 27692 15876 27748 15886
rect 27692 15874 27860 15876
rect 27692 15822 27694 15874
rect 27746 15822 27860 15874
rect 27692 15820 27860 15822
rect 27692 15810 27748 15820
rect 27692 15652 27748 15662
rect 27356 15538 27524 15540
rect 27356 15486 27358 15538
rect 27410 15486 27524 15538
rect 27356 15484 27524 15486
rect 27580 15540 27636 15550
rect 27356 15474 27412 15484
rect 27580 15446 27636 15484
rect 26348 15426 26628 15428
rect 26348 15374 26350 15426
rect 26402 15374 26628 15426
rect 26348 15372 26628 15374
rect 27692 15426 27748 15596
rect 27692 15374 27694 15426
rect 27746 15374 27748 15426
rect 26348 15362 26404 15372
rect 27692 15362 27748 15374
rect 27804 15316 27860 15820
rect 27916 15428 27972 16046
rect 28140 16100 28196 16110
rect 28252 16100 28308 17836
rect 28476 17890 28532 17948
rect 28476 17838 28478 17890
rect 28530 17838 28532 17890
rect 28476 16884 28532 17838
rect 28588 17892 28644 19854
rect 29260 18340 29316 18350
rect 29484 18340 29540 21534
rect 30318 21196 30582 21206
rect 30374 21140 30422 21196
rect 30478 21140 30526 21196
rect 30318 21130 30582 21140
rect 34476 20412 34740 20422
rect 34532 20356 34580 20412
rect 34636 20356 34684 20412
rect 34476 20346 34740 20356
rect 30318 19628 30582 19638
rect 30374 19572 30422 19628
rect 30478 19572 30526 19628
rect 30318 19562 30582 19572
rect 34476 18844 34740 18854
rect 34532 18788 34580 18844
rect 34636 18788 34684 18844
rect 34476 18778 34740 18788
rect 29316 18284 29652 18340
rect 29260 18246 29316 18284
rect 28588 17826 28644 17836
rect 29148 17778 29204 17790
rect 29148 17726 29150 17778
rect 29202 17726 29204 17778
rect 29148 17668 29204 17726
rect 29036 17612 29148 17668
rect 28924 17556 28980 17566
rect 28924 17106 28980 17500
rect 28924 17054 28926 17106
rect 28978 17054 28980 17106
rect 28924 17042 28980 17054
rect 29036 17108 29092 17612
rect 29148 17602 29204 17612
rect 29596 17668 29652 18284
rect 30318 18060 30582 18070
rect 30374 18004 30422 18060
rect 30478 18004 30526 18060
rect 30318 17994 30582 18004
rect 29036 17052 29428 17108
rect 29036 16994 29092 17052
rect 29036 16942 29038 16994
rect 29090 16942 29092 16994
rect 29036 16930 29092 16942
rect 28588 16884 28644 16894
rect 28476 16882 28980 16884
rect 28476 16830 28590 16882
rect 28642 16830 28980 16882
rect 28476 16828 28980 16830
rect 28140 16098 28308 16100
rect 28140 16046 28142 16098
rect 28194 16046 28308 16098
rect 28140 16044 28308 16046
rect 28364 16324 28420 16334
rect 28140 16034 28196 16044
rect 28364 15986 28420 16268
rect 28364 15934 28366 15986
rect 28418 15934 28420 15986
rect 28364 15922 28420 15934
rect 28476 15652 28532 16828
rect 28588 16818 28644 16828
rect 28924 16100 28980 16828
rect 29260 16882 29316 16894
rect 29260 16830 29262 16882
rect 29314 16830 29316 16882
rect 29260 16210 29316 16830
rect 29260 16158 29262 16210
rect 29314 16158 29316 16210
rect 29260 16146 29316 16158
rect 29148 16100 29204 16110
rect 28924 16098 29204 16100
rect 28924 16046 29150 16098
rect 29202 16046 29204 16098
rect 28924 16044 29204 16046
rect 29148 16034 29204 16044
rect 29372 16098 29428 17052
rect 29596 16882 29652 17612
rect 31388 17668 31444 17678
rect 31276 17556 31332 17566
rect 31276 17462 31332 17500
rect 29596 16830 29598 16882
rect 29650 16830 29652 16882
rect 29596 16818 29652 16830
rect 30380 16772 30436 16782
rect 30380 16678 30436 16716
rect 30318 16492 30582 16502
rect 30374 16436 30422 16492
rect 30478 16436 30526 16492
rect 30318 16426 30582 16436
rect 30716 16324 30772 16334
rect 29372 16046 29374 16098
rect 29426 16046 29428 16098
rect 28476 15586 28532 15596
rect 29372 15540 29428 16046
rect 29820 16100 29876 16110
rect 30044 16100 30100 16110
rect 29820 16098 30100 16100
rect 29820 16046 29822 16098
rect 29874 16046 30046 16098
rect 30098 16046 30100 16098
rect 29820 16044 30100 16046
rect 29820 16034 29876 16044
rect 29708 15540 29764 15550
rect 29372 15474 29428 15484
rect 29484 15484 29708 15540
rect 27916 15372 28308 15428
rect 27804 15260 27972 15316
rect 27916 15204 27972 15260
rect 27916 15148 28084 15204
rect 28028 14756 28084 15148
rect 27916 14700 28084 14756
rect 28252 14754 28308 15372
rect 28812 15426 28868 15438
rect 28812 15374 28814 15426
rect 28866 15374 28868 15426
rect 28252 14702 28254 14754
rect 28306 14702 28308 14754
rect 25788 14252 26180 14308
rect 27244 14530 27300 14542
rect 27244 14478 27246 14530
rect 27298 14478 27300 14530
rect 27244 14308 27300 14478
rect 23996 14140 24612 14196
rect 23660 13972 23716 13982
rect 24220 13972 24276 13982
rect 23548 13970 24276 13972
rect 23548 13918 23662 13970
rect 23714 13918 24222 13970
rect 24274 13918 24276 13970
rect 23548 13916 24276 13918
rect 23660 13906 23716 13916
rect 24220 13906 24276 13916
rect 23212 10546 23268 10556
rect 23548 13746 23604 13758
rect 23548 13694 23550 13746
rect 23602 13694 23604 13746
rect 22002 10220 22266 10230
rect 22058 10164 22106 10220
rect 22162 10164 22210 10220
rect 22002 10154 22266 10164
rect 21756 9938 21812 9950
rect 21756 9886 21758 9938
rect 21810 9886 21812 9938
rect 21420 8204 21588 8260
rect 21644 9716 21700 9726
rect 21420 6692 21476 8204
rect 21532 8036 21588 8046
rect 21644 8036 21700 9660
rect 21756 9154 21812 9886
rect 22092 9714 22148 9726
rect 22092 9662 22094 9714
rect 22146 9662 22148 9714
rect 21756 9102 21758 9154
rect 21810 9102 21812 9154
rect 21756 9090 21812 9102
rect 21868 9602 21924 9614
rect 21868 9550 21870 9602
rect 21922 9550 21924 9602
rect 21868 8932 21924 9550
rect 22092 9268 22148 9662
rect 22092 9202 22148 9212
rect 22876 9716 22932 9726
rect 21868 8484 21924 8876
rect 22876 9044 22932 9660
rect 22002 8652 22266 8662
rect 22058 8596 22106 8652
rect 22162 8596 22210 8652
rect 22002 8586 22266 8596
rect 21868 8428 22372 8484
rect 21532 8034 21700 8036
rect 21532 7982 21534 8034
rect 21586 7982 21700 8034
rect 21532 7980 21700 7982
rect 21756 8036 21812 8046
rect 21532 7970 21588 7980
rect 21644 7476 21700 7486
rect 21644 7362 21700 7420
rect 21644 7310 21646 7362
rect 21698 7310 21700 7362
rect 21644 7298 21700 7310
rect 21756 6916 21812 7980
rect 21980 7474 22036 8428
rect 22316 8372 22372 8428
rect 22316 8370 22708 8372
rect 22316 8318 22318 8370
rect 22370 8318 22708 8370
rect 22316 8316 22708 8318
rect 22316 8306 22372 8316
rect 21980 7422 21982 7474
rect 22034 7422 22036 7474
rect 21980 7410 22036 7422
rect 22092 8258 22148 8270
rect 22092 8206 22094 8258
rect 22146 8206 22148 8258
rect 22092 7476 22148 8206
rect 22428 7586 22484 7598
rect 22428 7534 22430 7586
rect 22482 7534 22484 7586
rect 22204 7476 22260 7486
rect 22092 7420 22204 7476
rect 22204 7382 22260 7420
rect 22002 7084 22266 7094
rect 22058 7028 22106 7084
rect 22162 7028 22210 7084
rect 22002 7018 22266 7028
rect 21420 6626 21476 6636
rect 21644 6860 21812 6916
rect 22092 6916 22148 6926
rect 21644 6244 21700 6860
rect 21868 6804 21924 6814
rect 21756 6692 21812 6702
rect 21756 6598 21812 6636
rect 21644 6188 21812 6244
rect 20972 6132 21028 6142
rect 21308 6132 21364 6142
rect 20860 6130 21252 6132
rect 20860 6078 20974 6130
rect 21026 6078 21252 6130
rect 20860 6076 21252 6078
rect 20860 4564 20916 6076
rect 20972 6066 21028 6076
rect 21196 5796 21252 6076
rect 21308 6018 21364 6076
rect 21308 5966 21310 6018
rect 21362 5966 21364 6018
rect 21308 5954 21364 5966
rect 21644 6020 21700 6030
rect 21644 5906 21700 5964
rect 21644 5854 21646 5906
rect 21698 5854 21700 5906
rect 21644 5842 21700 5854
rect 21756 5906 21812 6188
rect 21756 5854 21758 5906
rect 21810 5854 21812 5906
rect 21420 5796 21476 5806
rect 21196 5794 21476 5796
rect 21196 5742 21422 5794
rect 21474 5742 21476 5794
rect 21196 5740 21476 5742
rect 21420 5730 21476 5740
rect 21644 5236 21700 5246
rect 21644 5142 21700 5180
rect 20860 4498 20916 4508
rect 21532 5010 21588 5022
rect 21532 4958 21534 5010
rect 21586 4958 21588 5010
rect 19628 4286 19630 4338
rect 19682 4286 19684 4338
rect 19068 4226 19124 4238
rect 19068 4174 19070 4226
rect 19122 4174 19124 4226
rect 19068 3666 19124 4174
rect 19068 3614 19070 3666
rect 19122 3614 19124 3666
rect 19068 3602 19124 3614
rect 19628 3556 19684 4286
rect 20300 4228 20356 4238
rect 20300 4134 20356 4172
rect 21532 3666 21588 4958
rect 21756 4340 21812 5854
rect 21868 5348 21924 6748
rect 22092 6690 22148 6860
rect 22092 6638 22094 6690
rect 22146 6638 22148 6690
rect 22092 6626 22148 6638
rect 22316 6692 22372 6702
rect 22428 6692 22484 7534
rect 22316 6690 22484 6692
rect 22316 6638 22318 6690
rect 22370 6638 22484 6690
rect 22316 6636 22484 6638
rect 22316 6626 22372 6636
rect 22002 5516 22266 5526
rect 22058 5460 22106 5516
rect 22162 5460 22210 5516
rect 22002 5450 22266 5460
rect 21980 5348 22036 5358
rect 21868 5346 22036 5348
rect 21868 5294 21982 5346
rect 22034 5294 22036 5346
rect 21868 5292 22036 5294
rect 21980 5282 22036 5292
rect 21868 5122 21924 5134
rect 21868 5070 21870 5122
rect 21922 5070 21924 5122
rect 21868 4564 21924 5070
rect 21868 4498 21924 4508
rect 21756 4274 21812 4284
rect 22428 4226 22484 6636
rect 22540 7476 22596 7486
rect 22540 5794 22596 7420
rect 22652 5906 22708 8316
rect 22876 8260 22932 8988
rect 23548 8708 23604 13694
rect 23884 13748 23940 13758
rect 23884 13654 23940 13692
rect 24108 12962 24164 12974
rect 24108 12910 24110 12962
rect 24162 12910 24164 12962
rect 23660 12740 23716 12750
rect 23660 12290 23716 12684
rect 23660 12238 23662 12290
rect 23714 12238 23716 12290
rect 23660 12226 23716 12238
rect 24108 12180 24164 12910
rect 24332 12180 24388 12190
rect 24108 12178 24388 12180
rect 24108 12126 24334 12178
rect 24386 12126 24388 12178
rect 24108 12124 24388 12126
rect 24332 11396 24388 12124
rect 24444 11396 24500 11406
rect 24332 11394 24500 11396
rect 24332 11342 24446 11394
rect 24498 11342 24500 11394
rect 24332 11340 24500 11342
rect 24332 9716 24388 11340
rect 24444 11330 24500 11340
rect 24332 9650 24388 9660
rect 24556 9604 24612 14140
rect 25676 13972 25732 13982
rect 25676 13878 25732 13916
rect 25452 13860 25508 13870
rect 25452 13746 25508 13804
rect 25452 13694 25454 13746
rect 25506 13694 25508 13746
rect 25452 13682 25508 13694
rect 24780 13524 24836 13534
rect 24780 13074 24836 13468
rect 24780 13022 24782 13074
rect 24834 13022 24836 13074
rect 24780 13010 24836 13022
rect 25228 11284 25284 11294
rect 25228 11282 25732 11284
rect 25228 11230 25230 11282
rect 25282 11230 25732 11282
rect 25228 11228 25732 11230
rect 25228 11218 25284 11228
rect 25676 10498 25732 11228
rect 25788 10836 25844 14252
rect 27244 14242 27300 14252
rect 27468 14418 27524 14430
rect 27468 14366 27470 14418
rect 27522 14366 27524 14418
rect 26160 14140 26424 14150
rect 26216 14084 26264 14140
rect 26320 14084 26368 14140
rect 26160 14074 26424 14084
rect 26684 13972 26740 13982
rect 27020 13972 27076 13982
rect 26740 13916 26852 13972
rect 26684 13906 26740 13916
rect 26124 13748 26180 13758
rect 26124 13654 26180 13692
rect 26348 13746 26404 13758
rect 26348 13694 26350 13746
rect 26402 13694 26404 13746
rect 26348 13412 26404 13694
rect 26684 13746 26740 13758
rect 26684 13694 26686 13746
rect 26738 13694 26740 13746
rect 26460 13636 26516 13646
rect 26460 13542 26516 13580
rect 26348 13076 26404 13356
rect 26684 13300 26740 13694
rect 26348 13020 26628 13076
rect 26160 12572 26424 12582
rect 26216 12516 26264 12572
rect 26320 12516 26368 12572
rect 26160 12506 26424 12516
rect 26012 12178 26068 12190
rect 26012 12126 26014 12178
rect 26066 12126 26068 12178
rect 25788 10834 25956 10836
rect 25788 10782 25790 10834
rect 25842 10782 25956 10834
rect 25788 10780 25956 10782
rect 25788 10770 25844 10780
rect 25676 10446 25678 10498
rect 25730 10446 25732 10498
rect 25676 10434 25732 10446
rect 24668 9604 24724 9614
rect 24556 9548 24668 9604
rect 24668 9538 24724 9548
rect 25900 9380 25956 10780
rect 26012 10722 26068 12126
rect 26572 12178 26628 13020
rect 26572 12126 26574 12178
rect 26626 12126 26628 12178
rect 26572 12114 26628 12126
rect 26684 12066 26740 13244
rect 26684 12014 26686 12066
rect 26738 12014 26740 12066
rect 26684 12002 26740 12014
rect 26160 11004 26424 11014
rect 26216 10948 26264 11004
rect 26320 10948 26368 11004
rect 26160 10938 26424 10948
rect 26012 10670 26014 10722
rect 26066 10670 26068 10722
rect 26012 10658 26068 10670
rect 26160 9436 26424 9446
rect 26216 9380 26264 9436
rect 26320 9380 26368 9436
rect 25900 9324 26068 9380
rect 26160 9370 26424 9380
rect 24556 9268 24612 9278
rect 24332 9044 24388 9054
rect 23996 9042 24388 9044
rect 23996 8990 24334 9042
rect 24386 8990 24388 9042
rect 23996 8988 24388 8990
rect 23884 8932 23940 8942
rect 23884 8838 23940 8876
rect 23548 8652 23716 8708
rect 22988 8260 23044 8270
rect 22876 8258 23044 8260
rect 22876 8206 22990 8258
rect 23042 8206 23044 8258
rect 22876 8204 23044 8206
rect 22988 8194 23044 8204
rect 23324 8036 23380 8046
rect 23324 7586 23380 7980
rect 23324 7534 23326 7586
rect 23378 7534 23380 7586
rect 23324 7522 23380 7534
rect 23548 7586 23604 7598
rect 23548 7534 23550 7586
rect 23602 7534 23604 7586
rect 22652 5854 22654 5906
rect 22706 5854 22708 5906
rect 22652 5842 22708 5854
rect 22764 7474 22820 7486
rect 22764 7422 22766 7474
rect 22818 7422 22820 7474
rect 22540 5742 22542 5794
rect 22594 5742 22596 5794
rect 22540 5730 22596 5742
rect 22764 5122 22820 7422
rect 22988 7476 23044 7486
rect 22988 7382 23044 7420
rect 23436 7362 23492 7374
rect 23436 7310 23438 7362
rect 23490 7310 23492 7362
rect 23324 6916 23380 6926
rect 23212 6692 23268 6702
rect 23100 6690 23268 6692
rect 23100 6638 23214 6690
rect 23266 6638 23268 6690
rect 23100 6636 23268 6638
rect 22988 6580 23044 6590
rect 22988 6486 23044 6524
rect 22988 6020 23044 6030
rect 23100 6020 23156 6636
rect 23212 6626 23268 6636
rect 23044 5964 23156 6020
rect 22988 5926 23044 5964
rect 22764 5070 22766 5122
rect 22818 5070 22820 5122
rect 22764 5012 22820 5070
rect 22764 4946 22820 4956
rect 23324 5122 23380 6860
rect 23436 6804 23492 7310
rect 23548 6916 23604 7534
rect 23548 6850 23604 6860
rect 23660 6804 23716 8652
rect 23772 8372 23828 8382
rect 23996 8372 24052 8988
rect 24332 8978 24388 8988
rect 24556 9042 24612 9212
rect 26012 9268 26068 9324
rect 26236 9268 26292 9278
rect 26068 9266 26292 9268
rect 26068 9214 26238 9266
rect 26290 9214 26292 9266
rect 26068 9212 26292 9214
rect 26012 9174 26068 9212
rect 26236 9202 26292 9212
rect 26572 9268 26628 9278
rect 26796 9268 26852 13916
rect 27020 13746 27076 13916
rect 27020 13694 27022 13746
rect 27074 13694 27076 13746
rect 27020 13682 27076 13694
rect 27468 13748 27524 14366
rect 27244 13636 27300 13646
rect 27244 13542 27300 13580
rect 26908 13524 26964 13534
rect 26908 13430 26964 13468
rect 27356 13524 27412 13534
rect 27356 13430 27412 13468
rect 27468 13300 27524 13692
rect 27356 13244 27524 13300
rect 27580 14418 27636 14430
rect 27580 14366 27582 14418
rect 27634 14366 27636 14418
rect 27580 13412 27636 14366
rect 27804 14308 27860 14318
rect 27804 13636 27860 14252
rect 27804 13542 27860 13580
rect 26908 13076 26964 13086
rect 27356 13076 27412 13244
rect 26908 13074 27412 13076
rect 26908 13022 26910 13074
rect 26962 13022 27412 13074
rect 26908 13020 27412 13022
rect 26908 13010 26964 13020
rect 27356 12850 27412 13020
rect 27356 12798 27358 12850
rect 27410 12798 27412 12850
rect 27356 12786 27412 12798
rect 27468 12964 27524 12974
rect 27580 12964 27636 13356
rect 27468 12962 27636 12964
rect 27468 12910 27470 12962
rect 27522 12910 27636 12962
rect 27468 12908 27636 12910
rect 27132 12738 27188 12750
rect 27132 12686 27134 12738
rect 27186 12686 27188 12738
rect 27132 10836 27188 12686
rect 27356 11508 27412 11518
rect 27468 11508 27524 12908
rect 27356 11506 27524 11508
rect 27356 11454 27358 11506
rect 27410 11454 27524 11506
rect 27356 11452 27524 11454
rect 27356 11442 27412 11452
rect 27132 10770 27188 10780
rect 26908 10612 26964 10622
rect 27244 10612 27300 10622
rect 26964 10610 27300 10612
rect 26964 10558 27246 10610
rect 27298 10558 27300 10610
rect 26964 10556 27300 10558
rect 26908 9826 26964 10556
rect 27244 10546 27300 10556
rect 26908 9774 26910 9826
rect 26962 9774 26964 9826
rect 26908 9762 26964 9774
rect 27804 9604 27860 9614
rect 27132 9268 27188 9278
rect 26572 9266 27132 9268
rect 26572 9214 26574 9266
rect 26626 9214 27132 9266
rect 26572 9212 27132 9214
rect 26572 9202 26628 9212
rect 24556 8990 24558 9042
rect 24610 8990 24612 9042
rect 24556 8978 24612 8990
rect 27020 9042 27076 9054
rect 27020 8990 27022 9042
rect 27074 8990 27076 9042
rect 23772 8370 24052 8372
rect 23772 8318 23774 8370
rect 23826 8318 24052 8370
rect 23772 8316 24052 8318
rect 24220 8818 24276 8830
rect 24220 8766 24222 8818
rect 24274 8766 24276 8818
rect 23772 8306 23828 8316
rect 24108 7364 24164 7374
rect 23772 6804 23828 6814
rect 23660 6802 23828 6804
rect 23660 6750 23774 6802
rect 23826 6750 23828 6802
rect 23660 6748 23828 6750
rect 23436 6738 23492 6748
rect 23772 5908 23828 6748
rect 24108 6578 24164 7308
rect 24108 6526 24110 6578
rect 24162 6526 24164 6578
rect 24108 6514 24164 6526
rect 23772 5842 23828 5852
rect 24108 5684 24164 5694
rect 24220 5684 24276 8766
rect 27020 8428 27076 8990
rect 25900 8370 25956 8382
rect 25900 8318 25902 8370
rect 25954 8318 25956 8370
rect 25900 8260 25956 8318
rect 26908 8372 27076 8428
rect 26236 8260 26292 8270
rect 26908 8260 26964 8372
rect 25900 8258 26292 8260
rect 25900 8206 26238 8258
rect 26290 8206 26292 8258
rect 25900 8204 26292 8206
rect 25900 7586 25956 8204
rect 26236 8194 26292 8204
rect 26796 8204 26964 8260
rect 27132 8258 27188 9212
rect 27804 9154 27860 9548
rect 27804 9102 27806 9154
rect 27858 9102 27860 9154
rect 27804 9090 27860 9102
rect 27692 8260 27748 8270
rect 27132 8206 27134 8258
rect 27186 8206 27188 8258
rect 26572 8034 26628 8046
rect 26572 7982 26574 8034
rect 26626 7982 26628 8034
rect 26160 7868 26424 7878
rect 26216 7812 26264 7868
rect 26320 7812 26368 7868
rect 26160 7802 26424 7812
rect 25900 7534 25902 7586
rect 25954 7534 25956 7586
rect 25900 7522 25956 7534
rect 26012 7588 26068 7598
rect 26012 7474 26068 7532
rect 26012 7422 26014 7474
rect 26066 7422 26068 7474
rect 25676 7362 25732 7374
rect 25676 7310 25678 7362
rect 25730 7310 25732 7362
rect 25676 7252 25732 7310
rect 24780 6580 24836 6590
rect 24780 6486 24836 6524
rect 25676 6356 25732 7196
rect 25452 6300 25732 6356
rect 24444 6132 24500 6142
rect 24108 5682 24276 5684
rect 24108 5630 24110 5682
rect 24162 5630 24276 5682
rect 24108 5628 24276 5630
rect 24332 6076 24444 6132
rect 24332 5794 24388 6076
rect 24444 6066 24500 6076
rect 24444 5908 24500 5918
rect 24444 5814 24500 5852
rect 25340 5908 25396 5918
rect 25452 5908 25508 6300
rect 25676 6132 25732 6142
rect 25676 6018 25732 6076
rect 25676 5966 25678 6018
rect 25730 5966 25732 6018
rect 25676 5954 25732 5966
rect 25340 5906 25508 5908
rect 25340 5854 25342 5906
rect 25394 5854 25508 5906
rect 25340 5852 25508 5854
rect 25564 5908 25620 5918
rect 24332 5742 24334 5794
rect 24386 5742 24388 5794
rect 24108 5618 24164 5628
rect 24108 5460 24164 5470
rect 23324 5070 23326 5122
rect 23378 5070 23380 5122
rect 22428 4174 22430 4226
rect 22482 4174 22484 4226
rect 22002 3948 22266 3958
rect 22058 3892 22106 3948
rect 22162 3892 22210 3948
rect 22002 3882 22266 3892
rect 21532 3614 21534 3666
rect 21586 3614 21588 3666
rect 21532 3602 21588 3614
rect 19740 3556 19796 3566
rect 19628 3500 19740 3556
rect 19740 3462 19796 3500
rect 20748 3556 20804 3566
rect 20748 3462 20804 3500
rect 22428 3556 22484 4174
rect 22764 4564 22820 4574
rect 22764 3668 22820 4508
rect 23100 4340 23156 4350
rect 23100 4246 23156 4284
rect 23324 4226 23380 5070
rect 23772 5236 23828 5246
rect 23436 5012 23492 5022
rect 23492 4956 23604 5012
rect 23436 4946 23492 4956
rect 23324 4174 23326 4226
rect 23378 4174 23380 4226
rect 23324 4116 23380 4174
rect 23324 4050 23380 4060
rect 23548 3668 23604 4956
rect 23772 4338 23828 5180
rect 24108 5234 24164 5404
rect 24108 5182 24110 5234
rect 24162 5182 24164 5234
rect 24108 5170 24164 5182
rect 23772 4286 23774 4338
rect 23826 4286 23828 4338
rect 23772 4274 23828 4286
rect 24220 4340 24276 4350
rect 24332 4340 24388 5742
rect 25340 5460 25396 5852
rect 25564 5814 25620 5852
rect 25340 5394 25396 5404
rect 24220 4338 24388 4340
rect 24220 4286 24222 4338
rect 24274 4286 24388 4338
rect 24220 4284 24388 4286
rect 24220 4274 24276 4284
rect 23660 4228 23716 4238
rect 23660 4134 23716 4172
rect 25788 4228 25844 4238
rect 26012 4228 26068 7422
rect 26236 7476 26292 7486
rect 26236 7382 26292 7420
rect 26572 6804 26628 7982
rect 26796 7812 26852 8204
rect 27132 8194 27188 8206
rect 27468 8258 27748 8260
rect 27468 8206 27694 8258
rect 27746 8206 27748 8258
rect 27468 8204 27748 8206
rect 26908 8036 26964 8046
rect 26908 8034 27188 8036
rect 26908 7982 26910 8034
rect 26962 7982 27188 8034
rect 26908 7980 27188 7982
rect 26908 7970 26964 7980
rect 26796 7756 26964 7812
rect 26796 7476 26852 7486
rect 26684 7250 26740 7262
rect 26684 7198 26686 7250
rect 26738 7198 26740 7250
rect 26684 7140 26740 7198
rect 26684 7074 26740 7084
rect 26796 7028 26852 7420
rect 26796 6962 26852 6972
rect 26684 6804 26740 6814
rect 26572 6748 26684 6804
rect 26460 6692 26516 6702
rect 26460 6598 26516 6636
rect 26160 6300 26424 6310
rect 26216 6244 26264 6300
rect 26320 6244 26368 6300
rect 26160 6234 26424 6244
rect 26684 6020 26740 6748
rect 26908 6468 26964 7756
rect 27132 7476 27188 7980
rect 27468 7698 27524 8204
rect 27692 8194 27748 8204
rect 27468 7646 27470 7698
rect 27522 7646 27524 7698
rect 27468 7634 27524 7646
rect 27916 7586 27972 14700
rect 28028 14532 28084 14542
rect 28028 14438 28084 14476
rect 28252 13524 28308 14702
rect 28588 15314 28644 15326
rect 28588 15262 28590 15314
rect 28642 15262 28644 15314
rect 28588 15092 28644 15262
rect 28588 13860 28644 15036
rect 28812 14644 28868 15374
rect 29260 15428 29316 15466
rect 29260 15362 29316 15372
rect 29484 15426 29540 15484
rect 29708 15474 29764 15484
rect 29932 15538 29988 16044
rect 30044 16034 30100 16044
rect 30380 15874 30436 15886
rect 30380 15822 30382 15874
rect 30434 15822 30436 15874
rect 30380 15652 30436 15822
rect 30716 15652 30772 16268
rect 31388 16098 31444 17612
rect 31948 17668 32004 17678
rect 31948 17574 32004 17612
rect 34476 17276 34740 17286
rect 34532 17220 34580 17276
rect 34636 17220 34684 17276
rect 34476 17210 34740 17220
rect 33068 17108 33124 17118
rect 33068 17106 33460 17108
rect 33068 17054 33070 17106
rect 33122 17054 33460 17106
rect 33068 17052 33460 17054
rect 33068 17042 33124 17052
rect 33292 16882 33348 16894
rect 33292 16830 33294 16882
rect 33346 16830 33348 16882
rect 31948 16772 32004 16782
rect 31388 16046 31390 16098
rect 31442 16046 31444 16098
rect 31388 16034 31444 16046
rect 31724 16660 31780 16670
rect 30380 15596 30772 15652
rect 29932 15486 29934 15538
rect 29986 15486 29988 15538
rect 29932 15474 29988 15486
rect 29484 15374 29486 15426
rect 29538 15374 29540 15426
rect 29260 15202 29316 15214
rect 29260 15150 29262 15202
rect 29314 15150 29316 15202
rect 29260 14754 29316 15150
rect 29260 14702 29262 14754
rect 29314 14702 29316 14754
rect 29260 14690 29316 14702
rect 28812 14578 28868 14588
rect 29372 14532 29428 14542
rect 28588 13794 28644 13804
rect 29148 14530 29428 14532
rect 29148 14478 29374 14530
rect 29426 14478 29428 14530
rect 29148 14476 29428 14478
rect 28252 13458 28308 13468
rect 29148 13300 29204 14476
rect 29372 14466 29428 14476
rect 29484 14532 29540 15374
rect 30044 15428 30100 15438
rect 29820 15202 29876 15214
rect 29820 15150 29822 15202
rect 29874 15150 29876 15202
rect 29820 15092 29876 15150
rect 29820 15026 29876 15036
rect 29596 14644 29652 14654
rect 29596 14550 29652 14588
rect 29148 13186 29204 13244
rect 29148 13134 29150 13186
rect 29202 13134 29204 13186
rect 29148 13122 29204 13134
rect 29484 13186 29540 14476
rect 29708 14420 29764 14430
rect 29708 14418 29988 14420
rect 29708 14366 29710 14418
rect 29762 14366 29988 14418
rect 29708 14364 29988 14366
rect 29708 14354 29764 14364
rect 29932 13858 29988 14364
rect 29932 13806 29934 13858
rect 29986 13806 29988 13858
rect 29932 13794 29988 13806
rect 29484 13134 29486 13186
rect 29538 13134 29540 13186
rect 29484 13122 29540 13134
rect 29708 13636 29764 13646
rect 30044 13636 30100 15372
rect 30380 15426 30436 15438
rect 30380 15374 30382 15426
rect 30434 15374 30436 15426
rect 30380 15316 30436 15374
rect 30380 15250 30436 15260
rect 30492 15202 30548 15214
rect 30492 15150 30494 15202
rect 30546 15150 30548 15202
rect 30492 15092 30548 15150
rect 30604 15204 30660 15214
rect 30604 15110 30660 15148
rect 30492 15026 30548 15036
rect 30318 14924 30582 14934
rect 30374 14868 30422 14924
rect 30478 14868 30526 14924
rect 30318 14858 30582 14868
rect 30716 14756 30772 15596
rect 30940 15876 30996 15886
rect 30940 15426 30996 15820
rect 30940 15374 30942 15426
rect 30994 15374 30996 15426
rect 30940 15362 30996 15374
rect 31500 15428 31556 15438
rect 31052 15316 31108 15326
rect 31052 15222 31108 15260
rect 31388 15316 31444 15326
rect 31276 15092 31332 15102
rect 31164 15090 31332 15092
rect 31164 15038 31278 15090
rect 31330 15038 31332 15090
rect 31164 15036 31332 15038
rect 31164 14868 31220 15036
rect 31276 15026 31332 15036
rect 31388 14868 31444 15260
rect 31500 15314 31556 15372
rect 31724 15316 31780 16604
rect 31500 15262 31502 15314
rect 31554 15262 31556 15314
rect 31500 15250 31556 15262
rect 31612 15314 31780 15316
rect 31612 15262 31726 15314
rect 31778 15262 31780 15314
rect 31612 15260 31780 15262
rect 30604 14700 30772 14756
rect 30828 14812 31220 14868
rect 31276 14812 31444 14868
rect 30828 14754 30884 14812
rect 30828 14702 30830 14754
rect 30882 14702 30884 14754
rect 30604 14196 30660 14700
rect 30828 14690 30884 14702
rect 31164 14644 31220 14654
rect 31276 14644 31332 14812
rect 31164 14642 31332 14644
rect 31164 14590 31166 14642
rect 31218 14590 31332 14642
rect 31164 14588 31332 14590
rect 31164 14578 31220 14588
rect 30716 14420 30772 14430
rect 31276 14420 31332 14430
rect 30716 14418 31332 14420
rect 30716 14366 30718 14418
rect 30770 14366 31278 14418
rect 31330 14366 31332 14418
rect 30716 14364 31332 14366
rect 30716 14354 30772 14364
rect 30604 14140 30884 14196
rect 29764 13580 30100 13636
rect 30716 13746 30772 13758
rect 30716 13694 30718 13746
rect 30770 13694 30772 13746
rect 29708 13074 29764 13580
rect 30318 13356 30582 13366
rect 30374 13300 30422 13356
rect 30478 13300 30526 13356
rect 30318 13290 30582 13300
rect 29708 13022 29710 13074
rect 29762 13022 29764 13074
rect 29708 13010 29764 13022
rect 30716 12964 30772 13694
rect 30716 11844 30772 12908
rect 30318 11788 30582 11798
rect 30374 11732 30422 11788
rect 30478 11732 30526 11788
rect 30318 11722 30582 11732
rect 29148 11394 29204 11406
rect 29148 11342 29150 11394
rect 29202 11342 29204 11394
rect 29148 10388 29204 11342
rect 29484 11396 29540 11406
rect 29484 11394 29876 11396
rect 29484 11342 29486 11394
rect 29538 11342 29876 11394
rect 29484 11340 29876 11342
rect 29484 11330 29540 11340
rect 29596 11170 29652 11182
rect 29596 11118 29598 11170
rect 29650 11118 29652 11170
rect 29596 10388 29652 11118
rect 29148 10322 29204 10332
rect 29260 10332 29652 10388
rect 29708 11170 29764 11182
rect 29708 11118 29710 11170
rect 29762 11118 29764 11170
rect 29260 9826 29316 10332
rect 29596 10052 29652 10062
rect 29260 9774 29262 9826
rect 29314 9774 29316 9826
rect 29260 9762 29316 9774
rect 29484 9828 29540 9838
rect 29596 9828 29652 9996
rect 29484 9826 29652 9828
rect 29484 9774 29486 9826
rect 29538 9774 29652 9826
rect 29484 9772 29652 9774
rect 29484 9762 29540 9772
rect 28252 9602 28308 9614
rect 28252 9550 28254 9602
rect 28306 9550 28308 9602
rect 28252 9268 28308 9550
rect 28252 9202 28308 9212
rect 28588 9602 28644 9614
rect 28588 9550 28590 9602
rect 28642 9550 28644 9602
rect 28028 8932 28084 8942
rect 28028 8258 28084 8876
rect 28028 8206 28030 8258
rect 28082 8206 28084 8258
rect 28028 8194 28084 8206
rect 28140 8370 28196 8382
rect 28140 8318 28142 8370
rect 28194 8318 28196 8370
rect 28140 7698 28196 8318
rect 28140 7646 28142 7698
rect 28194 7646 28196 7698
rect 28140 7634 28196 7646
rect 28252 8034 28308 8046
rect 28252 7982 28254 8034
rect 28306 7982 28308 8034
rect 27916 7534 27918 7586
rect 27970 7534 27972 7586
rect 27916 7522 27972 7534
rect 28252 7588 28308 7982
rect 28252 7522 28308 7532
rect 27580 7476 27636 7486
rect 27132 7420 27524 7476
rect 27132 7252 27188 7262
rect 27132 7158 27188 7196
rect 27356 7250 27412 7262
rect 27356 7198 27358 7250
rect 27410 7198 27412 7250
rect 27020 7140 27076 7150
rect 27020 6916 27076 7084
rect 27132 6916 27188 6926
rect 27020 6914 27188 6916
rect 27020 6862 27134 6914
rect 27186 6862 27188 6914
rect 27020 6860 27188 6862
rect 27132 6850 27188 6860
rect 27356 6804 27412 7198
rect 27356 6738 27412 6748
rect 27244 6690 27300 6702
rect 27244 6638 27246 6690
rect 27298 6638 27300 6690
rect 26908 6412 27188 6468
rect 26684 5926 26740 5964
rect 26908 6020 26964 6030
rect 26964 5964 27076 6020
rect 26908 5954 26964 5964
rect 26124 5908 26180 5918
rect 26124 5814 26180 5852
rect 26460 5906 26516 5918
rect 26460 5854 26462 5906
rect 26514 5854 26516 5906
rect 26236 5684 26292 5694
rect 26236 5234 26292 5628
rect 26460 5460 26516 5854
rect 27020 5906 27076 5964
rect 27020 5854 27022 5906
rect 27074 5854 27076 5906
rect 27020 5842 27076 5854
rect 26908 5796 26964 5806
rect 26908 5702 26964 5740
rect 26460 5394 26516 5404
rect 26236 5182 26238 5234
rect 26290 5182 26292 5234
rect 26236 5170 26292 5182
rect 27020 5124 27076 5134
rect 27132 5124 27188 6412
rect 27244 5348 27300 6638
rect 27468 6690 27524 7420
rect 27580 7382 27636 7420
rect 28028 7364 28084 7374
rect 28028 7270 28084 7308
rect 27468 6638 27470 6690
rect 27522 6638 27524 6690
rect 27356 5684 27412 5694
rect 27356 5590 27412 5628
rect 27468 5682 27524 6638
rect 28140 7028 28196 7038
rect 28140 6690 28196 6972
rect 28588 6916 28644 9550
rect 29484 9604 29540 9614
rect 29484 9510 29540 9548
rect 29596 9044 29652 9772
rect 29596 8978 29652 8988
rect 29708 9826 29764 11118
rect 29820 11172 29876 11340
rect 30268 11394 30324 11406
rect 30268 11342 30270 11394
rect 30322 11342 30324 11394
rect 30044 11172 30100 11182
rect 29820 11170 30100 11172
rect 29820 11118 30046 11170
rect 30098 11118 30100 11170
rect 29820 11116 30100 11118
rect 30044 10164 30100 11116
rect 30268 10388 30324 11342
rect 30044 10098 30100 10108
rect 30156 10332 30324 10388
rect 30716 10722 30772 11788
rect 30716 10670 30718 10722
rect 30770 10670 30772 10722
rect 30044 9940 30100 9950
rect 29708 9774 29710 9826
rect 29762 9774 29764 9826
rect 29708 8260 29764 9774
rect 29820 9884 30044 9940
rect 29820 8428 29876 9884
rect 30044 9846 30100 9884
rect 30156 9940 30212 10332
rect 30318 10220 30582 10230
rect 30374 10164 30422 10220
rect 30478 10164 30526 10220
rect 30318 10154 30582 10164
rect 30716 10052 30772 10670
rect 30828 10388 30884 14140
rect 31276 13970 31332 14364
rect 31612 14418 31668 15260
rect 31724 15250 31780 15260
rect 31948 15092 32004 16716
rect 32508 16770 32564 16782
rect 32508 16718 32510 16770
rect 32562 16718 32564 16770
rect 32508 16660 32564 16718
rect 32508 16594 32564 16604
rect 33180 16770 33236 16782
rect 33180 16718 33182 16770
rect 33234 16718 33236 16770
rect 32060 15986 32116 15998
rect 33180 15988 33236 16718
rect 33292 16660 33348 16830
rect 33292 16594 33348 16604
rect 32060 15934 32062 15986
rect 32114 15934 32116 15986
rect 32060 15876 32116 15934
rect 32396 15932 33236 15988
rect 32060 15820 32340 15876
rect 32060 15540 32116 15550
rect 32060 15316 32116 15484
rect 32060 15314 32228 15316
rect 32060 15262 32062 15314
rect 32114 15262 32228 15314
rect 32060 15260 32228 15262
rect 32060 15250 32116 15260
rect 32060 15092 32116 15102
rect 31948 15090 32116 15092
rect 31948 15038 32062 15090
rect 32114 15038 32116 15090
rect 31948 15036 32116 15038
rect 32060 15026 32116 15036
rect 32172 14754 32228 15260
rect 32172 14702 32174 14754
rect 32226 14702 32228 14754
rect 32172 14690 32228 14702
rect 31612 14366 31614 14418
rect 31666 14366 31668 14418
rect 31612 14354 31668 14366
rect 31836 14530 31892 14542
rect 31836 14478 31838 14530
rect 31890 14478 31892 14530
rect 31276 13918 31278 13970
rect 31330 13918 31332 13970
rect 31276 13860 31332 13918
rect 31276 13804 31780 13860
rect 30828 10322 30884 10332
rect 31052 13522 31108 13534
rect 31052 13470 31054 13522
rect 31106 13470 31108 13522
rect 31052 11172 31108 13470
rect 31276 13074 31332 13804
rect 31724 13746 31780 13804
rect 31724 13694 31726 13746
rect 31778 13694 31780 13746
rect 31724 13682 31780 13694
rect 31500 13636 31556 13646
rect 31388 13524 31444 13534
rect 31388 13430 31444 13468
rect 31276 13022 31278 13074
rect 31330 13022 31332 13074
rect 31276 13010 31332 13022
rect 31500 12178 31556 13580
rect 31836 13524 31892 14478
rect 32284 14308 32340 15820
rect 32396 15426 32452 15932
rect 33404 15652 33460 17052
rect 33628 16882 33684 16894
rect 33628 16830 33630 16882
rect 33682 16830 33684 16882
rect 33628 16324 33684 16830
rect 33628 16258 33684 16268
rect 33180 15596 33460 15652
rect 34188 16210 34244 16222
rect 34188 16158 34190 16210
rect 34242 16158 34244 16210
rect 33068 15540 33124 15550
rect 33180 15540 33236 15596
rect 32396 15374 32398 15426
rect 32450 15374 32452 15426
rect 32396 15362 32452 15374
rect 32620 15538 33236 15540
rect 32620 15486 33070 15538
rect 33122 15486 33236 15538
rect 32620 15484 33236 15486
rect 32508 15204 32564 15214
rect 32396 15092 32452 15102
rect 32396 14530 32452 15036
rect 32396 14478 32398 14530
rect 32450 14478 32452 14530
rect 32396 14466 32452 14478
rect 32508 14532 32564 15148
rect 32620 14754 32676 15484
rect 33068 15474 33124 15484
rect 33628 15316 33684 15326
rect 33628 15222 33684 15260
rect 34188 15316 34244 16158
rect 34476 15708 34740 15718
rect 34532 15652 34580 15708
rect 34636 15652 34684 15708
rect 34476 15642 34740 15652
rect 34188 15250 34244 15260
rect 33404 15204 33460 15214
rect 32620 14702 32622 14754
rect 32674 14702 32676 14754
rect 32620 14690 32676 14702
rect 33180 15148 33404 15204
rect 32844 14532 32900 14542
rect 32508 14476 32676 14532
rect 32508 14308 32564 14318
rect 32284 14306 32564 14308
rect 32284 14254 32510 14306
rect 32562 14254 32564 14306
rect 32284 14252 32564 14254
rect 32508 14242 32564 14252
rect 32620 14084 32676 14476
rect 32284 14028 32676 14084
rect 32284 13970 32340 14028
rect 32284 13918 32286 13970
rect 32338 13918 32340 13970
rect 32284 13906 32340 13918
rect 32844 13636 32900 14476
rect 33180 13746 33236 15148
rect 33404 15110 33460 15148
rect 34476 14140 34740 14150
rect 34532 14084 34580 14140
rect 34636 14084 34684 14140
rect 34476 14074 34740 14084
rect 33628 13748 33684 13758
rect 33180 13694 33182 13746
rect 33234 13694 33236 13746
rect 33180 13682 33236 13694
rect 33404 13746 33684 13748
rect 33404 13694 33630 13746
rect 33682 13694 33684 13746
rect 33404 13692 33684 13694
rect 32844 13570 32900 13580
rect 31948 13524 32004 13534
rect 31500 12126 31502 12178
rect 31554 12126 31556 12178
rect 31500 12114 31556 12126
rect 31724 13522 32004 13524
rect 31724 13470 31950 13522
rect 32002 13470 32004 13522
rect 31724 13468 32004 13470
rect 31388 11954 31444 11966
rect 31388 11902 31390 11954
rect 31442 11902 31444 11954
rect 31276 11844 31332 11854
rect 31276 11394 31332 11788
rect 31388 11508 31444 11902
rect 31388 11442 31444 11452
rect 31724 11954 31780 13468
rect 31948 13458 32004 13468
rect 33292 13524 33348 13534
rect 33292 13430 33348 13468
rect 33404 13074 33460 13692
rect 33628 13682 33684 13692
rect 33516 13524 33572 13534
rect 33516 13430 33572 13468
rect 33404 13022 33406 13074
rect 33458 13022 33460 13074
rect 33404 13010 33460 13022
rect 34076 12964 34132 12974
rect 34076 12870 34132 12908
rect 34476 12572 34740 12582
rect 34532 12516 34580 12572
rect 34636 12516 34684 12572
rect 34476 12506 34740 12516
rect 31724 11902 31726 11954
rect 31778 11902 31780 11954
rect 31276 11342 31278 11394
rect 31330 11342 31332 11394
rect 31276 11330 31332 11342
rect 31724 11172 31780 11902
rect 31052 11116 31780 11172
rect 31836 11954 31892 11966
rect 31836 11902 31838 11954
rect 31890 11902 31892 11954
rect 30716 9986 30772 9996
rect 30828 10164 30884 10174
rect 30156 9884 30436 9940
rect 30156 9604 30212 9884
rect 30380 9826 30436 9884
rect 30380 9774 30382 9826
rect 30434 9774 30436 9826
rect 30380 9762 30436 9774
rect 30828 9826 30884 10108
rect 31052 10050 31108 11116
rect 31836 10388 31892 11902
rect 32060 11508 32116 11518
rect 34188 11508 34244 11518
rect 32060 11414 32116 11452
rect 33628 11506 34244 11508
rect 33628 11454 34190 11506
rect 34242 11454 34244 11506
rect 33628 11452 34244 11454
rect 33292 10722 33348 10734
rect 33292 10670 33294 10722
rect 33346 10670 33348 10722
rect 33180 10500 33236 10510
rect 31836 10322 31892 10332
rect 33068 10386 33124 10398
rect 33068 10334 33070 10386
rect 33122 10334 33124 10386
rect 31612 10164 31668 10174
rect 31052 9998 31054 10050
rect 31106 9998 31108 10050
rect 31052 9986 31108 9998
rect 31164 10052 31220 10062
rect 31164 9940 31220 9996
rect 31164 9884 31332 9940
rect 30828 9774 30830 9826
rect 30882 9774 30884 9826
rect 30268 9716 30324 9726
rect 30268 9622 30324 9660
rect 29932 9548 30212 9604
rect 29932 8930 29988 9548
rect 30380 9156 30436 9166
rect 30380 9154 30772 9156
rect 30380 9102 30382 9154
rect 30434 9102 30772 9154
rect 30380 9100 30772 9102
rect 30380 9090 30436 9100
rect 30268 9044 30324 9054
rect 29932 8878 29934 8930
rect 29986 8878 29988 8930
rect 29932 8866 29988 8878
rect 30044 9042 30324 9044
rect 30044 8990 30270 9042
rect 30322 8990 30324 9042
rect 30044 8988 30324 8990
rect 29820 8372 29988 8428
rect 29932 8278 29988 8316
rect 30044 8370 30100 8988
rect 30268 8978 30324 8988
rect 30604 8932 30660 8942
rect 30604 8838 30660 8876
rect 30318 8652 30582 8662
rect 30374 8596 30422 8652
rect 30478 8596 30526 8652
rect 30318 8586 30582 8596
rect 30716 8428 30772 9100
rect 30044 8318 30046 8370
rect 30098 8318 30100 8370
rect 30044 8306 30100 8318
rect 30380 8372 30436 8382
rect 30380 8278 30436 8316
rect 30492 8372 30772 8428
rect 30828 8428 30884 9774
rect 31276 9828 31332 9884
rect 31276 9826 31444 9828
rect 31276 9774 31278 9826
rect 31330 9774 31444 9826
rect 31276 9772 31444 9774
rect 31276 9762 31332 9772
rect 31164 9716 31220 9726
rect 31164 9156 31220 9660
rect 31164 9044 31220 9100
rect 31276 9044 31332 9054
rect 31164 9042 31332 9044
rect 31164 8990 31278 9042
rect 31330 8990 31332 9042
rect 31164 8988 31332 8990
rect 31276 8978 31332 8988
rect 31388 8484 31444 9772
rect 31276 8428 31444 8484
rect 30828 8372 30996 8428
rect 29708 8194 29764 8204
rect 29484 8148 29540 8158
rect 29484 7586 29540 8092
rect 30492 8148 30548 8372
rect 30492 8082 30548 8092
rect 30604 8260 30660 8270
rect 30940 8260 30996 8372
rect 30604 8258 30996 8260
rect 30604 8206 30606 8258
rect 30658 8206 30996 8258
rect 30604 8204 30996 8206
rect 31052 8260 31108 8270
rect 30268 7700 30324 7710
rect 30604 7700 30660 8204
rect 30940 8036 30996 8046
rect 31052 8036 31108 8204
rect 30940 8034 31108 8036
rect 30940 7982 30942 8034
rect 30994 7982 31108 8034
rect 30940 7980 31108 7982
rect 31276 8258 31332 8428
rect 31276 8206 31278 8258
rect 31330 8206 31332 8258
rect 30940 7970 30996 7980
rect 30268 7698 30660 7700
rect 30268 7646 30270 7698
rect 30322 7646 30660 7698
rect 30268 7644 30660 7646
rect 30268 7634 30324 7644
rect 29484 7534 29486 7586
rect 29538 7534 29540 7586
rect 29484 7522 29540 7534
rect 29260 7476 29316 7486
rect 29148 7420 29260 7476
rect 28588 6850 28644 6860
rect 28700 7140 28756 7150
rect 28140 6638 28142 6690
rect 28194 6638 28196 6690
rect 28140 6626 28196 6638
rect 27468 5630 27470 5682
rect 27522 5630 27524 5682
rect 27356 5348 27412 5358
rect 27244 5346 27412 5348
rect 27244 5294 27358 5346
rect 27410 5294 27412 5346
rect 27244 5292 27412 5294
rect 27356 5282 27412 5292
rect 27468 5236 27524 5630
rect 27468 5170 27524 5180
rect 27580 6578 27636 6590
rect 27580 6526 27582 6578
rect 27634 6526 27636 6578
rect 27356 5124 27412 5134
rect 27020 5122 27132 5124
rect 27020 5070 27022 5122
rect 27074 5070 27132 5122
rect 27020 5068 27132 5070
rect 27020 5058 27076 5068
rect 27132 5030 27188 5068
rect 27244 5122 27412 5124
rect 27244 5070 27358 5122
rect 27410 5070 27412 5122
rect 27244 5068 27412 5070
rect 27580 5124 27636 6526
rect 27916 6466 27972 6478
rect 27916 6414 27918 6466
rect 27970 6414 27972 6466
rect 27916 6020 27972 6414
rect 27916 5954 27972 5964
rect 28700 6018 28756 7084
rect 29148 6804 29204 7420
rect 29260 7382 29316 7420
rect 29596 7474 29652 7486
rect 29596 7422 29598 7474
rect 29650 7422 29652 7474
rect 29372 7140 29428 7150
rect 28700 5966 28702 6018
rect 28754 5966 28756 6018
rect 28700 5954 28756 5966
rect 29036 6802 29204 6804
rect 29036 6750 29150 6802
rect 29202 6750 29204 6802
rect 29036 6748 29204 6750
rect 27692 5908 27748 5918
rect 29036 5908 29092 6748
rect 29148 6738 29204 6748
rect 29260 6916 29316 6926
rect 27692 5346 27748 5852
rect 28924 5906 29092 5908
rect 28924 5854 29038 5906
rect 29090 5854 29092 5906
rect 28924 5852 29092 5854
rect 27804 5796 27860 5806
rect 27804 5702 27860 5740
rect 27692 5294 27694 5346
rect 27746 5294 27748 5346
rect 27692 5282 27748 5294
rect 28588 5124 28644 5134
rect 27580 5068 27972 5124
rect 27244 4900 27300 5068
rect 27356 5058 27412 5068
rect 26796 4844 27300 4900
rect 26160 4732 26424 4742
rect 26216 4676 26264 4732
rect 26320 4676 26368 4732
rect 26160 4666 26424 4676
rect 26796 4228 26852 4844
rect 27916 4450 27972 5068
rect 27916 4398 27918 4450
rect 27970 4398 27972 4450
rect 27916 4386 27972 4398
rect 28588 4338 28644 5068
rect 28588 4286 28590 4338
rect 28642 4286 28644 4338
rect 28588 4274 28644 4286
rect 25788 4226 26852 4228
rect 25788 4174 25790 4226
rect 25842 4174 26852 4226
rect 25788 4172 26852 4174
rect 28924 4228 28980 5852
rect 29036 5842 29092 5852
rect 29036 5682 29092 5694
rect 29036 5630 29038 5682
rect 29090 5630 29092 5682
rect 29036 5124 29092 5630
rect 29260 5346 29316 6860
rect 29372 6914 29428 7084
rect 29372 6862 29374 6914
rect 29426 6862 29428 6914
rect 29372 6850 29428 6862
rect 29596 6692 29652 7422
rect 29820 7474 29876 7486
rect 29820 7422 29822 7474
rect 29874 7422 29876 7474
rect 29820 7140 29876 7422
rect 30716 7252 30772 7262
rect 29820 7074 29876 7084
rect 30318 7084 30582 7094
rect 30374 7028 30422 7084
rect 30478 7028 30526 7084
rect 30318 7018 30582 7028
rect 29708 6804 29764 6814
rect 29708 6710 29764 6748
rect 30044 6804 30100 6814
rect 29596 6626 29652 6636
rect 29260 5294 29262 5346
rect 29314 5294 29316 5346
rect 29260 5282 29316 5294
rect 29820 6018 29876 6030
rect 29820 5966 29822 6018
rect 29874 5966 29876 6018
rect 29820 5908 29876 5966
rect 29484 5124 29540 5134
rect 29036 5122 29540 5124
rect 29036 5070 29486 5122
rect 29538 5070 29540 5122
rect 29036 5068 29540 5070
rect 29484 5058 29540 5068
rect 29708 5124 29764 5134
rect 29820 5124 29876 5852
rect 30044 5906 30100 6748
rect 30380 6804 30436 6814
rect 30380 6710 30436 6748
rect 30044 5854 30046 5906
rect 30098 5854 30100 5906
rect 30044 5842 30100 5854
rect 30156 6692 30212 6702
rect 30156 5684 30212 6636
rect 30716 6690 30772 7196
rect 30716 6638 30718 6690
rect 30770 6638 30772 6690
rect 30716 6626 30772 6638
rect 31052 6692 31108 6702
rect 31276 6692 31332 8206
rect 31500 8372 31556 8382
rect 31500 8148 31556 8316
rect 31500 8082 31556 8092
rect 31612 7474 31668 10108
rect 33068 10164 33124 10334
rect 33068 10098 33124 10108
rect 32060 9716 32116 9726
rect 32060 9714 33012 9716
rect 32060 9662 32062 9714
rect 32114 9662 33012 9714
rect 32060 9660 33012 9662
rect 32060 9650 32116 9660
rect 31836 9154 31892 9166
rect 31836 9102 31838 9154
rect 31890 9102 31892 9154
rect 31836 9044 31892 9102
rect 31836 8978 31892 8988
rect 32396 8820 32452 8830
rect 32060 8148 32116 8158
rect 31724 8146 32116 8148
rect 31724 8094 32062 8146
rect 32114 8094 32116 8146
rect 31724 8092 32116 8094
rect 31724 7698 31780 8092
rect 32060 8082 32116 8092
rect 31724 7646 31726 7698
rect 31778 7646 31780 7698
rect 31724 7634 31780 7646
rect 31612 7422 31614 7474
rect 31666 7422 31668 7474
rect 31612 7410 31668 7422
rect 31836 7476 31892 7486
rect 32284 7476 32340 7486
rect 31836 7474 32340 7476
rect 31836 7422 31838 7474
rect 31890 7422 32286 7474
rect 32338 7422 32340 7474
rect 31836 7420 32340 7422
rect 31836 7410 31892 7420
rect 32284 7410 32340 7420
rect 31388 7250 31444 7262
rect 31388 7198 31390 7250
rect 31442 7198 31444 7250
rect 31388 6916 31444 7198
rect 31388 6850 31444 6860
rect 31500 7252 31556 7262
rect 31052 6690 31332 6692
rect 31052 6638 31054 6690
rect 31106 6638 31332 6690
rect 31052 6636 31332 6638
rect 30940 6132 30996 6142
rect 30940 6020 30996 6076
rect 30828 6018 30996 6020
rect 30828 5966 30942 6018
rect 30994 5966 30996 6018
rect 30828 5964 30996 5966
rect 30604 5908 30660 5918
rect 30604 5814 30660 5852
rect 30716 5796 30772 5806
rect 30716 5702 30772 5740
rect 30156 5618 30212 5628
rect 30716 5572 30772 5582
rect 30318 5516 30582 5526
rect 30374 5460 30422 5516
rect 30478 5460 30526 5516
rect 30318 5450 30582 5460
rect 30716 5348 30772 5516
rect 30492 5292 30772 5348
rect 30492 5234 30548 5292
rect 30492 5182 30494 5234
rect 30546 5182 30548 5234
rect 30492 5170 30548 5182
rect 30268 5124 30324 5134
rect 29708 5122 30324 5124
rect 29708 5070 29710 5122
rect 29762 5070 30270 5122
rect 30322 5070 30324 5122
rect 29708 5068 30324 5070
rect 29708 5058 29764 5068
rect 30268 5058 30324 5068
rect 30716 5124 30772 5134
rect 30828 5124 30884 5964
rect 30940 5954 30996 5964
rect 30716 5122 30884 5124
rect 30716 5070 30718 5122
rect 30770 5070 30884 5122
rect 30716 5068 30884 5070
rect 30940 5348 30996 5358
rect 30940 5122 30996 5292
rect 30940 5070 30942 5122
rect 30994 5070 30996 5122
rect 30716 5058 30772 5068
rect 30940 5058 30996 5070
rect 31052 5124 31108 6636
rect 31164 5906 31220 5918
rect 31164 5854 31166 5906
rect 31218 5854 31220 5906
rect 31164 5460 31220 5854
rect 31500 5906 31556 7196
rect 32172 7252 32228 7262
rect 32172 7158 32228 7196
rect 31948 6916 32004 6926
rect 31500 5854 31502 5906
rect 31554 5854 31556 5906
rect 31500 5842 31556 5854
rect 31836 6578 31892 6590
rect 31836 6526 31838 6578
rect 31890 6526 31892 6578
rect 31724 5796 31780 5806
rect 31724 5702 31780 5740
rect 31836 5572 31892 6526
rect 31948 5906 32004 6860
rect 31948 5854 31950 5906
rect 32002 5854 32004 5906
rect 31948 5842 32004 5854
rect 31836 5506 31892 5516
rect 32060 5682 32116 5694
rect 32060 5630 32062 5682
rect 32114 5630 32116 5682
rect 31164 5394 31220 5404
rect 32060 5234 32116 5630
rect 32060 5182 32062 5234
rect 32114 5182 32116 5234
rect 32060 5170 32116 5182
rect 31276 5124 31332 5134
rect 31108 5122 31332 5124
rect 31108 5070 31278 5122
rect 31330 5070 31332 5122
rect 31108 5068 31332 5070
rect 31052 5058 31108 5068
rect 31276 5058 31332 5068
rect 31836 5124 31892 5134
rect 31892 5068 32004 5124
rect 31836 5058 31892 5068
rect 29596 4900 29652 4910
rect 29596 4806 29652 4844
rect 31164 4900 31220 4910
rect 31164 4450 31220 4844
rect 31164 4398 31166 4450
rect 31218 4398 31220 4450
rect 31164 4386 31220 4398
rect 31948 4338 32004 5068
rect 31948 4286 31950 4338
rect 32002 4286 32004 4338
rect 31948 4274 32004 4286
rect 29036 4228 29092 4238
rect 28924 4226 29092 4228
rect 28924 4174 29038 4226
rect 29090 4174 29092 4226
rect 28924 4172 29092 4174
rect 25788 4162 25844 4172
rect 29036 4162 29092 4172
rect 23996 4114 24052 4126
rect 23996 4062 23998 4114
rect 24050 4062 24052 4114
rect 23996 3892 24052 4062
rect 25228 4116 25284 4126
rect 23996 3836 24724 3892
rect 23660 3668 23716 3678
rect 23548 3666 23716 3668
rect 23548 3614 23662 3666
rect 23714 3614 23716 3666
rect 23548 3612 23716 3614
rect 22764 3602 22820 3612
rect 23660 3602 23716 3612
rect 24556 3668 24612 3678
rect 24556 3574 24612 3612
rect 24668 3666 24724 3836
rect 24668 3614 24670 3666
rect 24722 3614 24724 3666
rect 24668 3602 24724 3614
rect 22428 3490 22484 3500
rect 24892 3556 24948 3566
rect 24892 3462 24948 3500
rect 25228 3554 25284 4060
rect 30318 3948 30582 3958
rect 30374 3892 30422 3948
rect 30478 3892 30526 3948
rect 30318 3882 30582 3892
rect 32396 3668 32452 8764
rect 32508 8372 32564 8382
rect 32508 7474 32564 8316
rect 32956 7588 33012 9660
rect 33180 9266 33236 10444
rect 33292 9940 33348 10670
rect 33292 9874 33348 9884
rect 33404 10386 33460 10398
rect 33404 10334 33406 10386
rect 33458 10334 33460 10386
rect 33180 9214 33182 9266
rect 33234 9214 33236 9266
rect 33180 9202 33236 9214
rect 33068 9042 33124 9054
rect 33068 8990 33070 9042
rect 33122 8990 33124 9042
rect 33068 8428 33124 8990
rect 33292 9044 33348 9054
rect 33292 8950 33348 8988
rect 33404 8428 33460 10334
rect 33628 9156 33684 11452
rect 34188 11442 34244 11452
rect 34476 11004 34740 11014
rect 34532 10948 34580 11004
rect 34636 10948 34684 11004
rect 34476 10938 34740 10948
rect 33628 9062 33684 9100
rect 33740 10276 33796 10286
rect 33740 8428 33796 10220
rect 34188 9940 34244 9950
rect 34188 9846 34244 9884
rect 34476 9436 34740 9446
rect 34532 9380 34580 9436
rect 34636 9380 34684 9436
rect 34476 9370 34740 9380
rect 33068 8372 33236 8428
rect 33180 8260 33236 8372
rect 33068 7588 33124 7598
rect 32956 7586 33124 7588
rect 32956 7534 33070 7586
rect 33122 7534 33124 7586
rect 32956 7532 33124 7534
rect 33068 7522 33124 7532
rect 32508 7422 32510 7474
rect 32562 7422 32564 7474
rect 32508 7410 32564 7422
rect 33180 7476 33236 8204
rect 33292 8372 33460 8428
rect 33628 8372 33796 8428
rect 34188 8372 34244 8382
rect 33292 7476 33348 8372
rect 33404 7476 33460 7486
rect 33292 7474 33460 7476
rect 33292 7422 33406 7474
rect 33458 7422 33460 7474
rect 33292 7420 33460 7422
rect 33180 7410 33236 7420
rect 33404 7410 33460 7420
rect 33516 7476 33572 7486
rect 33516 7382 33572 7420
rect 33180 7250 33236 7262
rect 33180 7198 33182 7250
rect 33234 7198 33236 7250
rect 33180 6916 33236 7198
rect 33180 6850 33236 6860
rect 33292 6132 33348 6142
rect 33292 6038 33348 6076
rect 33068 5908 33124 5918
rect 33068 5814 33124 5852
rect 33628 5906 33684 8372
rect 34188 8278 34244 8316
rect 34476 7868 34740 7878
rect 34532 7812 34580 7868
rect 34636 7812 34684 7868
rect 34476 7802 34740 7812
rect 33964 6802 34020 6814
rect 33964 6750 33966 6802
rect 34018 6750 34020 6802
rect 33964 6132 34020 6750
rect 34476 6300 34740 6310
rect 34532 6244 34580 6300
rect 34636 6244 34684 6300
rect 34476 6234 34740 6244
rect 33628 5854 33630 5906
rect 33682 5854 33684 5906
rect 33628 5842 33684 5854
rect 33740 6076 33964 6132
rect 33180 5794 33236 5806
rect 33180 5742 33182 5794
rect 33234 5742 33236 5794
rect 33068 5684 33124 5694
rect 33068 4562 33124 5628
rect 33180 5348 33236 5742
rect 33180 5282 33236 5292
rect 33404 5460 33460 5470
rect 33068 4510 33070 4562
rect 33122 4510 33124 4562
rect 33068 4498 33124 4510
rect 33404 4338 33460 5404
rect 33404 4286 33406 4338
rect 33458 4286 33460 4338
rect 33404 4274 33460 4286
rect 33628 4340 33684 4350
rect 33740 4340 33796 6076
rect 33964 6066 34020 6076
rect 34188 5460 34244 5470
rect 34188 5234 34244 5404
rect 34188 5182 34190 5234
rect 34242 5182 34244 5234
rect 34188 5170 34244 5182
rect 34476 4732 34740 4742
rect 34532 4676 34580 4732
rect 34636 4676 34684 4732
rect 34476 4666 34740 4676
rect 33628 4338 33796 4340
rect 33628 4286 33630 4338
rect 33682 4286 33796 4338
rect 33628 4284 33796 4286
rect 33628 4274 33684 4284
rect 32956 3668 33012 3678
rect 32396 3666 33012 3668
rect 32396 3614 32958 3666
rect 33010 3614 33012 3666
rect 32396 3612 33012 3614
rect 25228 3502 25230 3554
rect 25282 3502 25284 3554
rect 25228 3490 25284 3502
rect 31612 3556 31668 3566
rect 31612 3554 32228 3556
rect 31612 3502 31614 3554
rect 31666 3502 32228 3554
rect 31612 3500 32228 3502
rect 31612 3490 31668 3500
rect 17948 2380 18340 2436
rect 25116 3444 25172 3454
rect 17948 800 18004 2380
rect 25116 800 25172 3388
rect 26908 3444 26964 3454
rect 26908 3350 26964 3388
rect 30044 3444 30100 3454
rect 30044 3350 30100 3388
rect 32172 3442 32228 3500
rect 32396 3554 32452 3612
rect 32956 3602 33012 3612
rect 32396 3502 32398 3554
rect 32450 3502 32452 3554
rect 32396 3490 32452 3502
rect 32172 3390 32174 3442
rect 32226 3390 32228 3442
rect 32172 3378 32228 3390
rect 32284 3444 32340 3454
rect 26160 3164 26424 3174
rect 26216 3108 26264 3164
rect 26320 3108 26368 3164
rect 26160 3098 26424 3108
rect 32284 800 32340 3388
rect 34476 3164 34740 3174
rect 34532 3108 34580 3164
rect 34636 3108 34684 3164
rect 34476 3098 34740 3108
rect 3584 0 3696 800
rect 10752 0 10864 800
rect 17920 0 18032 800
rect 25088 0 25200 800
rect 32256 0 32368 800
<< via2 >>
rect 5370 32170 5426 32172
rect 5370 32118 5372 32170
rect 5372 32118 5424 32170
rect 5424 32118 5426 32170
rect 5370 32116 5426 32118
rect 5474 32170 5530 32172
rect 5474 32118 5476 32170
rect 5476 32118 5528 32170
rect 5528 32118 5530 32170
rect 5474 32116 5530 32118
rect 5578 32170 5634 32172
rect 5578 32118 5580 32170
rect 5580 32118 5632 32170
rect 5632 32118 5634 32170
rect 5578 32116 5634 32118
rect 13686 32170 13742 32172
rect 13686 32118 13688 32170
rect 13688 32118 13740 32170
rect 13740 32118 13742 32170
rect 13686 32116 13742 32118
rect 13790 32170 13846 32172
rect 13790 32118 13792 32170
rect 13792 32118 13844 32170
rect 13844 32118 13846 32170
rect 13790 32116 13846 32118
rect 13894 32170 13950 32172
rect 13894 32118 13896 32170
rect 13896 32118 13948 32170
rect 13948 32118 13950 32170
rect 13894 32116 13950 32118
rect 22002 32170 22058 32172
rect 22002 32118 22004 32170
rect 22004 32118 22056 32170
rect 22056 32118 22058 32170
rect 22002 32116 22058 32118
rect 22106 32170 22162 32172
rect 22106 32118 22108 32170
rect 22108 32118 22160 32170
rect 22160 32118 22162 32170
rect 22106 32116 22162 32118
rect 22210 32170 22266 32172
rect 22210 32118 22212 32170
rect 22212 32118 22264 32170
rect 22264 32118 22266 32170
rect 22210 32116 22266 32118
rect 30318 32170 30374 32172
rect 30318 32118 30320 32170
rect 30320 32118 30372 32170
rect 30372 32118 30374 32170
rect 30318 32116 30374 32118
rect 30422 32170 30478 32172
rect 30422 32118 30424 32170
rect 30424 32118 30476 32170
rect 30476 32118 30478 32170
rect 30422 32116 30478 32118
rect 30526 32170 30582 32172
rect 30526 32118 30528 32170
rect 30528 32118 30580 32170
rect 30580 32118 30582 32170
rect 30526 32116 30582 32118
rect 9528 31386 9584 31388
rect 9528 31334 9530 31386
rect 9530 31334 9582 31386
rect 9582 31334 9584 31386
rect 9528 31332 9584 31334
rect 9632 31386 9688 31388
rect 9632 31334 9634 31386
rect 9634 31334 9686 31386
rect 9686 31334 9688 31386
rect 9632 31332 9688 31334
rect 9736 31386 9792 31388
rect 9736 31334 9738 31386
rect 9738 31334 9790 31386
rect 9790 31334 9792 31386
rect 9736 31332 9792 31334
rect 17844 31386 17900 31388
rect 17844 31334 17846 31386
rect 17846 31334 17898 31386
rect 17898 31334 17900 31386
rect 17844 31332 17900 31334
rect 17948 31386 18004 31388
rect 17948 31334 17950 31386
rect 17950 31334 18002 31386
rect 18002 31334 18004 31386
rect 17948 31332 18004 31334
rect 18052 31386 18108 31388
rect 18052 31334 18054 31386
rect 18054 31334 18106 31386
rect 18106 31334 18108 31386
rect 18052 31332 18108 31334
rect 26160 31386 26216 31388
rect 26160 31334 26162 31386
rect 26162 31334 26214 31386
rect 26214 31334 26216 31386
rect 26160 31332 26216 31334
rect 26264 31386 26320 31388
rect 26264 31334 26266 31386
rect 26266 31334 26318 31386
rect 26318 31334 26320 31386
rect 26264 31332 26320 31334
rect 26368 31386 26424 31388
rect 26368 31334 26370 31386
rect 26370 31334 26422 31386
rect 26422 31334 26424 31386
rect 26368 31332 26424 31334
rect 34476 31386 34532 31388
rect 34476 31334 34478 31386
rect 34478 31334 34530 31386
rect 34530 31334 34532 31386
rect 34476 31332 34532 31334
rect 34580 31386 34636 31388
rect 34580 31334 34582 31386
rect 34582 31334 34634 31386
rect 34634 31334 34636 31386
rect 34580 31332 34636 31334
rect 34684 31386 34740 31388
rect 34684 31334 34686 31386
rect 34686 31334 34738 31386
rect 34738 31334 34740 31386
rect 34684 31332 34740 31334
rect 5370 30602 5426 30604
rect 5370 30550 5372 30602
rect 5372 30550 5424 30602
rect 5424 30550 5426 30602
rect 5370 30548 5426 30550
rect 5474 30602 5530 30604
rect 5474 30550 5476 30602
rect 5476 30550 5528 30602
rect 5528 30550 5530 30602
rect 5474 30548 5530 30550
rect 5578 30602 5634 30604
rect 5578 30550 5580 30602
rect 5580 30550 5632 30602
rect 5632 30550 5634 30602
rect 5578 30548 5634 30550
rect 13686 30602 13742 30604
rect 13686 30550 13688 30602
rect 13688 30550 13740 30602
rect 13740 30550 13742 30602
rect 13686 30548 13742 30550
rect 13790 30602 13846 30604
rect 13790 30550 13792 30602
rect 13792 30550 13844 30602
rect 13844 30550 13846 30602
rect 13790 30548 13846 30550
rect 13894 30602 13950 30604
rect 13894 30550 13896 30602
rect 13896 30550 13948 30602
rect 13948 30550 13950 30602
rect 13894 30548 13950 30550
rect 22002 30602 22058 30604
rect 22002 30550 22004 30602
rect 22004 30550 22056 30602
rect 22056 30550 22058 30602
rect 22002 30548 22058 30550
rect 22106 30602 22162 30604
rect 22106 30550 22108 30602
rect 22108 30550 22160 30602
rect 22160 30550 22162 30602
rect 22106 30548 22162 30550
rect 22210 30602 22266 30604
rect 22210 30550 22212 30602
rect 22212 30550 22264 30602
rect 22264 30550 22266 30602
rect 22210 30548 22266 30550
rect 30318 30602 30374 30604
rect 30318 30550 30320 30602
rect 30320 30550 30372 30602
rect 30372 30550 30374 30602
rect 30318 30548 30374 30550
rect 30422 30602 30478 30604
rect 30422 30550 30424 30602
rect 30424 30550 30476 30602
rect 30476 30550 30478 30602
rect 30422 30548 30478 30550
rect 30526 30602 30582 30604
rect 30526 30550 30528 30602
rect 30528 30550 30580 30602
rect 30580 30550 30582 30602
rect 30526 30548 30582 30550
rect 9528 29818 9584 29820
rect 9528 29766 9530 29818
rect 9530 29766 9582 29818
rect 9582 29766 9584 29818
rect 9528 29764 9584 29766
rect 9632 29818 9688 29820
rect 9632 29766 9634 29818
rect 9634 29766 9686 29818
rect 9686 29766 9688 29818
rect 9632 29764 9688 29766
rect 9736 29818 9792 29820
rect 9736 29766 9738 29818
rect 9738 29766 9790 29818
rect 9790 29766 9792 29818
rect 9736 29764 9792 29766
rect 17844 29818 17900 29820
rect 17844 29766 17846 29818
rect 17846 29766 17898 29818
rect 17898 29766 17900 29818
rect 17844 29764 17900 29766
rect 17948 29818 18004 29820
rect 17948 29766 17950 29818
rect 17950 29766 18002 29818
rect 18002 29766 18004 29818
rect 17948 29764 18004 29766
rect 18052 29818 18108 29820
rect 18052 29766 18054 29818
rect 18054 29766 18106 29818
rect 18106 29766 18108 29818
rect 18052 29764 18108 29766
rect 26160 29818 26216 29820
rect 26160 29766 26162 29818
rect 26162 29766 26214 29818
rect 26214 29766 26216 29818
rect 26160 29764 26216 29766
rect 26264 29818 26320 29820
rect 26264 29766 26266 29818
rect 26266 29766 26318 29818
rect 26318 29766 26320 29818
rect 26264 29764 26320 29766
rect 26368 29818 26424 29820
rect 26368 29766 26370 29818
rect 26370 29766 26422 29818
rect 26422 29766 26424 29818
rect 26368 29764 26424 29766
rect 34476 29818 34532 29820
rect 34476 29766 34478 29818
rect 34478 29766 34530 29818
rect 34530 29766 34532 29818
rect 34476 29764 34532 29766
rect 34580 29818 34636 29820
rect 34580 29766 34582 29818
rect 34582 29766 34634 29818
rect 34634 29766 34636 29818
rect 34580 29764 34636 29766
rect 34684 29818 34740 29820
rect 34684 29766 34686 29818
rect 34686 29766 34738 29818
rect 34738 29766 34740 29818
rect 34684 29764 34740 29766
rect 5370 29034 5426 29036
rect 5370 28982 5372 29034
rect 5372 28982 5424 29034
rect 5424 28982 5426 29034
rect 5370 28980 5426 28982
rect 5474 29034 5530 29036
rect 5474 28982 5476 29034
rect 5476 28982 5528 29034
rect 5528 28982 5530 29034
rect 5474 28980 5530 28982
rect 5578 29034 5634 29036
rect 5578 28982 5580 29034
rect 5580 28982 5632 29034
rect 5632 28982 5634 29034
rect 5578 28980 5634 28982
rect 13686 29034 13742 29036
rect 13686 28982 13688 29034
rect 13688 28982 13740 29034
rect 13740 28982 13742 29034
rect 13686 28980 13742 28982
rect 13790 29034 13846 29036
rect 13790 28982 13792 29034
rect 13792 28982 13844 29034
rect 13844 28982 13846 29034
rect 13790 28980 13846 28982
rect 13894 29034 13950 29036
rect 13894 28982 13896 29034
rect 13896 28982 13948 29034
rect 13948 28982 13950 29034
rect 13894 28980 13950 28982
rect 22002 29034 22058 29036
rect 22002 28982 22004 29034
rect 22004 28982 22056 29034
rect 22056 28982 22058 29034
rect 22002 28980 22058 28982
rect 22106 29034 22162 29036
rect 22106 28982 22108 29034
rect 22108 28982 22160 29034
rect 22160 28982 22162 29034
rect 22106 28980 22162 28982
rect 22210 29034 22266 29036
rect 22210 28982 22212 29034
rect 22212 28982 22264 29034
rect 22264 28982 22266 29034
rect 22210 28980 22266 28982
rect 30318 29034 30374 29036
rect 30318 28982 30320 29034
rect 30320 28982 30372 29034
rect 30372 28982 30374 29034
rect 30318 28980 30374 28982
rect 30422 29034 30478 29036
rect 30422 28982 30424 29034
rect 30424 28982 30476 29034
rect 30476 28982 30478 29034
rect 30422 28980 30478 28982
rect 30526 29034 30582 29036
rect 30526 28982 30528 29034
rect 30528 28982 30580 29034
rect 30580 28982 30582 29034
rect 30526 28980 30582 28982
rect 2492 26348 2548 26404
rect 9528 28250 9584 28252
rect 9528 28198 9530 28250
rect 9530 28198 9582 28250
rect 9582 28198 9584 28250
rect 9528 28196 9584 28198
rect 9632 28250 9688 28252
rect 9632 28198 9634 28250
rect 9634 28198 9686 28250
rect 9686 28198 9688 28250
rect 9632 28196 9688 28198
rect 9736 28250 9792 28252
rect 9736 28198 9738 28250
rect 9738 28198 9790 28250
rect 9790 28198 9792 28250
rect 9736 28196 9792 28198
rect 8428 27804 8484 27860
rect 5370 27466 5426 27468
rect 5370 27414 5372 27466
rect 5372 27414 5424 27466
rect 5424 27414 5426 27466
rect 5370 27412 5426 27414
rect 5474 27466 5530 27468
rect 5474 27414 5476 27466
rect 5476 27414 5528 27466
rect 5528 27414 5530 27466
rect 5474 27412 5530 27414
rect 5578 27466 5634 27468
rect 5578 27414 5580 27466
rect 5580 27414 5632 27466
rect 5632 27414 5634 27466
rect 5578 27412 5634 27414
rect 5180 27244 5236 27300
rect 5852 27298 5908 27300
rect 5852 27246 5854 27298
rect 5854 27246 5906 27298
rect 5906 27246 5908 27298
rect 5852 27244 5908 27246
rect 5964 27074 6020 27076
rect 5964 27022 5966 27074
rect 5966 27022 6018 27074
rect 6018 27022 6020 27074
rect 5964 27020 6020 27022
rect 4956 26908 5012 26964
rect 3276 26348 3332 26404
rect 1820 25452 1876 25508
rect 2492 22258 2548 22260
rect 2492 22206 2494 22258
rect 2494 22206 2546 22258
rect 2546 22206 2548 22258
rect 2492 22204 2548 22206
rect 3276 24892 3332 24948
rect 4060 24834 4116 24836
rect 4060 24782 4062 24834
rect 4062 24782 4114 24834
rect 4114 24782 4116 24834
rect 4060 24780 4116 24782
rect 4620 25340 4676 25396
rect 5068 25340 5124 25396
rect 5180 26908 5236 26964
rect 5068 24780 5124 24836
rect 4620 24668 4676 24724
rect 5370 25898 5426 25900
rect 5370 25846 5372 25898
rect 5372 25846 5424 25898
rect 5424 25846 5426 25898
rect 5370 25844 5426 25846
rect 5474 25898 5530 25900
rect 5474 25846 5476 25898
rect 5476 25846 5528 25898
rect 5528 25846 5530 25898
rect 5474 25844 5530 25846
rect 5578 25898 5634 25900
rect 5578 25846 5580 25898
rect 5580 25846 5632 25898
rect 5632 25846 5634 25898
rect 5578 25844 5634 25846
rect 5852 25340 5908 25396
rect 5964 24780 6020 24836
rect 5628 24722 5684 24724
rect 5628 24670 5630 24722
rect 5630 24670 5682 24722
rect 5682 24670 5684 24722
rect 5628 24668 5684 24670
rect 4396 24444 4452 24500
rect 5370 24330 5426 24332
rect 5370 24278 5372 24330
rect 5372 24278 5424 24330
rect 5424 24278 5426 24330
rect 5370 24276 5426 24278
rect 5474 24330 5530 24332
rect 5474 24278 5476 24330
rect 5476 24278 5528 24330
rect 5528 24278 5530 24330
rect 5474 24276 5530 24278
rect 5578 24330 5634 24332
rect 5578 24278 5580 24330
rect 5580 24278 5632 24330
rect 5632 24278 5634 24330
rect 5578 24276 5634 24278
rect 4060 23548 4116 23604
rect 2828 23042 2884 23044
rect 2828 22990 2830 23042
rect 2830 22990 2882 23042
rect 2882 22990 2884 23042
rect 2828 22988 2884 22990
rect 4956 23212 5012 23268
rect 5404 23548 5460 23604
rect 6748 27074 6804 27076
rect 6748 27022 6750 27074
rect 6750 27022 6802 27074
rect 6802 27022 6804 27074
rect 6748 27020 6804 27022
rect 6300 26348 6356 26404
rect 6412 26908 6468 26964
rect 6188 24444 6244 24500
rect 6188 23212 6244 23268
rect 5370 22762 5426 22764
rect 5370 22710 5372 22762
rect 5372 22710 5424 22762
rect 5424 22710 5426 22762
rect 5370 22708 5426 22710
rect 5474 22762 5530 22764
rect 5474 22710 5476 22762
rect 5476 22710 5528 22762
rect 5528 22710 5530 22762
rect 5474 22708 5530 22710
rect 5578 22762 5634 22764
rect 5578 22710 5580 22762
rect 5580 22710 5632 22762
rect 5632 22710 5634 22762
rect 5578 22708 5634 22710
rect 3612 22316 3668 22372
rect 3948 21698 4004 21700
rect 3948 21646 3950 21698
rect 3950 21646 4002 21698
rect 4002 21646 4004 21698
rect 3948 21644 4004 21646
rect 5628 22258 5684 22260
rect 5628 22206 5630 22258
rect 5630 22206 5682 22258
rect 5682 22206 5684 22258
rect 5628 22204 5684 22206
rect 6076 22370 6132 22372
rect 6076 22318 6078 22370
rect 6078 22318 6130 22370
rect 6130 22318 6132 22370
rect 6076 22316 6132 22318
rect 4620 21698 4676 21700
rect 4620 21646 4622 21698
rect 4622 21646 4674 21698
rect 4674 21646 4676 21698
rect 4620 21644 4676 21646
rect 5404 21698 5460 21700
rect 5404 21646 5406 21698
rect 5406 21646 5458 21698
rect 5458 21646 5460 21698
rect 5404 21644 5460 21646
rect 3276 20802 3332 20804
rect 3276 20750 3278 20802
rect 3278 20750 3330 20802
rect 3330 20750 3332 20802
rect 3276 20748 3332 20750
rect 2380 20578 2436 20580
rect 2380 20526 2382 20578
rect 2382 20526 2434 20578
rect 2434 20526 2436 20578
rect 2380 20524 2436 20526
rect 2940 20578 2996 20580
rect 2940 20526 2942 20578
rect 2942 20526 2994 20578
rect 2994 20526 2996 20578
rect 2940 20524 2996 20526
rect 3388 20524 3444 20580
rect 5370 21194 5426 21196
rect 5370 21142 5372 21194
rect 5372 21142 5424 21194
rect 5424 21142 5426 21194
rect 5370 21140 5426 21142
rect 5474 21194 5530 21196
rect 5474 21142 5476 21194
rect 5476 21142 5528 21194
rect 5528 21142 5530 21194
rect 5474 21140 5530 21142
rect 5578 21194 5634 21196
rect 5578 21142 5580 21194
rect 5580 21142 5632 21194
rect 5632 21142 5634 21194
rect 5578 21140 5634 21142
rect 3948 20690 4004 20692
rect 3948 20638 3950 20690
rect 3950 20638 4002 20690
rect 4002 20638 4004 20690
rect 3948 20636 4004 20638
rect 4284 20578 4340 20580
rect 4284 20526 4286 20578
rect 4286 20526 4338 20578
rect 4338 20526 4340 20578
rect 4284 20524 4340 20526
rect 4396 20076 4452 20132
rect 3612 19964 3668 20020
rect 4508 19964 4564 20020
rect 4732 20748 4788 20804
rect 2604 19906 2660 19908
rect 2604 19854 2606 19906
rect 2606 19854 2658 19906
rect 2658 19854 2660 19906
rect 2604 19852 2660 19854
rect 4844 20636 4900 20692
rect 5068 20524 5124 20580
rect 6860 26962 6916 26964
rect 6860 26910 6862 26962
rect 6862 26910 6914 26962
rect 6914 26910 6916 26962
rect 6860 26908 6916 26910
rect 7308 26402 7364 26404
rect 7308 26350 7310 26402
rect 7310 26350 7362 26402
rect 7362 26350 7364 26402
rect 7308 26348 7364 26350
rect 6636 24780 6692 24836
rect 7084 25506 7140 25508
rect 7084 25454 7086 25506
rect 7086 25454 7138 25506
rect 7138 25454 7140 25506
rect 7084 25452 7140 25454
rect 6636 24444 6692 24500
rect 6636 23154 6692 23156
rect 6636 23102 6638 23154
rect 6638 23102 6690 23154
rect 6690 23102 6692 23154
rect 6636 23100 6692 23102
rect 8092 26460 8148 26516
rect 7420 25452 7476 25508
rect 9528 26682 9584 26684
rect 9528 26630 9530 26682
rect 9530 26630 9582 26682
rect 9582 26630 9584 26682
rect 9528 26628 9584 26630
rect 9632 26682 9688 26684
rect 9632 26630 9634 26682
rect 9634 26630 9686 26682
rect 9686 26630 9688 26682
rect 9632 26628 9688 26630
rect 9736 26682 9792 26684
rect 9736 26630 9738 26682
rect 9738 26630 9790 26682
rect 9790 26630 9792 26682
rect 9736 26628 9792 26630
rect 8876 26460 8932 26516
rect 7980 25452 8036 25508
rect 10220 27858 10276 27860
rect 10220 27806 10222 27858
rect 10222 27806 10274 27858
rect 10274 27806 10276 27858
rect 10220 27804 10276 27806
rect 11004 27746 11060 27748
rect 11004 27694 11006 27746
rect 11006 27694 11058 27746
rect 11058 27694 11060 27746
rect 11004 27692 11060 27694
rect 9528 25114 9584 25116
rect 9528 25062 9530 25114
rect 9530 25062 9582 25114
rect 9582 25062 9584 25114
rect 9528 25060 9584 25062
rect 9632 25114 9688 25116
rect 9632 25062 9634 25114
rect 9634 25062 9686 25114
rect 9686 25062 9688 25114
rect 9632 25060 9688 25062
rect 9736 25114 9792 25116
rect 9736 25062 9738 25114
rect 9738 25062 9790 25114
rect 9790 25062 9792 25114
rect 9736 25060 9792 25062
rect 7756 24108 7812 24164
rect 8876 24108 8932 24164
rect 6748 23042 6804 23044
rect 6748 22990 6750 23042
rect 6750 22990 6802 23042
rect 6802 22990 6804 23042
rect 6748 22988 6804 22990
rect 8988 23996 9044 24052
rect 9528 23546 9584 23548
rect 9528 23494 9530 23546
rect 9530 23494 9582 23546
rect 9582 23494 9584 23546
rect 9528 23492 9584 23494
rect 9632 23546 9688 23548
rect 9632 23494 9634 23546
rect 9634 23494 9686 23546
rect 9686 23494 9688 23546
rect 9632 23492 9688 23494
rect 9736 23546 9792 23548
rect 9736 23494 9738 23546
rect 9738 23494 9790 23546
rect 9790 23494 9792 23546
rect 9736 23492 9792 23494
rect 9996 24892 10052 24948
rect 17844 28250 17900 28252
rect 17844 28198 17846 28250
rect 17846 28198 17898 28250
rect 17898 28198 17900 28250
rect 17844 28196 17900 28198
rect 17948 28250 18004 28252
rect 17948 28198 17950 28250
rect 17950 28198 18002 28250
rect 18002 28198 18004 28250
rect 17948 28196 18004 28198
rect 18052 28250 18108 28252
rect 18052 28198 18054 28250
rect 18054 28198 18106 28250
rect 18106 28198 18108 28250
rect 18052 28196 18108 28198
rect 26160 28250 26216 28252
rect 26160 28198 26162 28250
rect 26162 28198 26214 28250
rect 26214 28198 26216 28250
rect 26160 28196 26216 28198
rect 26264 28250 26320 28252
rect 26264 28198 26266 28250
rect 26266 28198 26318 28250
rect 26318 28198 26320 28250
rect 26264 28196 26320 28198
rect 26368 28250 26424 28252
rect 26368 28198 26370 28250
rect 26370 28198 26422 28250
rect 26422 28198 26424 28250
rect 26368 28196 26424 28198
rect 34476 28250 34532 28252
rect 34476 28198 34478 28250
rect 34478 28198 34530 28250
rect 34530 28198 34532 28250
rect 34476 28196 34532 28198
rect 34580 28250 34636 28252
rect 34580 28198 34582 28250
rect 34582 28198 34634 28250
rect 34634 28198 34636 28250
rect 34580 28196 34636 28198
rect 34684 28250 34740 28252
rect 34684 28198 34686 28250
rect 34686 28198 34738 28250
rect 34738 28198 34740 28250
rect 34684 28196 34740 28198
rect 19292 27804 19348 27860
rect 12236 27692 12292 27748
rect 11004 25340 11060 25396
rect 10220 24332 10276 24388
rect 11116 24946 11172 24948
rect 11116 24894 11118 24946
rect 11118 24894 11170 24946
rect 11170 24894 11172 24946
rect 11116 24892 11172 24894
rect 11788 24780 11844 24836
rect 11116 24332 11172 24388
rect 11004 24050 11060 24052
rect 11004 23998 11006 24050
rect 11006 23998 11058 24050
rect 11058 23998 11060 24050
rect 11004 23996 11060 23998
rect 9996 23548 10052 23604
rect 11340 23772 11396 23828
rect 9996 23378 10052 23380
rect 9996 23326 9998 23378
rect 9998 23326 10050 23378
rect 10050 23326 10052 23378
rect 9996 23324 10052 23326
rect 7084 22428 7140 22484
rect 7868 22482 7924 22484
rect 7868 22430 7870 22482
rect 7870 22430 7922 22482
rect 7922 22430 7924 22482
rect 7868 22428 7924 22430
rect 8988 23042 9044 23044
rect 8988 22990 8990 23042
rect 8990 22990 9042 23042
rect 9042 22990 9044 23042
rect 8988 22988 9044 22990
rect 9884 22876 9940 22932
rect 8540 22204 8596 22260
rect 9528 21978 9584 21980
rect 9528 21926 9530 21978
rect 9530 21926 9582 21978
rect 9582 21926 9584 21978
rect 9528 21924 9584 21926
rect 9632 21978 9688 21980
rect 9632 21926 9634 21978
rect 9634 21926 9686 21978
rect 9686 21926 9688 21978
rect 9632 21924 9688 21926
rect 9736 21978 9792 21980
rect 9736 21926 9738 21978
rect 9738 21926 9790 21978
rect 9790 21926 9792 21978
rect 9736 21924 9792 21926
rect 11452 22930 11508 22932
rect 11452 22878 11454 22930
rect 11454 22878 11506 22930
rect 11506 22878 11508 22930
rect 11452 22876 11508 22878
rect 12460 26962 12516 26964
rect 12460 26910 12462 26962
rect 12462 26910 12514 26962
rect 12514 26910 12516 26962
rect 12460 26908 12516 26910
rect 12348 26290 12404 26292
rect 12348 26238 12350 26290
rect 12350 26238 12402 26290
rect 12402 26238 12404 26290
rect 12348 26236 12404 26238
rect 12348 25676 12404 25732
rect 12684 25564 12740 25620
rect 13686 27466 13742 27468
rect 13686 27414 13688 27466
rect 13688 27414 13740 27466
rect 13740 27414 13742 27466
rect 13686 27412 13742 27414
rect 13790 27466 13846 27468
rect 13790 27414 13792 27466
rect 13792 27414 13844 27466
rect 13844 27414 13846 27466
rect 13790 27412 13846 27414
rect 13894 27466 13950 27468
rect 13894 27414 13896 27466
rect 13896 27414 13948 27466
rect 13948 27414 13950 27466
rect 13894 27412 13950 27414
rect 13020 26236 13076 26292
rect 13132 27020 13188 27076
rect 14252 27074 14308 27076
rect 14252 27022 14254 27074
rect 14254 27022 14306 27074
rect 14306 27022 14308 27074
rect 14252 27020 14308 27022
rect 13686 25898 13742 25900
rect 13686 25846 13688 25898
rect 13688 25846 13740 25898
rect 13740 25846 13742 25898
rect 13686 25844 13742 25846
rect 13790 25898 13846 25900
rect 13790 25846 13792 25898
rect 13792 25846 13844 25898
rect 13844 25846 13846 25898
rect 13790 25844 13846 25846
rect 13894 25898 13950 25900
rect 13894 25846 13896 25898
rect 13896 25846 13948 25898
rect 13948 25846 13950 25898
rect 13894 25844 13950 25846
rect 14252 25676 14308 25732
rect 13580 25618 13636 25620
rect 13580 25566 13582 25618
rect 13582 25566 13634 25618
rect 13634 25566 13636 25618
rect 13580 25564 13636 25566
rect 14140 25564 14196 25620
rect 13020 25452 13076 25508
rect 13692 25506 13748 25508
rect 13692 25454 13694 25506
rect 13694 25454 13746 25506
rect 13746 25454 13748 25506
rect 13692 25452 13748 25454
rect 12012 24556 12068 24612
rect 12348 24892 12404 24948
rect 12236 24722 12292 24724
rect 12236 24670 12238 24722
rect 12238 24670 12290 24722
rect 12290 24670 12292 24722
rect 12236 24668 12292 24670
rect 12460 24610 12516 24612
rect 12460 24558 12462 24610
rect 12462 24558 12514 24610
rect 12514 24558 12516 24610
rect 12460 24556 12516 24558
rect 12124 24444 12180 24500
rect 11676 23996 11732 24052
rect 12684 24722 12740 24724
rect 12684 24670 12686 24722
rect 12686 24670 12738 24722
rect 12738 24670 12740 24722
rect 12684 24668 12740 24670
rect 13468 24780 13524 24836
rect 13244 24668 13300 24724
rect 11788 23660 11844 23716
rect 11676 23548 11732 23604
rect 10668 21756 10724 21812
rect 10780 21362 10836 21364
rect 10780 21310 10782 21362
rect 10782 21310 10834 21362
rect 10834 21310 10836 21362
rect 10780 21308 10836 21310
rect 7644 20802 7700 20804
rect 7644 20750 7646 20802
rect 7646 20750 7698 20802
rect 7698 20750 7700 20802
rect 7644 20748 7700 20750
rect 8204 20690 8260 20692
rect 8204 20638 8206 20690
rect 8206 20638 8258 20690
rect 8258 20638 8260 20690
rect 8204 20636 8260 20638
rect 5516 20076 5572 20132
rect 5292 20018 5348 20020
rect 5292 19966 5294 20018
rect 5294 19966 5346 20018
rect 5346 19966 5348 20018
rect 5292 19964 5348 19966
rect 5180 19906 5236 19908
rect 5180 19854 5182 19906
rect 5182 19854 5234 19906
rect 5234 19854 5236 19906
rect 5180 19852 5236 19854
rect 6748 19852 6804 19908
rect 5370 19626 5426 19628
rect 5370 19574 5372 19626
rect 5372 19574 5424 19626
rect 5424 19574 5426 19626
rect 5370 19572 5426 19574
rect 5474 19626 5530 19628
rect 5474 19574 5476 19626
rect 5476 19574 5528 19626
rect 5528 19574 5530 19626
rect 5474 19572 5530 19574
rect 5578 19626 5634 19628
rect 5578 19574 5580 19626
rect 5580 19574 5632 19626
rect 5632 19574 5634 19626
rect 5578 19572 5634 19574
rect 4956 19404 5012 19460
rect 4620 18396 4676 18452
rect 5628 18450 5684 18452
rect 5628 18398 5630 18450
rect 5630 18398 5682 18450
rect 5682 18398 5684 18450
rect 5628 18396 5684 18398
rect 5852 18284 5908 18340
rect 6300 18172 6356 18228
rect 6412 18396 6468 18452
rect 6636 18396 6692 18452
rect 5370 18058 5426 18060
rect 5370 18006 5372 18058
rect 5372 18006 5424 18058
rect 5424 18006 5426 18058
rect 5370 18004 5426 18006
rect 5474 18058 5530 18060
rect 5474 18006 5476 18058
rect 5476 18006 5528 18058
rect 5528 18006 5530 18058
rect 5474 18004 5530 18006
rect 5578 18058 5634 18060
rect 5578 18006 5580 18058
rect 5580 18006 5632 18058
rect 5632 18006 5634 18058
rect 5578 18004 5634 18006
rect 7420 19906 7476 19908
rect 7420 19854 7422 19906
rect 7422 19854 7474 19906
rect 7474 19854 7476 19906
rect 7420 19852 7476 19854
rect 6972 18732 7028 18788
rect 6860 18172 6916 18228
rect 1596 15148 1652 15204
rect 6188 17666 6244 17668
rect 6188 17614 6190 17666
rect 6190 17614 6242 17666
rect 6242 17614 6244 17666
rect 6188 17612 6244 17614
rect 1820 15036 1876 15092
rect 2268 15036 2324 15092
rect 2044 12124 2100 12180
rect 2940 14252 2996 14308
rect 3948 16882 4004 16884
rect 3948 16830 3950 16882
rect 3950 16830 4002 16882
rect 4002 16830 4004 16882
rect 3948 16828 4004 16830
rect 5068 16828 5124 16884
rect 5068 16604 5124 16660
rect 3276 15036 3332 15092
rect 5370 16490 5426 16492
rect 5370 16438 5372 16490
rect 5372 16438 5424 16490
rect 5424 16438 5426 16490
rect 5370 16436 5426 16438
rect 5474 16490 5530 16492
rect 5474 16438 5476 16490
rect 5476 16438 5528 16490
rect 5528 16438 5530 16490
rect 5474 16436 5530 16438
rect 5578 16490 5634 16492
rect 5578 16438 5580 16490
rect 5580 16438 5632 16490
rect 5632 16438 5634 16490
rect 5578 16436 5634 16438
rect 7084 18338 7140 18340
rect 7084 18286 7086 18338
rect 7086 18286 7138 18338
rect 7138 18286 7140 18338
rect 7084 18284 7140 18286
rect 7420 18674 7476 18676
rect 7420 18622 7422 18674
rect 7422 18622 7474 18674
rect 7474 18622 7476 18674
rect 7420 18620 7476 18622
rect 10780 20748 10836 20804
rect 9528 20410 9584 20412
rect 9528 20358 9530 20410
rect 9530 20358 9582 20410
rect 9582 20358 9584 20410
rect 9528 20356 9584 20358
rect 9632 20410 9688 20412
rect 9632 20358 9634 20410
rect 9634 20358 9686 20410
rect 9686 20358 9688 20410
rect 9632 20356 9688 20358
rect 9736 20410 9792 20412
rect 9736 20358 9738 20410
rect 9738 20358 9790 20410
rect 9790 20358 9792 20410
rect 9736 20356 9792 20358
rect 8204 20188 8260 20244
rect 10220 20188 10276 20244
rect 8876 19964 8932 20020
rect 9436 19964 9492 20020
rect 7980 19852 8036 19908
rect 8204 18732 8260 18788
rect 7308 18396 7364 18452
rect 7980 18562 8036 18564
rect 7980 18510 7982 18562
rect 7982 18510 8034 18562
rect 8034 18510 8036 18562
rect 7980 18508 8036 18510
rect 7420 17724 7476 17780
rect 7084 17666 7140 17668
rect 7084 17614 7086 17666
rect 7086 17614 7138 17666
rect 7138 17614 7140 17666
rect 7084 17612 7140 17614
rect 7420 17276 7476 17332
rect 7644 18284 7700 18340
rect 8092 18060 8148 18116
rect 8316 18284 8372 18340
rect 8204 17948 8260 18004
rect 8876 19740 8932 19796
rect 8988 19346 9044 19348
rect 8988 19294 8990 19346
rect 8990 19294 9042 19346
rect 9042 19294 9044 19346
rect 8988 19292 9044 19294
rect 9996 20018 10052 20020
rect 9996 19966 9998 20018
rect 9998 19966 10050 20018
rect 10050 19966 10052 20018
rect 9996 19964 10052 19966
rect 10444 19964 10500 20020
rect 9660 19906 9716 19908
rect 9660 19854 9662 19906
rect 9662 19854 9714 19906
rect 9714 19854 9716 19906
rect 9660 19852 9716 19854
rect 10220 19516 10276 19572
rect 9100 19068 9156 19124
rect 10668 19628 10724 19684
rect 11004 21644 11060 21700
rect 11340 21196 11396 21252
rect 12572 23884 12628 23940
rect 12796 23884 12852 23940
rect 12012 23826 12068 23828
rect 12012 23774 12014 23826
rect 12014 23774 12066 23826
rect 12066 23774 12068 23826
rect 12012 23772 12068 23774
rect 12684 23772 12740 23828
rect 12124 23324 12180 23380
rect 12124 21980 12180 22036
rect 12012 21756 12068 21812
rect 10556 19292 10612 19348
rect 10668 19180 10724 19236
rect 9772 18956 9828 19012
rect 9528 18842 9584 18844
rect 9528 18790 9530 18842
rect 9530 18790 9582 18842
rect 9582 18790 9584 18842
rect 9528 18788 9584 18790
rect 9632 18842 9688 18844
rect 9632 18790 9634 18842
rect 9634 18790 9686 18842
rect 9686 18790 9688 18842
rect 9632 18788 9688 18790
rect 9736 18842 9792 18844
rect 9736 18790 9738 18842
rect 9738 18790 9790 18842
rect 9790 18790 9792 18842
rect 9736 18788 9792 18790
rect 8428 17836 8484 17892
rect 7868 17666 7924 17668
rect 7868 17614 7870 17666
rect 7870 17614 7922 17666
rect 7922 17614 7924 17666
rect 7868 17612 7924 17614
rect 6748 16882 6804 16884
rect 6748 16830 6750 16882
rect 6750 16830 6802 16882
rect 6802 16830 6804 16882
rect 6748 16828 6804 16830
rect 7532 16882 7588 16884
rect 7532 16830 7534 16882
rect 7534 16830 7586 16882
rect 7586 16830 7588 16882
rect 7532 16828 7588 16830
rect 5370 14922 5426 14924
rect 5370 14870 5372 14922
rect 5372 14870 5424 14922
rect 5424 14870 5426 14922
rect 5370 14868 5426 14870
rect 5474 14922 5530 14924
rect 5474 14870 5476 14922
rect 5476 14870 5528 14922
rect 5528 14870 5530 14922
rect 5474 14868 5530 14870
rect 5578 14922 5634 14924
rect 5578 14870 5580 14922
rect 5580 14870 5632 14922
rect 5632 14870 5634 14922
rect 5578 14868 5634 14870
rect 4620 14642 4676 14644
rect 4620 14590 4622 14642
rect 4622 14590 4674 14642
rect 4674 14590 4676 14642
rect 4620 14588 4676 14590
rect 3276 14028 3332 14084
rect 3500 14252 3556 14308
rect 2492 13468 2548 13524
rect 2828 13020 2884 13076
rect 3388 12684 3444 12740
rect 5068 14028 5124 14084
rect 5628 14588 5684 14644
rect 5964 14306 6020 14308
rect 5964 14254 5966 14306
rect 5966 14254 6018 14306
rect 6018 14254 6020 14306
rect 5964 14252 6020 14254
rect 5964 14028 6020 14084
rect 5628 13580 5684 13636
rect 5068 13132 5124 13188
rect 2828 12178 2884 12180
rect 2828 12126 2830 12178
rect 2830 12126 2882 12178
rect 2882 12126 2884 12178
rect 2828 12124 2884 12126
rect 3612 12290 3668 12292
rect 3612 12238 3614 12290
rect 3614 12238 3666 12290
rect 3666 12238 3668 12290
rect 3612 12236 3668 12238
rect 3500 12178 3556 12180
rect 3500 12126 3502 12178
rect 3502 12126 3554 12178
rect 3554 12126 3556 12178
rect 3500 12124 3556 12126
rect 3948 11900 4004 11956
rect 3052 11506 3108 11508
rect 3052 11454 3054 11506
rect 3054 11454 3106 11506
rect 3106 11454 3108 11506
rect 3052 11452 3108 11454
rect 2156 11394 2212 11396
rect 2156 11342 2158 11394
rect 2158 11342 2210 11394
rect 2210 11342 2212 11394
rect 2156 11340 2212 11342
rect 2044 9100 2100 9156
rect 2604 11170 2660 11172
rect 2604 11118 2606 11170
rect 2606 11118 2658 11170
rect 2658 11118 2660 11170
rect 2604 11116 2660 11118
rect 2716 10050 2772 10052
rect 2716 9998 2718 10050
rect 2718 9998 2770 10050
rect 2770 9998 2772 10050
rect 2716 9996 2772 9998
rect 2156 8652 2212 8708
rect 2156 7308 2212 7364
rect 2604 9772 2660 9828
rect 2492 9154 2548 9156
rect 2492 9102 2494 9154
rect 2494 9102 2546 9154
rect 2546 9102 2548 9154
rect 2492 9100 2548 9102
rect 4508 12236 4564 12292
rect 3948 11564 4004 11620
rect 4396 12012 4452 12068
rect 4732 12738 4788 12740
rect 4732 12686 4734 12738
rect 4734 12686 4786 12738
rect 4786 12686 4788 12738
rect 4732 12684 4788 12686
rect 4620 11788 4676 11844
rect 4732 12178 4788 12180
rect 4732 12126 4734 12178
rect 4734 12126 4786 12178
rect 4786 12126 4788 12178
rect 4732 12124 4788 12126
rect 4956 12178 5012 12180
rect 4956 12126 4958 12178
rect 4958 12126 5010 12178
rect 5010 12126 5012 12178
rect 4956 12124 5012 12126
rect 4508 11676 4564 11732
rect 3500 11394 3556 11396
rect 3500 11342 3502 11394
rect 3502 11342 3554 11394
rect 3554 11342 3556 11394
rect 3500 11340 3556 11342
rect 3276 11004 3332 11060
rect 4284 11228 4340 11284
rect 3612 11116 3668 11172
rect 3276 9996 3332 10052
rect 3164 9826 3220 9828
rect 3164 9774 3166 9826
rect 3166 9774 3218 9826
rect 3218 9774 3220 9826
rect 3164 9772 3220 9774
rect 3052 9548 3108 9604
rect 2940 9212 2996 9268
rect 4284 10668 4340 10724
rect 4620 11282 4676 11284
rect 4620 11230 4622 11282
rect 4622 11230 4674 11282
rect 4674 11230 4676 11282
rect 4620 11228 4676 11230
rect 4396 10556 4452 10612
rect 3948 9996 4004 10052
rect 3500 9714 3556 9716
rect 3500 9662 3502 9714
rect 3502 9662 3554 9714
rect 3554 9662 3556 9714
rect 3500 9660 3556 9662
rect 3612 9602 3668 9604
rect 3612 9550 3614 9602
rect 3614 9550 3666 9602
rect 3666 9550 3668 9602
rect 3612 9548 3668 9550
rect 3500 9436 3556 9492
rect 2828 9154 2884 9156
rect 2828 9102 2830 9154
rect 2830 9102 2882 9154
rect 2882 9102 2884 9154
rect 2828 9100 2884 9102
rect 3612 8988 3668 9044
rect 2828 8146 2884 8148
rect 2828 8094 2830 8146
rect 2830 8094 2882 8146
rect 2882 8094 2884 8146
rect 2828 8092 2884 8094
rect 2492 7756 2548 7812
rect 3948 8988 4004 9044
rect 3612 8258 3668 8260
rect 3612 8206 3614 8258
rect 3614 8206 3666 8258
rect 3666 8206 3668 8258
rect 3612 8204 3668 8206
rect 3388 8092 3444 8148
rect 3276 7756 3332 7812
rect 2604 7308 2660 7364
rect 2716 5180 2772 5236
rect 2156 5122 2212 5124
rect 2156 5070 2158 5122
rect 2158 5070 2210 5122
rect 2210 5070 2212 5122
rect 2156 5068 2212 5070
rect 3500 7196 3556 7252
rect 3052 6188 3108 6244
rect 3164 6860 3220 6916
rect 3052 5628 3108 5684
rect 2828 5068 2884 5124
rect 3388 5068 3444 5124
rect 3836 8652 3892 8708
rect 4060 8316 4116 8372
rect 3948 7868 4004 7924
rect 3948 6972 4004 7028
rect 3836 6636 3892 6692
rect 4284 7868 4340 7924
rect 4172 7362 4228 7364
rect 4172 7310 4174 7362
rect 4174 7310 4226 7362
rect 4226 7310 4228 7362
rect 4172 7308 4228 7310
rect 4060 6636 4116 6692
rect 4396 8092 4452 8148
rect 4620 9660 4676 9716
rect 4956 11676 5012 11732
rect 5068 10610 5124 10612
rect 5068 10558 5070 10610
rect 5070 10558 5122 10610
rect 5122 10558 5124 10610
rect 5068 10556 5124 10558
rect 5068 10332 5124 10388
rect 5370 13354 5426 13356
rect 5370 13302 5372 13354
rect 5372 13302 5424 13354
rect 5424 13302 5426 13354
rect 5370 13300 5426 13302
rect 5474 13354 5530 13356
rect 5474 13302 5476 13354
rect 5476 13302 5528 13354
rect 5528 13302 5530 13354
rect 5474 13300 5530 13302
rect 5578 13354 5634 13356
rect 5578 13302 5580 13354
rect 5580 13302 5632 13354
rect 5632 13302 5634 13354
rect 5578 13300 5634 13302
rect 5628 12962 5684 12964
rect 5628 12910 5630 12962
rect 5630 12910 5682 12962
rect 5682 12910 5684 12962
rect 5628 12908 5684 12910
rect 5292 12684 5348 12740
rect 5628 12402 5684 12404
rect 5628 12350 5630 12402
rect 5630 12350 5682 12402
rect 5682 12350 5684 12402
rect 5628 12348 5684 12350
rect 5852 12124 5908 12180
rect 5370 11786 5426 11788
rect 5370 11734 5372 11786
rect 5372 11734 5424 11786
rect 5424 11734 5426 11786
rect 5370 11732 5426 11734
rect 5474 11786 5530 11788
rect 5474 11734 5476 11786
rect 5476 11734 5528 11786
rect 5528 11734 5530 11786
rect 5474 11732 5530 11734
rect 5578 11786 5634 11788
rect 5578 11734 5580 11786
rect 5580 11734 5632 11786
rect 5632 11734 5634 11786
rect 5578 11732 5634 11734
rect 5516 11394 5572 11396
rect 5516 11342 5518 11394
rect 5518 11342 5570 11394
rect 5570 11342 5572 11394
rect 5516 11340 5572 11342
rect 5852 11282 5908 11284
rect 5852 11230 5854 11282
rect 5854 11230 5906 11282
rect 5906 11230 5908 11282
rect 5852 11228 5908 11230
rect 5516 10332 5572 10388
rect 5370 10218 5426 10220
rect 5370 10166 5372 10218
rect 5372 10166 5424 10218
rect 5424 10166 5426 10218
rect 5370 10164 5426 10166
rect 5474 10218 5530 10220
rect 5474 10166 5476 10218
rect 5476 10166 5528 10218
rect 5528 10166 5530 10218
rect 5474 10164 5530 10166
rect 5578 10218 5634 10220
rect 5578 10166 5580 10218
rect 5580 10166 5632 10218
rect 5632 10166 5634 10218
rect 5578 10164 5634 10166
rect 4844 9436 4900 9492
rect 4620 9212 4676 9268
rect 4844 9212 4900 9268
rect 4508 7644 4564 7700
rect 4732 8204 4788 8260
rect 4732 7420 4788 7476
rect 4956 8258 5012 8260
rect 4956 8206 4958 8258
rect 4958 8206 5010 8258
rect 5010 8206 5012 8258
rect 4956 8204 5012 8206
rect 5628 9826 5684 9828
rect 5628 9774 5630 9826
rect 5630 9774 5682 9826
rect 5682 9774 5684 9826
rect 5628 9772 5684 9774
rect 5740 9436 5796 9492
rect 5516 8876 5572 8932
rect 5370 8650 5426 8652
rect 5370 8598 5372 8650
rect 5372 8598 5424 8650
rect 5424 8598 5426 8650
rect 5370 8596 5426 8598
rect 5474 8650 5530 8652
rect 5474 8598 5476 8650
rect 5476 8598 5528 8650
rect 5528 8598 5530 8650
rect 5474 8596 5530 8598
rect 5578 8650 5634 8652
rect 5578 8598 5580 8650
rect 5580 8598 5632 8650
rect 5632 8598 5634 8650
rect 5578 8596 5634 8598
rect 5628 8316 5684 8372
rect 5628 7980 5684 8036
rect 4844 6860 4900 6916
rect 5292 7474 5348 7476
rect 5292 7422 5294 7474
rect 5294 7422 5346 7474
rect 5346 7422 5348 7474
rect 5292 7420 5348 7422
rect 5852 8428 5908 8484
rect 5852 8258 5908 8260
rect 5852 8206 5854 8258
rect 5854 8206 5906 8258
rect 5906 8206 5908 8258
rect 5852 8204 5908 8206
rect 5740 7474 5796 7476
rect 5740 7422 5742 7474
rect 5742 7422 5794 7474
rect 5794 7422 5796 7474
rect 5740 7420 5796 7422
rect 5370 7082 5426 7084
rect 5370 7030 5372 7082
rect 5372 7030 5424 7082
rect 5424 7030 5426 7082
rect 5370 7028 5426 7030
rect 5474 7082 5530 7084
rect 5474 7030 5476 7082
rect 5476 7030 5528 7082
rect 5528 7030 5530 7082
rect 5474 7028 5530 7030
rect 5578 7082 5634 7084
rect 5578 7030 5580 7082
rect 5580 7030 5632 7082
rect 5632 7030 5634 7082
rect 5578 7028 5634 7030
rect 4732 6748 4788 6804
rect 4956 6690 5012 6692
rect 4956 6638 4958 6690
rect 4958 6638 5010 6690
rect 5010 6638 5012 6690
rect 4956 6636 5012 6638
rect 5628 6690 5684 6692
rect 5628 6638 5630 6690
rect 5630 6638 5682 6690
rect 5682 6638 5684 6690
rect 5628 6636 5684 6638
rect 5852 6636 5908 6692
rect 5068 6578 5124 6580
rect 5068 6526 5070 6578
rect 5070 6526 5122 6578
rect 5122 6526 5124 6578
rect 5068 6524 5124 6526
rect 5852 6300 5908 6356
rect 4620 6188 4676 6244
rect 5516 6130 5572 6132
rect 5516 6078 5518 6130
rect 5518 6078 5570 6130
rect 5570 6078 5572 6130
rect 5516 6076 5572 6078
rect 4508 5964 4564 6020
rect 4284 5180 4340 5236
rect 3612 4732 3668 4788
rect 5852 6018 5908 6020
rect 5852 5966 5854 6018
rect 5854 5966 5906 6018
rect 5906 5966 5908 6018
rect 5852 5964 5908 5966
rect 5370 5514 5426 5516
rect 5370 5462 5372 5514
rect 5372 5462 5424 5514
rect 5424 5462 5426 5514
rect 5370 5460 5426 5462
rect 5474 5514 5530 5516
rect 5474 5462 5476 5514
rect 5476 5462 5528 5514
rect 5528 5462 5530 5514
rect 5474 5460 5530 5462
rect 5578 5514 5634 5516
rect 5578 5462 5580 5514
rect 5580 5462 5632 5514
rect 5632 5462 5634 5514
rect 5578 5460 5634 5462
rect 6860 14252 6916 14308
rect 6076 12236 6132 12292
rect 6076 11900 6132 11956
rect 6076 11004 6132 11060
rect 6412 13356 6468 13412
rect 6412 13132 6468 13188
rect 8876 18562 8932 18564
rect 8876 18510 8878 18562
rect 8878 18510 8930 18562
rect 8930 18510 8932 18562
rect 8876 18508 8932 18510
rect 8876 18226 8932 18228
rect 8876 18174 8878 18226
rect 8878 18174 8930 18226
rect 8930 18174 8932 18226
rect 8876 18172 8932 18174
rect 8540 17612 8596 17668
rect 8204 17500 8260 17556
rect 9100 17500 9156 17556
rect 9660 18562 9716 18564
rect 9660 18510 9662 18562
rect 9662 18510 9714 18562
rect 9714 18510 9716 18562
rect 9660 18508 9716 18510
rect 9884 18284 9940 18340
rect 10556 19122 10612 19124
rect 10556 19070 10558 19122
rect 10558 19070 10610 19122
rect 10610 19070 10612 19122
rect 10556 19068 10612 19070
rect 10556 18620 10612 18676
rect 10108 18226 10164 18228
rect 10108 18174 10110 18226
rect 10110 18174 10162 18226
rect 10162 18174 10164 18226
rect 10108 18172 10164 18174
rect 9660 17948 9716 18004
rect 9548 17890 9604 17892
rect 9548 17838 9550 17890
rect 9550 17838 9602 17890
rect 9602 17838 9604 17890
rect 9548 17836 9604 17838
rect 10556 18450 10612 18452
rect 10556 18398 10558 18450
rect 10558 18398 10610 18450
rect 10610 18398 10612 18450
rect 10556 18396 10612 18398
rect 11452 20690 11508 20692
rect 11452 20638 11454 20690
rect 11454 20638 11506 20690
rect 11506 20638 11508 20690
rect 11452 20636 11508 20638
rect 11340 20076 11396 20132
rect 12348 21868 12404 21924
rect 12348 21532 12404 21588
rect 12572 23042 12628 23044
rect 12572 22990 12574 23042
rect 12574 22990 12626 23042
rect 12626 22990 12628 23042
rect 12572 22988 12628 22990
rect 12684 22876 12740 22932
rect 12460 21420 12516 21476
rect 12684 22316 12740 22372
rect 12348 20748 12404 20804
rect 12572 21308 12628 21364
rect 12908 23436 12964 23492
rect 17500 27074 17556 27076
rect 17500 27022 17502 27074
rect 17502 27022 17554 27074
rect 17554 27022 17556 27074
rect 17500 27020 17556 27022
rect 14700 25506 14756 25508
rect 14700 25454 14702 25506
rect 14702 25454 14754 25506
rect 14754 25454 14756 25506
rect 14700 25452 14756 25454
rect 14588 24722 14644 24724
rect 14588 24670 14590 24722
rect 14590 24670 14642 24722
rect 14642 24670 14644 24722
rect 14588 24668 14644 24670
rect 14140 24610 14196 24612
rect 14140 24558 14142 24610
rect 14142 24558 14194 24610
rect 14194 24558 14196 24610
rect 14140 24556 14196 24558
rect 13686 24330 13742 24332
rect 13686 24278 13688 24330
rect 13688 24278 13740 24330
rect 13740 24278 13742 24330
rect 13686 24276 13742 24278
rect 13790 24330 13846 24332
rect 13790 24278 13792 24330
rect 13792 24278 13844 24330
rect 13844 24278 13846 24330
rect 13790 24276 13846 24278
rect 13894 24330 13950 24332
rect 13894 24278 13896 24330
rect 13896 24278 13948 24330
rect 13948 24278 13950 24330
rect 13894 24276 13950 24278
rect 13580 23772 13636 23828
rect 13468 23548 13524 23604
rect 13132 23212 13188 23268
rect 12908 22092 12964 22148
rect 12796 21532 12852 21588
rect 13020 21980 13076 22036
rect 13692 23714 13748 23716
rect 13692 23662 13694 23714
rect 13694 23662 13746 23714
rect 13746 23662 13748 23714
rect 13692 23660 13748 23662
rect 14140 24332 14196 24388
rect 14924 25394 14980 25396
rect 14924 25342 14926 25394
rect 14926 25342 14978 25394
rect 14978 25342 14980 25394
rect 14924 25340 14980 25342
rect 15484 25506 15540 25508
rect 15484 25454 15486 25506
rect 15486 25454 15538 25506
rect 15538 25454 15540 25506
rect 15484 25452 15540 25454
rect 15260 25116 15316 25172
rect 16268 26124 16324 26180
rect 16268 25394 16324 25396
rect 16268 25342 16270 25394
rect 16270 25342 16322 25394
rect 16322 25342 16324 25394
rect 16268 25340 16324 25342
rect 15708 25116 15764 25172
rect 16380 25116 16436 25172
rect 16604 25282 16660 25284
rect 16604 25230 16606 25282
rect 16606 25230 16658 25282
rect 16658 25230 16660 25282
rect 16604 25228 16660 25230
rect 17612 26908 17668 26964
rect 17500 26236 17556 26292
rect 17844 26682 17900 26684
rect 17844 26630 17846 26682
rect 17846 26630 17898 26682
rect 17898 26630 17900 26682
rect 17844 26628 17900 26630
rect 17948 26682 18004 26684
rect 17948 26630 17950 26682
rect 17950 26630 18002 26682
rect 18002 26630 18004 26682
rect 17948 26628 18004 26630
rect 18052 26682 18108 26684
rect 18052 26630 18054 26682
rect 18054 26630 18106 26682
rect 18106 26630 18108 26682
rect 18052 26628 18108 26630
rect 18284 26908 18340 26964
rect 19068 26402 19124 26404
rect 19068 26350 19070 26402
rect 19070 26350 19122 26402
rect 19122 26350 19124 26402
rect 19068 26348 19124 26350
rect 18844 26124 18900 26180
rect 19516 27132 19572 27188
rect 19516 25564 19572 25620
rect 18844 25452 18900 25508
rect 16940 25228 16996 25284
rect 17500 25228 17556 25284
rect 15260 24332 15316 24388
rect 14028 23772 14084 23828
rect 13916 23714 13972 23716
rect 13916 23662 13918 23714
rect 13918 23662 13970 23714
rect 13970 23662 13972 23714
rect 13916 23660 13972 23662
rect 13916 23436 13972 23492
rect 13916 22876 13972 22932
rect 13686 22762 13742 22764
rect 13686 22710 13688 22762
rect 13688 22710 13740 22762
rect 13740 22710 13742 22762
rect 13686 22708 13742 22710
rect 13790 22762 13846 22764
rect 13790 22710 13792 22762
rect 13792 22710 13844 22762
rect 13844 22710 13846 22762
rect 13790 22708 13846 22710
rect 13894 22762 13950 22764
rect 13894 22710 13896 22762
rect 13896 22710 13948 22762
rect 13948 22710 13950 22762
rect 13894 22708 13950 22710
rect 14476 23548 14532 23604
rect 13468 22316 13524 22372
rect 14364 22876 14420 22932
rect 13580 22204 13636 22260
rect 13468 21698 13524 21700
rect 13468 21646 13470 21698
rect 13470 21646 13522 21698
rect 13522 21646 13524 21698
rect 13468 21644 13524 21646
rect 12684 21026 12740 21028
rect 12684 20974 12686 21026
rect 12686 20974 12738 21026
rect 12738 20974 12740 21026
rect 12684 20972 12740 20974
rect 12684 20690 12740 20692
rect 12684 20638 12686 20690
rect 12686 20638 12738 20690
rect 12738 20638 12740 20690
rect 12684 20636 12740 20638
rect 12796 20524 12852 20580
rect 12124 20188 12180 20244
rect 10780 18956 10836 19012
rect 10220 17666 10276 17668
rect 10220 17614 10222 17666
rect 10222 17614 10274 17666
rect 10274 17614 10276 17666
rect 10220 17612 10276 17614
rect 11116 19180 11172 19236
rect 11452 18732 11508 18788
rect 11340 18508 11396 18564
rect 11004 18172 11060 18228
rect 10668 17554 10724 17556
rect 10668 17502 10670 17554
rect 10670 17502 10722 17554
rect 10722 17502 10724 17554
rect 10668 17500 10724 17502
rect 9772 17442 9828 17444
rect 9772 17390 9774 17442
rect 9774 17390 9826 17442
rect 9826 17390 9828 17442
rect 9772 17388 9828 17390
rect 9528 17274 9584 17276
rect 9528 17222 9530 17274
rect 9530 17222 9582 17274
rect 9582 17222 9584 17274
rect 9528 17220 9584 17222
rect 9632 17274 9688 17276
rect 9632 17222 9634 17274
rect 9634 17222 9686 17274
rect 9686 17222 9688 17274
rect 9632 17220 9688 17222
rect 9736 17274 9792 17276
rect 9736 17222 9738 17274
rect 9738 17222 9790 17274
rect 9790 17222 9792 17274
rect 9736 17220 9792 17222
rect 9884 17276 9940 17332
rect 11452 18396 11508 18452
rect 13686 21194 13742 21196
rect 13686 21142 13688 21194
rect 13688 21142 13740 21194
rect 13740 21142 13742 21194
rect 13686 21140 13742 21142
rect 13790 21194 13846 21196
rect 13790 21142 13792 21194
rect 13792 21142 13844 21194
rect 13844 21142 13846 21194
rect 13790 21140 13846 21142
rect 13894 21194 13950 21196
rect 13894 21142 13896 21194
rect 13896 21142 13948 21194
rect 13948 21142 13950 21194
rect 13894 21140 13950 21142
rect 14476 21756 14532 21812
rect 14588 22988 14644 23044
rect 13020 20076 13076 20132
rect 12572 19964 12628 20020
rect 12572 19628 12628 19684
rect 12236 19346 12292 19348
rect 12236 19294 12238 19346
rect 12238 19294 12290 19346
rect 12290 19294 12292 19346
rect 12236 19292 12292 19294
rect 11900 18620 11956 18676
rect 12124 18508 12180 18564
rect 11900 18396 11956 18452
rect 12348 18338 12404 18340
rect 12348 18286 12350 18338
rect 12350 18286 12402 18338
rect 12402 18286 12404 18338
rect 12348 18284 12404 18286
rect 11788 18172 11844 18228
rect 13580 20578 13636 20580
rect 13580 20526 13582 20578
rect 13582 20526 13634 20578
rect 13634 20526 13636 20578
rect 13580 20524 13636 20526
rect 14364 20748 14420 20804
rect 14140 20524 14196 20580
rect 13580 20076 13636 20132
rect 14252 20130 14308 20132
rect 14252 20078 14254 20130
rect 14254 20078 14306 20130
rect 14306 20078 14308 20130
rect 14252 20076 14308 20078
rect 13356 19292 13412 19348
rect 14700 23660 14756 23716
rect 14812 23266 14868 23268
rect 14812 23214 14814 23266
rect 14814 23214 14866 23266
rect 14866 23214 14868 23266
rect 14812 23212 14868 23214
rect 14924 22988 14980 23044
rect 14700 21868 14756 21924
rect 15036 22092 15092 22148
rect 14812 21698 14868 21700
rect 14812 21646 14814 21698
rect 14814 21646 14866 21698
rect 14866 21646 14868 21698
rect 14812 21644 14868 21646
rect 15372 23996 15428 24052
rect 15596 23884 15652 23940
rect 15372 23436 15428 23492
rect 15932 23772 15988 23828
rect 17164 23826 17220 23828
rect 17164 23774 17166 23826
rect 17166 23774 17218 23826
rect 17218 23774 17220 23826
rect 17164 23772 17220 23774
rect 17388 23378 17444 23380
rect 17388 23326 17390 23378
rect 17390 23326 17442 23378
rect 17442 23326 17444 23378
rect 17388 23324 17444 23326
rect 15820 23266 15876 23268
rect 15820 23214 15822 23266
rect 15822 23214 15874 23266
rect 15874 23214 15876 23266
rect 15820 23212 15876 23214
rect 16044 22876 16100 22932
rect 15260 21868 15316 21924
rect 15708 21810 15764 21812
rect 15708 21758 15710 21810
rect 15710 21758 15762 21810
rect 15762 21758 15764 21810
rect 15708 21756 15764 21758
rect 15372 21474 15428 21476
rect 15372 21422 15374 21474
rect 15374 21422 15426 21474
rect 15426 21422 15428 21474
rect 15372 21420 15428 21422
rect 15484 20972 15540 21028
rect 15596 21420 15652 21476
rect 14028 19852 14084 19908
rect 12908 18172 12964 18228
rect 12796 18060 12852 18116
rect 11116 17442 11172 17444
rect 11116 17390 11118 17442
rect 11118 17390 11170 17442
rect 11170 17390 11172 17442
rect 11116 17388 11172 17390
rect 11228 17276 11284 17332
rect 10444 17052 10500 17108
rect 10780 16828 10836 16884
rect 12124 16882 12180 16884
rect 12124 16830 12126 16882
rect 12126 16830 12178 16882
rect 12178 16830 12180 16882
rect 12124 16828 12180 16830
rect 12908 16828 12964 16884
rect 12236 16716 12292 16772
rect 12796 16156 12852 16212
rect 13686 19626 13742 19628
rect 13686 19574 13688 19626
rect 13688 19574 13740 19626
rect 13740 19574 13742 19626
rect 13686 19572 13742 19574
rect 13790 19626 13846 19628
rect 13790 19574 13792 19626
rect 13792 19574 13844 19626
rect 13844 19574 13846 19626
rect 13790 19572 13846 19574
rect 13894 19626 13950 19628
rect 13894 19574 13896 19626
rect 13896 19574 13948 19626
rect 13948 19574 13950 19626
rect 13894 19572 13950 19574
rect 14700 19740 14756 19796
rect 13916 19404 13972 19460
rect 14028 18450 14084 18452
rect 14028 18398 14030 18450
rect 14030 18398 14082 18450
rect 14082 18398 14084 18450
rect 14028 18396 14084 18398
rect 14700 18338 14756 18340
rect 14700 18286 14702 18338
rect 14702 18286 14754 18338
rect 14754 18286 14756 18338
rect 14700 18284 14756 18286
rect 13686 18058 13742 18060
rect 13686 18006 13688 18058
rect 13688 18006 13740 18058
rect 13740 18006 13742 18058
rect 13686 18004 13742 18006
rect 13790 18058 13846 18060
rect 13790 18006 13792 18058
rect 13792 18006 13844 18058
rect 13844 18006 13846 18058
rect 13790 18004 13846 18006
rect 13894 18058 13950 18060
rect 13894 18006 13896 18058
rect 13896 18006 13948 18058
rect 13948 18006 13950 18058
rect 13894 18004 13950 18006
rect 14364 17500 14420 17556
rect 14140 16828 14196 16884
rect 14028 16770 14084 16772
rect 14028 16718 14030 16770
rect 14030 16718 14082 16770
rect 14082 16718 14084 16770
rect 14028 16716 14084 16718
rect 13916 16604 13972 16660
rect 13686 16490 13742 16492
rect 13686 16438 13688 16490
rect 13688 16438 13740 16490
rect 13740 16438 13742 16490
rect 13686 16436 13742 16438
rect 13790 16490 13846 16492
rect 13790 16438 13792 16490
rect 13792 16438 13844 16490
rect 13844 16438 13846 16490
rect 13790 16436 13846 16438
rect 13894 16490 13950 16492
rect 13894 16438 13896 16490
rect 13896 16438 13948 16490
rect 13948 16438 13950 16490
rect 13894 16436 13950 16438
rect 13692 16210 13748 16212
rect 13692 16158 13694 16210
rect 13694 16158 13746 16210
rect 13746 16158 13748 16210
rect 13692 16156 13748 16158
rect 14140 15986 14196 15988
rect 14140 15934 14142 15986
rect 14142 15934 14194 15986
rect 14194 15934 14196 15986
rect 14140 15932 14196 15934
rect 15260 19852 15316 19908
rect 16828 21810 16884 21812
rect 16828 21758 16830 21810
rect 16830 21758 16882 21810
rect 16882 21758 16884 21810
rect 16828 21756 16884 21758
rect 16492 21308 16548 21364
rect 15820 20914 15876 20916
rect 15820 20862 15822 20914
rect 15822 20862 15874 20914
rect 15874 20862 15876 20914
rect 15820 20860 15876 20862
rect 16716 20860 16772 20916
rect 16044 20802 16100 20804
rect 16044 20750 16046 20802
rect 16046 20750 16098 20802
rect 16098 20750 16100 20802
rect 16044 20748 16100 20750
rect 17844 25114 17900 25116
rect 17844 25062 17846 25114
rect 17846 25062 17898 25114
rect 17898 25062 17900 25114
rect 17844 25060 17900 25062
rect 17948 25114 18004 25116
rect 17948 25062 17950 25114
rect 17950 25062 18002 25114
rect 18002 25062 18004 25114
rect 17948 25060 18004 25062
rect 18052 25114 18108 25116
rect 18052 25062 18054 25114
rect 18054 25062 18106 25114
rect 18106 25062 18108 25114
rect 18052 25060 18108 25062
rect 19516 25394 19572 25396
rect 19516 25342 19518 25394
rect 19518 25342 19570 25394
rect 19570 25342 19572 25394
rect 19516 25340 19572 25342
rect 19292 25228 19348 25284
rect 18172 24834 18228 24836
rect 18172 24782 18174 24834
rect 18174 24782 18226 24834
rect 18226 24782 18228 24834
rect 18172 24780 18228 24782
rect 17844 23546 17900 23548
rect 17844 23494 17846 23546
rect 17846 23494 17898 23546
rect 17898 23494 17900 23546
rect 17844 23492 17900 23494
rect 17948 23546 18004 23548
rect 17948 23494 17950 23546
rect 17950 23494 18002 23546
rect 18002 23494 18004 23546
rect 17948 23492 18004 23494
rect 18052 23546 18108 23548
rect 18052 23494 18054 23546
rect 18054 23494 18106 23546
rect 18106 23494 18108 23546
rect 18052 23492 18108 23494
rect 17836 23324 17892 23380
rect 17724 23042 17780 23044
rect 17724 22990 17726 23042
rect 17726 22990 17778 23042
rect 17778 22990 17780 23042
rect 17724 22988 17780 22990
rect 18284 23660 18340 23716
rect 18172 23100 18228 23156
rect 19292 23660 19348 23716
rect 19068 23378 19124 23380
rect 19068 23326 19070 23378
rect 19070 23326 19122 23378
rect 19122 23326 19124 23378
rect 19068 23324 19124 23326
rect 17844 21978 17900 21980
rect 17844 21926 17846 21978
rect 17846 21926 17898 21978
rect 17898 21926 17900 21978
rect 17844 21924 17900 21926
rect 17948 21978 18004 21980
rect 17948 21926 17950 21978
rect 17950 21926 18002 21978
rect 18002 21926 18004 21978
rect 17948 21924 18004 21926
rect 18052 21978 18108 21980
rect 18052 21926 18054 21978
rect 18054 21926 18106 21978
rect 18106 21926 18108 21978
rect 18052 21924 18108 21926
rect 17612 21474 17668 21476
rect 17612 21422 17614 21474
rect 17614 21422 17666 21474
rect 17666 21422 17668 21474
rect 17612 21420 17668 21422
rect 18172 21420 18228 21476
rect 17500 20412 17556 20468
rect 16940 20076 16996 20132
rect 16380 19964 16436 20020
rect 14812 16268 14868 16324
rect 16604 19852 16660 19908
rect 15932 19740 15988 19796
rect 14700 15932 14756 15988
rect 9528 15706 9584 15708
rect 9528 15654 9530 15706
rect 9530 15654 9582 15706
rect 9582 15654 9584 15706
rect 9528 15652 9584 15654
rect 9632 15706 9688 15708
rect 9632 15654 9634 15706
rect 9634 15654 9686 15706
rect 9686 15654 9688 15706
rect 9632 15652 9688 15654
rect 9736 15706 9792 15708
rect 9736 15654 9738 15706
rect 9738 15654 9790 15706
rect 9790 15654 9792 15706
rect 9736 15652 9792 15654
rect 11228 15314 11284 15316
rect 11228 15262 11230 15314
rect 11230 15262 11282 15314
rect 11282 15262 11284 15314
rect 11228 15260 11284 15262
rect 13468 15260 13524 15316
rect 8988 15036 9044 15092
rect 7756 13916 7812 13972
rect 9996 15036 10052 15092
rect 12684 14252 12740 14308
rect 8428 14028 8484 14084
rect 9528 14138 9584 14140
rect 9528 14086 9530 14138
rect 9530 14086 9582 14138
rect 9582 14086 9584 14138
rect 9528 14084 9584 14086
rect 9632 14138 9688 14140
rect 9632 14086 9634 14138
rect 9634 14086 9686 14138
rect 9686 14086 9688 14138
rect 9632 14084 9688 14086
rect 9736 14138 9792 14140
rect 9736 14086 9738 14138
rect 9738 14086 9790 14138
rect 9790 14086 9792 14138
rect 9736 14084 9792 14086
rect 6972 13692 7028 13748
rect 6636 13468 6692 13524
rect 6748 12962 6804 12964
rect 6748 12910 6750 12962
rect 6750 12910 6802 12962
rect 6802 12910 6804 12962
rect 6748 12908 6804 12910
rect 6860 12738 6916 12740
rect 6860 12686 6862 12738
rect 6862 12686 6914 12738
rect 6914 12686 6916 12738
rect 6860 12684 6916 12686
rect 6412 12402 6468 12404
rect 6412 12350 6414 12402
rect 6414 12350 6466 12402
rect 6466 12350 6468 12402
rect 6412 12348 6468 12350
rect 6636 12348 6692 12404
rect 6300 11394 6356 11396
rect 6300 11342 6302 11394
rect 6302 11342 6354 11394
rect 6354 11342 6356 11394
rect 6300 11340 6356 11342
rect 6748 12290 6804 12292
rect 6748 12238 6750 12290
rect 6750 12238 6802 12290
rect 6802 12238 6804 12290
rect 6748 12236 6804 12238
rect 7084 13132 7140 13188
rect 7756 13132 7812 13188
rect 7420 13074 7476 13076
rect 7420 13022 7422 13074
rect 7422 13022 7474 13074
rect 7474 13022 7476 13074
rect 7420 13020 7476 13022
rect 7196 12684 7252 12740
rect 7084 12402 7140 12404
rect 7084 12350 7086 12402
rect 7086 12350 7138 12402
rect 7138 12350 7140 12402
rect 7084 12348 7140 12350
rect 6972 11564 7028 11620
rect 7084 11394 7140 11396
rect 7084 11342 7086 11394
rect 7086 11342 7138 11394
rect 7138 11342 7140 11394
rect 7084 11340 7140 11342
rect 7532 12348 7588 12404
rect 7308 12236 7364 12292
rect 7420 11676 7476 11732
rect 11900 13916 11956 13972
rect 10556 13858 10612 13860
rect 10556 13806 10558 13858
rect 10558 13806 10610 13858
rect 10610 13806 10612 13858
rect 10556 13804 10612 13806
rect 10332 13746 10388 13748
rect 10332 13694 10334 13746
rect 10334 13694 10386 13746
rect 10386 13694 10388 13746
rect 10332 13692 10388 13694
rect 10108 13468 10164 13524
rect 8652 13356 8708 13412
rect 8428 12908 8484 12964
rect 8540 13020 8596 13076
rect 9528 12570 9584 12572
rect 9528 12518 9530 12570
rect 9530 12518 9582 12570
rect 9582 12518 9584 12570
rect 9528 12516 9584 12518
rect 9632 12570 9688 12572
rect 9632 12518 9634 12570
rect 9634 12518 9686 12570
rect 9686 12518 9688 12570
rect 9632 12516 9688 12518
rect 9736 12570 9792 12572
rect 9736 12518 9738 12570
rect 9738 12518 9790 12570
rect 9790 12518 9792 12570
rect 9736 12516 9792 12518
rect 9884 12402 9940 12404
rect 9884 12350 9886 12402
rect 9886 12350 9938 12402
rect 9938 12350 9940 12402
rect 9884 12348 9940 12350
rect 11788 13858 11844 13860
rect 11788 13806 11790 13858
rect 11790 13806 11842 13858
rect 11842 13806 11844 13858
rect 11788 13804 11844 13806
rect 11900 13020 11956 13076
rect 12124 13692 12180 13748
rect 12236 13468 12292 13524
rect 11004 12684 11060 12740
rect 10892 12348 10948 12404
rect 8988 12290 9044 12292
rect 8988 12238 8990 12290
rect 8990 12238 9042 12290
rect 9042 12238 9044 12290
rect 8988 12236 9044 12238
rect 7980 12012 8036 12068
rect 7868 11676 7924 11732
rect 7420 11282 7476 11284
rect 7420 11230 7422 11282
rect 7422 11230 7474 11282
rect 7474 11230 7476 11282
rect 7420 11228 7476 11230
rect 6300 10556 6356 10612
rect 6300 9884 6356 9940
rect 6188 9714 6244 9716
rect 6188 9662 6190 9714
rect 6190 9662 6242 9714
rect 6242 9662 6244 9714
rect 6188 9660 6244 9662
rect 6860 9266 6916 9268
rect 6860 9214 6862 9266
rect 6862 9214 6914 9266
rect 6914 9214 6916 9266
rect 6860 9212 6916 9214
rect 6412 9042 6468 9044
rect 6412 8990 6414 9042
rect 6414 8990 6466 9042
rect 6466 8990 6468 9042
rect 6412 8988 6468 8990
rect 6636 9042 6692 9044
rect 6636 8990 6638 9042
rect 6638 8990 6690 9042
rect 6690 8990 6692 9042
rect 6636 8988 6692 8990
rect 6524 8930 6580 8932
rect 6524 8878 6526 8930
rect 6526 8878 6578 8930
rect 6578 8878 6580 8930
rect 6524 8876 6580 8878
rect 6524 8146 6580 8148
rect 6524 8094 6526 8146
rect 6526 8094 6578 8146
rect 6578 8094 6580 8146
rect 6524 8092 6580 8094
rect 7196 9996 7252 10052
rect 6972 8204 7028 8260
rect 7084 8428 7140 8484
rect 7868 11282 7924 11284
rect 7868 11230 7870 11282
rect 7870 11230 7922 11282
rect 7922 11230 7924 11282
rect 7868 11228 7924 11230
rect 8316 11676 8372 11732
rect 7868 10892 7924 10948
rect 7532 9996 7588 10052
rect 8092 10556 8148 10612
rect 8204 10444 8260 10500
rect 7868 9772 7924 9828
rect 10556 12290 10612 12292
rect 10556 12238 10558 12290
rect 10558 12238 10610 12290
rect 10610 12238 10612 12290
rect 10556 12236 10612 12238
rect 8652 11618 8708 11620
rect 8652 11566 8654 11618
rect 8654 11566 8706 11618
rect 8706 11566 8708 11618
rect 8652 11564 8708 11566
rect 8876 11618 8932 11620
rect 8876 11566 8878 11618
rect 8878 11566 8930 11618
rect 8930 11566 8932 11618
rect 8876 11564 8932 11566
rect 8876 11004 8932 11060
rect 8988 10892 9044 10948
rect 9100 11340 9156 11396
rect 10668 11506 10724 11508
rect 10668 11454 10670 11506
rect 10670 11454 10722 11506
rect 10722 11454 10724 11506
rect 10668 11452 10724 11454
rect 10444 11394 10500 11396
rect 10444 11342 10446 11394
rect 10446 11342 10498 11394
rect 10498 11342 10500 11394
rect 10444 11340 10500 11342
rect 9660 11282 9716 11284
rect 9660 11230 9662 11282
rect 9662 11230 9714 11282
rect 9714 11230 9716 11282
rect 9660 11228 9716 11230
rect 9548 11116 9604 11172
rect 9528 11002 9584 11004
rect 9528 10950 9530 11002
rect 9530 10950 9582 11002
rect 9582 10950 9584 11002
rect 9528 10948 9584 10950
rect 9632 11002 9688 11004
rect 9632 10950 9634 11002
rect 9634 10950 9686 11002
rect 9686 10950 9688 11002
rect 9632 10948 9688 10950
rect 9736 11002 9792 11004
rect 9736 10950 9738 11002
rect 9738 10950 9790 11002
rect 9790 10950 9792 11002
rect 9736 10948 9792 10950
rect 10780 11228 10836 11284
rect 9324 10668 9380 10724
rect 8204 9436 8260 9492
rect 9212 10050 9268 10052
rect 9212 9998 9214 10050
rect 9214 9998 9266 10050
rect 9266 9998 9268 10050
rect 9212 9996 9268 9998
rect 7756 9154 7812 9156
rect 7756 9102 7758 9154
rect 7758 9102 7810 9154
rect 7810 9102 7812 9154
rect 7756 9100 7812 9102
rect 8540 9660 8596 9716
rect 7644 8764 7700 8820
rect 7308 8652 7364 8708
rect 7308 8428 7364 8484
rect 6860 7868 6916 7924
rect 6076 7644 6132 7700
rect 6860 7698 6916 7700
rect 6860 7646 6862 7698
rect 6862 7646 6914 7698
rect 6914 7646 6916 7698
rect 6860 7644 6916 7646
rect 6188 7420 6244 7476
rect 6188 6972 6244 7028
rect 6076 6636 6132 6692
rect 6412 6690 6468 6692
rect 6412 6638 6414 6690
rect 6414 6638 6466 6690
rect 6466 6638 6468 6690
rect 6412 6636 6468 6638
rect 6188 6412 6244 6468
rect 6972 7308 7028 7364
rect 6636 6636 6692 6692
rect 6524 6300 6580 6356
rect 6300 5740 6356 5796
rect 4844 5122 4900 5124
rect 4844 5070 4846 5122
rect 4846 5070 4898 5122
rect 4898 5070 4900 5122
rect 4844 5068 4900 5070
rect 4956 5180 5012 5236
rect 4396 4732 4452 4788
rect 4732 4562 4788 4564
rect 4732 4510 4734 4562
rect 4734 4510 4786 4562
rect 4786 4510 4788 4562
rect 4732 4508 4788 4510
rect 5516 5068 5572 5124
rect 5068 4844 5124 4900
rect 5180 4450 5236 4452
rect 5180 4398 5182 4450
rect 5182 4398 5234 4450
rect 5234 4398 5236 4450
rect 5180 4396 5236 4398
rect 1820 4338 1876 4340
rect 1820 4286 1822 4338
rect 1822 4286 1874 4338
rect 1874 4286 1876 4338
rect 1820 4284 1876 4286
rect 5740 4508 5796 4564
rect 1596 4172 1652 4228
rect 3612 4172 3668 4228
rect 5740 4172 5796 4228
rect 5964 5122 6020 5124
rect 5964 5070 5966 5122
rect 5966 5070 6018 5122
rect 6018 5070 6020 5122
rect 5964 5068 6020 5070
rect 6188 4898 6244 4900
rect 6188 4846 6190 4898
rect 6190 4846 6242 4898
rect 6242 4846 6244 4898
rect 6188 4844 6244 4846
rect 6860 6300 6916 6356
rect 7084 6412 7140 6468
rect 7196 7474 7252 7476
rect 7196 7422 7198 7474
rect 7198 7422 7250 7474
rect 7250 7422 7252 7474
rect 7196 7420 7252 7422
rect 7868 7644 7924 7700
rect 7756 6802 7812 6804
rect 7756 6750 7758 6802
rect 7758 6750 7810 6802
rect 7810 6750 7812 6802
rect 7756 6748 7812 6750
rect 7644 6690 7700 6692
rect 7644 6638 7646 6690
rect 7646 6638 7698 6690
rect 7698 6638 7700 6690
rect 7644 6636 7700 6638
rect 7980 6636 8036 6692
rect 7980 6300 8036 6356
rect 8204 7308 8260 7364
rect 9324 9884 9380 9940
rect 9996 10668 10052 10724
rect 9548 10610 9604 10612
rect 9548 10558 9550 10610
rect 9550 10558 9602 10610
rect 9602 10558 9604 10610
rect 9548 10556 9604 10558
rect 9548 9996 9604 10052
rect 9548 9826 9604 9828
rect 9548 9774 9550 9826
rect 9550 9774 9602 9826
rect 9602 9774 9604 9826
rect 9548 9772 9604 9774
rect 8988 8988 9044 9044
rect 8092 6412 8148 6468
rect 7644 6130 7700 6132
rect 7644 6078 7646 6130
rect 7646 6078 7698 6130
rect 7698 6078 7700 6130
rect 7644 6076 7700 6078
rect 6972 5964 7028 6020
rect 6860 5740 6916 5796
rect 6636 4956 6692 5012
rect 5852 4284 5908 4340
rect 5370 3946 5426 3948
rect 5370 3894 5372 3946
rect 5372 3894 5424 3946
rect 5424 3894 5426 3946
rect 5370 3892 5426 3894
rect 5474 3946 5530 3948
rect 5474 3894 5476 3946
rect 5476 3894 5528 3946
rect 5528 3894 5530 3946
rect 5474 3892 5530 3894
rect 5578 3946 5634 3948
rect 5578 3894 5580 3946
rect 5580 3894 5632 3946
rect 5632 3894 5634 3946
rect 5578 3892 5634 3894
rect 6748 4732 6804 4788
rect 6636 4284 6692 4340
rect 6860 4450 6916 4452
rect 6860 4398 6862 4450
rect 6862 4398 6914 4450
rect 6914 4398 6916 4450
rect 6860 4396 6916 4398
rect 7196 4620 7252 4676
rect 7308 5516 7364 5572
rect 7084 4562 7140 4564
rect 7084 4510 7086 4562
rect 7086 4510 7138 4562
rect 7138 4510 7140 4562
rect 7084 4508 7140 4510
rect 7980 6130 8036 6132
rect 7980 6078 7982 6130
rect 7982 6078 8034 6130
rect 8034 6078 8036 6130
rect 7980 6076 8036 6078
rect 7868 5852 7924 5908
rect 8204 6188 8260 6244
rect 8652 6300 8708 6356
rect 8428 5852 8484 5908
rect 8540 6188 8596 6244
rect 7532 4732 7588 4788
rect 7420 4450 7476 4452
rect 7420 4398 7422 4450
rect 7422 4398 7474 4450
rect 7474 4398 7476 4450
rect 7420 4396 7476 4398
rect 7868 4732 7924 4788
rect 8204 4956 8260 5012
rect 7756 4562 7812 4564
rect 7756 4510 7758 4562
rect 7758 4510 7810 4562
rect 7810 4510 7812 4562
rect 7756 4508 7812 4510
rect 6860 4172 6916 4228
rect 6748 3724 6804 3780
rect 8316 4284 8372 4340
rect 9100 9436 9156 9492
rect 8876 7698 8932 7700
rect 8876 7646 8878 7698
rect 8878 7646 8930 7698
rect 8930 7646 8932 7698
rect 8876 7644 8932 7646
rect 8876 7250 8932 7252
rect 8876 7198 8878 7250
rect 8878 7198 8930 7250
rect 8930 7198 8932 7250
rect 8876 7196 8932 7198
rect 8988 6412 9044 6468
rect 8876 6188 8932 6244
rect 8764 6076 8820 6132
rect 8876 5964 8932 6020
rect 9528 9434 9584 9436
rect 9528 9382 9530 9434
rect 9530 9382 9582 9434
rect 9582 9382 9584 9434
rect 9528 9380 9584 9382
rect 9632 9434 9688 9436
rect 9632 9382 9634 9434
rect 9634 9382 9686 9434
rect 9686 9382 9688 9434
rect 9632 9380 9688 9382
rect 9736 9434 9792 9436
rect 9736 9382 9738 9434
rect 9738 9382 9790 9434
rect 9790 9382 9792 9434
rect 9736 9380 9792 9382
rect 10220 10498 10276 10500
rect 10220 10446 10222 10498
rect 10222 10446 10274 10498
rect 10274 10446 10276 10498
rect 10220 10444 10276 10446
rect 10668 10332 10724 10388
rect 9884 9324 9940 9380
rect 11116 11564 11172 11620
rect 11116 10108 11172 10164
rect 10668 9884 10724 9940
rect 10444 9660 10500 9716
rect 9660 9212 9716 9268
rect 9548 8764 9604 8820
rect 10108 8988 10164 9044
rect 9884 8316 9940 8372
rect 9772 8092 9828 8148
rect 11340 12738 11396 12740
rect 11340 12686 11342 12738
rect 11342 12686 11394 12738
rect 11394 12686 11396 12738
rect 11340 12684 11396 12686
rect 12012 12738 12068 12740
rect 12012 12686 12014 12738
rect 12014 12686 12066 12738
rect 12066 12686 12068 12738
rect 12012 12684 12068 12686
rect 11228 9884 11284 9940
rect 11340 11676 11396 11732
rect 10780 9660 10836 9716
rect 10556 8428 10612 8484
rect 10108 7980 10164 8036
rect 9528 7866 9584 7868
rect 9528 7814 9530 7866
rect 9530 7814 9582 7866
rect 9582 7814 9584 7866
rect 9528 7812 9584 7814
rect 9632 7866 9688 7868
rect 9632 7814 9634 7866
rect 9634 7814 9686 7866
rect 9686 7814 9688 7866
rect 9632 7812 9688 7814
rect 9736 7866 9792 7868
rect 9736 7814 9738 7866
rect 9738 7814 9790 7866
rect 9790 7814 9792 7866
rect 9736 7812 9792 7814
rect 9996 7644 10052 7700
rect 9212 7196 9268 7252
rect 10668 9212 10724 9268
rect 10332 7532 10388 7588
rect 11452 9996 11508 10052
rect 11900 9884 11956 9940
rect 11452 9212 11508 9268
rect 11788 9660 11844 9716
rect 11340 8316 11396 8372
rect 11452 8764 11508 8820
rect 11004 7532 11060 7588
rect 10220 7196 10276 7252
rect 9660 6748 9716 6804
rect 9884 6972 9940 7028
rect 9212 5964 9268 6020
rect 9528 6298 9584 6300
rect 9528 6246 9530 6298
rect 9530 6246 9582 6298
rect 9582 6246 9584 6298
rect 9528 6244 9584 6246
rect 9632 6298 9688 6300
rect 9632 6246 9634 6298
rect 9634 6246 9686 6298
rect 9686 6246 9688 6298
rect 9632 6244 9688 6246
rect 9736 6298 9792 6300
rect 9736 6246 9738 6298
rect 9738 6246 9790 6298
rect 9790 6246 9792 6298
rect 9736 6244 9792 6246
rect 9436 5852 9492 5908
rect 9324 5628 9380 5684
rect 8652 5292 8708 5348
rect 8876 5180 8932 5236
rect 8652 4844 8708 4900
rect 8988 4732 9044 4788
rect 8652 4450 8708 4452
rect 8652 4398 8654 4450
rect 8654 4398 8706 4450
rect 8706 4398 8708 4450
rect 8652 4396 8708 4398
rect 9436 5010 9492 5012
rect 9436 4958 9438 5010
rect 9438 4958 9490 5010
rect 9490 4958 9492 5010
rect 9436 4956 9492 4958
rect 10892 7196 10948 7252
rect 10220 6076 10276 6132
rect 10780 5292 10836 5348
rect 10892 5234 10948 5236
rect 10892 5182 10894 5234
rect 10894 5182 10946 5234
rect 10946 5182 10948 5234
rect 10892 5180 10948 5182
rect 12572 12962 12628 12964
rect 12572 12910 12574 12962
rect 12574 12910 12626 12962
rect 12626 12910 12628 12962
rect 12572 12908 12628 12910
rect 14812 15820 14868 15876
rect 14700 15426 14756 15428
rect 14700 15374 14702 15426
rect 14702 15374 14754 15426
rect 14754 15374 14756 15426
rect 14700 15372 14756 15374
rect 14028 15260 14084 15316
rect 13686 14922 13742 14924
rect 13686 14870 13688 14922
rect 13688 14870 13740 14922
rect 13740 14870 13742 14922
rect 13686 14868 13742 14870
rect 13790 14922 13846 14924
rect 13790 14870 13792 14922
rect 13792 14870 13844 14922
rect 13844 14870 13846 14922
rect 13790 14868 13846 14870
rect 13894 14922 13950 14924
rect 13894 14870 13896 14922
rect 13896 14870 13948 14922
rect 13948 14870 13950 14922
rect 13894 14868 13950 14870
rect 13580 14306 13636 14308
rect 13580 14254 13582 14306
rect 13582 14254 13634 14306
rect 13634 14254 13636 14306
rect 13580 14252 13636 14254
rect 13686 13354 13742 13356
rect 13686 13302 13688 13354
rect 13688 13302 13740 13354
rect 13740 13302 13742 13354
rect 13686 13300 13742 13302
rect 13790 13354 13846 13356
rect 13790 13302 13792 13354
rect 13792 13302 13844 13354
rect 13844 13302 13846 13354
rect 13790 13300 13846 13302
rect 13894 13354 13950 13356
rect 13894 13302 13896 13354
rect 13896 13302 13948 13354
rect 13948 13302 13950 13354
rect 13894 13300 13950 13302
rect 13804 12850 13860 12852
rect 13804 12798 13806 12850
rect 13806 12798 13858 12850
rect 13858 12798 13860 12850
rect 13804 12796 13860 12798
rect 14140 12850 14196 12852
rect 14140 12798 14142 12850
rect 14142 12798 14194 12850
rect 14194 12798 14196 12850
rect 14140 12796 14196 12798
rect 16828 18508 16884 18564
rect 16044 18284 16100 18340
rect 16492 18284 16548 18340
rect 15932 16994 15988 16996
rect 15932 16942 15934 16994
rect 15934 16942 15986 16994
rect 15986 16942 15988 16994
rect 15932 16940 15988 16942
rect 15260 16828 15316 16884
rect 15260 16658 15316 16660
rect 15260 16606 15262 16658
rect 15262 16606 15314 16658
rect 15314 16606 15316 16658
rect 15260 16604 15316 16606
rect 15260 16044 15316 16100
rect 15148 15986 15204 15988
rect 15148 15934 15150 15986
rect 15150 15934 15202 15986
rect 15202 15934 15204 15986
rect 15148 15932 15204 15934
rect 15148 15708 15204 15764
rect 16156 17500 16212 17556
rect 16716 16994 16772 16996
rect 16716 16942 16718 16994
rect 16718 16942 16770 16994
rect 16770 16942 16772 16994
rect 16716 16940 16772 16942
rect 15484 15820 15540 15876
rect 15260 15314 15316 15316
rect 15260 15262 15262 15314
rect 15262 15262 15314 15314
rect 15314 15262 15316 15314
rect 15260 15260 15316 15262
rect 15708 15708 15764 15764
rect 15596 15372 15652 15428
rect 14924 12796 14980 12852
rect 15596 14140 15652 14196
rect 16492 16604 16548 16660
rect 15932 16380 15988 16436
rect 16044 15986 16100 15988
rect 16044 15934 16046 15986
rect 16046 15934 16098 15986
rect 16098 15934 16100 15986
rect 16044 15932 16100 15934
rect 16380 15932 16436 15988
rect 17724 20690 17780 20692
rect 17724 20638 17726 20690
rect 17726 20638 17778 20690
rect 17778 20638 17780 20690
rect 17724 20636 17780 20638
rect 17388 19346 17444 19348
rect 17388 19294 17390 19346
rect 17390 19294 17442 19346
rect 17442 19294 17444 19346
rect 17388 19292 17444 19294
rect 17500 18508 17556 18564
rect 17500 18338 17556 18340
rect 17500 18286 17502 18338
rect 17502 18286 17554 18338
rect 17554 18286 17556 18338
rect 17500 18284 17556 18286
rect 17836 20524 17892 20580
rect 17844 20410 17900 20412
rect 17844 20358 17846 20410
rect 17846 20358 17898 20410
rect 17898 20358 17900 20410
rect 17844 20356 17900 20358
rect 17948 20410 18004 20412
rect 17948 20358 17950 20410
rect 17950 20358 18002 20410
rect 18002 20358 18004 20410
rect 17948 20356 18004 20358
rect 18052 20410 18108 20412
rect 18052 20358 18054 20410
rect 18054 20358 18106 20410
rect 18106 20358 18108 20410
rect 18052 20356 18108 20358
rect 18172 20018 18228 20020
rect 18172 19966 18174 20018
rect 18174 19966 18226 20018
rect 18226 19966 18228 20018
rect 18172 19964 18228 19966
rect 17948 19740 18004 19796
rect 18060 19628 18116 19684
rect 17844 18842 17900 18844
rect 17844 18790 17846 18842
rect 17846 18790 17898 18842
rect 17898 18790 17900 18842
rect 17844 18788 17900 18790
rect 17948 18842 18004 18844
rect 17948 18790 17950 18842
rect 17950 18790 18002 18842
rect 18002 18790 18004 18842
rect 17948 18788 18004 18790
rect 18052 18842 18108 18844
rect 18052 18790 18054 18842
rect 18054 18790 18106 18842
rect 18106 18790 18108 18842
rect 18052 18788 18108 18790
rect 18060 18172 18116 18228
rect 17164 17500 17220 17556
rect 17164 17276 17220 17332
rect 17052 17052 17108 17108
rect 16716 16658 16772 16660
rect 16716 16606 16718 16658
rect 16718 16606 16770 16658
rect 16770 16606 16772 16658
rect 16716 16604 16772 16606
rect 17052 16268 17108 16324
rect 15820 14588 15876 14644
rect 16156 14700 16212 14756
rect 16716 15932 16772 15988
rect 16940 15986 16996 15988
rect 16940 15934 16942 15986
rect 16942 15934 16994 15986
rect 16994 15934 16996 15986
rect 16940 15932 16996 15934
rect 17836 17500 17892 17556
rect 18172 17500 18228 17556
rect 17724 17442 17780 17444
rect 17724 17390 17726 17442
rect 17726 17390 17778 17442
rect 17778 17390 17780 17442
rect 17724 17388 17780 17390
rect 17612 17276 17668 17332
rect 17844 17274 17900 17276
rect 17844 17222 17846 17274
rect 17846 17222 17898 17274
rect 17898 17222 17900 17274
rect 17844 17220 17900 17222
rect 17948 17274 18004 17276
rect 17948 17222 17950 17274
rect 17950 17222 18002 17274
rect 18002 17222 18004 17274
rect 17948 17220 18004 17222
rect 18052 17274 18108 17276
rect 18052 17222 18054 17274
rect 18054 17222 18106 17274
rect 18106 17222 18108 17274
rect 18052 17220 18108 17222
rect 17948 17052 18004 17108
rect 17276 16828 17332 16884
rect 17612 16716 17668 16772
rect 17836 16940 17892 16996
rect 18956 23212 19012 23268
rect 18732 22988 18788 23044
rect 18396 21756 18452 21812
rect 18732 21980 18788 22036
rect 18844 23100 18900 23156
rect 20300 27858 20356 27860
rect 20300 27806 20302 27858
rect 20302 27806 20354 27858
rect 20354 27806 20356 27858
rect 20300 27804 20356 27806
rect 19516 23154 19572 23156
rect 19516 23102 19518 23154
rect 19518 23102 19570 23154
rect 19570 23102 19572 23154
rect 19516 23100 19572 23102
rect 19740 26290 19796 26292
rect 19740 26238 19742 26290
rect 19742 26238 19794 26290
rect 19794 26238 19796 26290
rect 19740 26236 19796 26238
rect 20300 26348 20356 26404
rect 22002 27466 22058 27468
rect 22002 27414 22004 27466
rect 22004 27414 22056 27466
rect 22056 27414 22058 27466
rect 22002 27412 22058 27414
rect 22106 27466 22162 27468
rect 22106 27414 22108 27466
rect 22108 27414 22160 27466
rect 22160 27414 22162 27466
rect 22106 27412 22162 27414
rect 22210 27466 22266 27468
rect 22210 27414 22212 27466
rect 22212 27414 22264 27466
rect 22264 27414 22266 27466
rect 22210 27412 22266 27414
rect 30318 27466 30374 27468
rect 30318 27414 30320 27466
rect 30320 27414 30372 27466
rect 30372 27414 30374 27466
rect 30318 27412 30374 27414
rect 30422 27466 30478 27468
rect 30422 27414 30424 27466
rect 30424 27414 30476 27466
rect 30476 27414 30478 27466
rect 30422 27412 30478 27414
rect 30526 27466 30582 27468
rect 30526 27414 30528 27466
rect 30528 27414 30580 27466
rect 30580 27414 30582 27466
rect 30526 27412 30582 27414
rect 20636 27132 20692 27188
rect 20636 26962 20692 26964
rect 20636 26910 20638 26962
rect 20638 26910 20690 26962
rect 20690 26910 20692 26962
rect 20636 26908 20692 26910
rect 20300 25676 20356 25732
rect 20524 25564 20580 25620
rect 19852 25506 19908 25508
rect 19852 25454 19854 25506
rect 19854 25454 19906 25506
rect 19906 25454 19908 25506
rect 19852 25452 19908 25454
rect 20076 25506 20132 25508
rect 20076 25454 20078 25506
rect 20078 25454 20130 25506
rect 20130 25454 20132 25506
rect 20076 25452 20132 25454
rect 26160 26682 26216 26684
rect 26160 26630 26162 26682
rect 26162 26630 26214 26682
rect 26214 26630 26216 26682
rect 26160 26628 26216 26630
rect 26264 26682 26320 26684
rect 26264 26630 26266 26682
rect 26266 26630 26318 26682
rect 26318 26630 26320 26682
rect 26264 26628 26320 26630
rect 26368 26682 26424 26684
rect 26368 26630 26370 26682
rect 26370 26630 26422 26682
rect 26422 26630 26424 26682
rect 26368 26628 26424 26630
rect 34476 26682 34532 26684
rect 34476 26630 34478 26682
rect 34478 26630 34530 26682
rect 34530 26630 34532 26682
rect 34476 26628 34532 26630
rect 34580 26682 34636 26684
rect 34580 26630 34582 26682
rect 34582 26630 34634 26682
rect 34634 26630 34636 26682
rect 34580 26628 34636 26630
rect 34684 26682 34740 26684
rect 34684 26630 34686 26682
rect 34686 26630 34738 26682
rect 34738 26630 34740 26682
rect 34684 26628 34740 26630
rect 22002 25898 22058 25900
rect 22002 25846 22004 25898
rect 22004 25846 22056 25898
rect 22056 25846 22058 25898
rect 22002 25844 22058 25846
rect 22106 25898 22162 25900
rect 22106 25846 22108 25898
rect 22108 25846 22160 25898
rect 22160 25846 22162 25898
rect 22106 25844 22162 25846
rect 22210 25898 22266 25900
rect 22210 25846 22212 25898
rect 22212 25846 22264 25898
rect 22264 25846 22266 25898
rect 22210 25844 22266 25846
rect 21980 25564 22036 25620
rect 20748 25452 20804 25508
rect 21644 25506 21700 25508
rect 21644 25454 21646 25506
rect 21646 25454 21698 25506
rect 21698 25454 21700 25506
rect 21644 25452 21700 25454
rect 20860 25340 20916 25396
rect 21756 25340 21812 25396
rect 20188 24556 20244 24612
rect 19740 23100 19796 23156
rect 19516 22876 19572 22932
rect 20300 23266 20356 23268
rect 20300 23214 20302 23266
rect 20302 23214 20354 23266
rect 20354 23214 20356 23266
rect 20300 23212 20356 23214
rect 19292 21980 19348 22036
rect 19628 21644 19684 21700
rect 18396 19852 18452 19908
rect 18508 19628 18564 19684
rect 18396 19346 18452 19348
rect 18396 19294 18398 19346
rect 18398 19294 18450 19346
rect 18450 19294 18452 19346
rect 18396 19292 18452 19294
rect 19068 20018 19124 20020
rect 19068 19966 19070 20018
rect 19070 19966 19122 20018
rect 19122 19966 19124 20018
rect 19068 19964 19124 19966
rect 18844 19740 18900 19796
rect 19740 21308 19796 21364
rect 19516 19964 19572 20020
rect 20300 22370 20356 22372
rect 20300 22318 20302 22370
rect 20302 22318 20354 22370
rect 20354 22318 20356 22370
rect 20300 22316 20356 22318
rect 19964 22092 20020 22148
rect 19964 21810 20020 21812
rect 19964 21758 19966 21810
rect 19966 21758 20018 21810
rect 20018 21758 20020 21810
rect 19964 21756 20020 21758
rect 20300 21308 20356 21364
rect 20300 20018 20356 20020
rect 20300 19966 20302 20018
rect 20302 19966 20354 20018
rect 20354 19966 20356 20018
rect 20300 19964 20356 19966
rect 18844 18620 18900 18676
rect 18732 18450 18788 18452
rect 18732 18398 18734 18450
rect 18734 18398 18786 18450
rect 18786 18398 18788 18450
rect 18732 18396 18788 18398
rect 18956 17554 19012 17556
rect 18956 17502 18958 17554
rect 18958 17502 19010 17554
rect 19010 17502 19012 17554
rect 18956 17500 19012 17502
rect 18396 17442 18452 17444
rect 18396 17390 18398 17442
rect 18398 17390 18450 17442
rect 18450 17390 18452 17442
rect 18396 17388 18452 17390
rect 19068 17442 19124 17444
rect 19068 17390 19070 17442
rect 19070 17390 19122 17442
rect 19122 17390 19124 17442
rect 19068 17388 19124 17390
rect 18508 16770 18564 16772
rect 18508 16718 18510 16770
rect 18510 16718 18562 16770
rect 18562 16718 18564 16770
rect 18508 16716 18564 16718
rect 19068 16604 19124 16660
rect 17948 16322 18004 16324
rect 17948 16270 17950 16322
rect 17950 16270 18002 16322
rect 18002 16270 18004 16322
rect 17948 16268 18004 16270
rect 16828 15708 16884 15764
rect 16604 14700 16660 14756
rect 17276 15036 17332 15092
rect 16380 14476 16436 14532
rect 16492 14642 16548 14644
rect 16492 14590 16494 14642
rect 16494 14590 16546 14642
rect 16546 14590 16548 14642
rect 16492 14588 16548 14590
rect 15820 14140 15876 14196
rect 13686 11786 13742 11788
rect 13686 11734 13688 11786
rect 13688 11734 13740 11786
rect 13740 11734 13742 11786
rect 13686 11732 13742 11734
rect 13790 11786 13846 11788
rect 13790 11734 13792 11786
rect 13792 11734 13844 11786
rect 13844 11734 13846 11786
rect 13790 11732 13846 11734
rect 13894 11786 13950 11788
rect 13894 11734 13896 11786
rect 13896 11734 13948 11786
rect 13948 11734 13950 11786
rect 13894 11732 13950 11734
rect 14252 11506 14308 11508
rect 14252 11454 14254 11506
rect 14254 11454 14306 11506
rect 14306 11454 14308 11506
rect 14252 11452 14308 11454
rect 13020 11228 13076 11284
rect 12348 10332 12404 10388
rect 17052 14530 17108 14532
rect 17052 14478 17054 14530
rect 17054 14478 17106 14530
rect 17106 14478 17108 14530
rect 17052 14476 17108 14478
rect 17388 14530 17444 14532
rect 17388 14478 17390 14530
rect 17390 14478 17442 14530
rect 17442 14478 17444 14530
rect 17388 14476 17444 14478
rect 16492 13804 16548 13860
rect 17276 14252 17332 14308
rect 15372 13074 15428 13076
rect 15372 13022 15374 13074
rect 15374 13022 15426 13074
rect 15426 13022 15428 13074
rect 15372 13020 15428 13022
rect 17388 14140 17444 14196
rect 16380 13020 16436 13076
rect 18284 15874 18340 15876
rect 18284 15822 18286 15874
rect 18286 15822 18338 15874
rect 18338 15822 18340 15874
rect 18284 15820 18340 15822
rect 17844 15706 17900 15708
rect 17844 15654 17846 15706
rect 17846 15654 17898 15706
rect 17898 15654 17900 15706
rect 17844 15652 17900 15654
rect 17948 15706 18004 15708
rect 17948 15654 17950 15706
rect 17950 15654 18002 15706
rect 18002 15654 18004 15706
rect 17948 15652 18004 15654
rect 18052 15706 18108 15708
rect 18052 15654 18054 15706
rect 18054 15654 18106 15706
rect 18106 15654 18108 15706
rect 18052 15652 18108 15654
rect 17836 15260 17892 15316
rect 17948 15148 18004 15204
rect 18620 16044 18676 16100
rect 18508 15986 18564 15988
rect 18508 15934 18510 15986
rect 18510 15934 18562 15986
rect 18562 15934 18564 15986
rect 18508 15932 18564 15934
rect 17844 14138 17900 14140
rect 17844 14086 17846 14138
rect 17846 14086 17898 14138
rect 17898 14086 17900 14138
rect 17844 14084 17900 14086
rect 17948 14138 18004 14140
rect 17948 14086 17950 14138
rect 17950 14086 18002 14138
rect 18002 14086 18004 14138
rect 17948 14084 18004 14086
rect 18052 14138 18108 14140
rect 18052 14086 18054 14138
rect 18054 14086 18106 14138
rect 18106 14086 18108 14138
rect 18052 14084 18108 14086
rect 17724 13746 17780 13748
rect 17724 13694 17726 13746
rect 17726 13694 17778 13746
rect 17778 13694 17780 13746
rect 17724 13692 17780 13694
rect 16492 10780 16548 10836
rect 13468 10332 13524 10388
rect 14924 10332 14980 10388
rect 13686 10218 13742 10220
rect 13686 10166 13688 10218
rect 13688 10166 13740 10218
rect 13740 10166 13742 10218
rect 13686 10164 13742 10166
rect 13790 10218 13846 10220
rect 13790 10166 13792 10218
rect 13792 10166 13844 10218
rect 13844 10166 13846 10218
rect 13790 10164 13846 10166
rect 13894 10218 13950 10220
rect 13894 10166 13896 10218
rect 13896 10166 13948 10218
rect 13948 10166 13950 10218
rect 13894 10164 13950 10166
rect 12236 9884 12292 9940
rect 12012 9602 12068 9604
rect 12012 9550 12014 9602
rect 12014 9550 12066 9602
rect 12066 9550 12068 9602
rect 12012 9548 12068 9550
rect 12348 9548 12404 9604
rect 11900 8764 11956 8820
rect 12236 8652 12292 8708
rect 11788 8540 11844 8596
rect 12236 8146 12292 8148
rect 12236 8094 12238 8146
rect 12238 8094 12290 8146
rect 12290 8094 12292 8146
rect 12236 8092 12292 8094
rect 14476 9938 14532 9940
rect 14476 9886 14478 9938
rect 14478 9886 14530 9938
rect 14530 9886 14532 9938
rect 14476 9884 14532 9886
rect 12908 9826 12964 9828
rect 12908 9774 12910 9826
rect 12910 9774 12962 9826
rect 12962 9774 12964 9826
rect 12908 9772 12964 9774
rect 13580 9602 13636 9604
rect 13580 9550 13582 9602
rect 13582 9550 13634 9602
rect 13634 9550 13636 9602
rect 13580 9548 13636 9550
rect 13804 9660 13860 9716
rect 14028 9548 14084 9604
rect 12572 9436 12628 9492
rect 12572 8482 12628 8484
rect 12572 8430 12574 8482
rect 12574 8430 12626 8482
rect 12626 8430 12628 8482
rect 12572 8428 12628 8430
rect 13692 9436 13748 9492
rect 12908 8652 12964 8708
rect 12908 8428 12964 8484
rect 12796 8370 12852 8372
rect 12796 8318 12798 8370
rect 12798 8318 12850 8370
rect 12850 8318 12852 8370
rect 12796 8316 12852 8318
rect 12684 8092 12740 8148
rect 11228 7308 11284 7364
rect 9528 4730 9584 4732
rect 9528 4678 9530 4730
rect 9530 4678 9582 4730
rect 9582 4678 9584 4730
rect 9528 4676 9584 4678
rect 9632 4730 9688 4732
rect 9632 4678 9634 4730
rect 9634 4678 9686 4730
rect 9686 4678 9688 4730
rect 9632 4676 9688 4678
rect 9736 4730 9792 4732
rect 9736 4678 9738 4730
rect 9738 4678 9790 4730
rect 9790 4678 9792 4730
rect 9736 4676 9792 4678
rect 9100 4508 9156 4564
rect 9772 4508 9828 4564
rect 11340 4562 11396 4564
rect 11340 4510 11342 4562
rect 11342 4510 11394 4562
rect 11394 4510 11396 4562
rect 11340 4508 11396 4510
rect 11676 7474 11732 7476
rect 11676 7422 11678 7474
rect 11678 7422 11730 7474
rect 11730 7422 11732 7474
rect 11676 7420 11732 7422
rect 11564 6466 11620 6468
rect 11564 6414 11566 6466
rect 11566 6414 11618 6466
rect 11618 6414 11620 6466
rect 11564 6412 11620 6414
rect 12012 7474 12068 7476
rect 12012 7422 12014 7474
rect 12014 7422 12066 7474
rect 12066 7422 12068 7474
rect 12012 7420 12068 7422
rect 12796 7250 12852 7252
rect 12796 7198 12798 7250
rect 12798 7198 12850 7250
rect 12850 7198 12852 7250
rect 12796 7196 12852 7198
rect 12012 6860 12068 6916
rect 12572 6860 12628 6916
rect 12460 6748 12516 6804
rect 11900 5740 11956 5796
rect 11788 5122 11844 5124
rect 11788 5070 11790 5122
rect 11790 5070 11842 5122
rect 11842 5070 11844 5122
rect 11788 5068 11844 5070
rect 11564 4844 11620 4900
rect 12124 5292 12180 5348
rect 12124 4508 12180 4564
rect 11452 4396 11508 4452
rect 8988 3612 9044 3668
rect 10220 3666 10276 3668
rect 10220 3614 10222 3666
rect 10222 3614 10274 3666
rect 10274 3614 10276 3666
rect 10220 3612 10276 3614
rect 9548 3554 9604 3556
rect 9548 3502 9550 3554
rect 9550 3502 9602 3554
rect 9602 3502 9604 3554
rect 9548 3500 9604 3502
rect 9528 3162 9584 3164
rect 9528 3110 9530 3162
rect 9530 3110 9582 3162
rect 9582 3110 9584 3162
rect 9528 3108 9584 3110
rect 9632 3162 9688 3164
rect 9632 3110 9634 3162
rect 9634 3110 9686 3162
rect 9686 3110 9688 3162
rect 9632 3108 9688 3110
rect 9736 3162 9792 3164
rect 9736 3110 9738 3162
rect 9738 3110 9790 3162
rect 9790 3110 9792 3162
rect 9736 3108 9792 3110
rect 12908 6860 12964 6916
rect 12684 6524 12740 6580
rect 13132 7980 13188 8036
rect 13356 8764 13412 8820
rect 13686 8650 13742 8652
rect 13686 8598 13688 8650
rect 13688 8598 13740 8650
rect 13740 8598 13742 8650
rect 13686 8596 13742 8598
rect 13790 8650 13846 8652
rect 13790 8598 13792 8650
rect 13792 8598 13844 8650
rect 13844 8598 13846 8650
rect 13790 8596 13846 8598
rect 13894 8650 13950 8652
rect 13894 8598 13896 8650
rect 13896 8598 13948 8650
rect 13948 8598 13950 8650
rect 13894 8596 13950 8598
rect 13244 7644 13300 7700
rect 14140 7980 14196 8036
rect 14140 7532 14196 7588
rect 13132 6524 13188 6580
rect 13020 6188 13076 6244
rect 14364 7644 14420 7700
rect 13916 7362 13972 7364
rect 13916 7310 13918 7362
rect 13918 7310 13970 7362
rect 13970 7310 13972 7362
rect 13916 7308 13972 7310
rect 13686 7082 13742 7084
rect 13686 7030 13688 7082
rect 13688 7030 13740 7082
rect 13740 7030 13742 7082
rect 13686 7028 13742 7030
rect 13790 7082 13846 7084
rect 13790 7030 13792 7082
rect 13792 7030 13844 7082
rect 13844 7030 13846 7082
rect 13790 7028 13846 7030
rect 13894 7082 13950 7084
rect 13894 7030 13896 7082
rect 13896 7030 13948 7082
rect 13948 7030 13950 7082
rect 13894 7028 13950 7030
rect 14364 6748 14420 6804
rect 13356 6690 13412 6692
rect 13356 6638 13358 6690
rect 13358 6638 13410 6690
rect 13410 6638 13412 6690
rect 13356 6636 13412 6638
rect 13804 6578 13860 6580
rect 13804 6526 13806 6578
rect 13806 6526 13858 6578
rect 13858 6526 13860 6578
rect 13804 6524 13860 6526
rect 13244 6412 13300 6468
rect 13692 6130 13748 6132
rect 13692 6078 13694 6130
rect 13694 6078 13746 6130
rect 13746 6078 13748 6130
rect 13692 6076 13748 6078
rect 14252 6188 14308 6244
rect 12684 5068 12740 5124
rect 13686 5514 13742 5516
rect 13686 5462 13688 5514
rect 13688 5462 13740 5514
rect 13740 5462 13742 5514
rect 13686 5460 13742 5462
rect 13790 5514 13846 5516
rect 13790 5462 13792 5514
rect 13792 5462 13844 5514
rect 13844 5462 13846 5514
rect 13790 5460 13846 5462
rect 13894 5514 13950 5516
rect 13894 5462 13896 5514
rect 13896 5462 13948 5514
rect 13948 5462 13950 5514
rect 13894 5460 13950 5462
rect 13580 5346 13636 5348
rect 13580 5294 13582 5346
rect 13582 5294 13634 5346
rect 13634 5294 13636 5346
rect 13580 5292 13636 5294
rect 13244 5068 13300 5124
rect 13916 5122 13972 5124
rect 13916 5070 13918 5122
rect 13918 5070 13970 5122
rect 13970 5070 13972 5122
rect 13916 5068 13972 5070
rect 15036 9660 15092 9716
rect 15036 9042 15092 9044
rect 15036 8990 15038 9042
rect 15038 8990 15090 9042
rect 15090 8990 15092 9042
rect 15036 8988 15092 8990
rect 14924 8146 14980 8148
rect 14924 8094 14926 8146
rect 14926 8094 14978 8146
rect 14978 8094 14980 8146
rect 14924 8092 14980 8094
rect 14588 6690 14644 6692
rect 14588 6638 14590 6690
rect 14590 6638 14642 6690
rect 14642 6638 14644 6690
rect 14588 6636 14644 6638
rect 15372 8428 15428 8484
rect 16604 10610 16660 10612
rect 16604 10558 16606 10610
rect 16606 10558 16658 10610
rect 16658 10558 16660 10610
rect 16604 10556 16660 10558
rect 16268 10108 16324 10164
rect 16268 9154 16324 9156
rect 16268 9102 16270 9154
rect 16270 9102 16322 9154
rect 16322 9102 16324 9154
rect 16268 9100 16324 9102
rect 16268 8316 16324 8372
rect 16492 8204 16548 8260
rect 15708 7532 15764 7588
rect 15484 7474 15540 7476
rect 15484 7422 15486 7474
rect 15486 7422 15538 7474
rect 15538 7422 15540 7474
rect 15484 7420 15540 7422
rect 15260 7084 15316 7140
rect 14476 5852 14532 5908
rect 14588 5794 14644 5796
rect 14588 5742 14590 5794
rect 14590 5742 14642 5794
rect 14642 5742 14644 5794
rect 14588 5740 14644 5742
rect 14588 5292 14644 5348
rect 14028 5010 14084 5012
rect 14028 4958 14030 5010
rect 14030 4958 14082 5010
rect 14082 4958 14084 5010
rect 14028 4956 14084 4958
rect 13468 4508 13524 4564
rect 13356 4450 13412 4452
rect 13356 4398 13358 4450
rect 13358 4398 13410 4450
rect 13410 4398 13412 4450
rect 13356 4396 13412 4398
rect 12572 4338 12628 4340
rect 12572 4286 12574 4338
rect 12574 4286 12626 4338
rect 12626 4286 12628 4338
rect 12572 4284 12628 4286
rect 15596 5852 15652 5908
rect 15484 5516 15540 5572
rect 15036 4284 15092 4340
rect 15260 4956 15316 5012
rect 14140 4172 14196 4228
rect 13686 3946 13742 3948
rect 13686 3894 13688 3946
rect 13688 3894 13740 3946
rect 13740 3894 13742 3946
rect 13686 3892 13742 3894
rect 13790 3946 13846 3948
rect 13790 3894 13792 3946
rect 13792 3894 13844 3946
rect 13844 3894 13846 3946
rect 13790 3892 13846 3894
rect 13894 3946 13950 3948
rect 13894 3894 13896 3946
rect 13896 3894 13948 3946
rect 13948 3894 13950 3946
rect 13894 3892 13950 3894
rect 14924 3778 14980 3780
rect 14924 3726 14926 3778
rect 14926 3726 14978 3778
rect 14978 3726 14980 3778
rect 14924 3724 14980 3726
rect 16044 7532 16100 7588
rect 16156 7308 16212 7364
rect 16044 5292 16100 5348
rect 16044 4844 16100 4900
rect 17612 12236 17668 12292
rect 17388 11116 17444 11172
rect 17388 10834 17444 10836
rect 17388 10782 17390 10834
rect 17390 10782 17442 10834
rect 17442 10782 17444 10834
rect 17388 10780 17444 10782
rect 17948 13804 18004 13860
rect 18396 13970 18452 13972
rect 18396 13918 18398 13970
rect 18398 13918 18450 13970
rect 18450 13918 18452 13970
rect 18396 13916 18452 13918
rect 18172 13804 18228 13860
rect 17948 12908 18004 12964
rect 18844 15874 18900 15876
rect 18844 15822 18846 15874
rect 18846 15822 18898 15874
rect 18898 15822 18900 15874
rect 18844 15820 18900 15822
rect 19964 19292 20020 19348
rect 22652 25452 22708 25508
rect 22876 25676 22932 25732
rect 22540 25340 22596 25396
rect 22764 24892 22820 24948
rect 23100 25618 23156 25620
rect 23100 25566 23102 25618
rect 23102 25566 23154 25618
rect 23154 25566 23156 25618
rect 23100 25564 23156 25566
rect 22988 25228 23044 25284
rect 23548 25340 23604 25396
rect 23212 24892 23268 24948
rect 23100 24668 23156 24724
rect 21980 24444 22036 24500
rect 22002 24330 22058 24332
rect 22002 24278 22004 24330
rect 22004 24278 22056 24330
rect 22056 24278 22058 24330
rect 22002 24276 22058 24278
rect 22106 24330 22162 24332
rect 22106 24278 22108 24330
rect 22108 24278 22160 24330
rect 22160 24278 22162 24330
rect 22106 24276 22162 24278
rect 22210 24330 22266 24332
rect 22210 24278 22212 24330
rect 22212 24278 22264 24330
rect 22264 24278 22266 24330
rect 22210 24276 22266 24278
rect 21084 22316 21140 22372
rect 20636 22258 20692 22260
rect 20636 22206 20638 22258
rect 20638 22206 20690 22258
rect 20690 22206 20692 22258
rect 20636 22204 20692 22206
rect 20636 21698 20692 21700
rect 20636 21646 20638 21698
rect 20638 21646 20690 21698
rect 20690 21646 20692 21698
rect 20636 21644 20692 21646
rect 20524 21532 20580 21588
rect 21308 21868 21364 21924
rect 23212 24444 23268 24500
rect 22002 22762 22058 22764
rect 22002 22710 22004 22762
rect 22004 22710 22056 22762
rect 22056 22710 22058 22762
rect 22002 22708 22058 22710
rect 22106 22762 22162 22764
rect 22106 22710 22108 22762
rect 22108 22710 22160 22762
rect 22160 22710 22162 22762
rect 22106 22708 22162 22710
rect 22210 22762 22266 22764
rect 22210 22710 22212 22762
rect 22212 22710 22264 22762
rect 22264 22710 22266 22762
rect 22210 22708 22266 22710
rect 22092 22258 22148 22260
rect 22092 22206 22094 22258
rect 22094 22206 22146 22258
rect 22146 22206 22148 22258
rect 22092 22204 22148 22206
rect 21980 21868 22036 21924
rect 21756 21698 21812 21700
rect 21756 21646 21758 21698
rect 21758 21646 21810 21698
rect 21810 21646 21812 21698
rect 21756 21644 21812 21646
rect 20860 21420 20916 21476
rect 21756 21420 21812 21476
rect 22876 21756 22932 21812
rect 22092 21644 22148 21700
rect 22540 21698 22596 21700
rect 22540 21646 22542 21698
rect 22542 21646 22594 21698
rect 22594 21646 22596 21698
rect 22540 21644 22596 21646
rect 22428 21586 22484 21588
rect 22428 21534 22430 21586
rect 22430 21534 22482 21586
rect 22482 21534 22484 21586
rect 22428 21532 22484 21534
rect 21308 20636 21364 20692
rect 22652 21308 22708 21364
rect 22002 21194 22058 21196
rect 22002 21142 22004 21194
rect 22004 21142 22056 21194
rect 22056 21142 22058 21194
rect 22002 21140 22058 21142
rect 22106 21194 22162 21196
rect 22106 21142 22108 21194
rect 22108 21142 22160 21194
rect 22160 21142 22162 21194
rect 22106 21140 22162 21142
rect 22210 21194 22266 21196
rect 22210 21142 22212 21194
rect 22212 21142 22264 21194
rect 22264 21142 22266 21194
rect 22210 21140 22266 21142
rect 21868 20748 21924 20804
rect 21196 19906 21252 19908
rect 21196 19854 21198 19906
rect 21198 19854 21250 19906
rect 21250 19854 21252 19906
rect 21196 19852 21252 19854
rect 20412 19292 20468 19348
rect 20636 17388 20692 17444
rect 21868 19852 21924 19908
rect 22002 19626 22058 19628
rect 22002 19574 22004 19626
rect 22004 19574 22056 19626
rect 22056 19574 22058 19626
rect 22002 19572 22058 19574
rect 22106 19626 22162 19628
rect 22106 19574 22108 19626
rect 22108 19574 22160 19626
rect 22160 19574 22162 19626
rect 22106 19572 22162 19574
rect 22210 19626 22266 19628
rect 22210 19574 22212 19626
rect 22212 19574 22264 19626
rect 22264 19574 22266 19626
rect 22210 19572 22266 19574
rect 21644 18620 21700 18676
rect 22652 18674 22708 18676
rect 22652 18622 22654 18674
rect 22654 18622 22706 18674
rect 22706 18622 22708 18674
rect 22652 18620 22708 18622
rect 23100 20802 23156 20804
rect 23100 20750 23102 20802
rect 23102 20750 23154 20802
rect 23154 20750 23156 20802
rect 23100 20748 23156 20750
rect 22092 18284 22148 18340
rect 21644 16156 21700 16212
rect 21756 16044 21812 16100
rect 19404 13858 19460 13860
rect 19404 13806 19406 13858
rect 19406 13806 19458 13858
rect 19458 13806 19460 13858
rect 19404 13804 19460 13806
rect 18732 13746 18788 13748
rect 18732 13694 18734 13746
rect 18734 13694 18786 13746
rect 18786 13694 18788 13746
rect 18732 13692 18788 13694
rect 19068 13746 19124 13748
rect 19068 13694 19070 13746
rect 19070 13694 19122 13746
rect 19122 13694 19124 13746
rect 19068 13692 19124 13694
rect 19628 13916 19684 13972
rect 19516 13468 19572 13524
rect 18172 12684 18228 12740
rect 17844 12570 17900 12572
rect 17844 12518 17846 12570
rect 17846 12518 17898 12570
rect 17898 12518 17900 12570
rect 17844 12516 17900 12518
rect 17948 12570 18004 12572
rect 17948 12518 17950 12570
rect 17950 12518 18002 12570
rect 18002 12518 18004 12570
rect 17948 12516 18004 12518
rect 18052 12570 18108 12572
rect 18052 12518 18054 12570
rect 18054 12518 18106 12570
rect 18106 12518 18108 12570
rect 18052 12516 18108 12518
rect 18508 12348 18564 12404
rect 18396 12236 18452 12292
rect 17500 10668 17556 10724
rect 17724 11116 17780 11172
rect 17844 11002 17900 11004
rect 17844 10950 17846 11002
rect 17846 10950 17898 11002
rect 17898 10950 17900 11002
rect 17844 10948 17900 10950
rect 17948 11002 18004 11004
rect 17948 10950 17950 11002
rect 17950 10950 18002 11002
rect 18002 10950 18004 11002
rect 17948 10948 18004 10950
rect 18052 11002 18108 11004
rect 18052 10950 18054 11002
rect 18054 10950 18106 11002
rect 18106 10950 18108 11002
rect 18052 10948 18108 10950
rect 18284 10780 18340 10836
rect 18396 10668 18452 10724
rect 17836 10498 17892 10500
rect 17836 10446 17838 10498
rect 17838 10446 17890 10498
rect 17890 10446 17892 10498
rect 17836 10444 17892 10446
rect 17276 10108 17332 10164
rect 19068 13132 19124 13188
rect 18844 12962 18900 12964
rect 18844 12910 18846 12962
rect 18846 12910 18898 12962
rect 18898 12910 18900 12962
rect 18844 12908 18900 12910
rect 18732 12012 18788 12068
rect 19292 12572 19348 12628
rect 19404 12236 19460 12292
rect 19404 12012 19460 12068
rect 18732 10668 18788 10724
rect 16940 9772 16996 9828
rect 17836 9826 17892 9828
rect 17836 9774 17838 9826
rect 17838 9774 17890 9826
rect 17890 9774 17892 9826
rect 17836 9772 17892 9774
rect 17844 9434 17900 9436
rect 17844 9382 17846 9434
rect 17846 9382 17898 9434
rect 17898 9382 17900 9434
rect 17844 9380 17900 9382
rect 17948 9434 18004 9436
rect 17948 9382 17950 9434
rect 17950 9382 18002 9434
rect 18002 9382 18004 9434
rect 17948 9380 18004 9382
rect 18052 9434 18108 9436
rect 18052 9382 18054 9434
rect 18054 9382 18106 9434
rect 18106 9382 18108 9434
rect 18052 9380 18108 9382
rect 17276 9154 17332 9156
rect 17276 9102 17278 9154
rect 17278 9102 17330 9154
rect 17330 9102 17332 9154
rect 17276 9100 17332 9102
rect 18060 9100 18116 9156
rect 16716 7644 16772 7700
rect 16492 7474 16548 7476
rect 16492 7422 16494 7474
rect 16494 7422 16546 7474
rect 16546 7422 16548 7474
rect 16492 7420 16548 7422
rect 16268 7084 16324 7140
rect 17844 7866 17900 7868
rect 17844 7814 17846 7866
rect 17846 7814 17898 7866
rect 17898 7814 17900 7866
rect 17844 7812 17900 7814
rect 17948 7866 18004 7868
rect 17948 7814 17950 7866
rect 17950 7814 18002 7866
rect 18002 7814 18004 7866
rect 17948 7812 18004 7814
rect 18052 7866 18108 7868
rect 18052 7814 18054 7866
rect 18054 7814 18106 7866
rect 18106 7814 18108 7866
rect 18052 7812 18108 7814
rect 17164 6412 17220 6468
rect 17276 6636 17332 6692
rect 16156 4508 16212 4564
rect 16604 5628 16660 5684
rect 17388 7084 17444 7140
rect 18620 9714 18676 9716
rect 18620 9662 18622 9714
rect 18622 9662 18674 9714
rect 18674 9662 18676 9714
rect 18620 9660 18676 9662
rect 18508 8204 18564 8260
rect 22876 18396 22932 18452
rect 22002 18058 22058 18060
rect 22002 18006 22004 18058
rect 22004 18006 22056 18058
rect 22056 18006 22058 18058
rect 22002 18004 22058 18006
rect 22106 18058 22162 18060
rect 22106 18006 22108 18058
rect 22108 18006 22160 18058
rect 22160 18006 22162 18058
rect 22106 18004 22162 18006
rect 22210 18058 22266 18060
rect 22210 18006 22212 18058
rect 22212 18006 22264 18058
rect 22264 18006 22266 18058
rect 22210 18004 22266 18006
rect 22002 16490 22058 16492
rect 22002 16438 22004 16490
rect 22004 16438 22056 16490
rect 22056 16438 22058 16490
rect 22002 16436 22058 16438
rect 22106 16490 22162 16492
rect 22106 16438 22108 16490
rect 22108 16438 22160 16490
rect 22160 16438 22162 16490
rect 22106 16436 22162 16438
rect 22210 16490 22266 16492
rect 22210 16438 22212 16490
rect 22212 16438 22264 16490
rect 22264 16438 22266 16490
rect 22210 16436 22266 16438
rect 22428 16098 22484 16100
rect 22428 16046 22430 16098
rect 22430 16046 22482 16098
rect 22482 16046 22484 16098
rect 22428 16044 22484 16046
rect 21756 15148 21812 15204
rect 22652 15986 22708 15988
rect 22652 15934 22654 15986
rect 22654 15934 22706 15986
rect 22706 15934 22708 15986
rect 22652 15932 22708 15934
rect 23772 25228 23828 25284
rect 24556 25564 24612 25620
rect 23660 24946 23716 24948
rect 23660 24894 23662 24946
rect 23662 24894 23714 24946
rect 23714 24894 23716 24946
rect 23660 24892 23716 24894
rect 23884 24722 23940 24724
rect 23884 24670 23886 24722
rect 23886 24670 23938 24722
rect 23938 24670 23940 24722
rect 23884 24668 23940 24670
rect 24444 24722 24500 24724
rect 24444 24670 24446 24722
rect 24446 24670 24498 24722
rect 24498 24670 24500 24722
rect 24444 24668 24500 24670
rect 25452 25228 25508 25284
rect 25564 25340 25620 25396
rect 30318 25898 30374 25900
rect 30318 25846 30320 25898
rect 30320 25846 30372 25898
rect 30372 25846 30374 25898
rect 30318 25844 30374 25846
rect 30422 25898 30478 25900
rect 30422 25846 30424 25898
rect 30424 25846 30476 25898
rect 30476 25846 30478 25898
rect 30422 25844 30478 25846
rect 30526 25898 30582 25900
rect 30526 25846 30528 25898
rect 30528 25846 30580 25898
rect 30580 25846 30582 25898
rect 30526 25844 30582 25846
rect 26348 25564 26404 25620
rect 25788 25228 25844 25284
rect 25116 24444 25172 24500
rect 25228 23324 25284 23380
rect 25676 23772 25732 23828
rect 24332 23212 24388 23268
rect 24444 23154 24500 23156
rect 24444 23102 24446 23154
rect 24446 23102 24498 23154
rect 24498 23102 24500 23154
rect 24444 23100 24500 23102
rect 24668 22764 24724 22820
rect 25116 23212 25172 23268
rect 25788 23660 25844 23716
rect 25228 22370 25284 22372
rect 25228 22318 25230 22370
rect 25230 22318 25282 22370
rect 25282 22318 25284 22370
rect 25228 22316 25284 22318
rect 24220 21698 24276 21700
rect 24220 21646 24222 21698
rect 24222 21646 24274 21698
rect 24274 21646 24276 21698
rect 24220 21644 24276 21646
rect 25676 21644 25732 21700
rect 24444 21586 24500 21588
rect 24444 21534 24446 21586
rect 24446 21534 24498 21586
rect 24498 21534 24500 21586
rect 24444 21532 24500 21534
rect 24108 21420 24164 21476
rect 23324 18674 23380 18676
rect 23324 18622 23326 18674
rect 23326 18622 23378 18674
rect 23378 18622 23380 18674
rect 23324 18620 23380 18622
rect 23996 20076 24052 20132
rect 24668 21474 24724 21476
rect 24668 21422 24670 21474
rect 24670 21422 24722 21474
rect 24722 21422 24724 21474
rect 24668 21420 24724 21422
rect 24556 20748 24612 20804
rect 22988 18172 23044 18228
rect 23436 16210 23492 16212
rect 23436 16158 23438 16210
rect 23438 16158 23490 16210
rect 23490 16158 23492 16210
rect 23436 16156 23492 16158
rect 22876 15426 22932 15428
rect 22876 15374 22878 15426
rect 22878 15374 22930 15426
rect 22930 15374 22932 15426
rect 22876 15372 22932 15374
rect 19852 13132 19908 13188
rect 20076 14418 20132 14420
rect 20076 14366 20078 14418
rect 20078 14366 20130 14418
rect 20130 14366 20132 14418
rect 20076 14364 20132 14366
rect 19740 12738 19796 12740
rect 19740 12686 19742 12738
rect 19742 12686 19794 12738
rect 19794 12686 19796 12738
rect 19740 12684 19796 12686
rect 19852 12572 19908 12628
rect 20188 13916 20244 13972
rect 20076 13746 20132 13748
rect 20076 13694 20078 13746
rect 20078 13694 20130 13746
rect 20130 13694 20132 13746
rect 20076 13692 20132 13694
rect 20524 14306 20580 14308
rect 20524 14254 20526 14306
rect 20526 14254 20578 14306
rect 20578 14254 20580 14306
rect 20524 14252 20580 14254
rect 20300 13186 20356 13188
rect 20300 13134 20302 13186
rect 20302 13134 20354 13186
rect 20354 13134 20356 13186
rect 20300 13132 20356 13134
rect 20076 13074 20132 13076
rect 20076 13022 20078 13074
rect 20078 13022 20130 13074
rect 20130 13022 20132 13074
rect 20076 13020 20132 13022
rect 21532 14588 21588 14644
rect 22876 15148 22932 15204
rect 21420 14252 21476 14308
rect 21420 13580 21476 13636
rect 21308 13522 21364 13524
rect 21308 13470 21310 13522
rect 21310 13470 21362 13522
rect 21362 13470 21364 13522
rect 21308 13468 21364 13470
rect 20748 13020 20804 13076
rect 20524 12962 20580 12964
rect 20524 12910 20526 12962
rect 20526 12910 20578 12962
rect 20578 12910 20580 12962
rect 20524 12908 20580 12910
rect 20972 12684 21028 12740
rect 19628 11676 19684 11732
rect 18844 10556 18900 10612
rect 19852 11564 19908 11620
rect 19964 12348 20020 12404
rect 20636 12402 20692 12404
rect 20636 12350 20638 12402
rect 20638 12350 20690 12402
rect 20690 12350 20692 12402
rect 20636 12348 20692 12350
rect 20076 11676 20132 11732
rect 20412 11618 20468 11620
rect 20412 11566 20414 11618
rect 20414 11566 20466 11618
rect 20466 11566 20468 11618
rect 20412 11564 20468 11566
rect 21308 11676 21364 11732
rect 18844 9660 18900 9716
rect 18956 10444 19012 10500
rect 19292 10108 19348 10164
rect 22002 14922 22058 14924
rect 22002 14870 22004 14922
rect 22004 14870 22056 14922
rect 22056 14870 22058 14922
rect 22002 14868 22058 14870
rect 22106 14922 22162 14924
rect 22106 14870 22108 14922
rect 22108 14870 22160 14922
rect 22160 14870 22162 14922
rect 22106 14868 22162 14870
rect 22210 14922 22266 14924
rect 22210 14870 22212 14922
rect 22212 14870 22264 14922
rect 22264 14870 22266 14922
rect 22210 14868 22266 14870
rect 22204 14364 22260 14420
rect 21980 13522 22036 13524
rect 21980 13470 21982 13522
rect 21982 13470 22034 13522
rect 22034 13470 22036 13522
rect 21980 13468 22036 13470
rect 22002 13354 22058 13356
rect 22002 13302 22004 13354
rect 22004 13302 22056 13354
rect 22056 13302 22058 13354
rect 22002 13300 22058 13302
rect 22106 13354 22162 13356
rect 22106 13302 22108 13354
rect 22108 13302 22160 13354
rect 22160 13302 22162 13354
rect 22106 13300 22162 13302
rect 22210 13354 22266 13356
rect 22210 13302 22212 13354
rect 22212 13302 22264 13354
rect 22264 13302 22266 13354
rect 22210 13300 22266 13302
rect 22092 13186 22148 13188
rect 22092 13134 22094 13186
rect 22094 13134 22146 13186
rect 22146 13134 22148 13186
rect 22092 13132 22148 13134
rect 22652 13132 22708 13188
rect 22988 13468 23044 13524
rect 22316 13074 22372 13076
rect 22316 13022 22318 13074
rect 22318 13022 22370 13074
rect 22370 13022 22372 13074
rect 22316 13020 22372 13022
rect 21868 12962 21924 12964
rect 21868 12910 21870 12962
rect 21870 12910 21922 12962
rect 21922 12910 21924 12962
rect 21868 12908 21924 12910
rect 21644 12850 21700 12852
rect 21644 12798 21646 12850
rect 21646 12798 21698 12850
rect 21698 12798 21700 12850
rect 21644 12796 21700 12798
rect 22428 12738 22484 12740
rect 22428 12686 22430 12738
rect 22430 12686 22482 12738
rect 22482 12686 22484 12738
rect 22428 12684 22484 12686
rect 21532 11452 21588 11508
rect 22002 11786 22058 11788
rect 22002 11734 22004 11786
rect 22004 11734 22056 11786
rect 22056 11734 22058 11786
rect 22002 11732 22058 11734
rect 22106 11786 22162 11788
rect 22106 11734 22108 11786
rect 22108 11734 22160 11786
rect 22160 11734 22162 11786
rect 22106 11732 22162 11734
rect 22210 11786 22266 11788
rect 22210 11734 22212 11786
rect 22212 11734 22264 11786
rect 22264 11734 22266 11786
rect 22210 11732 22266 11734
rect 22876 12850 22932 12852
rect 22876 12798 22878 12850
rect 22878 12798 22930 12850
rect 22930 12798 22932 12850
rect 22876 12796 22932 12798
rect 22876 11506 22932 11508
rect 22876 11454 22878 11506
rect 22878 11454 22930 11506
rect 22930 11454 22932 11506
rect 22876 11452 22932 11454
rect 21532 10780 21588 10836
rect 19852 9884 19908 9940
rect 18844 9154 18900 9156
rect 18844 9102 18846 9154
rect 18846 9102 18898 9154
rect 18898 9102 18900 9154
rect 18844 9100 18900 9102
rect 20412 9938 20468 9940
rect 20412 9886 20414 9938
rect 20414 9886 20466 9938
rect 20466 9886 20468 9938
rect 20412 9884 20468 9886
rect 19068 8876 19124 8932
rect 18732 8316 18788 8372
rect 19628 8316 19684 8372
rect 17724 6412 17780 6468
rect 17276 5628 17332 5684
rect 18732 6466 18788 6468
rect 18732 6414 18734 6466
rect 18734 6414 18786 6466
rect 18786 6414 18788 6466
rect 18732 6412 18788 6414
rect 17844 6298 17900 6300
rect 17844 6246 17846 6298
rect 17846 6246 17898 6298
rect 17898 6246 17900 6298
rect 17844 6244 17900 6246
rect 17948 6298 18004 6300
rect 17948 6246 17950 6298
rect 17950 6246 18002 6298
rect 18002 6246 18004 6298
rect 17948 6244 18004 6246
rect 18052 6298 18108 6300
rect 18052 6246 18054 6298
rect 18054 6246 18106 6298
rect 18106 6246 18108 6298
rect 18052 6244 18108 6246
rect 17724 5740 17780 5796
rect 16940 5068 16996 5124
rect 17836 5516 17892 5572
rect 18284 5180 18340 5236
rect 18172 5122 18228 5124
rect 18172 5070 18174 5122
rect 18174 5070 18226 5122
rect 18226 5070 18228 5122
rect 18172 5068 18228 5070
rect 17844 4730 17900 4732
rect 17844 4678 17846 4730
rect 17846 4678 17898 4730
rect 17898 4678 17900 4730
rect 17844 4676 17900 4678
rect 17948 4730 18004 4732
rect 17948 4678 17950 4730
rect 17950 4678 18002 4730
rect 18002 4678 18004 4730
rect 17948 4676 18004 4678
rect 18052 4730 18108 4732
rect 18052 4678 18054 4730
rect 18054 4678 18106 4730
rect 18106 4678 18108 4730
rect 18052 4676 18108 4678
rect 17500 4562 17556 4564
rect 17500 4510 17502 4562
rect 17502 4510 17554 4562
rect 17554 4510 17556 4562
rect 17500 4508 17556 4510
rect 12572 3500 12628 3556
rect 17844 3162 17900 3164
rect 17844 3110 17846 3162
rect 17846 3110 17898 3162
rect 17898 3110 17900 3162
rect 17844 3108 17900 3110
rect 17948 3162 18004 3164
rect 17948 3110 17950 3162
rect 17950 3110 18002 3162
rect 18002 3110 18004 3162
rect 17948 3108 18004 3110
rect 18052 3162 18108 3164
rect 18052 3110 18054 3162
rect 18054 3110 18106 3162
rect 18106 3110 18108 3162
rect 18052 3108 18108 3110
rect 18620 4562 18676 4564
rect 18620 4510 18622 4562
rect 18622 4510 18674 4562
rect 18674 4510 18676 4562
rect 18620 4508 18676 4510
rect 19068 8204 19124 8260
rect 19516 6076 19572 6132
rect 19292 5906 19348 5908
rect 19292 5854 19294 5906
rect 19294 5854 19346 5906
rect 19346 5854 19348 5906
rect 19292 5852 19348 5854
rect 18956 5516 19012 5572
rect 19180 5234 19236 5236
rect 19180 5182 19182 5234
rect 19182 5182 19234 5234
rect 19234 5182 19236 5234
rect 19180 5180 19236 5182
rect 18844 5068 18900 5124
rect 19180 4508 19236 4564
rect 21420 9714 21476 9716
rect 21420 9662 21422 9714
rect 21422 9662 21474 9714
rect 21474 9662 21476 9714
rect 21420 9660 21476 9662
rect 20972 9042 21028 9044
rect 20972 8990 20974 9042
rect 20974 8990 21026 9042
rect 21026 8990 21028 9042
rect 20972 8988 21028 8990
rect 20972 8428 21028 8484
rect 22316 10610 22372 10612
rect 22316 10558 22318 10610
rect 22318 10558 22370 10610
rect 22370 10558 22372 10610
rect 22316 10556 22372 10558
rect 23436 14642 23492 14644
rect 23436 14590 23438 14642
rect 23438 14590 23490 14642
rect 23490 14590 23492 14642
rect 23436 14588 23492 14590
rect 23660 18284 23716 18340
rect 25900 21420 25956 21476
rect 25900 20914 25956 20916
rect 25900 20862 25902 20914
rect 25902 20862 25954 20914
rect 25954 20862 25956 20914
rect 25900 20860 25956 20862
rect 25676 20188 25732 20244
rect 26460 25340 26516 25396
rect 26160 25114 26216 25116
rect 26160 25062 26162 25114
rect 26162 25062 26214 25114
rect 26214 25062 26216 25114
rect 26160 25060 26216 25062
rect 26264 25114 26320 25116
rect 26264 25062 26266 25114
rect 26266 25062 26318 25114
rect 26318 25062 26320 25114
rect 26264 25060 26320 25062
rect 26368 25114 26424 25116
rect 26368 25062 26370 25114
rect 26370 25062 26422 25114
rect 26422 25062 26424 25114
rect 26368 25060 26424 25062
rect 26348 24668 26404 24724
rect 27244 25282 27300 25284
rect 27244 25230 27246 25282
rect 27246 25230 27298 25282
rect 27298 25230 27300 25282
rect 27244 25228 27300 25230
rect 34476 25114 34532 25116
rect 34476 25062 34478 25114
rect 34478 25062 34530 25114
rect 34530 25062 34532 25114
rect 34476 25060 34532 25062
rect 34580 25114 34636 25116
rect 34580 25062 34582 25114
rect 34582 25062 34634 25114
rect 34634 25062 34636 25114
rect 34580 25060 34636 25062
rect 34684 25114 34740 25116
rect 34684 25062 34686 25114
rect 34686 25062 34738 25114
rect 34738 25062 34740 25114
rect 34684 25060 34740 25062
rect 26124 23996 26180 24052
rect 26684 23996 26740 24052
rect 26684 23826 26740 23828
rect 26684 23774 26686 23826
rect 26686 23774 26738 23826
rect 26738 23774 26740 23826
rect 26684 23772 26740 23774
rect 26348 23714 26404 23716
rect 26348 23662 26350 23714
rect 26350 23662 26402 23714
rect 26402 23662 26404 23714
rect 26348 23660 26404 23662
rect 26160 23546 26216 23548
rect 26160 23494 26162 23546
rect 26162 23494 26214 23546
rect 26214 23494 26216 23546
rect 26160 23492 26216 23494
rect 26264 23546 26320 23548
rect 26264 23494 26266 23546
rect 26266 23494 26318 23546
rect 26318 23494 26320 23546
rect 26264 23492 26320 23494
rect 26368 23546 26424 23548
rect 26368 23494 26370 23546
rect 26370 23494 26422 23546
rect 26422 23494 26424 23546
rect 26368 23492 26424 23494
rect 26348 23324 26404 23380
rect 26124 23154 26180 23156
rect 26124 23102 26126 23154
rect 26126 23102 26178 23154
rect 26178 23102 26180 23154
rect 26124 23100 26180 23102
rect 26908 23714 26964 23716
rect 26908 23662 26910 23714
rect 26910 23662 26962 23714
rect 26962 23662 26964 23714
rect 26908 23660 26964 23662
rect 27020 23212 27076 23268
rect 29148 23266 29204 23268
rect 29148 23214 29150 23266
rect 29150 23214 29202 23266
rect 29202 23214 29204 23266
rect 29148 23212 29204 23214
rect 30318 24330 30374 24332
rect 30318 24278 30320 24330
rect 30320 24278 30372 24330
rect 30372 24278 30374 24330
rect 30318 24276 30374 24278
rect 30422 24330 30478 24332
rect 30422 24278 30424 24330
rect 30424 24278 30476 24330
rect 30476 24278 30478 24330
rect 30422 24276 30478 24278
rect 30526 24330 30582 24332
rect 30526 24278 30528 24330
rect 30528 24278 30580 24330
rect 30580 24278 30582 24330
rect 30526 24276 30582 24278
rect 34476 23546 34532 23548
rect 34476 23494 34478 23546
rect 34478 23494 34530 23546
rect 34530 23494 34532 23546
rect 34476 23492 34532 23494
rect 34580 23546 34636 23548
rect 34580 23494 34582 23546
rect 34582 23494 34634 23546
rect 34634 23494 34636 23546
rect 34580 23492 34636 23494
rect 34684 23546 34740 23548
rect 34684 23494 34686 23546
rect 34686 23494 34738 23546
rect 34738 23494 34740 23546
rect 34684 23492 34740 23494
rect 26908 23100 26964 23156
rect 26348 22370 26404 22372
rect 26348 22318 26350 22370
rect 26350 22318 26402 22370
rect 26402 22318 26404 22370
rect 26348 22316 26404 22318
rect 26908 22764 26964 22820
rect 27020 22316 27076 22372
rect 26572 22146 26628 22148
rect 26572 22094 26574 22146
rect 26574 22094 26626 22146
rect 26626 22094 26628 22146
rect 26572 22092 26628 22094
rect 26160 21978 26216 21980
rect 26160 21926 26162 21978
rect 26162 21926 26214 21978
rect 26214 21926 26216 21978
rect 26160 21924 26216 21926
rect 26264 21978 26320 21980
rect 26264 21926 26266 21978
rect 26266 21926 26318 21978
rect 26318 21926 26320 21978
rect 26264 21924 26320 21926
rect 26368 21978 26424 21980
rect 26368 21926 26370 21978
rect 26370 21926 26422 21978
rect 26422 21926 26424 21978
rect 26368 21924 26424 21926
rect 26796 22092 26852 22148
rect 26124 21698 26180 21700
rect 26124 21646 26126 21698
rect 26126 21646 26178 21698
rect 26178 21646 26180 21698
rect 26124 21644 26180 21646
rect 26124 21362 26180 21364
rect 26124 21310 26126 21362
rect 26126 21310 26178 21362
rect 26178 21310 26180 21362
rect 26124 21308 26180 21310
rect 26012 20748 26068 20804
rect 26572 21532 26628 21588
rect 26684 20860 26740 20916
rect 27468 22092 27524 22148
rect 27580 21308 27636 21364
rect 30318 22762 30374 22764
rect 30318 22710 30320 22762
rect 30320 22710 30372 22762
rect 30372 22710 30374 22762
rect 30318 22708 30374 22710
rect 30422 22762 30478 22764
rect 30422 22710 30424 22762
rect 30424 22710 30476 22762
rect 30476 22710 30478 22762
rect 30422 22708 30478 22710
rect 30526 22762 30582 22764
rect 30526 22710 30528 22762
rect 30528 22710 30580 22762
rect 30580 22710 30582 22762
rect 30526 22708 30582 22710
rect 34476 21978 34532 21980
rect 34476 21926 34478 21978
rect 34478 21926 34530 21978
rect 34530 21926 34532 21978
rect 34476 21924 34532 21926
rect 34580 21978 34636 21980
rect 34580 21926 34582 21978
rect 34582 21926 34634 21978
rect 34634 21926 34636 21978
rect 34580 21924 34636 21926
rect 34684 21978 34740 21980
rect 34684 21926 34686 21978
rect 34686 21926 34738 21978
rect 34738 21926 34740 21978
rect 34684 21924 34740 21926
rect 28028 20914 28084 20916
rect 28028 20862 28030 20914
rect 28030 20862 28082 20914
rect 28082 20862 28084 20914
rect 28028 20860 28084 20862
rect 28700 20860 28756 20916
rect 26160 20410 26216 20412
rect 26160 20358 26162 20410
rect 26162 20358 26214 20410
rect 26214 20358 26216 20410
rect 26160 20356 26216 20358
rect 26264 20410 26320 20412
rect 26264 20358 26266 20410
rect 26266 20358 26318 20410
rect 26318 20358 26320 20410
rect 26264 20356 26320 20358
rect 26368 20410 26424 20412
rect 26368 20358 26370 20410
rect 26370 20358 26422 20410
rect 26422 20358 26424 20410
rect 26368 20356 26424 20358
rect 26572 20076 26628 20132
rect 26160 18842 26216 18844
rect 26160 18790 26162 18842
rect 26162 18790 26214 18842
rect 26214 18790 26216 18842
rect 26160 18788 26216 18790
rect 26264 18842 26320 18844
rect 26264 18790 26266 18842
rect 26266 18790 26318 18842
rect 26318 18790 26320 18842
rect 26264 18788 26320 18790
rect 26368 18842 26424 18844
rect 26368 18790 26370 18842
rect 26370 18790 26422 18842
rect 26422 18790 26424 18842
rect 26368 18788 26424 18790
rect 26236 18450 26292 18452
rect 26236 18398 26238 18450
rect 26238 18398 26290 18450
rect 26290 18398 26292 18450
rect 26236 18396 26292 18398
rect 25676 18284 25732 18340
rect 23660 16098 23716 16100
rect 23660 16046 23662 16098
rect 23662 16046 23714 16098
rect 23714 16046 23716 16098
rect 23660 16044 23716 16046
rect 27244 18450 27300 18452
rect 27244 18398 27246 18450
rect 27246 18398 27298 18450
rect 27298 18398 27300 18450
rect 27244 18396 27300 18398
rect 26684 17948 26740 18004
rect 26236 17890 26292 17892
rect 26236 17838 26238 17890
rect 26238 17838 26290 17890
rect 26290 17838 26292 17890
rect 26236 17836 26292 17838
rect 24332 15986 24388 15988
rect 24332 15934 24334 15986
rect 24334 15934 24386 15986
rect 24386 15934 24388 15986
rect 24332 15932 24388 15934
rect 26012 17554 26068 17556
rect 26012 17502 26014 17554
rect 26014 17502 26066 17554
rect 26066 17502 26068 17554
rect 26012 17500 26068 17502
rect 26160 17274 26216 17276
rect 26160 17222 26162 17274
rect 26162 17222 26214 17274
rect 26214 17222 26216 17274
rect 26160 17220 26216 17222
rect 26264 17274 26320 17276
rect 26264 17222 26266 17274
rect 26266 17222 26318 17274
rect 26318 17222 26320 17274
rect 26264 17220 26320 17222
rect 26368 17274 26424 17276
rect 26368 17222 26370 17274
rect 26370 17222 26422 17274
rect 26422 17222 26424 17274
rect 26368 17220 26424 17222
rect 25900 16044 25956 16100
rect 24556 15148 24612 15204
rect 26160 15706 26216 15708
rect 26160 15654 26162 15706
rect 26162 15654 26214 15706
rect 26214 15654 26216 15706
rect 26160 15652 26216 15654
rect 26264 15706 26320 15708
rect 26264 15654 26266 15706
rect 26266 15654 26318 15706
rect 26318 15654 26320 15706
rect 26264 15652 26320 15654
rect 26368 15706 26424 15708
rect 26368 15654 26370 15706
rect 26370 15654 26422 15706
rect 26422 15654 26424 15706
rect 26368 15652 26424 15654
rect 28476 17948 28532 18004
rect 27916 17836 27972 17892
rect 28140 17836 28196 17892
rect 27244 16716 27300 16772
rect 26908 16156 26964 16212
rect 27020 16098 27076 16100
rect 27020 16046 27022 16098
rect 27022 16046 27074 16098
rect 27074 16046 27076 16098
rect 27020 16044 27076 16046
rect 27356 15874 27412 15876
rect 27356 15822 27358 15874
rect 27358 15822 27410 15874
rect 27410 15822 27412 15874
rect 27356 15820 27412 15822
rect 27580 16716 27636 16772
rect 28140 16770 28196 16772
rect 28140 16718 28142 16770
rect 28142 16718 28194 16770
rect 28194 16718 28196 16770
rect 28140 16716 28196 16718
rect 28028 16210 28084 16212
rect 28028 16158 28030 16210
rect 28030 16158 28082 16210
rect 28082 16158 28084 16210
rect 28028 16156 28084 16158
rect 27692 15596 27748 15652
rect 27580 15538 27636 15540
rect 27580 15486 27582 15538
rect 27582 15486 27634 15538
rect 27634 15486 27636 15538
rect 27580 15484 27636 15486
rect 30318 21194 30374 21196
rect 30318 21142 30320 21194
rect 30320 21142 30372 21194
rect 30372 21142 30374 21194
rect 30318 21140 30374 21142
rect 30422 21194 30478 21196
rect 30422 21142 30424 21194
rect 30424 21142 30476 21194
rect 30476 21142 30478 21194
rect 30422 21140 30478 21142
rect 30526 21194 30582 21196
rect 30526 21142 30528 21194
rect 30528 21142 30580 21194
rect 30580 21142 30582 21194
rect 30526 21140 30582 21142
rect 34476 20410 34532 20412
rect 34476 20358 34478 20410
rect 34478 20358 34530 20410
rect 34530 20358 34532 20410
rect 34476 20356 34532 20358
rect 34580 20410 34636 20412
rect 34580 20358 34582 20410
rect 34582 20358 34634 20410
rect 34634 20358 34636 20410
rect 34580 20356 34636 20358
rect 34684 20410 34740 20412
rect 34684 20358 34686 20410
rect 34686 20358 34738 20410
rect 34738 20358 34740 20410
rect 34684 20356 34740 20358
rect 30318 19626 30374 19628
rect 30318 19574 30320 19626
rect 30320 19574 30372 19626
rect 30372 19574 30374 19626
rect 30318 19572 30374 19574
rect 30422 19626 30478 19628
rect 30422 19574 30424 19626
rect 30424 19574 30476 19626
rect 30476 19574 30478 19626
rect 30422 19572 30478 19574
rect 30526 19626 30582 19628
rect 30526 19574 30528 19626
rect 30528 19574 30580 19626
rect 30580 19574 30582 19626
rect 30526 19572 30582 19574
rect 34476 18842 34532 18844
rect 34476 18790 34478 18842
rect 34478 18790 34530 18842
rect 34530 18790 34532 18842
rect 34476 18788 34532 18790
rect 34580 18842 34636 18844
rect 34580 18790 34582 18842
rect 34582 18790 34634 18842
rect 34634 18790 34636 18842
rect 34580 18788 34636 18790
rect 34684 18842 34740 18844
rect 34684 18790 34686 18842
rect 34686 18790 34738 18842
rect 34738 18790 34740 18842
rect 34684 18788 34740 18790
rect 29260 18338 29316 18340
rect 29260 18286 29262 18338
rect 29262 18286 29314 18338
rect 29314 18286 29316 18338
rect 29260 18284 29316 18286
rect 28588 17836 28644 17892
rect 29148 17612 29204 17668
rect 28924 17500 28980 17556
rect 30318 18058 30374 18060
rect 30318 18006 30320 18058
rect 30320 18006 30372 18058
rect 30372 18006 30374 18058
rect 30318 18004 30374 18006
rect 30422 18058 30478 18060
rect 30422 18006 30424 18058
rect 30424 18006 30476 18058
rect 30476 18006 30478 18058
rect 30422 18004 30478 18006
rect 30526 18058 30582 18060
rect 30526 18006 30528 18058
rect 30528 18006 30580 18058
rect 30580 18006 30582 18058
rect 30526 18004 30582 18006
rect 29596 17612 29652 17668
rect 28364 16268 28420 16324
rect 31388 17612 31444 17668
rect 31276 17554 31332 17556
rect 31276 17502 31278 17554
rect 31278 17502 31330 17554
rect 31330 17502 31332 17554
rect 31276 17500 31332 17502
rect 30380 16770 30436 16772
rect 30380 16718 30382 16770
rect 30382 16718 30434 16770
rect 30434 16718 30436 16770
rect 30380 16716 30436 16718
rect 30318 16490 30374 16492
rect 30318 16438 30320 16490
rect 30320 16438 30372 16490
rect 30372 16438 30374 16490
rect 30318 16436 30374 16438
rect 30422 16490 30478 16492
rect 30422 16438 30424 16490
rect 30424 16438 30476 16490
rect 30476 16438 30478 16490
rect 30422 16436 30478 16438
rect 30526 16490 30582 16492
rect 30526 16438 30528 16490
rect 30528 16438 30580 16490
rect 30580 16438 30582 16490
rect 30526 16436 30582 16438
rect 30716 16268 30772 16324
rect 28476 15596 28532 15652
rect 29372 15484 29428 15540
rect 29708 15484 29764 15540
rect 27244 14252 27300 14308
rect 23212 10556 23268 10612
rect 22002 10218 22058 10220
rect 22002 10166 22004 10218
rect 22004 10166 22056 10218
rect 22056 10166 22058 10218
rect 22002 10164 22058 10166
rect 22106 10218 22162 10220
rect 22106 10166 22108 10218
rect 22108 10166 22160 10218
rect 22160 10166 22162 10218
rect 22106 10164 22162 10166
rect 22210 10218 22266 10220
rect 22210 10166 22212 10218
rect 22212 10166 22264 10218
rect 22264 10166 22266 10218
rect 22210 10164 22266 10166
rect 21644 9660 21700 9716
rect 22092 9212 22148 9268
rect 22876 9714 22932 9716
rect 22876 9662 22878 9714
rect 22878 9662 22930 9714
rect 22930 9662 22932 9714
rect 22876 9660 22932 9662
rect 21868 8876 21924 8932
rect 22876 8988 22932 9044
rect 22002 8650 22058 8652
rect 22002 8598 22004 8650
rect 22004 8598 22056 8650
rect 22056 8598 22058 8650
rect 22002 8596 22058 8598
rect 22106 8650 22162 8652
rect 22106 8598 22108 8650
rect 22108 8598 22160 8650
rect 22160 8598 22162 8650
rect 22106 8596 22162 8598
rect 22210 8650 22266 8652
rect 22210 8598 22212 8650
rect 22212 8598 22264 8650
rect 22264 8598 22266 8650
rect 22210 8596 22266 8598
rect 21756 8034 21812 8036
rect 21756 7982 21758 8034
rect 21758 7982 21810 8034
rect 21810 7982 21812 8034
rect 21756 7980 21812 7982
rect 21644 7420 21700 7476
rect 22204 7474 22260 7476
rect 22204 7422 22206 7474
rect 22206 7422 22258 7474
rect 22258 7422 22260 7474
rect 22204 7420 22260 7422
rect 22002 7082 22058 7084
rect 22002 7030 22004 7082
rect 22004 7030 22056 7082
rect 22056 7030 22058 7082
rect 22002 7028 22058 7030
rect 22106 7082 22162 7084
rect 22106 7030 22108 7082
rect 22108 7030 22160 7082
rect 22160 7030 22162 7082
rect 22106 7028 22162 7030
rect 22210 7082 22266 7084
rect 22210 7030 22212 7082
rect 22212 7030 22264 7082
rect 22264 7030 22266 7082
rect 22210 7028 22266 7030
rect 21420 6636 21476 6692
rect 22092 6860 22148 6916
rect 21868 6748 21924 6804
rect 21756 6690 21812 6692
rect 21756 6638 21758 6690
rect 21758 6638 21810 6690
rect 21810 6638 21812 6690
rect 21756 6636 21812 6638
rect 21308 6076 21364 6132
rect 21644 5964 21700 6020
rect 21644 5234 21700 5236
rect 21644 5182 21646 5234
rect 21646 5182 21698 5234
rect 21698 5182 21700 5234
rect 21644 5180 21700 5182
rect 20860 4508 20916 4564
rect 20300 4226 20356 4228
rect 20300 4174 20302 4226
rect 20302 4174 20354 4226
rect 20354 4174 20356 4226
rect 20300 4172 20356 4174
rect 22002 5514 22058 5516
rect 22002 5462 22004 5514
rect 22004 5462 22056 5514
rect 22056 5462 22058 5514
rect 22002 5460 22058 5462
rect 22106 5514 22162 5516
rect 22106 5462 22108 5514
rect 22108 5462 22160 5514
rect 22160 5462 22162 5514
rect 22106 5460 22162 5462
rect 22210 5514 22266 5516
rect 22210 5462 22212 5514
rect 22212 5462 22264 5514
rect 22264 5462 22266 5514
rect 22210 5460 22266 5462
rect 21868 4508 21924 4564
rect 21756 4284 21812 4340
rect 22540 7420 22596 7476
rect 23884 13746 23940 13748
rect 23884 13694 23886 13746
rect 23886 13694 23938 13746
rect 23938 13694 23940 13746
rect 23884 13692 23940 13694
rect 23660 12684 23716 12740
rect 24332 9660 24388 9716
rect 25676 13970 25732 13972
rect 25676 13918 25678 13970
rect 25678 13918 25730 13970
rect 25730 13918 25732 13970
rect 25676 13916 25732 13918
rect 25452 13804 25508 13860
rect 24780 13468 24836 13524
rect 26160 14138 26216 14140
rect 26160 14086 26162 14138
rect 26162 14086 26214 14138
rect 26214 14086 26216 14138
rect 26160 14084 26216 14086
rect 26264 14138 26320 14140
rect 26264 14086 26266 14138
rect 26266 14086 26318 14138
rect 26318 14086 26320 14138
rect 26264 14084 26320 14086
rect 26368 14138 26424 14140
rect 26368 14086 26370 14138
rect 26370 14086 26422 14138
rect 26422 14086 26424 14138
rect 26368 14084 26424 14086
rect 26684 13916 26740 13972
rect 26124 13746 26180 13748
rect 26124 13694 26126 13746
rect 26126 13694 26178 13746
rect 26178 13694 26180 13746
rect 26124 13692 26180 13694
rect 26460 13634 26516 13636
rect 26460 13582 26462 13634
rect 26462 13582 26514 13634
rect 26514 13582 26516 13634
rect 26460 13580 26516 13582
rect 26348 13356 26404 13412
rect 26684 13244 26740 13300
rect 26160 12570 26216 12572
rect 26160 12518 26162 12570
rect 26162 12518 26214 12570
rect 26214 12518 26216 12570
rect 26160 12516 26216 12518
rect 26264 12570 26320 12572
rect 26264 12518 26266 12570
rect 26266 12518 26318 12570
rect 26318 12518 26320 12570
rect 26264 12516 26320 12518
rect 26368 12570 26424 12572
rect 26368 12518 26370 12570
rect 26370 12518 26422 12570
rect 26422 12518 26424 12570
rect 26368 12516 26424 12518
rect 24668 9548 24724 9604
rect 26160 11002 26216 11004
rect 26160 10950 26162 11002
rect 26162 10950 26214 11002
rect 26214 10950 26216 11002
rect 26160 10948 26216 10950
rect 26264 11002 26320 11004
rect 26264 10950 26266 11002
rect 26266 10950 26318 11002
rect 26318 10950 26320 11002
rect 26264 10948 26320 10950
rect 26368 11002 26424 11004
rect 26368 10950 26370 11002
rect 26370 10950 26422 11002
rect 26422 10950 26424 11002
rect 26368 10948 26424 10950
rect 26160 9434 26216 9436
rect 26160 9382 26162 9434
rect 26162 9382 26214 9434
rect 26214 9382 26216 9434
rect 26160 9380 26216 9382
rect 26264 9434 26320 9436
rect 26264 9382 26266 9434
rect 26266 9382 26318 9434
rect 26318 9382 26320 9434
rect 26264 9380 26320 9382
rect 26368 9434 26424 9436
rect 26368 9382 26370 9434
rect 26370 9382 26422 9434
rect 26422 9382 26424 9434
rect 26368 9380 26424 9382
rect 24556 9212 24612 9268
rect 23884 8930 23940 8932
rect 23884 8878 23886 8930
rect 23886 8878 23938 8930
rect 23938 8878 23940 8930
rect 23884 8876 23940 8878
rect 23324 7980 23380 8036
rect 22988 7474 23044 7476
rect 22988 7422 22990 7474
rect 22990 7422 23042 7474
rect 23042 7422 23044 7474
rect 22988 7420 23044 7422
rect 23324 6860 23380 6916
rect 22988 6578 23044 6580
rect 22988 6526 22990 6578
rect 22990 6526 23042 6578
rect 23042 6526 23044 6578
rect 22988 6524 23044 6526
rect 22988 6018 23044 6020
rect 22988 5966 22990 6018
rect 22990 5966 23042 6018
rect 23042 5966 23044 6018
rect 22988 5964 23044 5966
rect 22764 4956 22820 5012
rect 23548 6860 23604 6916
rect 23436 6748 23492 6804
rect 26012 9212 26068 9268
rect 27020 13916 27076 13972
rect 27468 13692 27524 13748
rect 27244 13634 27300 13636
rect 27244 13582 27246 13634
rect 27246 13582 27298 13634
rect 27298 13582 27300 13634
rect 27244 13580 27300 13582
rect 26908 13522 26964 13524
rect 26908 13470 26910 13522
rect 26910 13470 26962 13522
rect 26962 13470 26964 13522
rect 26908 13468 26964 13470
rect 27356 13522 27412 13524
rect 27356 13470 27358 13522
rect 27358 13470 27410 13522
rect 27410 13470 27412 13522
rect 27356 13468 27412 13470
rect 27804 14252 27860 14308
rect 27804 13634 27860 13636
rect 27804 13582 27806 13634
rect 27806 13582 27858 13634
rect 27858 13582 27860 13634
rect 27804 13580 27860 13582
rect 27580 13356 27636 13412
rect 27132 10780 27188 10836
rect 26908 10610 26964 10612
rect 26908 10558 26910 10610
rect 26910 10558 26962 10610
rect 26962 10558 26964 10610
rect 26908 10556 26964 10558
rect 27804 9548 27860 9604
rect 27132 9212 27188 9268
rect 24108 7308 24164 7364
rect 23772 5852 23828 5908
rect 26160 7866 26216 7868
rect 26160 7814 26162 7866
rect 26162 7814 26214 7866
rect 26214 7814 26216 7866
rect 26160 7812 26216 7814
rect 26264 7866 26320 7868
rect 26264 7814 26266 7866
rect 26266 7814 26318 7866
rect 26318 7814 26320 7866
rect 26264 7812 26320 7814
rect 26368 7866 26424 7868
rect 26368 7814 26370 7866
rect 26370 7814 26422 7866
rect 26422 7814 26424 7866
rect 26368 7812 26424 7814
rect 26012 7532 26068 7588
rect 25676 7196 25732 7252
rect 24780 6578 24836 6580
rect 24780 6526 24782 6578
rect 24782 6526 24834 6578
rect 24834 6526 24836 6578
rect 24780 6524 24836 6526
rect 24444 6076 24500 6132
rect 24444 5906 24500 5908
rect 24444 5854 24446 5906
rect 24446 5854 24498 5906
rect 24498 5854 24500 5906
rect 24444 5852 24500 5854
rect 25676 6076 25732 6132
rect 25564 5906 25620 5908
rect 25564 5854 25566 5906
rect 25566 5854 25618 5906
rect 25618 5854 25620 5906
rect 25564 5852 25620 5854
rect 24108 5404 24164 5460
rect 22002 3946 22058 3948
rect 22002 3894 22004 3946
rect 22004 3894 22056 3946
rect 22056 3894 22058 3946
rect 22002 3892 22058 3894
rect 22106 3946 22162 3948
rect 22106 3894 22108 3946
rect 22108 3894 22160 3946
rect 22160 3894 22162 3946
rect 22106 3892 22162 3894
rect 22210 3946 22266 3948
rect 22210 3894 22212 3946
rect 22212 3894 22264 3946
rect 22264 3894 22266 3946
rect 22210 3892 22266 3894
rect 19740 3554 19796 3556
rect 19740 3502 19742 3554
rect 19742 3502 19794 3554
rect 19794 3502 19796 3554
rect 19740 3500 19796 3502
rect 20748 3554 20804 3556
rect 20748 3502 20750 3554
rect 20750 3502 20802 3554
rect 20802 3502 20804 3554
rect 20748 3500 20804 3502
rect 22764 4562 22820 4564
rect 22764 4510 22766 4562
rect 22766 4510 22818 4562
rect 22818 4510 22820 4562
rect 22764 4508 22820 4510
rect 23100 4338 23156 4340
rect 23100 4286 23102 4338
rect 23102 4286 23154 4338
rect 23154 4286 23156 4338
rect 23100 4284 23156 4286
rect 23772 5180 23828 5236
rect 23436 4956 23492 5012
rect 23324 4060 23380 4116
rect 22764 3612 22820 3668
rect 25340 5404 25396 5460
rect 23660 4226 23716 4228
rect 23660 4174 23662 4226
rect 23662 4174 23714 4226
rect 23714 4174 23716 4226
rect 23660 4172 23716 4174
rect 26236 7474 26292 7476
rect 26236 7422 26238 7474
rect 26238 7422 26290 7474
rect 26290 7422 26292 7474
rect 26236 7420 26292 7422
rect 26796 7420 26852 7476
rect 26684 7084 26740 7140
rect 26796 6972 26852 7028
rect 26684 6748 26740 6804
rect 26460 6690 26516 6692
rect 26460 6638 26462 6690
rect 26462 6638 26514 6690
rect 26514 6638 26516 6690
rect 26460 6636 26516 6638
rect 26160 6298 26216 6300
rect 26160 6246 26162 6298
rect 26162 6246 26214 6298
rect 26214 6246 26216 6298
rect 26160 6244 26216 6246
rect 26264 6298 26320 6300
rect 26264 6246 26266 6298
rect 26266 6246 26318 6298
rect 26318 6246 26320 6298
rect 26264 6244 26320 6246
rect 26368 6298 26424 6300
rect 26368 6246 26370 6298
rect 26370 6246 26422 6298
rect 26422 6246 26424 6298
rect 26368 6244 26424 6246
rect 28028 14530 28084 14532
rect 28028 14478 28030 14530
rect 28030 14478 28082 14530
rect 28082 14478 28084 14530
rect 28028 14476 28084 14478
rect 28588 15036 28644 15092
rect 29260 15426 29316 15428
rect 29260 15374 29262 15426
rect 29262 15374 29314 15426
rect 29314 15374 29316 15426
rect 29260 15372 29316 15374
rect 31948 17666 32004 17668
rect 31948 17614 31950 17666
rect 31950 17614 32002 17666
rect 32002 17614 32004 17666
rect 31948 17612 32004 17614
rect 34476 17274 34532 17276
rect 34476 17222 34478 17274
rect 34478 17222 34530 17274
rect 34530 17222 34532 17274
rect 34476 17220 34532 17222
rect 34580 17274 34636 17276
rect 34580 17222 34582 17274
rect 34582 17222 34634 17274
rect 34634 17222 34636 17274
rect 34580 17220 34636 17222
rect 34684 17274 34740 17276
rect 34684 17222 34686 17274
rect 34686 17222 34738 17274
rect 34738 17222 34740 17274
rect 34684 17220 34740 17222
rect 31948 16716 32004 16772
rect 31724 16604 31780 16660
rect 28812 14588 28868 14644
rect 28588 13804 28644 13860
rect 28252 13468 28308 13524
rect 30044 15372 30100 15428
rect 29820 15036 29876 15092
rect 29596 14642 29652 14644
rect 29596 14590 29598 14642
rect 29598 14590 29650 14642
rect 29650 14590 29652 14642
rect 29596 14588 29652 14590
rect 29484 14476 29540 14532
rect 29148 13244 29204 13300
rect 30380 15260 30436 15316
rect 30604 15202 30660 15204
rect 30604 15150 30606 15202
rect 30606 15150 30658 15202
rect 30658 15150 30660 15202
rect 30604 15148 30660 15150
rect 30492 15036 30548 15092
rect 30318 14922 30374 14924
rect 30318 14870 30320 14922
rect 30320 14870 30372 14922
rect 30372 14870 30374 14922
rect 30318 14868 30374 14870
rect 30422 14922 30478 14924
rect 30422 14870 30424 14922
rect 30424 14870 30476 14922
rect 30476 14870 30478 14922
rect 30422 14868 30478 14870
rect 30526 14922 30582 14924
rect 30526 14870 30528 14922
rect 30528 14870 30580 14922
rect 30580 14870 30582 14922
rect 30526 14868 30582 14870
rect 30940 15820 30996 15876
rect 31500 15372 31556 15428
rect 31052 15314 31108 15316
rect 31052 15262 31054 15314
rect 31054 15262 31106 15314
rect 31106 15262 31108 15314
rect 31052 15260 31108 15262
rect 31388 15260 31444 15316
rect 29708 13580 29764 13636
rect 30318 13354 30374 13356
rect 30318 13302 30320 13354
rect 30320 13302 30372 13354
rect 30372 13302 30374 13354
rect 30318 13300 30374 13302
rect 30422 13354 30478 13356
rect 30422 13302 30424 13354
rect 30424 13302 30476 13354
rect 30476 13302 30478 13354
rect 30422 13300 30478 13302
rect 30526 13354 30582 13356
rect 30526 13302 30528 13354
rect 30528 13302 30580 13354
rect 30580 13302 30582 13354
rect 30526 13300 30582 13302
rect 30716 12908 30772 12964
rect 30318 11786 30374 11788
rect 30318 11734 30320 11786
rect 30320 11734 30372 11786
rect 30372 11734 30374 11786
rect 30318 11732 30374 11734
rect 30422 11786 30478 11788
rect 30422 11734 30424 11786
rect 30424 11734 30476 11786
rect 30476 11734 30478 11786
rect 30422 11732 30478 11734
rect 30526 11786 30582 11788
rect 30526 11734 30528 11786
rect 30528 11734 30580 11786
rect 30580 11734 30582 11786
rect 30526 11732 30582 11734
rect 30716 11788 30772 11844
rect 29148 10332 29204 10388
rect 29596 9996 29652 10052
rect 28252 9212 28308 9268
rect 28028 8876 28084 8932
rect 28252 7532 28308 7588
rect 27132 7250 27188 7252
rect 27132 7198 27134 7250
rect 27134 7198 27186 7250
rect 27186 7198 27188 7250
rect 27132 7196 27188 7198
rect 27020 7084 27076 7140
rect 27356 6748 27412 6804
rect 26684 6018 26740 6020
rect 26684 5966 26686 6018
rect 26686 5966 26738 6018
rect 26738 5966 26740 6018
rect 26684 5964 26740 5966
rect 26908 5964 26964 6020
rect 26124 5906 26180 5908
rect 26124 5854 26126 5906
rect 26126 5854 26178 5906
rect 26178 5854 26180 5906
rect 26124 5852 26180 5854
rect 26236 5628 26292 5684
rect 26908 5794 26964 5796
rect 26908 5742 26910 5794
rect 26910 5742 26962 5794
rect 26962 5742 26964 5794
rect 26908 5740 26964 5742
rect 26460 5404 26516 5460
rect 27580 7474 27636 7476
rect 27580 7422 27582 7474
rect 27582 7422 27634 7474
rect 27634 7422 27636 7474
rect 27580 7420 27636 7422
rect 28028 7362 28084 7364
rect 28028 7310 28030 7362
rect 28030 7310 28082 7362
rect 28082 7310 28084 7362
rect 28028 7308 28084 7310
rect 27356 5682 27412 5684
rect 27356 5630 27358 5682
rect 27358 5630 27410 5682
rect 27410 5630 27412 5682
rect 27356 5628 27412 5630
rect 28140 6972 28196 7028
rect 29484 9602 29540 9604
rect 29484 9550 29486 9602
rect 29486 9550 29538 9602
rect 29538 9550 29540 9602
rect 29484 9548 29540 9550
rect 29596 8988 29652 9044
rect 30044 10108 30100 10164
rect 30044 9938 30100 9940
rect 30044 9886 30046 9938
rect 30046 9886 30098 9938
rect 30098 9886 30100 9938
rect 30044 9884 30100 9886
rect 30318 10218 30374 10220
rect 30318 10166 30320 10218
rect 30320 10166 30372 10218
rect 30372 10166 30374 10218
rect 30318 10164 30374 10166
rect 30422 10218 30478 10220
rect 30422 10166 30424 10218
rect 30424 10166 30476 10218
rect 30476 10166 30478 10218
rect 30422 10164 30478 10166
rect 30526 10218 30582 10220
rect 30526 10166 30528 10218
rect 30528 10166 30580 10218
rect 30580 10166 30582 10218
rect 30526 10164 30582 10166
rect 32508 16604 32564 16660
rect 33292 16604 33348 16660
rect 32060 15484 32116 15540
rect 30828 10332 30884 10388
rect 31500 13580 31556 13636
rect 31388 13522 31444 13524
rect 31388 13470 31390 13522
rect 31390 13470 31442 13522
rect 31442 13470 31444 13522
rect 31388 13468 31444 13470
rect 33628 16268 33684 16324
rect 32508 15148 32564 15204
rect 32396 15036 32452 15092
rect 33628 15314 33684 15316
rect 33628 15262 33630 15314
rect 33630 15262 33682 15314
rect 33682 15262 33684 15314
rect 33628 15260 33684 15262
rect 34476 15706 34532 15708
rect 34476 15654 34478 15706
rect 34478 15654 34530 15706
rect 34530 15654 34532 15706
rect 34476 15652 34532 15654
rect 34580 15706 34636 15708
rect 34580 15654 34582 15706
rect 34582 15654 34634 15706
rect 34634 15654 34636 15706
rect 34580 15652 34636 15654
rect 34684 15706 34740 15708
rect 34684 15654 34686 15706
rect 34686 15654 34738 15706
rect 34738 15654 34740 15706
rect 34684 15652 34740 15654
rect 34188 15260 34244 15316
rect 33404 15202 33460 15204
rect 33404 15150 33406 15202
rect 33406 15150 33458 15202
rect 33458 15150 33460 15202
rect 33404 15148 33460 15150
rect 32844 14530 32900 14532
rect 32844 14478 32846 14530
rect 32846 14478 32898 14530
rect 32898 14478 32900 14530
rect 32844 14476 32900 14478
rect 34476 14138 34532 14140
rect 34476 14086 34478 14138
rect 34478 14086 34530 14138
rect 34530 14086 34532 14138
rect 34476 14084 34532 14086
rect 34580 14138 34636 14140
rect 34580 14086 34582 14138
rect 34582 14086 34634 14138
rect 34634 14086 34636 14138
rect 34580 14084 34636 14086
rect 34684 14138 34740 14140
rect 34684 14086 34686 14138
rect 34686 14086 34738 14138
rect 34738 14086 34740 14138
rect 34684 14084 34740 14086
rect 32844 13580 32900 13636
rect 31276 11788 31332 11844
rect 31388 11452 31444 11508
rect 33292 13522 33348 13524
rect 33292 13470 33294 13522
rect 33294 13470 33346 13522
rect 33346 13470 33348 13522
rect 33292 13468 33348 13470
rect 33516 13522 33572 13524
rect 33516 13470 33518 13522
rect 33518 13470 33570 13522
rect 33570 13470 33572 13522
rect 33516 13468 33572 13470
rect 34076 12962 34132 12964
rect 34076 12910 34078 12962
rect 34078 12910 34130 12962
rect 34130 12910 34132 12962
rect 34076 12908 34132 12910
rect 34476 12570 34532 12572
rect 34476 12518 34478 12570
rect 34478 12518 34530 12570
rect 34530 12518 34532 12570
rect 34476 12516 34532 12518
rect 34580 12570 34636 12572
rect 34580 12518 34582 12570
rect 34582 12518 34634 12570
rect 34634 12518 34636 12570
rect 34580 12516 34636 12518
rect 34684 12570 34740 12572
rect 34684 12518 34686 12570
rect 34686 12518 34738 12570
rect 34738 12518 34740 12570
rect 34684 12516 34740 12518
rect 30716 9996 30772 10052
rect 30828 10108 30884 10164
rect 32060 11506 32116 11508
rect 32060 11454 32062 11506
rect 32062 11454 32114 11506
rect 32114 11454 32116 11506
rect 32060 11452 32116 11454
rect 33180 10444 33236 10500
rect 31836 10332 31892 10388
rect 31612 10108 31668 10164
rect 31164 9996 31220 10052
rect 30268 9714 30324 9716
rect 30268 9662 30270 9714
rect 30270 9662 30322 9714
rect 30322 9662 30324 9714
rect 30268 9660 30324 9662
rect 29932 8370 29988 8372
rect 29932 8318 29934 8370
rect 29934 8318 29986 8370
rect 29986 8318 29988 8370
rect 29932 8316 29988 8318
rect 30604 8930 30660 8932
rect 30604 8878 30606 8930
rect 30606 8878 30658 8930
rect 30658 8878 30660 8930
rect 30604 8876 30660 8878
rect 30318 8650 30374 8652
rect 30318 8598 30320 8650
rect 30320 8598 30372 8650
rect 30372 8598 30374 8650
rect 30318 8596 30374 8598
rect 30422 8650 30478 8652
rect 30422 8598 30424 8650
rect 30424 8598 30476 8650
rect 30476 8598 30478 8650
rect 30422 8596 30478 8598
rect 30526 8650 30582 8652
rect 30526 8598 30528 8650
rect 30528 8598 30580 8650
rect 30580 8598 30582 8650
rect 30526 8596 30582 8598
rect 30380 8370 30436 8372
rect 30380 8318 30382 8370
rect 30382 8318 30434 8370
rect 30434 8318 30436 8370
rect 30380 8316 30436 8318
rect 31164 9660 31220 9716
rect 31164 9100 31220 9156
rect 29708 8204 29764 8260
rect 29484 8092 29540 8148
rect 30492 8092 30548 8148
rect 31052 8204 31108 8260
rect 29260 7474 29316 7476
rect 29260 7422 29262 7474
rect 29262 7422 29314 7474
rect 29314 7422 29316 7474
rect 29260 7420 29316 7422
rect 28588 6860 28644 6916
rect 28700 7084 28756 7140
rect 27468 5180 27524 5236
rect 27132 5068 27188 5124
rect 27916 5964 27972 6020
rect 29372 7084 29428 7140
rect 29260 6860 29316 6916
rect 27692 5906 27748 5908
rect 27692 5854 27694 5906
rect 27694 5854 27746 5906
rect 27746 5854 27748 5906
rect 27692 5852 27748 5854
rect 27804 5794 27860 5796
rect 27804 5742 27806 5794
rect 27806 5742 27858 5794
rect 27858 5742 27860 5794
rect 27804 5740 27860 5742
rect 26160 4730 26216 4732
rect 26160 4678 26162 4730
rect 26162 4678 26214 4730
rect 26214 4678 26216 4730
rect 26160 4676 26216 4678
rect 26264 4730 26320 4732
rect 26264 4678 26266 4730
rect 26266 4678 26318 4730
rect 26318 4678 26320 4730
rect 26264 4676 26320 4678
rect 26368 4730 26424 4732
rect 26368 4678 26370 4730
rect 26370 4678 26422 4730
rect 26422 4678 26424 4730
rect 26368 4676 26424 4678
rect 28588 5068 28644 5124
rect 29820 7084 29876 7140
rect 30716 7196 30772 7252
rect 30318 7082 30374 7084
rect 30318 7030 30320 7082
rect 30320 7030 30372 7082
rect 30372 7030 30374 7082
rect 30318 7028 30374 7030
rect 30422 7082 30478 7084
rect 30422 7030 30424 7082
rect 30424 7030 30476 7082
rect 30476 7030 30478 7082
rect 30422 7028 30478 7030
rect 30526 7082 30582 7084
rect 30526 7030 30528 7082
rect 30528 7030 30580 7082
rect 30580 7030 30582 7082
rect 30526 7028 30582 7030
rect 29708 6802 29764 6804
rect 29708 6750 29710 6802
rect 29710 6750 29762 6802
rect 29762 6750 29764 6802
rect 29708 6748 29764 6750
rect 30044 6748 30100 6804
rect 29596 6636 29652 6692
rect 29820 5852 29876 5908
rect 30380 6802 30436 6804
rect 30380 6750 30382 6802
rect 30382 6750 30434 6802
rect 30434 6750 30436 6802
rect 30380 6748 30436 6750
rect 30156 6690 30212 6692
rect 30156 6638 30158 6690
rect 30158 6638 30210 6690
rect 30210 6638 30212 6690
rect 30156 6636 30212 6638
rect 31500 8316 31556 8372
rect 31500 8092 31556 8148
rect 33068 10108 33124 10164
rect 31836 8988 31892 9044
rect 32396 8764 32452 8820
rect 31388 6860 31444 6916
rect 31500 7196 31556 7252
rect 30940 6076 30996 6132
rect 30604 5906 30660 5908
rect 30604 5854 30606 5906
rect 30606 5854 30658 5906
rect 30658 5854 30660 5906
rect 30604 5852 30660 5854
rect 30716 5794 30772 5796
rect 30716 5742 30718 5794
rect 30718 5742 30770 5794
rect 30770 5742 30772 5794
rect 30716 5740 30772 5742
rect 30156 5628 30212 5684
rect 30318 5514 30374 5516
rect 30318 5462 30320 5514
rect 30320 5462 30372 5514
rect 30372 5462 30374 5514
rect 30318 5460 30374 5462
rect 30422 5514 30478 5516
rect 30422 5462 30424 5514
rect 30424 5462 30476 5514
rect 30476 5462 30478 5514
rect 30422 5460 30478 5462
rect 30526 5514 30582 5516
rect 30526 5462 30528 5514
rect 30528 5462 30580 5514
rect 30580 5462 30582 5514
rect 30526 5460 30582 5462
rect 30716 5516 30772 5572
rect 30940 5292 30996 5348
rect 32172 7250 32228 7252
rect 32172 7198 32174 7250
rect 32174 7198 32226 7250
rect 32226 7198 32228 7250
rect 32172 7196 32228 7198
rect 31948 6860 32004 6916
rect 31724 5794 31780 5796
rect 31724 5742 31726 5794
rect 31726 5742 31778 5794
rect 31778 5742 31780 5794
rect 31724 5740 31780 5742
rect 31836 5516 31892 5572
rect 31164 5404 31220 5460
rect 31052 5068 31108 5124
rect 31836 5068 31892 5124
rect 29596 4898 29652 4900
rect 29596 4846 29598 4898
rect 29598 4846 29650 4898
rect 29650 4846 29652 4898
rect 29596 4844 29652 4846
rect 31164 4844 31220 4900
rect 25228 4060 25284 4116
rect 24556 3666 24612 3668
rect 24556 3614 24558 3666
rect 24558 3614 24610 3666
rect 24610 3614 24612 3666
rect 24556 3612 24612 3614
rect 22428 3500 22484 3556
rect 24892 3554 24948 3556
rect 24892 3502 24894 3554
rect 24894 3502 24946 3554
rect 24946 3502 24948 3554
rect 24892 3500 24948 3502
rect 30318 3946 30374 3948
rect 30318 3894 30320 3946
rect 30320 3894 30372 3946
rect 30372 3894 30374 3946
rect 30318 3892 30374 3894
rect 30422 3946 30478 3948
rect 30422 3894 30424 3946
rect 30424 3894 30476 3946
rect 30476 3894 30478 3946
rect 30422 3892 30478 3894
rect 30526 3946 30582 3948
rect 30526 3894 30528 3946
rect 30528 3894 30580 3946
rect 30580 3894 30582 3946
rect 30526 3892 30582 3894
rect 32508 8316 32564 8372
rect 33292 9884 33348 9940
rect 33292 9042 33348 9044
rect 33292 8990 33294 9042
rect 33294 8990 33346 9042
rect 33346 8990 33348 9042
rect 33292 8988 33348 8990
rect 34476 11002 34532 11004
rect 34476 10950 34478 11002
rect 34478 10950 34530 11002
rect 34530 10950 34532 11002
rect 34476 10948 34532 10950
rect 34580 11002 34636 11004
rect 34580 10950 34582 11002
rect 34582 10950 34634 11002
rect 34634 10950 34636 11002
rect 34580 10948 34636 10950
rect 34684 11002 34740 11004
rect 34684 10950 34686 11002
rect 34686 10950 34738 11002
rect 34738 10950 34740 11002
rect 34684 10948 34740 10950
rect 33628 9154 33684 9156
rect 33628 9102 33630 9154
rect 33630 9102 33682 9154
rect 33682 9102 33684 9154
rect 33628 9100 33684 9102
rect 33740 10220 33796 10276
rect 34188 9938 34244 9940
rect 34188 9886 34190 9938
rect 34190 9886 34242 9938
rect 34242 9886 34244 9938
rect 34188 9884 34244 9886
rect 34476 9434 34532 9436
rect 34476 9382 34478 9434
rect 34478 9382 34530 9434
rect 34530 9382 34532 9434
rect 34476 9380 34532 9382
rect 34580 9434 34636 9436
rect 34580 9382 34582 9434
rect 34582 9382 34634 9434
rect 34634 9382 34636 9434
rect 34580 9380 34636 9382
rect 34684 9434 34740 9436
rect 34684 9382 34686 9434
rect 34686 9382 34738 9434
rect 34738 9382 34740 9434
rect 34684 9380 34740 9382
rect 33180 8204 33236 8260
rect 33180 7420 33236 7476
rect 33516 7474 33572 7476
rect 33516 7422 33518 7474
rect 33518 7422 33570 7474
rect 33570 7422 33572 7474
rect 33516 7420 33572 7422
rect 33180 6860 33236 6916
rect 33292 6130 33348 6132
rect 33292 6078 33294 6130
rect 33294 6078 33346 6130
rect 33346 6078 33348 6130
rect 33292 6076 33348 6078
rect 33068 5906 33124 5908
rect 33068 5854 33070 5906
rect 33070 5854 33122 5906
rect 33122 5854 33124 5906
rect 33068 5852 33124 5854
rect 34188 8370 34244 8372
rect 34188 8318 34190 8370
rect 34190 8318 34242 8370
rect 34242 8318 34244 8370
rect 34188 8316 34244 8318
rect 34476 7866 34532 7868
rect 34476 7814 34478 7866
rect 34478 7814 34530 7866
rect 34530 7814 34532 7866
rect 34476 7812 34532 7814
rect 34580 7866 34636 7868
rect 34580 7814 34582 7866
rect 34582 7814 34634 7866
rect 34634 7814 34636 7866
rect 34580 7812 34636 7814
rect 34684 7866 34740 7868
rect 34684 7814 34686 7866
rect 34686 7814 34738 7866
rect 34738 7814 34740 7866
rect 34684 7812 34740 7814
rect 34476 6298 34532 6300
rect 34476 6246 34478 6298
rect 34478 6246 34530 6298
rect 34530 6246 34532 6298
rect 34476 6244 34532 6246
rect 34580 6298 34636 6300
rect 34580 6246 34582 6298
rect 34582 6246 34634 6298
rect 34634 6246 34636 6298
rect 34580 6244 34636 6246
rect 34684 6298 34740 6300
rect 34684 6246 34686 6298
rect 34686 6246 34738 6298
rect 34738 6246 34740 6298
rect 34684 6244 34740 6246
rect 33964 6076 34020 6132
rect 33068 5628 33124 5684
rect 33180 5292 33236 5348
rect 33404 5404 33460 5460
rect 34188 5404 34244 5460
rect 34476 4730 34532 4732
rect 34476 4678 34478 4730
rect 34478 4678 34530 4730
rect 34530 4678 34532 4730
rect 34476 4676 34532 4678
rect 34580 4730 34636 4732
rect 34580 4678 34582 4730
rect 34582 4678 34634 4730
rect 34634 4678 34636 4730
rect 34580 4676 34636 4678
rect 34684 4730 34740 4732
rect 34684 4678 34686 4730
rect 34686 4678 34738 4730
rect 34738 4678 34740 4730
rect 34684 4676 34740 4678
rect 25116 3388 25172 3444
rect 26908 3442 26964 3444
rect 26908 3390 26910 3442
rect 26910 3390 26962 3442
rect 26962 3390 26964 3442
rect 26908 3388 26964 3390
rect 30044 3442 30100 3444
rect 30044 3390 30046 3442
rect 30046 3390 30098 3442
rect 30098 3390 30100 3442
rect 30044 3388 30100 3390
rect 32284 3388 32340 3444
rect 26160 3162 26216 3164
rect 26160 3110 26162 3162
rect 26162 3110 26214 3162
rect 26214 3110 26216 3162
rect 26160 3108 26216 3110
rect 26264 3162 26320 3164
rect 26264 3110 26266 3162
rect 26266 3110 26318 3162
rect 26318 3110 26320 3162
rect 26264 3108 26320 3110
rect 26368 3162 26424 3164
rect 26368 3110 26370 3162
rect 26370 3110 26422 3162
rect 26422 3110 26424 3162
rect 26368 3108 26424 3110
rect 34476 3162 34532 3164
rect 34476 3110 34478 3162
rect 34478 3110 34530 3162
rect 34530 3110 34532 3162
rect 34476 3108 34532 3110
rect 34580 3162 34636 3164
rect 34580 3110 34582 3162
rect 34582 3110 34634 3162
rect 34634 3110 34636 3162
rect 34580 3108 34636 3110
rect 34684 3162 34740 3164
rect 34684 3110 34686 3162
rect 34686 3110 34738 3162
rect 34738 3110 34740 3162
rect 34684 3108 34740 3110
<< metal3 >>
rect 5360 32116 5370 32172
rect 5426 32116 5474 32172
rect 5530 32116 5578 32172
rect 5634 32116 5644 32172
rect 13676 32116 13686 32172
rect 13742 32116 13790 32172
rect 13846 32116 13894 32172
rect 13950 32116 13960 32172
rect 21992 32116 22002 32172
rect 22058 32116 22106 32172
rect 22162 32116 22210 32172
rect 22266 32116 22276 32172
rect 30308 32116 30318 32172
rect 30374 32116 30422 32172
rect 30478 32116 30526 32172
rect 30582 32116 30592 32172
rect 9518 31332 9528 31388
rect 9584 31332 9632 31388
rect 9688 31332 9736 31388
rect 9792 31332 9802 31388
rect 17834 31332 17844 31388
rect 17900 31332 17948 31388
rect 18004 31332 18052 31388
rect 18108 31332 18118 31388
rect 26150 31332 26160 31388
rect 26216 31332 26264 31388
rect 26320 31332 26368 31388
rect 26424 31332 26434 31388
rect 34466 31332 34476 31388
rect 34532 31332 34580 31388
rect 34636 31332 34684 31388
rect 34740 31332 34750 31388
rect 5360 30548 5370 30604
rect 5426 30548 5474 30604
rect 5530 30548 5578 30604
rect 5634 30548 5644 30604
rect 13676 30548 13686 30604
rect 13742 30548 13790 30604
rect 13846 30548 13894 30604
rect 13950 30548 13960 30604
rect 21992 30548 22002 30604
rect 22058 30548 22106 30604
rect 22162 30548 22210 30604
rect 22266 30548 22276 30604
rect 30308 30548 30318 30604
rect 30374 30548 30422 30604
rect 30478 30548 30526 30604
rect 30582 30548 30592 30604
rect 9518 29764 9528 29820
rect 9584 29764 9632 29820
rect 9688 29764 9736 29820
rect 9792 29764 9802 29820
rect 17834 29764 17844 29820
rect 17900 29764 17948 29820
rect 18004 29764 18052 29820
rect 18108 29764 18118 29820
rect 26150 29764 26160 29820
rect 26216 29764 26264 29820
rect 26320 29764 26368 29820
rect 26424 29764 26434 29820
rect 34466 29764 34476 29820
rect 34532 29764 34580 29820
rect 34636 29764 34684 29820
rect 34740 29764 34750 29820
rect 5360 28980 5370 29036
rect 5426 28980 5474 29036
rect 5530 28980 5578 29036
rect 5634 28980 5644 29036
rect 13676 28980 13686 29036
rect 13742 28980 13790 29036
rect 13846 28980 13894 29036
rect 13950 28980 13960 29036
rect 21992 28980 22002 29036
rect 22058 28980 22106 29036
rect 22162 28980 22210 29036
rect 22266 28980 22276 29036
rect 30308 28980 30318 29036
rect 30374 28980 30422 29036
rect 30478 28980 30526 29036
rect 30582 28980 30592 29036
rect 9518 28196 9528 28252
rect 9584 28196 9632 28252
rect 9688 28196 9736 28252
rect 9792 28196 9802 28252
rect 17834 28196 17844 28252
rect 17900 28196 17948 28252
rect 18004 28196 18052 28252
rect 18108 28196 18118 28252
rect 26150 28196 26160 28252
rect 26216 28196 26264 28252
rect 26320 28196 26368 28252
rect 26424 28196 26434 28252
rect 34466 28196 34476 28252
rect 34532 28196 34580 28252
rect 34636 28196 34684 28252
rect 34740 28196 34750 28252
rect 8418 27804 8428 27860
rect 8484 27804 10220 27860
rect 10276 27804 10286 27860
rect 19282 27804 19292 27860
rect 19348 27804 20300 27860
rect 20356 27804 20366 27860
rect 10994 27692 11004 27748
rect 11060 27692 12236 27748
rect 12292 27692 12302 27748
rect 5360 27412 5370 27468
rect 5426 27412 5474 27468
rect 5530 27412 5578 27468
rect 5634 27412 5644 27468
rect 13676 27412 13686 27468
rect 13742 27412 13790 27468
rect 13846 27412 13894 27468
rect 13950 27412 13960 27468
rect 21992 27412 22002 27468
rect 22058 27412 22106 27468
rect 22162 27412 22210 27468
rect 22266 27412 22276 27468
rect 30308 27412 30318 27468
rect 30374 27412 30422 27468
rect 30478 27412 30526 27468
rect 30582 27412 30592 27468
rect 5170 27244 5180 27300
rect 5236 27244 5852 27300
rect 5908 27244 5918 27300
rect 5180 27076 5236 27244
rect 17724 27132 19516 27188
rect 19572 27132 20636 27188
rect 20692 27132 20702 27188
rect 4956 27020 5236 27076
rect 5954 27020 5964 27076
rect 6020 27020 6748 27076
rect 6804 27020 6814 27076
rect 13122 27020 13132 27076
rect 13188 27020 14252 27076
rect 14308 27020 17500 27076
rect 17556 27020 17566 27076
rect 4956 26964 5012 27020
rect 17724 26964 17780 27132
rect 4946 26908 4956 26964
rect 5012 26908 5022 26964
rect 5170 26908 5180 26964
rect 5236 26908 6412 26964
rect 6468 26908 6860 26964
rect 6916 26908 6926 26964
rect 12450 26908 12460 26964
rect 12516 26908 17612 26964
rect 17668 26908 17780 26964
rect 18274 26908 18284 26964
rect 18340 26908 20636 26964
rect 20692 26908 20702 26964
rect 9518 26628 9528 26684
rect 9584 26628 9632 26684
rect 9688 26628 9736 26684
rect 9792 26628 9802 26684
rect 17834 26628 17844 26684
rect 17900 26628 17948 26684
rect 18004 26628 18052 26684
rect 18108 26628 18118 26684
rect 26150 26628 26160 26684
rect 26216 26628 26264 26684
rect 26320 26628 26368 26684
rect 26424 26628 26434 26684
rect 34466 26628 34476 26684
rect 34532 26628 34580 26684
rect 34636 26628 34684 26684
rect 34740 26628 34750 26684
rect 8082 26460 8092 26516
rect 8148 26460 8876 26516
rect 8932 26460 8942 26516
rect 2482 26348 2492 26404
rect 2548 26348 3276 26404
rect 3332 26348 3342 26404
rect 6290 26348 6300 26404
rect 6356 26348 7308 26404
rect 7364 26348 7374 26404
rect 19058 26348 19068 26404
rect 19124 26348 20300 26404
rect 20356 26348 20366 26404
rect 12338 26236 12348 26292
rect 12404 26236 13020 26292
rect 13076 26236 13086 26292
rect 17490 26236 17500 26292
rect 17556 26236 19740 26292
rect 19796 26236 19806 26292
rect 16258 26124 16268 26180
rect 16324 26124 18844 26180
rect 18900 26124 18910 26180
rect 5360 25844 5370 25900
rect 5426 25844 5474 25900
rect 5530 25844 5578 25900
rect 5634 25844 5644 25900
rect 13676 25844 13686 25900
rect 13742 25844 13790 25900
rect 13846 25844 13894 25900
rect 13950 25844 13960 25900
rect 21992 25844 22002 25900
rect 22058 25844 22106 25900
rect 22162 25844 22210 25900
rect 22266 25844 22276 25900
rect 30308 25844 30318 25900
rect 30374 25844 30422 25900
rect 30478 25844 30526 25900
rect 30582 25844 30592 25900
rect 12338 25676 12348 25732
rect 12404 25676 14252 25732
rect 14308 25676 14318 25732
rect 20290 25676 20300 25732
rect 20356 25676 22876 25732
rect 22932 25676 22942 25732
rect 12674 25564 12684 25620
rect 12740 25564 13580 25620
rect 13636 25564 13646 25620
rect 14130 25564 14140 25620
rect 14196 25564 16660 25620
rect 19506 25564 19516 25620
rect 19572 25564 20524 25620
rect 20580 25564 21980 25620
rect 22036 25564 22046 25620
rect 23090 25564 23100 25620
rect 23156 25564 24556 25620
rect 24612 25564 26348 25620
rect 26404 25564 26414 25620
rect 1810 25452 1820 25508
rect 1876 25452 7084 25508
rect 7140 25452 7420 25508
rect 7476 25452 7980 25508
rect 8036 25452 8046 25508
rect 13010 25452 13020 25508
rect 13076 25452 13692 25508
rect 13748 25452 13758 25508
rect 14690 25452 14700 25508
rect 14756 25452 15484 25508
rect 15540 25452 15550 25508
rect 14700 25396 14756 25452
rect 4610 25340 4620 25396
rect 4676 25340 5068 25396
rect 5124 25340 5852 25396
rect 5908 25340 5918 25396
rect 10994 25340 11004 25396
rect 11060 25340 14756 25396
rect 14914 25340 14924 25396
rect 14980 25340 16268 25396
rect 16324 25340 16334 25396
rect 16604 25284 16660 25564
rect 18834 25452 18844 25508
rect 18900 25452 19852 25508
rect 19908 25452 19918 25508
rect 20066 25452 20076 25508
rect 20132 25452 20748 25508
rect 20804 25452 21644 25508
rect 21700 25452 22652 25508
rect 22708 25452 22718 25508
rect 19506 25340 19516 25396
rect 19572 25340 20860 25396
rect 20916 25340 21756 25396
rect 21812 25340 21822 25396
rect 22530 25340 22540 25396
rect 22596 25340 23548 25396
rect 23604 25340 23614 25396
rect 25554 25340 25564 25396
rect 25620 25340 26460 25396
rect 26516 25340 26526 25396
rect 16594 25228 16604 25284
rect 16660 25228 16940 25284
rect 16996 25228 17500 25284
rect 17556 25228 17566 25284
rect 19282 25228 19292 25284
rect 19348 25228 22988 25284
rect 23044 25228 23772 25284
rect 23828 25228 23838 25284
rect 25442 25228 25452 25284
rect 25508 25228 25788 25284
rect 25844 25228 26796 25284
rect 26852 25228 27244 25284
rect 27300 25228 27310 25284
rect 15250 25116 15260 25172
rect 15316 25116 15708 25172
rect 15764 25116 16380 25172
rect 16436 25116 16446 25172
rect 9518 25060 9528 25116
rect 9584 25060 9632 25116
rect 9688 25060 9736 25116
rect 9792 25060 9802 25116
rect 17834 25060 17844 25116
rect 17900 25060 17948 25116
rect 18004 25060 18052 25116
rect 18108 25060 18118 25116
rect 26150 25060 26160 25116
rect 26216 25060 26264 25116
rect 26320 25060 26368 25116
rect 26424 25060 26434 25116
rect 34466 25060 34476 25116
rect 34532 25060 34580 25116
rect 34636 25060 34684 25116
rect 34740 25060 34750 25116
rect 3266 24892 3276 24948
rect 3332 24836 3388 24948
rect 9986 24892 9996 24948
rect 10052 24892 11116 24948
rect 11172 24892 11182 24948
rect 12338 24892 12348 24948
rect 12404 24892 12852 24948
rect 22754 24892 22764 24948
rect 22820 24892 23212 24948
rect 23268 24892 23660 24948
rect 23716 24892 23726 24948
rect 12796 24836 12852 24892
rect 3332 24780 4060 24836
rect 4116 24780 4126 24836
rect 5058 24780 5068 24836
rect 5124 24780 5964 24836
rect 6020 24780 6636 24836
rect 6692 24780 6702 24836
rect 11778 24780 11788 24836
rect 11844 24780 12516 24836
rect 12786 24780 12796 24836
rect 12852 24780 12862 24836
rect 13458 24780 13468 24836
rect 13524 24780 18172 24836
rect 18228 24780 18238 24836
rect 12460 24724 12516 24780
rect 4610 24668 4620 24724
rect 4676 24668 5628 24724
rect 5684 24668 5694 24724
rect 12198 24668 12236 24724
rect 12292 24668 12302 24724
rect 12460 24668 12684 24724
rect 12740 24668 13244 24724
rect 13300 24668 13310 24724
rect 13458 24668 13468 24724
rect 13524 24668 14588 24724
rect 14644 24668 14654 24724
rect 23090 24668 23100 24724
rect 23156 24668 23884 24724
rect 23940 24668 23950 24724
rect 24434 24668 24444 24724
rect 24500 24668 26348 24724
rect 26404 24668 26414 24724
rect 12002 24556 12012 24612
rect 12068 24556 12460 24612
rect 12516 24556 12526 24612
rect 14130 24556 14140 24612
rect 14196 24556 20188 24612
rect 20244 24556 20254 24612
rect 4386 24444 4396 24500
rect 4452 24444 6188 24500
rect 6244 24444 6636 24500
rect 6692 24444 6702 24500
rect 12114 24444 12124 24500
rect 12180 24444 12348 24500
rect 12404 24444 12414 24500
rect 21970 24444 21980 24500
rect 22036 24444 23212 24500
rect 23268 24444 25116 24500
rect 25172 24444 25182 24500
rect 10210 24332 10220 24388
rect 10276 24332 11116 24388
rect 11172 24332 11182 24388
rect 14130 24332 14140 24388
rect 14196 24332 15260 24388
rect 15316 24332 15326 24388
rect 5360 24276 5370 24332
rect 5426 24276 5474 24332
rect 5530 24276 5578 24332
rect 5634 24276 5644 24332
rect 13676 24276 13686 24332
rect 13742 24276 13790 24332
rect 13846 24276 13894 24332
rect 13950 24276 13960 24332
rect 21992 24276 22002 24332
rect 22058 24276 22106 24332
rect 22162 24276 22210 24332
rect 22266 24276 22276 24332
rect 30308 24276 30318 24332
rect 30374 24276 30422 24332
rect 30478 24276 30526 24332
rect 30582 24276 30592 24332
rect 7746 24108 7756 24164
rect 7812 24108 8876 24164
rect 8932 24108 8942 24164
rect 8978 23996 8988 24052
rect 9044 23996 11004 24052
rect 11060 23996 11070 24052
rect 11666 23996 11676 24052
rect 11732 23996 15372 24052
rect 15428 23996 15438 24052
rect 26114 23996 26124 24052
rect 26180 23996 26684 24052
rect 26740 23996 26750 24052
rect 12226 23884 12236 23940
rect 12292 23884 12572 23940
rect 12628 23884 12638 23940
rect 12786 23884 12796 23940
rect 12852 23884 12890 23940
rect 14700 23884 15596 23940
rect 15652 23884 15662 23940
rect 11330 23772 11340 23828
rect 11396 23772 12012 23828
rect 12068 23772 12078 23828
rect 12338 23772 12348 23828
rect 12404 23772 12684 23828
rect 12740 23772 12750 23828
rect 13570 23772 13580 23828
rect 13636 23772 14028 23828
rect 14084 23772 14094 23828
rect 14700 23716 14756 23884
rect 15922 23772 15932 23828
rect 15988 23772 17164 23828
rect 17220 23772 17230 23828
rect 25666 23772 25676 23828
rect 25732 23772 26684 23828
rect 26740 23772 26750 23828
rect 11778 23660 11788 23716
rect 11844 23660 13692 23716
rect 13748 23660 13758 23716
rect 13906 23660 13916 23716
rect 13972 23660 14700 23716
rect 14756 23660 14766 23716
rect 15092 23660 18284 23716
rect 18340 23660 19292 23716
rect 19348 23660 19358 23716
rect 25778 23660 25788 23716
rect 25844 23660 26348 23716
rect 26404 23660 26908 23716
rect 26964 23660 26974 23716
rect 4050 23548 4060 23604
rect 4116 23548 5404 23604
rect 5460 23548 5470 23604
rect 9986 23548 9996 23604
rect 10052 23548 11676 23604
rect 11732 23548 13468 23604
rect 13524 23548 14476 23604
rect 14532 23548 14542 23604
rect 9518 23492 9528 23548
rect 9584 23492 9632 23548
rect 9688 23492 9736 23548
rect 9792 23492 9802 23548
rect 15092 23492 15148 23660
rect 17834 23492 17844 23548
rect 17900 23492 17948 23548
rect 18004 23492 18052 23548
rect 18108 23492 18118 23548
rect 26150 23492 26160 23548
rect 26216 23492 26264 23548
rect 26320 23492 26368 23548
rect 26424 23492 26434 23548
rect 34466 23492 34476 23548
rect 34532 23492 34580 23548
rect 34636 23492 34684 23548
rect 34740 23492 34750 23548
rect 12898 23436 12908 23492
rect 12964 23436 13916 23492
rect 13972 23436 15148 23492
rect 15362 23436 15372 23492
rect 15428 23436 17668 23492
rect 17612 23380 17668 23436
rect 9986 23324 9996 23380
rect 10052 23324 12124 23380
rect 12180 23324 12190 23380
rect 14578 23324 14588 23380
rect 14644 23324 17388 23380
rect 17444 23324 17454 23380
rect 17612 23324 17836 23380
rect 17892 23324 19068 23380
rect 19124 23324 19134 23380
rect 25218 23324 25228 23380
rect 25284 23324 26348 23380
rect 26404 23324 26414 23380
rect 12124 23268 12180 23324
rect 4946 23212 4956 23268
rect 5012 23212 6188 23268
rect 6244 23212 6254 23268
rect 12124 23212 13132 23268
rect 13188 23212 14812 23268
rect 14868 23212 15820 23268
rect 15876 23212 15886 23268
rect 18946 23212 18956 23268
rect 19012 23212 20300 23268
rect 20356 23212 20366 23268
rect 24322 23212 24332 23268
rect 24388 23212 25116 23268
rect 25172 23212 26908 23268
rect 27010 23212 27020 23268
rect 27076 23212 29148 23268
rect 29204 23212 29214 23268
rect 6626 23100 6636 23156
rect 6692 23100 14588 23156
rect 14644 23100 14654 23156
rect 18162 23100 18172 23156
rect 18228 23100 18844 23156
rect 18900 23100 19516 23156
rect 19572 23100 19740 23156
rect 19796 23100 19806 23156
rect 24434 23100 24444 23156
rect 24500 23100 26124 23156
rect 26180 23100 26190 23156
rect 26852 23100 26908 23212
rect 26964 23100 26974 23156
rect 2818 22988 2828 23044
rect 2884 22988 6748 23044
rect 6804 22988 6814 23044
rect 8978 22988 8988 23044
rect 9044 22988 12572 23044
rect 12628 22988 12638 23044
rect 14578 22988 14588 23044
rect 14644 22988 14924 23044
rect 14980 22988 14990 23044
rect 17714 22988 17724 23044
rect 17780 22988 18732 23044
rect 18788 22988 18798 23044
rect 9874 22876 9884 22932
rect 9940 22876 11452 22932
rect 11508 22876 12684 22932
rect 12740 22876 12750 22932
rect 13906 22876 13916 22932
rect 13972 22876 14364 22932
rect 14420 22876 14430 22932
rect 16034 22876 16044 22932
rect 16100 22876 19516 22932
rect 19572 22876 19582 22932
rect 24658 22764 24668 22820
rect 24724 22764 26796 22820
rect 26852 22764 26908 22820
rect 26964 22764 26974 22820
rect 5360 22708 5370 22764
rect 5426 22708 5474 22764
rect 5530 22708 5578 22764
rect 5634 22708 5644 22764
rect 13676 22708 13686 22764
rect 13742 22708 13790 22764
rect 13846 22708 13894 22764
rect 13950 22708 13960 22764
rect 21992 22708 22002 22764
rect 22058 22708 22106 22764
rect 22162 22708 22210 22764
rect 22266 22708 22276 22764
rect 30308 22708 30318 22764
rect 30374 22708 30422 22764
rect 30478 22708 30526 22764
rect 30582 22708 30592 22764
rect 7074 22428 7084 22484
rect 7140 22428 7868 22484
rect 7924 22428 7934 22484
rect 3602 22316 3612 22372
rect 3668 22316 6076 22372
rect 6132 22316 6142 22372
rect 12674 22316 12684 22372
rect 12740 22316 13468 22372
rect 13524 22316 13534 22372
rect 20290 22316 20300 22372
rect 20356 22316 21084 22372
rect 21140 22316 25228 22372
rect 25284 22316 25294 22372
rect 26338 22316 26348 22372
rect 26404 22316 27020 22372
rect 27076 22316 27086 22372
rect 2482 22204 2492 22260
rect 2548 22204 5628 22260
rect 5684 22204 5694 22260
rect 8530 22204 8540 22260
rect 8596 22204 13580 22260
rect 13636 22204 13646 22260
rect 20626 22204 20636 22260
rect 20692 22204 22092 22260
rect 22148 22204 22158 22260
rect 12898 22092 12908 22148
rect 12964 22092 15036 22148
rect 15092 22092 19964 22148
rect 20020 22092 20030 22148
rect 26562 22092 26572 22148
rect 26628 22092 26796 22148
rect 26852 22092 27468 22148
rect 27524 22092 27534 22148
rect 12114 21980 12124 22036
rect 12180 21980 13020 22036
rect 13076 21980 13086 22036
rect 18722 21980 18732 22036
rect 18788 21980 19292 22036
rect 19348 21980 19358 22036
rect 9518 21924 9528 21980
rect 9584 21924 9632 21980
rect 9688 21924 9736 21980
rect 9792 21924 9802 21980
rect 17834 21924 17844 21980
rect 17900 21924 17948 21980
rect 18004 21924 18052 21980
rect 18108 21924 18118 21980
rect 26150 21924 26160 21980
rect 26216 21924 26264 21980
rect 26320 21924 26368 21980
rect 26424 21924 26434 21980
rect 34466 21924 34476 21980
rect 34532 21924 34580 21980
rect 34636 21924 34684 21980
rect 34740 21924 34750 21980
rect 12338 21868 12348 21924
rect 12404 21868 12414 21924
rect 14690 21868 14700 21924
rect 14756 21868 15260 21924
rect 15316 21868 15932 21924
rect 15988 21868 15998 21924
rect 21298 21868 21308 21924
rect 21364 21868 21980 21924
rect 22036 21868 22046 21924
rect 10658 21756 10668 21812
rect 10724 21756 12012 21812
rect 12068 21756 12078 21812
rect 12348 21700 12404 21868
rect 14466 21756 14476 21812
rect 14532 21756 15708 21812
rect 15764 21756 15774 21812
rect 16818 21756 16828 21812
rect 16884 21756 18396 21812
rect 18452 21756 18462 21812
rect 19954 21756 19964 21812
rect 20020 21756 22876 21812
rect 22932 21756 22942 21812
rect 3938 21644 3948 21700
rect 4004 21644 4620 21700
rect 4676 21644 5404 21700
rect 5460 21644 5470 21700
rect 10994 21644 11004 21700
rect 11060 21644 12404 21700
rect 13458 21644 13468 21700
rect 13524 21644 14812 21700
rect 14868 21644 14878 21700
rect 19618 21644 19628 21700
rect 19684 21644 20636 21700
rect 20692 21644 21756 21700
rect 21812 21644 21822 21700
rect 22082 21644 22092 21700
rect 22148 21644 22540 21700
rect 22596 21644 24220 21700
rect 24276 21644 24286 21700
rect 25666 21644 25676 21700
rect 25732 21644 26124 21700
rect 26180 21644 26190 21700
rect 12338 21532 12348 21588
rect 12404 21532 12796 21588
rect 12852 21532 12862 21588
rect 20514 21532 20524 21588
rect 20580 21532 22428 21588
rect 22484 21532 22494 21588
rect 24434 21532 24444 21588
rect 24500 21532 26572 21588
rect 26628 21532 26638 21588
rect 12450 21420 12460 21476
rect 12516 21420 15372 21476
rect 15428 21420 15438 21476
rect 15586 21420 15596 21476
rect 15652 21420 17612 21476
rect 17668 21420 18172 21476
rect 18228 21420 20692 21476
rect 20850 21420 20860 21476
rect 20916 21420 21756 21476
rect 21812 21420 24108 21476
rect 24164 21420 24174 21476
rect 24658 21420 24668 21476
rect 24724 21420 25900 21476
rect 25956 21420 25966 21476
rect 20636 21364 20692 21420
rect 10770 21308 10780 21364
rect 10836 21308 12572 21364
rect 12628 21308 12638 21364
rect 12796 21308 16492 21364
rect 16548 21308 19740 21364
rect 19796 21308 20300 21364
rect 20356 21308 20366 21364
rect 20636 21308 22652 21364
rect 22708 21308 22718 21364
rect 26114 21308 26124 21364
rect 26180 21308 27580 21364
rect 27636 21308 27646 21364
rect 12796 21252 12852 21308
rect 11330 21196 11340 21252
rect 11396 21196 12852 21252
rect 5360 21140 5370 21196
rect 5426 21140 5474 21196
rect 5530 21140 5578 21196
rect 5634 21140 5644 21196
rect 13676 21140 13686 21196
rect 13742 21140 13790 21196
rect 13846 21140 13894 21196
rect 13950 21140 13960 21196
rect 21992 21140 22002 21196
rect 22058 21140 22106 21196
rect 22162 21140 22210 21196
rect 22266 21140 22276 21196
rect 30308 21140 30318 21196
rect 30374 21140 30422 21196
rect 30478 21140 30526 21196
rect 30582 21140 30592 21196
rect 12674 20972 12684 21028
rect 12740 20972 15484 21028
rect 15540 20972 15550 21028
rect 15810 20860 15820 20916
rect 15876 20860 16716 20916
rect 16772 20860 16782 20916
rect 25890 20860 25900 20916
rect 25956 20860 26684 20916
rect 26740 20860 26750 20916
rect 28018 20860 28028 20916
rect 28084 20860 28700 20916
rect 28756 20860 28766 20916
rect 3266 20748 3276 20804
rect 3332 20748 4732 20804
rect 4788 20748 7644 20804
rect 7700 20748 7710 20804
rect 10770 20748 10780 20804
rect 10836 20748 12348 20804
rect 12404 20748 12414 20804
rect 14354 20748 14364 20804
rect 14420 20748 16044 20804
rect 16100 20748 16110 20804
rect 21858 20748 21868 20804
rect 21924 20748 23100 20804
rect 23156 20748 24556 20804
rect 24612 20748 26012 20804
rect 26068 20748 26078 20804
rect 14364 20692 14420 20748
rect 3938 20636 3948 20692
rect 4004 20636 4844 20692
rect 4900 20636 8204 20692
rect 8260 20636 8270 20692
rect 11442 20636 11452 20692
rect 11508 20636 12684 20692
rect 12740 20636 14420 20692
rect 17714 20636 17724 20692
rect 17780 20636 21308 20692
rect 21364 20636 21374 20692
rect 2370 20524 2380 20580
rect 2436 20524 2940 20580
rect 2996 20524 3388 20580
rect 3444 20524 4284 20580
rect 4340 20524 5068 20580
rect 5124 20524 5134 20580
rect 12786 20524 12796 20580
rect 12852 20524 13580 20580
rect 13636 20524 14140 20580
rect 14196 20524 14206 20580
rect 17500 20524 17836 20580
rect 17892 20524 17902 20580
rect 17500 20468 17556 20524
rect 17490 20412 17500 20468
rect 17556 20412 17566 20468
rect 9518 20356 9528 20412
rect 9584 20356 9632 20412
rect 9688 20356 9736 20412
rect 9792 20356 9802 20412
rect 17834 20356 17844 20412
rect 17900 20356 17948 20412
rect 18004 20356 18052 20412
rect 18108 20356 18118 20412
rect 26150 20356 26160 20412
rect 26216 20356 26264 20412
rect 26320 20356 26368 20412
rect 26424 20356 26434 20412
rect 34466 20356 34476 20412
rect 34532 20356 34580 20412
rect 34636 20356 34684 20412
rect 34740 20356 34750 20412
rect 8194 20188 8204 20244
rect 8260 20188 10220 20244
rect 10276 20188 10286 20244
rect 12114 20188 12124 20244
rect 12180 20188 12190 20244
rect 17836 20188 25676 20244
rect 25732 20188 25742 20244
rect 12124 20132 12180 20188
rect 17836 20132 17892 20188
rect 4386 20076 4396 20132
rect 4452 20076 5516 20132
rect 5572 20076 5582 20132
rect 11330 20076 11340 20132
rect 11396 20076 12180 20132
rect 13010 20076 13020 20132
rect 13076 20076 13580 20132
rect 13636 20076 14252 20132
rect 14308 20076 14318 20132
rect 16930 20076 16940 20132
rect 16996 20076 17892 20132
rect 23986 20076 23996 20132
rect 24052 20076 26572 20132
rect 26628 20076 26638 20132
rect 3602 19964 3612 20020
rect 3668 19964 4508 20020
rect 4564 19964 5292 20020
rect 5348 19964 5358 20020
rect 7420 19964 8876 20020
rect 8932 19964 9436 20020
rect 9492 19964 9502 20020
rect 9986 19964 9996 20020
rect 10052 19964 10444 20020
rect 10500 19964 12572 20020
rect 12628 19964 12638 20020
rect 16370 19964 16380 20020
rect 16436 19964 18172 20020
rect 18228 19964 19068 20020
rect 19124 19964 19134 20020
rect 19506 19964 19516 20020
rect 19572 19964 20300 20020
rect 20356 19964 20366 20020
rect 7420 19908 7476 19964
rect 2594 19852 2604 19908
rect 2660 19852 5180 19908
rect 5236 19852 5246 19908
rect 6738 19852 6748 19908
rect 6804 19852 7420 19908
rect 7476 19852 7486 19908
rect 7970 19852 7980 19908
rect 8036 19852 9660 19908
rect 9716 19852 9726 19908
rect 9996 19796 10052 19964
rect 14018 19852 14028 19908
rect 14084 19852 15260 19908
rect 15316 19852 16604 19908
rect 16660 19852 18396 19908
rect 18452 19852 18462 19908
rect 21186 19852 21196 19908
rect 21252 19852 21868 19908
rect 21924 19852 21934 19908
rect 8866 19740 8876 19796
rect 8932 19740 10052 19796
rect 14690 19740 14700 19796
rect 14756 19740 15932 19796
rect 15988 19740 15998 19796
rect 17938 19740 17948 19796
rect 18004 19740 18844 19796
rect 18900 19740 18910 19796
rect 10658 19628 10668 19684
rect 10724 19628 12572 19684
rect 12628 19628 12638 19684
rect 13458 19628 13468 19684
rect 13524 19628 13534 19684
rect 18050 19628 18060 19684
rect 18116 19628 18508 19684
rect 18564 19628 18574 19684
rect 5360 19572 5370 19628
rect 5426 19572 5474 19628
rect 5530 19572 5578 19628
rect 5634 19572 5644 19628
rect 13468 19572 13524 19628
rect 13676 19572 13686 19628
rect 13742 19572 13790 19628
rect 13846 19572 13894 19628
rect 13950 19572 13960 19628
rect 21992 19572 22002 19628
rect 22058 19572 22106 19628
rect 22162 19572 22210 19628
rect 22266 19572 22276 19628
rect 30308 19572 30318 19628
rect 30374 19572 30422 19628
rect 30478 19572 30526 19628
rect 30582 19572 30592 19628
rect 10210 19516 10220 19572
rect 10276 19516 13524 19572
rect 4946 19404 4956 19460
rect 5012 19404 13916 19460
rect 13972 19404 13982 19460
rect 8978 19292 8988 19348
rect 9044 19292 10556 19348
rect 10612 19292 10622 19348
rect 12226 19292 12236 19348
rect 12292 19292 13356 19348
rect 13412 19292 13422 19348
rect 17378 19292 17388 19348
rect 17444 19292 18396 19348
rect 18452 19292 19964 19348
rect 20020 19292 20412 19348
rect 20468 19292 20478 19348
rect 10658 19180 10668 19236
rect 10724 19180 11116 19236
rect 11172 19180 11182 19236
rect 9090 19068 9100 19124
rect 9156 19068 10556 19124
rect 10612 19068 10622 19124
rect 9762 18956 9772 19012
rect 9828 18956 10780 19012
rect 10836 18956 10846 19012
rect 9518 18788 9528 18844
rect 9584 18788 9632 18844
rect 9688 18788 9736 18844
rect 9792 18788 9802 18844
rect 17834 18788 17844 18844
rect 17900 18788 17948 18844
rect 18004 18788 18052 18844
rect 18108 18788 18118 18844
rect 26150 18788 26160 18844
rect 26216 18788 26264 18844
rect 26320 18788 26368 18844
rect 26424 18788 26434 18844
rect 34466 18788 34476 18844
rect 34532 18788 34580 18844
rect 34636 18788 34684 18844
rect 34740 18788 34750 18844
rect 6962 18732 6972 18788
rect 7028 18732 8204 18788
rect 8260 18732 8270 18788
rect 10332 18732 11452 18788
rect 11508 18732 11518 18788
rect 10332 18676 10388 18732
rect 7410 18620 7420 18676
rect 7476 18620 10388 18676
rect 10546 18620 10556 18676
rect 10612 18620 11900 18676
rect 11956 18620 11966 18676
rect 18834 18620 18844 18676
rect 18900 18620 21644 18676
rect 21700 18620 21710 18676
rect 22642 18620 22652 18676
rect 22708 18620 23324 18676
rect 23380 18620 23390 18676
rect 7970 18508 7980 18564
rect 8036 18508 8876 18564
rect 8932 18508 8942 18564
rect 9100 18508 9660 18564
rect 9716 18508 9726 18564
rect 10556 18508 11340 18564
rect 11396 18508 12124 18564
rect 12180 18508 12190 18564
rect 16818 18508 16828 18564
rect 16884 18508 17500 18564
rect 17556 18508 17566 18564
rect 9100 18452 9156 18508
rect 10556 18452 10612 18508
rect 4610 18396 4620 18452
rect 4676 18396 5628 18452
rect 5684 18396 6412 18452
rect 6468 18396 6478 18452
rect 6626 18396 6636 18452
rect 6692 18396 7308 18452
rect 7364 18396 9156 18452
rect 10546 18396 10556 18452
rect 10612 18396 10622 18452
rect 11442 18396 11452 18452
rect 11508 18396 11900 18452
rect 11956 18396 11966 18452
rect 14018 18396 14028 18452
rect 14084 18396 18732 18452
rect 18788 18396 18798 18452
rect 22866 18396 22876 18452
rect 22932 18396 26236 18452
rect 26292 18396 27244 18452
rect 27300 18396 27310 18452
rect 5842 18284 5852 18340
rect 5908 18284 7084 18340
rect 7140 18284 7644 18340
rect 7700 18284 8316 18340
rect 8372 18284 8382 18340
rect 9874 18284 9884 18340
rect 9940 18284 12348 18340
rect 12404 18284 12414 18340
rect 14690 18284 14700 18340
rect 14756 18284 16044 18340
rect 16100 18284 16110 18340
rect 16482 18284 16492 18340
rect 16548 18284 17500 18340
rect 17556 18284 17566 18340
rect 22082 18284 22092 18340
rect 22148 18284 23660 18340
rect 23716 18284 23726 18340
rect 25666 18284 25676 18340
rect 25732 18284 29260 18340
rect 29316 18284 29326 18340
rect 6290 18172 6300 18228
rect 6356 18172 6860 18228
rect 6916 18172 6926 18228
rect 8866 18172 8876 18228
rect 8932 18172 10108 18228
rect 10164 18172 10174 18228
rect 10994 18172 11004 18228
rect 11060 18172 11788 18228
rect 11844 18172 12908 18228
rect 12964 18172 12974 18228
rect 18050 18172 18060 18228
rect 18116 18172 22988 18228
rect 23044 18172 23054 18228
rect 8082 18060 8092 18116
rect 8148 18060 12796 18116
rect 12852 18060 12862 18116
rect 5360 18004 5370 18060
rect 5426 18004 5474 18060
rect 5530 18004 5578 18060
rect 5634 18004 5644 18060
rect 13676 18004 13686 18060
rect 13742 18004 13790 18060
rect 13846 18004 13894 18060
rect 13950 18004 13960 18060
rect 21992 18004 22002 18060
rect 22058 18004 22106 18060
rect 22162 18004 22210 18060
rect 22266 18004 22276 18060
rect 30308 18004 30318 18060
rect 30374 18004 30422 18060
rect 30478 18004 30526 18060
rect 30582 18004 30592 18060
rect 8194 17948 8204 18004
rect 8260 17948 9660 18004
rect 9716 17948 9726 18004
rect 26674 17948 26684 18004
rect 26740 17948 28476 18004
rect 28532 17948 28542 18004
rect 8418 17836 8428 17892
rect 8484 17836 9548 17892
rect 9604 17836 9614 17892
rect 26226 17836 26236 17892
rect 26292 17836 27916 17892
rect 27972 17836 28140 17892
rect 28196 17836 28588 17892
rect 28644 17836 28654 17892
rect 7410 17724 7420 17780
rect 7476 17724 8260 17780
rect 6178 17612 6188 17668
rect 6244 17612 7084 17668
rect 7140 17612 7868 17668
rect 7924 17612 7934 17668
rect 8204 17556 8260 17724
rect 8530 17612 8540 17668
rect 8596 17612 10220 17668
rect 10276 17612 10286 17668
rect 26852 17612 29148 17668
rect 29204 17612 29214 17668
rect 29586 17612 29596 17668
rect 29652 17612 31388 17668
rect 31444 17612 31948 17668
rect 32004 17612 32014 17668
rect 26852 17556 26908 17612
rect 8194 17500 8204 17556
rect 8260 17500 8270 17556
rect 9090 17500 9100 17556
rect 9156 17500 10668 17556
rect 10724 17500 10734 17556
rect 14354 17500 14364 17556
rect 14420 17500 16156 17556
rect 16212 17500 17164 17556
rect 17220 17500 17836 17556
rect 17892 17500 17902 17556
rect 18162 17500 18172 17556
rect 18228 17500 18956 17556
rect 19012 17500 19022 17556
rect 26002 17500 26012 17556
rect 26068 17500 26908 17556
rect 28914 17500 28924 17556
rect 28980 17500 31276 17556
rect 31332 17500 31342 17556
rect 9762 17388 9772 17444
rect 9828 17388 11116 17444
rect 11172 17388 11182 17444
rect 17714 17388 17724 17444
rect 17780 17388 18396 17444
rect 18452 17388 18462 17444
rect 19058 17388 19068 17444
rect 19124 17388 20636 17444
rect 20692 17388 20702 17444
rect 7410 17276 7420 17332
rect 7476 17276 7486 17332
rect 9874 17276 9884 17332
rect 9940 17276 11228 17332
rect 11284 17276 11294 17332
rect 17154 17276 17164 17332
rect 17220 17276 17612 17332
rect 17668 17276 17678 17332
rect 7420 17108 7476 17276
rect 9518 17220 9528 17276
rect 9584 17220 9632 17276
rect 9688 17220 9736 17276
rect 9792 17220 9802 17276
rect 17834 17220 17844 17276
rect 17900 17220 17948 17276
rect 18004 17220 18052 17276
rect 18108 17220 18118 17276
rect 26150 17220 26160 17276
rect 26216 17220 26264 17276
rect 26320 17220 26368 17276
rect 26424 17220 26434 17276
rect 34466 17220 34476 17276
rect 34532 17220 34580 17276
rect 34636 17220 34684 17276
rect 34740 17220 34750 17276
rect 7420 17052 10444 17108
rect 10500 17052 10510 17108
rect 17042 17052 17052 17108
rect 17108 17052 17948 17108
rect 18004 17052 18014 17108
rect 15092 16940 15932 16996
rect 15988 16940 16716 16996
rect 16772 16940 17836 16996
rect 17892 16940 17902 16996
rect 15092 16884 15148 16940
rect 3938 16828 3948 16884
rect 4004 16828 5068 16884
rect 5124 16828 5134 16884
rect 5292 16828 6748 16884
rect 6804 16828 7532 16884
rect 7588 16828 7598 16884
rect 10770 16828 10780 16884
rect 10836 16828 12124 16884
rect 12180 16828 12190 16884
rect 12898 16828 12908 16884
rect 12964 16828 14140 16884
rect 14196 16828 15148 16884
rect 15250 16828 15260 16884
rect 15316 16828 17276 16884
rect 17332 16828 17342 16884
rect 5292 16772 5348 16828
rect 5068 16716 5348 16772
rect 12226 16716 12236 16772
rect 12292 16716 14028 16772
rect 14084 16716 14094 16772
rect 16492 16716 17612 16772
rect 17668 16716 18508 16772
rect 18564 16716 18574 16772
rect 27234 16716 27244 16772
rect 27300 16716 27580 16772
rect 27636 16716 28140 16772
rect 28196 16716 28206 16772
rect 30370 16716 30380 16772
rect 30436 16716 31948 16772
rect 32004 16716 32014 16772
rect 5068 16660 5124 16716
rect 16492 16660 16548 16716
rect 5058 16604 5068 16660
rect 5124 16604 5134 16660
rect 13906 16604 13916 16660
rect 13972 16604 15260 16660
rect 15316 16604 15326 16660
rect 16482 16604 16492 16660
rect 16548 16604 16558 16660
rect 16706 16604 16716 16660
rect 16772 16604 19068 16660
rect 19124 16604 19134 16660
rect 31714 16604 31724 16660
rect 31780 16604 32508 16660
rect 32564 16604 33292 16660
rect 33348 16604 33358 16660
rect 5360 16436 5370 16492
rect 5426 16436 5474 16492
rect 5530 16436 5578 16492
rect 5634 16436 5644 16492
rect 13676 16436 13686 16492
rect 13742 16436 13790 16492
rect 13846 16436 13894 16492
rect 13950 16436 13960 16492
rect 21992 16436 22002 16492
rect 22058 16436 22106 16492
rect 22162 16436 22210 16492
rect 22266 16436 22276 16492
rect 30308 16436 30318 16492
rect 30374 16436 30422 16492
rect 30478 16436 30526 16492
rect 30582 16436 30592 16492
rect 15894 16380 15932 16436
rect 15988 16380 15998 16436
rect 14802 16268 14812 16324
rect 14868 16268 14878 16324
rect 17042 16268 17052 16324
rect 17108 16268 17948 16324
rect 18004 16268 18014 16324
rect 28354 16268 28364 16324
rect 28420 16268 30716 16324
rect 30772 16268 33628 16324
rect 33684 16268 33694 16324
rect 12786 16156 12796 16212
rect 12852 16156 13692 16212
rect 13748 16156 13758 16212
rect 14812 16100 14868 16268
rect 21634 16156 21644 16212
rect 21700 16156 23436 16212
rect 23492 16156 23502 16212
rect 26898 16156 26908 16212
rect 26964 16156 28028 16212
rect 28084 16156 28094 16212
rect 14812 16044 15260 16100
rect 15316 16044 18620 16100
rect 18676 16044 18686 16100
rect 21746 16044 21756 16100
rect 21812 16044 22428 16100
rect 22484 16044 23660 16100
rect 23716 16044 23726 16100
rect 25890 16044 25900 16100
rect 25956 16044 27020 16100
rect 27076 16044 27086 16100
rect 14130 15932 14140 15988
rect 14196 15932 14700 15988
rect 14756 15932 14766 15988
rect 15138 15932 15148 15988
rect 15204 15932 16044 15988
rect 16100 15932 16110 15988
rect 16370 15932 16380 15988
rect 16436 15932 16716 15988
rect 16772 15932 16782 15988
rect 16930 15932 16940 15988
rect 16996 15932 18508 15988
rect 18564 15932 18574 15988
rect 22642 15932 22652 15988
rect 22708 15932 24332 15988
rect 24388 15932 24398 15988
rect 14802 15820 14812 15876
rect 14868 15820 15484 15876
rect 15540 15820 15550 15876
rect 18274 15820 18284 15876
rect 18340 15820 18844 15876
rect 18900 15820 18910 15876
rect 27346 15820 27356 15876
rect 27412 15820 30940 15876
rect 30996 15820 31006 15876
rect 15138 15708 15148 15764
rect 15204 15708 15708 15764
rect 15764 15708 16828 15764
rect 16884 15708 16894 15764
rect 9518 15652 9528 15708
rect 9584 15652 9632 15708
rect 9688 15652 9736 15708
rect 9792 15652 9802 15708
rect 17834 15652 17844 15708
rect 17900 15652 17948 15708
rect 18004 15652 18052 15708
rect 18108 15652 18118 15708
rect 26150 15652 26160 15708
rect 26216 15652 26264 15708
rect 26320 15652 26368 15708
rect 26424 15652 26434 15708
rect 34466 15652 34476 15708
rect 34532 15652 34580 15708
rect 34636 15652 34684 15708
rect 34740 15652 34750 15708
rect 27682 15596 27692 15652
rect 27748 15596 28476 15652
rect 28532 15596 28542 15652
rect 27570 15484 27580 15540
rect 27636 15484 29372 15540
rect 29428 15484 29438 15540
rect 29698 15484 29708 15540
rect 29764 15484 32060 15540
rect 32116 15484 32126 15540
rect 14690 15372 14700 15428
rect 14756 15372 15596 15428
rect 15652 15372 15662 15428
rect 20132 15372 22876 15428
rect 22932 15372 22942 15428
rect 29250 15372 29260 15428
rect 29316 15372 30044 15428
rect 30100 15372 31500 15428
rect 31556 15372 31566 15428
rect 11218 15260 11228 15316
rect 11284 15260 13468 15316
rect 13524 15260 13534 15316
rect 14018 15260 14028 15316
rect 14084 15260 15260 15316
rect 15316 15260 17836 15316
rect 17892 15260 17902 15316
rect 1586 15148 1596 15204
rect 1652 15148 17948 15204
rect 18004 15148 18014 15204
rect 20132 15092 20188 15372
rect 30370 15260 30380 15316
rect 30436 15260 31052 15316
rect 31108 15260 31388 15316
rect 31444 15260 33628 15316
rect 33684 15260 34188 15316
rect 34244 15260 34254 15316
rect 21746 15148 21756 15204
rect 21812 15148 22876 15204
rect 22932 15148 24556 15204
rect 24612 15148 24622 15204
rect 30594 15148 30604 15204
rect 30660 15148 32508 15204
rect 32564 15148 33404 15204
rect 33460 15148 33470 15204
rect 1810 15036 1820 15092
rect 1876 15036 2268 15092
rect 2324 15036 3276 15092
rect 3332 15036 3342 15092
rect 8978 15036 8988 15092
rect 9044 15036 9996 15092
rect 10052 15036 10062 15092
rect 17266 15036 17276 15092
rect 17332 15036 20188 15092
rect 28578 15036 28588 15092
rect 28644 15036 29820 15092
rect 29876 15036 29886 15092
rect 30482 15036 30492 15092
rect 30548 15036 32396 15092
rect 32452 15036 32462 15092
rect 5360 14868 5370 14924
rect 5426 14868 5474 14924
rect 5530 14868 5578 14924
rect 5634 14868 5644 14924
rect 13676 14868 13686 14924
rect 13742 14868 13790 14924
rect 13846 14868 13894 14924
rect 13950 14868 13960 14924
rect 21992 14868 22002 14924
rect 22058 14868 22106 14924
rect 22162 14868 22210 14924
rect 22266 14868 22276 14924
rect 30308 14868 30318 14924
rect 30374 14868 30422 14924
rect 30478 14868 30526 14924
rect 30582 14868 30592 14924
rect 16146 14700 16156 14756
rect 16212 14700 16604 14756
rect 16660 14700 16670 14756
rect 4610 14588 4620 14644
rect 4676 14588 5628 14644
rect 5684 14588 5694 14644
rect 15810 14588 15820 14644
rect 15876 14588 16492 14644
rect 16548 14588 16558 14644
rect 21522 14588 21532 14644
rect 21588 14588 23436 14644
rect 23492 14588 23502 14644
rect 28802 14588 28812 14644
rect 28868 14588 29596 14644
rect 29652 14588 31948 14644
rect 31892 14532 31948 14588
rect 16370 14476 16380 14532
rect 16436 14476 17052 14532
rect 17108 14476 17388 14532
rect 17444 14476 17454 14532
rect 28018 14476 28028 14532
rect 28084 14476 29484 14532
rect 29540 14476 29550 14532
rect 31892 14476 32844 14532
rect 32900 14476 32910 14532
rect 20066 14364 20076 14420
rect 20132 14364 22204 14420
rect 22260 14364 22270 14420
rect 2930 14252 2940 14308
rect 2996 14252 3500 14308
rect 3556 14252 3566 14308
rect 5954 14252 5964 14308
rect 6020 14252 6860 14308
rect 6916 14252 6926 14308
rect 12674 14252 12684 14308
rect 12740 14252 13580 14308
rect 13636 14252 17276 14308
rect 17332 14252 17342 14308
rect 20514 14252 20524 14308
rect 20580 14252 21420 14308
rect 21476 14252 21486 14308
rect 27234 14252 27244 14308
rect 27300 14252 27804 14308
rect 27860 14252 27870 14308
rect 15586 14140 15596 14196
rect 15652 14140 15820 14196
rect 15876 14140 17388 14196
rect 17444 14140 17454 14196
rect 9518 14084 9528 14140
rect 9584 14084 9632 14140
rect 9688 14084 9736 14140
rect 9792 14084 9802 14140
rect 17834 14084 17844 14140
rect 17900 14084 17948 14140
rect 18004 14084 18052 14140
rect 18108 14084 18118 14140
rect 26150 14084 26160 14140
rect 26216 14084 26264 14140
rect 26320 14084 26368 14140
rect 26424 14084 26434 14140
rect 34466 14084 34476 14140
rect 34532 14084 34580 14140
rect 34636 14084 34684 14140
rect 34740 14084 34750 14140
rect 3266 14028 3276 14084
rect 3332 14028 5068 14084
rect 5124 14028 5964 14084
rect 6020 14028 8428 14084
rect 8484 14028 8494 14084
rect 7746 13916 7756 13972
rect 7812 13916 11900 13972
rect 11956 13916 11966 13972
rect 18386 13916 18396 13972
rect 18452 13916 19628 13972
rect 19684 13916 20188 13972
rect 20244 13916 20254 13972
rect 25666 13916 25676 13972
rect 25732 13916 26684 13972
rect 26740 13916 27020 13972
rect 27076 13916 27086 13972
rect 10546 13804 10556 13860
rect 10612 13804 11788 13860
rect 11844 13804 11854 13860
rect 16482 13804 16492 13860
rect 16548 13804 17948 13860
rect 18004 13804 18014 13860
rect 18162 13804 18172 13860
rect 18228 13804 19404 13860
rect 19460 13804 19470 13860
rect 25442 13804 25452 13860
rect 25508 13804 28588 13860
rect 28644 13804 28654 13860
rect 25452 13748 25508 13804
rect 6962 13692 6972 13748
rect 7028 13692 10332 13748
rect 10388 13692 12124 13748
rect 12180 13692 12190 13748
rect 17714 13692 17724 13748
rect 17780 13692 18732 13748
rect 18788 13692 18798 13748
rect 19058 13692 19068 13748
rect 19124 13692 20076 13748
rect 20132 13692 20142 13748
rect 23874 13692 23884 13748
rect 23940 13692 25508 13748
rect 26114 13692 26124 13748
rect 26180 13692 27468 13748
rect 27524 13692 27534 13748
rect 5618 13580 5628 13636
rect 5684 13580 10164 13636
rect 21410 13580 21420 13636
rect 21476 13580 22036 13636
rect 26450 13580 26460 13636
rect 26516 13580 27244 13636
rect 27300 13580 27310 13636
rect 27794 13580 27804 13636
rect 27860 13580 29708 13636
rect 29764 13580 29774 13636
rect 31490 13580 31500 13636
rect 31556 13580 32844 13636
rect 32900 13580 33572 13636
rect 10108 13524 10164 13580
rect 21980 13524 22036 13580
rect 33516 13524 33572 13580
rect 2482 13468 2492 13524
rect 2548 13468 6636 13524
rect 6692 13468 6702 13524
rect 10098 13468 10108 13524
rect 10164 13468 12236 13524
rect 12292 13468 12302 13524
rect 19506 13468 19516 13524
rect 19572 13468 21308 13524
rect 21364 13468 21374 13524
rect 21970 13468 21980 13524
rect 22036 13468 22988 13524
rect 23044 13468 23054 13524
rect 24770 13468 24780 13524
rect 24836 13468 26908 13524
rect 26964 13468 26974 13524
rect 27346 13468 27356 13524
rect 27412 13468 28252 13524
rect 28308 13468 28318 13524
rect 31378 13468 31388 13524
rect 31444 13468 33292 13524
rect 33348 13468 33358 13524
rect 33506 13468 33516 13524
rect 33572 13468 33582 13524
rect 5740 13356 6412 13412
rect 6468 13356 8652 13412
rect 8708 13356 8718 13412
rect 26338 13356 26348 13412
rect 26404 13356 27580 13412
rect 27636 13356 27646 13412
rect 5360 13300 5370 13356
rect 5426 13300 5474 13356
rect 5530 13300 5578 13356
rect 5634 13300 5644 13356
rect 5740 13188 5796 13356
rect 13676 13300 13686 13356
rect 13742 13300 13790 13356
rect 13846 13300 13894 13356
rect 13950 13300 13960 13356
rect 21992 13300 22002 13356
rect 22058 13300 22106 13356
rect 22162 13300 22210 13356
rect 22266 13300 22276 13356
rect 30308 13300 30318 13356
rect 30374 13300 30422 13356
rect 30478 13300 30526 13356
rect 30582 13300 30592 13356
rect 26674 13244 26684 13300
rect 26740 13244 29148 13300
rect 29204 13244 29214 13300
rect 5058 13132 5068 13188
rect 5124 13132 5796 13188
rect 6402 13132 6412 13188
rect 6468 13132 7084 13188
rect 7140 13132 7756 13188
rect 7812 13132 7822 13188
rect 19058 13132 19068 13188
rect 19124 13132 19852 13188
rect 19908 13132 19918 13188
rect 20290 13132 20300 13188
rect 20356 13132 22092 13188
rect 22148 13132 22652 13188
rect 22708 13132 22718 13188
rect 2818 13020 2828 13076
rect 2884 13020 7420 13076
rect 7476 13020 8540 13076
rect 8596 13020 8606 13076
rect 11890 13020 11900 13076
rect 11956 13020 15372 13076
rect 15428 13020 16380 13076
rect 16436 13020 16446 13076
rect 20066 13020 20076 13076
rect 20132 13020 20748 13076
rect 20804 13020 22316 13076
rect 22372 13020 22382 13076
rect 5618 12908 5628 12964
rect 5684 12908 6748 12964
rect 6804 12908 6814 12964
rect 8418 12908 8428 12964
rect 8484 12908 12572 12964
rect 12628 12908 12638 12964
rect 17938 12908 17948 12964
rect 18004 12908 18844 12964
rect 18900 12908 18910 12964
rect 20514 12908 20524 12964
rect 20580 12908 21868 12964
rect 21924 12908 21934 12964
rect 30706 12908 30716 12964
rect 30772 12908 34076 12964
rect 34132 12908 34142 12964
rect 11004 12796 13804 12852
rect 13860 12796 13870 12852
rect 14130 12796 14140 12852
rect 14196 12796 14924 12852
rect 14980 12796 14990 12852
rect 11004 12740 11060 12796
rect 20972 12740 21028 12908
rect 21634 12796 21644 12852
rect 21700 12796 22876 12852
rect 22932 12796 22942 12852
rect 3378 12684 3388 12740
rect 3444 12684 4732 12740
rect 4788 12684 5292 12740
rect 5348 12684 5358 12740
rect 6850 12684 6860 12740
rect 6916 12684 7196 12740
rect 7252 12684 11004 12740
rect 11060 12684 11070 12740
rect 11330 12684 11340 12740
rect 11396 12684 12012 12740
rect 12068 12684 12078 12740
rect 18162 12684 18172 12740
rect 18228 12684 19740 12740
rect 19796 12684 19806 12740
rect 20962 12684 20972 12740
rect 21028 12684 21038 12740
rect 22418 12684 22428 12740
rect 22484 12684 23660 12740
rect 23716 12684 23726 12740
rect 19282 12572 19292 12628
rect 19348 12572 19852 12628
rect 19908 12572 19918 12628
rect 9518 12516 9528 12572
rect 9584 12516 9632 12572
rect 9688 12516 9736 12572
rect 9792 12516 9802 12572
rect 17834 12516 17844 12572
rect 17900 12516 17948 12572
rect 18004 12516 18052 12572
rect 18108 12516 18118 12572
rect 26150 12516 26160 12572
rect 26216 12516 26264 12572
rect 26320 12516 26368 12572
rect 26424 12516 26434 12572
rect 34466 12516 34476 12572
rect 34532 12516 34580 12572
rect 34636 12516 34684 12572
rect 34740 12516 34750 12572
rect 5618 12348 5628 12404
rect 5684 12348 6412 12404
rect 6468 12348 6478 12404
rect 6626 12348 6636 12404
rect 6692 12348 7084 12404
rect 7140 12348 7150 12404
rect 7522 12348 7532 12404
rect 7588 12348 9884 12404
rect 9940 12348 10892 12404
rect 10948 12348 10958 12404
rect 18498 12348 18508 12404
rect 18564 12348 19964 12404
rect 20020 12348 20636 12404
rect 20692 12348 20702 12404
rect 3602 12236 3612 12292
rect 3668 12236 4508 12292
rect 4564 12236 6076 12292
rect 6132 12236 6142 12292
rect 6738 12236 6748 12292
rect 6804 12236 7308 12292
rect 7364 12236 7374 12292
rect 8978 12236 8988 12292
rect 9044 12236 10556 12292
rect 10612 12236 10622 12292
rect 17602 12236 17612 12292
rect 17668 12236 18396 12292
rect 18452 12236 19404 12292
rect 19460 12236 19470 12292
rect 2034 12124 2044 12180
rect 2100 12124 2828 12180
rect 2884 12124 2894 12180
rect 3490 12124 3500 12180
rect 3556 12124 4732 12180
rect 4788 12124 4798 12180
rect 4946 12124 4956 12180
rect 5012 12124 5852 12180
rect 5908 12124 5918 12180
rect 4386 12012 4396 12068
rect 4452 12012 7980 12068
rect 8036 12012 8046 12068
rect 18722 12012 18732 12068
rect 18788 12012 19404 12068
rect 19460 12012 19470 12068
rect 3938 11900 3948 11956
rect 4004 11900 6076 11956
rect 6132 11900 6142 11956
rect 4582 11788 4620 11844
rect 4676 11788 4686 11844
rect 30706 11788 30716 11844
rect 30772 11788 31276 11844
rect 31332 11788 31342 11844
rect 5360 11732 5370 11788
rect 5426 11732 5474 11788
rect 5530 11732 5578 11788
rect 5634 11732 5644 11788
rect 13676 11732 13686 11788
rect 13742 11732 13790 11788
rect 13846 11732 13894 11788
rect 13950 11732 13960 11788
rect 21992 11732 22002 11788
rect 22058 11732 22106 11788
rect 22162 11732 22210 11788
rect 22266 11732 22276 11788
rect 30308 11732 30318 11788
rect 30374 11732 30422 11788
rect 30478 11732 30526 11788
rect 30582 11732 30592 11788
rect 4498 11676 4508 11732
rect 4564 11676 4956 11732
rect 5012 11676 5022 11732
rect 7410 11676 7420 11732
rect 7476 11676 7868 11732
rect 7924 11676 8316 11732
rect 8372 11676 11340 11732
rect 11396 11676 11406 11732
rect 19618 11676 19628 11732
rect 19684 11676 20076 11732
rect 20132 11676 21308 11732
rect 21364 11676 21374 11732
rect 3938 11564 3948 11620
rect 4004 11564 4732 11620
rect 4788 11564 4798 11620
rect 6962 11564 6972 11620
rect 7028 11564 8652 11620
rect 8708 11564 8718 11620
rect 8866 11564 8876 11620
rect 8932 11564 11116 11620
rect 11172 11564 11182 11620
rect 19842 11564 19852 11620
rect 19908 11564 20412 11620
rect 20468 11564 20478 11620
rect 3042 11452 3052 11508
rect 3108 11452 5572 11508
rect 10658 11452 10668 11508
rect 10724 11452 14252 11508
rect 14308 11452 14318 11508
rect 21522 11452 21532 11508
rect 21588 11452 22876 11508
rect 22932 11452 22942 11508
rect 31378 11452 31388 11508
rect 31444 11452 32060 11508
rect 32116 11452 32126 11508
rect 5516 11396 5572 11452
rect 2146 11340 2156 11396
rect 2212 11340 3500 11396
rect 3556 11340 3566 11396
rect 5506 11340 5516 11396
rect 5572 11340 5582 11396
rect 6290 11340 6300 11396
rect 6356 11340 7084 11396
rect 7140 11340 7150 11396
rect 9090 11340 9100 11396
rect 9156 11340 10444 11396
rect 10500 11340 10510 11396
rect 4274 11228 4284 11284
rect 4340 11228 4620 11284
rect 4676 11228 4686 11284
rect 5842 11228 5852 11284
rect 5908 11228 7420 11284
rect 7476 11228 7486 11284
rect 7858 11228 7868 11284
rect 7924 11228 9660 11284
rect 9716 11228 9726 11284
rect 10770 11228 10780 11284
rect 10836 11228 13020 11284
rect 13076 11228 13086 11284
rect 2594 11116 2604 11172
rect 2660 11116 3612 11172
rect 3668 11116 3678 11172
rect 8876 11116 9548 11172
rect 9604 11116 9614 11172
rect 17378 11116 17388 11172
rect 17444 11116 17724 11172
rect 17780 11116 17790 11172
rect 8876 11060 8932 11116
rect 3266 11004 3276 11060
rect 3332 11004 6076 11060
rect 6132 11004 8876 11060
rect 8932 11004 8942 11060
rect 9518 10948 9528 11004
rect 9584 10948 9632 11004
rect 9688 10948 9736 11004
rect 9792 10948 9802 11004
rect 17834 10948 17844 11004
rect 17900 10948 17948 11004
rect 18004 10948 18052 11004
rect 18108 10948 18118 11004
rect 26150 10948 26160 11004
rect 26216 10948 26264 11004
rect 26320 10948 26368 11004
rect 26424 10948 26434 11004
rect 34466 10948 34476 11004
rect 34532 10948 34580 11004
rect 34636 10948 34684 11004
rect 34740 10948 34750 11004
rect 7858 10892 7868 10948
rect 7924 10892 8988 10948
rect 9044 10892 9054 10948
rect 16482 10780 16492 10836
rect 16548 10780 17388 10836
rect 17444 10780 18284 10836
rect 18340 10780 18350 10836
rect 21522 10780 21532 10836
rect 21588 10780 27132 10836
rect 27188 10780 27198 10836
rect 4274 10668 4284 10724
rect 4340 10668 9324 10724
rect 9380 10668 9996 10724
rect 10052 10668 10062 10724
rect 17490 10668 17500 10724
rect 17556 10668 18396 10724
rect 18452 10668 18732 10724
rect 18788 10668 18798 10724
rect 4386 10556 4396 10612
rect 4452 10556 5068 10612
rect 5124 10556 6300 10612
rect 6356 10556 6366 10612
rect 8082 10556 8092 10612
rect 8148 10556 9548 10612
rect 9604 10556 9614 10612
rect 16594 10556 16604 10612
rect 16660 10556 18844 10612
rect 18900 10556 18910 10612
rect 22306 10556 22316 10612
rect 22372 10556 23212 10612
rect 23268 10556 26908 10612
rect 26964 10556 26974 10612
rect 8194 10444 8204 10500
rect 8260 10444 10220 10500
rect 10276 10444 10286 10500
rect 17826 10444 17836 10500
rect 17892 10444 18956 10500
rect 19012 10444 19022 10500
rect 31892 10444 33180 10500
rect 33236 10444 33246 10500
rect 5058 10332 5068 10388
rect 5124 10332 5516 10388
rect 5572 10332 5582 10388
rect 9314 10332 9324 10388
rect 9380 10332 10668 10388
rect 10724 10332 10734 10388
rect 12338 10332 12348 10388
rect 12404 10332 13468 10388
rect 13524 10332 14924 10388
rect 14980 10332 14990 10388
rect 29138 10332 29148 10388
rect 29204 10332 30828 10388
rect 30884 10332 30894 10388
rect 31826 10332 31836 10388
rect 31892 10332 31948 10444
rect 30716 10276 30772 10332
rect 30716 10220 33740 10276
rect 33796 10220 33806 10276
rect 5360 10164 5370 10220
rect 5426 10164 5474 10220
rect 5530 10164 5578 10220
rect 5634 10164 5644 10220
rect 13676 10164 13686 10220
rect 13742 10164 13790 10220
rect 13846 10164 13894 10220
rect 13950 10164 13960 10220
rect 21992 10164 22002 10220
rect 22058 10164 22106 10220
rect 22162 10164 22210 10220
rect 22266 10164 22276 10220
rect 30308 10164 30318 10220
rect 30374 10164 30422 10220
rect 30478 10164 30526 10220
rect 30582 10164 30592 10220
rect 9874 10108 9884 10164
rect 9940 10108 11116 10164
rect 11172 10108 11182 10164
rect 16258 10108 16268 10164
rect 16324 10108 17276 10164
rect 17332 10108 19292 10164
rect 19348 10108 19358 10164
rect 30034 10108 30044 10164
rect 30100 10108 30110 10164
rect 30818 10108 30828 10164
rect 30884 10108 31612 10164
rect 31668 10108 33068 10164
rect 33124 10108 33134 10164
rect 30044 10052 30100 10108
rect 2706 9996 2716 10052
rect 2772 9996 3276 10052
rect 3332 9996 3948 10052
rect 4004 9996 4014 10052
rect 4610 9996 4620 10052
rect 4676 9996 7196 10052
rect 7252 9996 7262 10052
rect 7522 9996 7532 10052
rect 7588 9996 9212 10052
rect 9268 9996 9278 10052
rect 9538 9996 9548 10052
rect 9604 9996 11452 10052
rect 11508 9996 11518 10052
rect 29586 9996 29596 10052
rect 29652 9996 30100 10052
rect 30706 9996 30716 10052
rect 30772 9996 31164 10052
rect 31220 9996 31230 10052
rect 6262 9884 6300 9940
rect 6356 9884 6366 9940
rect 9314 9884 9324 9940
rect 9380 9884 10668 9940
rect 10724 9884 10734 9940
rect 11218 9884 11228 9940
rect 11284 9884 11900 9940
rect 11956 9884 11966 9940
rect 12226 9884 12236 9940
rect 12292 9884 14476 9940
rect 14532 9884 14542 9940
rect 19842 9884 19852 9940
rect 19908 9884 20412 9940
rect 20468 9884 20478 9940
rect 30034 9884 30044 9940
rect 30100 9884 33292 9940
rect 33348 9884 34188 9940
rect 34244 9884 34254 9940
rect 2594 9772 2604 9828
rect 2660 9772 3164 9828
rect 3220 9772 5628 9828
rect 5684 9772 5694 9828
rect 7858 9772 7868 9828
rect 7924 9772 9548 9828
rect 9604 9772 9614 9828
rect 12898 9772 12908 9828
rect 12964 9772 16940 9828
rect 16996 9772 17836 9828
rect 17892 9772 17902 9828
rect 3490 9660 3500 9716
rect 3556 9660 4620 9716
rect 4676 9660 4686 9716
rect 6178 9660 6188 9716
rect 6244 9660 8540 9716
rect 8596 9660 8606 9716
rect 10434 9660 10444 9716
rect 10500 9660 10780 9716
rect 10836 9660 10846 9716
rect 11778 9660 11788 9716
rect 11844 9660 13804 9716
rect 13860 9660 15036 9716
rect 15092 9660 15102 9716
rect 18610 9660 18620 9716
rect 18676 9660 18844 9716
rect 18900 9660 21420 9716
rect 21476 9660 21644 9716
rect 21700 9660 21710 9716
rect 22866 9660 22876 9716
rect 22932 9660 24332 9716
rect 24388 9660 24398 9716
rect 30258 9660 30268 9716
rect 30324 9660 31164 9716
rect 31220 9660 31230 9716
rect 3042 9548 3052 9604
rect 3108 9548 3612 9604
rect 3668 9548 3678 9604
rect 4722 9548 4732 9604
rect 4788 9548 12012 9604
rect 12068 9548 12078 9604
rect 12338 9548 12348 9604
rect 12404 9548 13580 9604
rect 13636 9548 14028 9604
rect 14084 9548 14094 9604
rect 24658 9548 24668 9604
rect 24724 9548 26964 9604
rect 27794 9548 27804 9604
rect 27860 9548 29484 9604
rect 29540 9548 29550 9604
rect 12012 9492 12068 9548
rect 3490 9436 3500 9492
rect 3556 9436 4844 9492
rect 4900 9436 5740 9492
rect 5796 9436 5806 9492
rect 8194 9436 8204 9492
rect 8260 9436 9100 9492
rect 9156 9436 9166 9492
rect 12012 9436 12572 9492
rect 12628 9436 13692 9492
rect 13748 9436 13758 9492
rect 9518 9380 9528 9436
rect 9584 9380 9632 9436
rect 9688 9380 9736 9436
rect 9792 9380 9802 9436
rect 17834 9380 17844 9436
rect 17900 9380 17948 9436
rect 18004 9380 18052 9436
rect 18108 9380 18118 9436
rect 26150 9380 26160 9436
rect 26216 9380 26264 9436
rect 26320 9380 26368 9436
rect 26424 9380 26434 9436
rect 9874 9324 9884 9380
rect 9940 9324 9950 9380
rect 9884 9268 9940 9324
rect 2930 9212 2940 9268
rect 2996 9212 4620 9268
rect 4676 9212 4686 9268
rect 4834 9212 4844 9268
rect 4900 9212 6860 9268
rect 6916 9212 6926 9268
rect 9650 9212 9660 9268
rect 9716 9212 9940 9268
rect 10658 9212 10668 9268
rect 10724 9212 11452 9268
rect 11508 9212 11518 9268
rect 22082 9212 22092 9268
rect 22148 9212 24556 9268
rect 24612 9212 26012 9268
rect 26068 9212 26078 9268
rect 2034 9100 2044 9156
rect 2100 9100 2492 9156
rect 2548 9100 2558 9156
rect 2818 9100 2828 9156
rect 2884 9100 3388 9156
rect 3332 9044 3388 9100
rect 6412 9100 7756 9156
rect 7812 9100 7822 9156
rect 16258 9100 16268 9156
rect 16324 9100 17276 9156
rect 17332 9100 17342 9156
rect 18050 9100 18060 9156
rect 18116 9100 18844 9156
rect 18900 9100 18910 9156
rect 6412 9044 6468 9100
rect 3332 8988 3612 9044
rect 3668 8988 3678 9044
rect 3938 8988 3948 9044
rect 4004 8988 6412 9044
rect 6468 8988 6478 9044
rect 6626 8988 6636 9044
rect 6692 8988 8428 9044
rect 8484 8988 8494 9044
rect 8978 8988 8988 9044
rect 9044 8988 10108 9044
rect 10164 8988 10174 9044
rect 15026 8988 15036 9044
rect 15092 8932 15148 9044
rect 20962 8988 20972 9044
rect 21028 8988 22876 9044
rect 22932 8988 22942 9044
rect 5506 8876 5516 8932
rect 5572 8876 6524 8932
rect 6580 8876 6590 8932
rect 15092 8876 19068 8932
rect 19124 8876 19134 8932
rect 21858 8876 21868 8932
rect 21924 8876 23884 8932
rect 23940 8876 23950 8932
rect 26908 8820 26964 9548
rect 34466 9380 34476 9436
rect 34532 9380 34580 9436
rect 34636 9380 34684 9436
rect 34740 9380 34750 9436
rect 27122 9212 27132 9268
rect 27188 9212 28252 9268
rect 28308 9212 28318 9268
rect 31154 9100 31164 9156
rect 31220 9100 33628 9156
rect 33684 9100 33694 9156
rect 29586 8988 29596 9044
rect 29652 8988 31836 9044
rect 31892 8988 33292 9044
rect 33348 8988 33358 9044
rect 28018 8876 28028 8932
rect 28084 8876 30604 8932
rect 30660 8876 30670 8932
rect 7074 8764 7084 8820
rect 7140 8764 7644 8820
rect 7700 8764 9548 8820
rect 9604 8764 9614 8820
rect 11442 8764 11452 8820
rect 11508 8764 11900 8820
rect 11956 8764 13356 8820
rect 13412 8764 13422 8820
rect 26908 8764 32396 8820
rect 32452 8764 32462 8820
rect 2146 8652 2156 8708
rect 2212 8652 3836 8708
rect 3892 8652 3902 8708
rect 7298 8652 7308 8708
rect 7364 8652 12236 8708
rect 12292 8652 12908 8708
rect 12964 8652 12974 8708
rect 5360 8596 5370 8652
rect 5426 8596 5474 8652
rect 5530 8596 5578 8652
rect 5634 8596 5644 8652
rect 13676 8596 13686 8652
rect 13742 8596 13790 8652
rect 13846 8596 13894 8652
rect 13950 8596 13960 8652
rect 21992 8596 22002 8652
rect 22058 8596 22106 8652
rect 22162 8596 22210 8652
rect 22266 8596 22276 8652
rect 30308 8596 30318 8652
rect 30374 8596 30422 8652
rect 30478 8596 30526 8652
rect 30582 8596 30592 8652
rect 11778 8540 11788 8596
rect 11844 8540 12292 8596
rect 5842 8428 5852 8484
rect 5908 8428 7084 8484
rect 7140 8428 7150 8484
rect 7298 8428 7308 8484
rect 7364 8428 7402 8484
rect 9660 8428 10556 8484
rect 10612 8428 10622 8484
rect 9660 8372 9716 8428
rect 4050 8316 4060 8372
rect 4116 8316 5628 8372
rect 5684 8316 9716 8372
rect 9874 8316 9884 8372
rect 9940 8316 11340 8372
rect 11396 8316 11406 8372
rect 3602 8204 3612 8260
rect 3668 8204 4732 8260
rect 4788 8204 4798 8260
rect 4946 8204 4956 8260
rect 5012 8204 5852 8260
rect 5908 8204 5918 8260
rect 6934 8204 6972 8260
rect 7028 8204 7038 8260
rect 12236 8148 12292 8540
rect 12562 8428 12572 8484
rect 12628 8428 12908 8484
rect 12964 8428 15372 8484
rect 15428 8428 15438 8484
rect 20962 8428 20972 8484
rect 21028 8428 21038 8484
rect 20972 8372 21028 8428
rect 12786 8316 12796 8372
rect 12852 8316 16268 8372
rect 16324 8316 16334 8372
rect 18722 8316 18732 8372
rect 18788 8316 19628 8372
rect 19684 8316 21028 8372
rect 29922 8316 29932 8372
rect 29988 8316 30380 8372
rect 30436 8316 30446 8372
rect 31490 8316 31500 8372
rect 31556 8316 32508 8372
rect 32564 8316 34188 8372
rect 34244 8316 34254 8372
rect 16482 8204 16492 8260
rect 16548 8204 18508 8260
rect 18564 8204 19068 8260
rect 19124 8204 19134 8260
rect 29698 8204 29708 8260
rect 29764 8204 31052 8260
rect 31108 8204 33180 8260
rect 33236 8204 33246 8260
rect 2818 8092 2828 8148
rect 2884 8092 3388 8148
rect 3444 8092 3454 8148
rect 4386 8092 4396 8148
rect 4452 8092 6524 8148
rect 6580 8092 6590 8148
rect 9762 8092 9772 8148
rect 9828 8092 9996 8148
rect 10052 8092 10062 8148
rect 12226 8092 12236 8148
rect 12292 8092 12302 8148
rect 12674 8092 12684 8148
rect 12740 8092 14924 8148
rect 14980 8092 14990 8148
rect 29474 8092 29484 8148
rect 29540 8092 30492 8148
rect 30548 8092 31500 8148
rect 31556 8092 31566 8148
rect 3332 7924 3388 8092
rect 5618 7980 5628 8036
rect 5684 7980 5740 8036
rect 5796 7980 10108 8036
rect 10164 7980 10174 8036
rect 13122 7980 13132 8036
rect 13188 7980 14140 8036
rect 14196 7980 14206 8036
rect 21746 7980 21756 8036
rect 21812 7980 23324 8036
rect 23380 7980 23390 8036
rect 3332 7868 3948 7924
rect 4004 7868 4014 7924
rect 4274 7868 4284 7924
rect 4340 7868 6860 7924
rect 6916 7868 9324 7924
rect 9380 7868 9390 7924
rect 9518 7812 9528 7868
rect 9584 7812 9632 7868
rect 9688 7812 9736 7868
rect 9792 7812 9802 7868
rect 17834 7812 17844 7868
rect 17900 7812 17948 7868
rect 18004 7812 18052 7868
rect 18108 7812 18118 7868
rect 26150 7812 26160 7868
rect 26216 7812 26264 7868
rect 26320 7812 26368 7868
rect 26424 7812 26434 7868
rect 34466 7812 34476 7868
rect 34532 7812 34580 7868
rect 34636 7812 34684 7868
rect 34740 7812 34750 7868
rect 2482 7756 2492 7812
rect 2548 7756 3276 7812
rect 3332 7588 3388 7812
rect 4498 7644 4508 7700
rect 4564 7644 6076 7700
rect 6132 7644 6142 7700
rect 6850 7644 6860 7700
rect 6916 7644 7868 7700
rect 7924 7644 7934 7700
rect 8866 7644 8876 7700
rect 8932 7644 9996 7700
rect 10052 7644 10062 7700
rect 13234 7644 13244 7700
rect 13300 7644 14364 7700
rect 14420 7644 16716 7700
rect 16772 7644 16782 7700
rect 3332 7532 10332 7588
rect 10388 7532 11004 7588
rect 11060 7532 11070 7588
rect 14130 7532 14140 7588
rect 14196 7532 15708 7588
rect 15764 7532 16044 7588
rect 16100 7532 16110 7588
rect 26002 7532 26012 7588
rect 26068 7532 28252 7588
rect 28308 7532 28318 7588
rect 4722 7420 4732 7476
rect 4788 7420 5292 7476
rect 5348 7420 5358 7476
rect 5730 7420 5740 7476
rect 5796 7420 6188 7476
rect 6244 7420 6254 7476
rect 7186 7420 7196 7476
rect 7252 7420 11676 7476
rect 11732 7420 11742 7476
rect 12002 7420 12012 7476
rect 12068 7420 15484 7476
rect 15540 7420 15550 7476
rect 16482 7420 16492 7476
rect 16548 7420 16558 7476
rect 21634 7420 21644 7476
rect 21700 7420 22204 7476
rect 22260 7420 22540 7476
rect 22596 7420 22606 7476
rect 22978 7420 22988 7476
rect 23044 7420 26236 7476
rect 26292 7420 26796 7476
rect 26852 7420 26862 7476
rect 27570 7420 27580 7476
rect 27636 7420 29260 7476
rect 29316 7420 29326 7476
rect 33170 7420 33180 7476
rect 33236 7420 33516 7476
rect 33572 7420 33582 7476
rect 16492 7364 16548 7420
rect 2146 7308 2156 7364
rect 2212 7308 2604 7364
rect 2660 7308 4172 7364
rect 4228 7308 4238 7364
rect 6962 7308 6972 7364
rect 7028 7308 8204 7364
rect 8260 7308 9996 7364
rect 10052 7308 11228 7364
rect 11284 7308 11294 7364
rect 13906 7308 13916 7364
rect 13972 7308 16156 7364
rect 16212 7308 16548 7364
rect 24098 7308 24108 7364
rect 24164 7308 28028 7364
rect 28084 7308 28094 7364
rect 3490 7196 3500 7252
rect 3556 7196 8876 7252
rect 8932 7196 9212 7252
rect 9268 7196 9278 7252
rect 10210 7196 10220 7252
rect 10276 7196 10892 7252
rect 10948 7196 12796 7252
rect 12852 7196 12862 7252
rect 25666 7196 25676 7252
rect 25732 7196 27132 7252
rect 27188 7196 27198 7252
rect 30706 7196 30716 7252
rect 30772 7196 31500 7252
rect 31556 7196 32172 7252
rect 32228 7196 32238 7252
rect 15250 7084 15260 7140
rect 15316 7084 16268 7140
rect 16324 7084 17388 7140
rect 17444 7084 17454 7140
rect 26674 7084 26684 7140
rect 26740 7084 27020 7140
rect 27076 7084 28700 7140
rect 28756 7084 29372 7140
rect 29428 7084 29820 7140
rect 29876 7084 29886 7140
rect 5360 7028 5370 7084
rect 5426 7028 5474 7084
rect 5530 7028 5578 7084
rect 5634 7028 5644 7084
rect 13676 7028 13686 7084
rect 13742 7028 13790 7084
rect 13846 7028 13894 7084
rect 13950 7028 13960 7084
rect 3938 6972 3948 7028
rect 4004 6972 5124 7028
rect 6178 6972 6188 7028
rect 6244 6972 9884 7028
rect 9940 6972 9950 7028
rect 5068 6916 5124 6972
rect 15260 6916 15316 7084
rect 21992 7028 22002 7084
rect 22058 7028 22106 7084
rect 22162 7028 22210 7084
rect 22266 7028 22276 7084
rect 30308 7028 30318 7084
rect 30374 7028 30422 7084
rect 30478 7028 30526 7084
rect 30582 7028 30592 7084
rect 26786 6972 26796 7028
rect 26852 6972 28140 7028
rect 28196 6972 28206 7028
rect 3154 6860 3164 6916
rect 3220 6860 4844 6916
rect 4900 6860 4910 6916
rect 5068 6860 12012 6916
rect 12068 6860 12078 6916
rect 12236 6860 12572 6916
rect 12628 6860 12638 6916
rect 12898 6860 12908 6916
rect 12964 6860 15316 6916
rect 22082 6860 22092 6916
rect 22148 6860 23324 6916
rect 23380 6860 23548 6916
rect 23604 6860 23614 6916
rect 28578 6860 28588 6916
rect 28644 6860 29260 6916
rect 29316 6860 31388 6916
rect 31444 6860 31948 6916
rect 32004 6860 33180 6916
rect 33236 6860 33246 6916
rect 12236 6804 12292 6860
rect 4722 6748 4732 6804
rect 4788 6748 7756 6804
rect 7812 6748 7822 6804
rect 8764 6748 9660 6804
rect 9716 6748 12292 6804
rect 12450 6748 12460 6804
rect 12516 6748 14364 6804
rect 14420 6748 14430 6804
rect 21858 6748 21868 6804
rect 21924 6748 23436 6804
rect 23492 6748 23502 6804
rect 26674 6748 26684 6804
rect 26740 6748 27356 6804
rect 27412 6748 27422 6804
rect 29698 6748 29708 6804
rect 29764 6748 30044 6804
rect 30100 6748 30380 6804
rect 30436 6748 30446 6804
rect 8764 6692 8820 6748
rect 3826 6636 3836 6692
rect 3892 6636 3902 6692
rect 4050 6636 4060 6692
rect 4116 6636 4956 6692
rect 5012 6636 5628 6692
rect 5684 6636 5694 6692
rect 5842 6636 5852 6692
rect 5908 6636 6076 6692
rect 6132 6636 6412 6692
rect 6468 6636 6478 6692
rect 6626 6636 6636 6692
rect 6692 6636 7420 6692
rect 7476 6636 7644 6692
rect 7700 6636 7710 6692
rect 7970 6636 7980 6692
rect 8036 6636 8820 6692
rect 9212 6636 13356 6692
rect 13412 6636 13422 6692
rect 14578 6636 14588 6692
rect 14644 6636 17276 6692
rect 17332 6636 17342 6692
rect 21410 6636 21420 6692
rect 21476 6636 21756 6692
rect 21812 6636 21822 6692
rect 26450 6636 26460 6692
rect 26516 6636 29596 6692
rect 29652 6636 30156 6692
rect 30212 6636 30222 6692
rect 3836 6468 3892 6636
rect 9212 6580 9268 6636
rect 5058 6524 5068 6580
rect 5124 6524 9268 6580
rect 12674 6524 12684 6580
rect 12740 6524 13132 6580
rect 13188 6524 13804 6580
rect 13860 6524 13870 6580
rect 22978 6524 22988 6580
rect 23044 6524 24780 6580
rect 24836 6524 24846 6580
rect 3836 6412 6188 6468
rect 6244 6412 7084 6468
rect 7140 6412 8092 6468
rect 8148 6412 8158 6468
rect 8316 6356 8372 6524
rect 8978 6412 8988 6468
rect 9044 6412 11564 6468
rect 11620 6412 11630 6468
rect 13234 6412 13244 6468
rect 13300 6412 17164 6468
rect 17220 6412 17230 6468
rect 17714 6412 17724 6468
rect 17780 6412 18732 6468
rect 18788 6412 18798 6468
rect 5842 6300 5852 6356
rect 5908 6300 6524 6356
rect 6580 6300 6590 6356
rect 6850 6300 6860 6356
rect 6916 6300 7308 6356
rect 7364 6300 7374 6356
rect 7522 6300 7532 6356
rect 7588 6300 7980 6356
rect 8036 6300 8046 6356
rect 8316 6300 8652 6356
rect 8708 6300 8718 6356
rect 9518 6244 9528 6300
rect 9584 6244 9632 6300
rect 9688 6244 9736 6300
rect 9792 6244 9802 6300
rect 17834 6244 17844 6300
rect 17900 6244 17948 6300
rect 18004 6244 18052 6300
rect 18108 6244 18118 6300
rect 26150 6244 26160 6300
rect 26216 6244 26264 6300
rect 26320 6244 26368 6300
rect 26424 6244 26434 6300
rect 34466 6244 34476 6300
rect 34532 6244 34580 6300
rect 34636 6244 34684 6300
rect 34740 6244 34750 6300
rect 3042 6188 3052 6244
rect 3108 6188 3388 6244
rect 4610 6188 4620 6244
rect 4676 6188 8204 6244
rect 8260 6188 8270 6244
rect 8530 6188 8540 6244
rect 8596 6188 8876 6244
rect 8932 6188 9380 6244
rect 13010 6188 13020 6244
rect 13076 6188 14252 6244
rect 14308 6188 14318 6244
rect 3332 5908 3388 6188
rect 9324 6132 9380 6188
rect 5506 6076 5516 6132
rect 5572 6076 7644 6132
rect 7700 6076 7710 6132
rect 7970 6076 7980 6132
rect 8036 6076 8764 6132
rect 8820 6076 8830 6132
rect 9324 6076 10220 6132
rect 10276 6076 13692 6132
rect 13748 6076 13758 6132
rect 19506 6076 19516 6132
rect 19572 6076 21308 6132
rect 21364 6076 21374 6132
rect 24434 6076 24444 6132
rect 24500 6076 25676 6132
rect 25732 6076 26964 6132
rect 30930 6076 30940 6132
rect 30996 6076 33292 6132
rect 33348 6076 33964 6132
rect 34020 6076 34030 6132
rect 7644 6020 7700 6076
rect 26908 6020 26964 6076
rect 4498 5964 4508 6020
rect 4564 5964 5852 6020
rect 5908 5964 6972 6020
rect 7028 5964 7038 6020
rect 7644 5964 8876 6020
rect 8932 5964 9212 6020
rect 9268 5964 9278 6020
rect 21634 5964 21644 6020
rect 21700 5964 22988 6020
rect 23044 5964 23054 6020
rect 25564 5964 26684 6020
rect 26740 5964 26750 6020
rect 26898 5964 26908 6020
rect 26964 5964 27916 6020
rect 27972 5964 27982 6020
rect 25564 5908 25620 5964
rect 3332 5852 7868 5908
rect 7924 5852 8428 5908
rect 8484 5852 8494 5908
rect 9314 5852 9324 5908
rect 9380 5852 9436 5908
rect 9492 5852 9502 5908
rect 14466 5852 14476 5908
rect 14532 5852 15596 5908
rect 15652 5852 15662 5908
rect 19282 5852 19292 5908
rect 19348 5852 23772 5908
rect 23828 5852 23838 5908
rect 24434 5852 24444 5908
rect 24500 5852 25564 5908
rect 25620 5852 25630 5908
rect 26114 5852 26124 5908
rect 26180 5852 27692 5908
rect 27748 5852 27758 5908
rect 29810 5852 29820 5908
rect 29876 5852 30604 5908
rect 30660 5852 33068 5908
rect 33124 5852 33134 5908
rect 6262 5740 6300 5796
rect 6356 5740 6366 5796
rect 6850 5740 6860 5796
rect 6916 5740 6972 5796
rect 7028 5740 11900 5796
rect 11956 5740 11966 5796
rect 14578 5740 14588 5796
rect 14644 5740 17724 5796
rect 17780 5740 17790 5796
rect 26898 5740 26908 5796
rect 26964 5740 27804 5796
rect 27860 5740 27870 5796
rect 30706 5740 30716 5796
rect 30772 5740 31724 5796
rect 31780 5740 31790 5796
rect 3042 5628 3052 5684
rect 3108 5628 9324 5684
rect 9380 5628 9390 5684
rect 16594 5628 16604 5684
rect 16660 5628 17276 5684
rect 17332 5628 17342 5684
rect 26226 5628 26236 5684
rect 26292 5628 27356 5684
rect 27412 5628 27422 5684
rect 30146 5628 30156 5684
rect 30212 5628 33068 5684
rect 33124 5628 33134 5684
rect 7298 5516 7308 5572
rect 7364 5516 7420 5572
rect 7476 5516 7486 5572
rect 15474 5516 15484 5572
rect 15540 5516 17836 5572
rect 17892 5516 18956 5572
rect 19012 5516 19022 5572
rect 30706 5516 30716 5572
rect 30772 5516 31836 5572
rect 31892 5516 31902 5572
rect 5360 5460 5370 5516
rect 5426 5460 5474 5516
rect 5530 5460 5578 5516
rect 5634 5460 5644 5516
rect 13676 5460 13686 5516
rect 13742 5460 13790 5516
rect 13846 5460 13894 5516
rect 13950 5460 13960 5516
rect 21992 5460 22002 5516
rect 22058 5460 22106 5516
rect 22162 5460 22210 5516
rect 22266 5460 22276 5516
rect 30308 5460 30318 5516
rect 30374 5460 30422 5516
rect 30478 5460 30526 5516
rect 30582 5460 30592 5516
rect 24098 5404 24108 5460
rect 24164 5404 25340 5460
rect 25396 5404 26460 5460
rect 26516 5404 26526 5460
rect 31154 5404 31164 5460
rect 31220 5404 33404 5460
rect 33460 5404 34188 5460
rect 34244 5404 34254 5460
rect 8642 5292 8652 5348
rect 8708 5292 10780 5348
rect 10836 5292 12124 5348
rect 12180 5292 12190 5348
rect 13570 5292 13580 5348
rect 13636 5292 14588 5348
rect 14644 5292 14654 5348
rect 15092 5292 16044 5348
rect 16100 5292 16110 5348
rect 30930 5292 30940 5348
rect 30996 5292 33180 5348
rect 33236 5292 33246 5348
rect 15092 5236 15148 5292
rect 2706 5180 2716 5236
rect 2772 5180 4284 5236
rect 4340 5180 4956 5236
rect 5012 5180 5022 5236
rect 8866 5180 8876 5236
rect 8932 5180 10892 5236
rect 10948 5180 15148 5236
rect 18274 5180 18284 5236
rect 18340 5180 19180 5236
rect 19236 5180 19246 5236
rect 21634 5180 21644 5236
rect 21700 5180 23772 5236
rect 23828 5180 27468 5236
rect 27524 5180 27534 5236
rect 2146 5068 2156 5124
rect 2212 5068 2828 5124
rect 2884 5068 3388 5124
rect 3444 5068 3454 5124
rect 4834 5068 4844 5124
rect 4900 5068 5516 5124
rect 5572 5068 5964 5124
rect 6020 5068 6030 5124
rect 11778 5068 11788 5124
rect 11844 5068 12684 5124
rect 12740 5068 12750 5124
rect 13234 5068 13244 5124
rect 13300 5068 13916 5124
rect 13972 5068 13982 5124
rect 16930 5068 16940 5124
rect 16996 5068 18172 5124
rect 18228 5068 18844 5124
rect 18900 5068 18910 5124
rect 27122 5068 27132 5124
rect 27188 5068 28588 5124
rect 28644 5068 31052 5124
rect 31108 5068 31836 5124
rect 31892 5068 31902 5124
rect 6626 4956 6636 5012
rect 6692 4956 8204 5012
rect 8260 4956 8270 5012
rect 8418 4956 8428 5012
rect 8484 4956 9436 5012
rect 9492 4956 9502 5012
rect 14018 4956 14028 5012
rect 14084 4956 15260 5012
rect 15316 4956 15326 5012
rect 22754 4956 22764 5012
rect 22820 4956 23436 5012
rect 23492 4956 23502 5012
rect 5058 4844 5068 4900
rect 5124 4844 6188 4900
rect 6244 4844 8652 4900
rect 8708 4844 8718 4900
rect 11554 4844 11564 4900
rect 11620 4844 16044 4900
rect 16100 4844 16110 4900
rect 29586 4844 29596 4900
rect 29652 4844 31164 4900
rect 31220 4844 31230 4900
rect 3602 4732 3612 4788
rect 3668 4732 4396 4788
rect 4452 4732 6748 4788
rect 6804 4732 6814 4788
rect 7494 4732 7532 4788
rect 7588 4732 7598 4788
rect 7858 4732 7868 4788
rect 7924 4732 8988 4788
rect 9044 4732 9054 4788
rect 9518 4676 9528 4732
rect 9584 4676 9632 4732
rect 9688 4676 9736 4732
rect 9792 4676 9802 4732
rect 17834 4676 17844 4732
rect 17900 4676 17948 4732
rect 18004 4676 18052 4732
rect 18108 4676 18118 4732
rect 26150 4676 26160 4732
rect 26216 4676 26264 4732
rect 26320 4676 26368 4732
rect 26424 4676 26434 4732
rect 34466 4676 34476 4732
rect 34532 4676 34580 4732
rect 34636 4676 34684 4732
rect 34740 4676 34750 4732
rect 7186 4620 7196 4676
rect 7252 4620 9380 4676
rect 9324 4564 9380 4620
rect 4694 4508 4732 4564
rect 4788 4508 4798 4564
rect 5702 4508 5740 4564
rect 5796 4508 5806 4564
rect 7046 4508 7084 4564
rect 7140 4508 7150 4564
rect 7746 4508 7756 4564
rect 7812 4508 9100 4564
rect 9156 4508 9166 4564
rect 9324 4508 9772 4564
rect 9828 4508 9838 4564
rect 11330 4508 11340 4564
rect 11396 4508 12124 4564
rect 12180 4508 13468 4564
rect 13524 4508 13534 4564
rect 16146 4508 16156 4564
rect 16212 4508 17500 4564
rect 17556 4508 17566 4564
rect 18610 4508 18620 4564
rect 18676 4508 19180 4564
rect 19236 4508 20860 4564
rect 20916 4508 20926 4564
rect 21858 4508 21868 4564
rect 21924 4508 22764 4564
rect 22820 4508 22830 4564
rect 5170 4396 5180 4452
rect 5236 4396 6860 4452
rect 6916 4396 6926 4452
rect 7410 4396 7420 4452
rect 7476 4396 8652 4452
rect 8708 4396 8718 4452
rect 11442 4396 11452 4452
rect 11508 4396 13356 4452
rect 13412 4396 13422 4452
rect 7420 4340 7476 4396
rect 11452 4340 11508 4396
rect 1810 4284 1820 4340
rect 1876 4284 5852 4340
rect 5908 4284 5918 4340
rect 6626 4284 6636 4340
rect 6692 4284 7476 4340
rect 8306 4284 8316 4340
rect 8372 4284 11508 4340
rect 12562 4284 12572 4340
rect 12628 4284 15036 4340
rect 15092 4284 15102 4340
rect 21746 4284 21756 4340
rect 21812 4284 23100 4340
rect 23156 4284 23166 4340
rect 1586 4172 1596 4228
rect 1652 4172 3612 4228
rect 3668 4172 3678 4228
rect 5730 4172 5740 4228
rect 5796 4172 6860 4228
rect 6916 4172 14140 4228
rect 14196 4172 14206 4228
rect 20290 4172 20300 4228
rect 20356 4172 23660 4228
rect 23716 4172 23726 4228
rect 23314 4060 23324 4116
rect 23380 4060 25228 4116
rect 25284 4060 25294 4116
rect 5360 3892 5370 3948
rect 5426 3892 5474 3948
rect 5530 3892 5578 3948
rect 5634 3892 5644 3948
rect 13676 3892 13686 3948
rect 13742 3892 13790 3948
rect 13846 3892 13894 3948
rect 13950 3892 13960 3948
rect 21992 3892 22002 3948
rect 22058 3892 22106 3948
rect 22162 3892 22210 3948
rect 22266 3892 22276 3948
rect 30308 3892 30318 3948
rect 30374 3892 30422 3948
rect 30478 3892 30526 3948
rect 30582 3892 30592 3948
rect 6738 3724 6748 3780
rect 6804 3724 14924 3780
rect 14980 3724 14990 3780
rect 8978 3612 8988 3668
rect 9044 3612 10220 3668
rect 10276 3612 10286 3668
rect 22754 3612 22764 3668
rect 22820 3612 24556 3668
rect 24612 3612 24622 3668
rect 9538 3500 9548 3556
rect 9604 3500 12572 3556
rect 12628 3500 12638 3556
rect 19730 3500 19740 3556
rect 19796 3500 20748 3556
rect 20804 3500 20814 3556
rect 22418 3500 22428 3556
rect 22484 3500 24892 3556
rect 24948 3500 24958 3556
rect 25106 3388 25116 3444
rect 25172 3388 26908 3444
rect 26964 3388 26974 3444
rect 30034 3388 30044 3444
rect 30100 3388 32284 3444
rect 32340 3388 32350 3444
rect 9518 3108 9528 3164
rect 9584 3108 9632 3164
rect 9688 3108 9736 3164
rect 9792 3108 9802 3164
rect 17834 3108 17844 3164
rect 17900 3108 17948 3164
rect 18004 3108 18052 3164
rect 18108 3108 18118 3164
rect 26150 3108 26160 3164
rect 26216 3108 26264 3164
rect 26320 3108 26368 3164
rect 26424 3108 26434 3164
rect 34466 3108 34476 3164
rect 34532 3108 34580 3164
rect 34636 3108 34684 3164
rect 34740 3108 34750 3164
<< via3 >>
rect 5370 32116 5426 32172
rect 5474 32116 5530 32172
rect 5578 32116 5634 32172
rect 13686 32116 13742 32172
rect 13790 32116 13846 32172
rect 13894 32116 13950 32172
rect 22002 32116 22058 32172
rect 22106 32116 22162 32172
rect 22210 32116 22266 32172
rect 30318 32116 30374 32172
rect 30422 32116 30478 32172
rect 30526 32116 30582 32172
rect 9528 31332 9584 31388
rect 9632 31332 9688 31388
rect 9736 31332 9792 31388
rect 17844 31332 17900 31388
rect 17948 31332 18004 31388
rect 18052 31332 18108 31388
rect 26160 31332 26216 31388
rect 26264 31332 26320 31388
rect 26368 31332 26424 31388
rect 34476 31332 34532 31388
rect 34580 31332 34636 31388
rect 34684 31332 34740 31388
rect 5370 30548 5426 30604
rect 5474 30548 5530 30604
rect 5578 30548 5634 30604
rect 13686 30548 13742 30604
rect 13790 30548 13846 30604
rect 13894 30548 13950 30604
rect 22002 30548 22058 30604
rect 22106 30548 22162 30604
rect 22210 30548 22266 30604
rect 30318 30548 30374 30604
rect 30422 30548 30478 30604
rect 30526 30548 30582 30604
rect 9528 29764 9584 29820
rect 9632 29764 9688 29820
rect 9736 29764 9792 29820
rect 17844 29764 17900 29820
rect 17948 29764 18004 29820
rect 18052 29764 18108 29820
rect 26160 29764 26216 29820
rect 26264 29764 26320 29820
rect 26368 29764 26424 29820
rect 34476 29764 34532 29820
rect 34580 29764 34636 29820
rect 34684 29764 34740 29820
rect 5370 28980 5426 29036
rect 5474 28980 5530 29036
rect 5578 28980 5634 29036
rect 13686 28980 13742 29036
rect 13790 28980 13846 29036
rect 13894 28980 13950 29036
rect 22002 28980 22058 29036
rect 22106 28980 22162 29036
rect 22210 28980 22266 29036
rect 30318 28980 30374 29036
rect 30422 28980 30478 29036
rect 30526 28980 30582 29036
rect 9528 28196 9584 28252
rect 9632 28196 9688 28252
rect 9736 28196 9792 28252
rect 17844 28196 17900 28252
rect 17948 28196 18004 28252
rect 18052 28196 18108 28252
rect 26160 28196 26216 28252
rect 26264 28196 26320 28252
rect 26368 28196 26424 28252
rect 34476 28196 34532 28252
rect 34580 28196 34636 28252
rect 34684 28196 34740 28252
rect 5370 27412 5426 27468
rect 5474 27412 5530 27468
rect 5578 27412 5634 27468
rect 13686 27412 13742 27468
rect 13790 27412 13846 27468
rect 13894 27412 13950 27468
rect 22002 27412 22058 27468
rect 22106 27412 22162 27468
rect 22210 27412 22266 27468
rect 30318 27412 30374 27468
rect 30422 27412 30478 27468
rect 30526 27412 30582 27468
rect 9528 26628 9584 26684
rect 9632 26628 9688 26684
rect 9736 26628 9792 26684
rect 17844 26628 17900 26684
rect 17948 26628 18004 26684
rect 18052 26628 18108 26684
rect 26160 26628 26216 26684
rect 26264 26628 26320 26684
rect 26368 26628 26424 26684
rect 34476 26628 34532 26684
rect 34580 26628 34636 26684
rect 34684 26628 34740 26684
rect 5370 25844 5426 25900
rect 5474 25844 5530 25900
rect 5578 25844 5634 25900
rect 13686 25844 13742 25900
rect 13790 25844 13846 25900
rect 13894 25844 13950 25900
rect 22002 25844 22058 25900
rect 22106 25844 22162 25900
rect 22210 25844 22266 25900
rect 30318 25844 30374 25900
rect 30422 25844 30478 25900
rect 30526 25844 30582 25900
rect 26796 25228 26852 25284
rect 9528 25060 9584 25116
rect 9632 25060 9688 25116
rect 9736 25060 9792 25116
rect 17844 25060 17900 25116
rect 17948 25060 18004 25116
rect 18052 25060 18108 25116
rect 26160 25060 26216 25116
rect 26264 25060 26320 25116
rect 26368 25060 26424 25116
rect 34476 25060 34532 25116
rect 34580 25060 34636 25116
rect 34684 25060 34740 25116
rect 12796 24780 12852 24836
rect 12236 24668 12292 24724
rect 13468 24668 13524 24724
rect 12348 24444 12404 24500
rect 5370 24276 5426 24332
rect 5474 24276 5530 24332
rect 5578 24276 5634 24332
rect 13686 24276 13742 24332
rect 13790 24276 13846 24332
rect 13894 24276 13950 24332
rect 22002 24276 22058 24332
rect 22106 24276 22162 24332
rect 22210 24276 22266 24332
rect 30318 24276 30374 24332
rect 30422 24276 30478 24332
rect 30526 24276 30582 24332
rect 12236 23884 12292 23940
rect 12796 23884 12852 23940
rect 12348 23772 12404 23828
rect 9528 23492 9584 23548
rect 9632 23492 9688 23548
rect 9736 23492 9792 23548
rect 17844 23492 17900 23548
rect 17948 23492 18004 23548
rect 18052 23492 18108 23548
rect 26160 23492 26216 23548
rect 26264 23492 26320 23548
rect 26368 23492 26424 23548
rect 34476 23492 34532 23548
rect 34580 23492 34636 23548
rect 34684 23492 34740 23548
rect 14588 23324 14644 23380
rect 14588 23100 14644 23156
rect 26796 22764 26852 22820
rect 5370 22708 5426 22764
rect 5474 22708 5530 22764
rect 5578 22708 5634 22764
rect 13686 22708 13742 22764
rect 13790 22708 13846 22764
rect 13894 22708 13950 22764
rect 22002 22708 22058 22764
rect 22106 22708 22162 22764
rect 22210 22708 22266 22764
rect 30318 22708 30374 22764
rect 30422 22708 30478 22764
rect 30526 22708 30582 22764
rect 9528 21924 9584 21980
rect 9632 21924 9688 21980
rect 9736 21924 9792 21980
rect 17844 21924 17900 21980
rect 17948 21924 18004 21980
rect 18052 21924 18108 21980
rect 26160 21924 26216 21980
rect 26264 21924 26320 21980
rect 26368 21924 26424 21980
rect 34476 21924 34532 21980
rect 34580 21924 34636 21980
rect 34684 21924 34740 21980
rect 15932 21868 15988 21924
rect 5370 21140 5426 21196
rect 5474 21140 5530 21196
rect 5578 21140 5634 21196
rect 13686 21140 13742 21196
rect 13790 21140 13846 21196
rect 13894 21140 13950 21196
rect 22002 21140 22058 21196
rect 22106 21140 22162 21196
rect 22210 21140 22266 21196
rect 30318 21140 30374 21196
rect 30422 21140 30478 21196
rect 30526 21140 30582 21196
rect 9528 20356 9584 20412
rect 9632 20356 9688 20412
rect 9736 20356 9792 20412
rect 17844 20356 17900 20412
rect 17948 20356 18004 20412
rect 18052 20356 18108 20412
rect 26160 20356 26216 20412
rect 26264 20356 26320 20412
rect 26368 20356 26424 20412
rect 34476 20356 34532 20412
rect 34580 20356 34636 20412
rect 34684 20356 34740 20412
rect 13468 19628 13524 19684
rect 5370 19572 5426 19628
rect 5474 19572 5530 19628
rect 5578 19572 5634 19628
rect 13686 19572 13742 19628
rect 13790 19572 13846 19628
rect 13894 19572 13950 19628
rect 22002 19572 22058 19628
rect 22106 19572 22162 19628
rect 22210 19572 22266 19628
rect 30318 19572 30374 19628
rect 30422 19572 30478 19628
rect 30526 19572 30582 19628
rect 9528 18788 9584 18844
rect 9632 18788 9688 18844
rect 9736 18788 9792 18844
rect 17844 18788 17900 18844
rect 17948 18788 18004 18844
rect 18052 18788 18108 18844
rect 26160 18788 26216 18844
rect 26264 18788 26320 18844
rect 26368 18788 26424 18844
rect 34476 18788 34532 18844
rect 34580 18788 34636 18844
rect 34684 18788 34740 18844
rect 5370 18004 5426 18060
rect 5474 18004 5530 18060
rect 5578 18004 5634 18060
rect 13686 18004 13742 18060
rect 13790 18004 13846 18060
rect 13894 18004 13950 18060
rect 22002 18004 22058 18060
rect 22106 18004 22162 18060
rect 22210 18004 22266 18060
rect 30318 18004 30374 18060
rect 30422 18004 30478 18060
rect 30526 18004 30582 18060
rect 9528 17220 9584 17276
rect 9632 17220 9688 17276
rect 9736 17220 9792 17276
rect 17844 17220 17900 17276
rect 17948 17220 18004 17276
rect 18052 17220 18108 17276
rect 26160 17220 26216 17276
rect 26264 17220 26320 17276
rect 26368 17220 26424 17276
rect 34476 17220 34532 17276
rect 34580 17220 34636 17276
rect 34684 17220 34740 17276
rect 5370 16436 5426 16492
rect 5474 16436 5530 16492
rect 5578 16436 5634 16492
rect 13686 16436 13742 16492
rect 13790 16436 13846 16492
rect 13894 16436 13950 16492
rect 22002 16436 22058 16492
rect 22106 16436 22162 16492
rect 22210 16436 22266 16492
rect 30318 16436 30374 16492
rect 30422 16436 30478 16492
rect 30526 16436 30582 16492
rect 15932 16380 15988 16436
rect 9528 15652 9584 15708
rect 9632 15652 9688 15708
rect 9736 15652 9792 15708
rect 17844 15652 17900 15708
rect 17948 15652 18004 15708
rect 18052 15652 18108 15708
rect 26160 15652 26216 15708
rect 26264 15652 26320 15708
rect 26368 15652 26424 15708
rect 34476 15652 34532 15708
rect 34580 15652 34636 15708
rect 34684 15652 34740 15708
rect 5370 14868 5426 14924
rect 5474 14868 5530 14924
rect 5578 14868 5634 14924
rect 13686 14868 13742 14924
rect 13790 14868 13846 14924
rect 13894 14868 13950 14924
rect 22002 14868 22058 14924
rect 22106 14868 22162 14924
rect 22210 14868 22266 14924
rect 30318 14868 30374 14924
rect 30422 14868 30478 14924
rect 30526 14868 30582 14924
rect 9528 14084 9584 14140
rect 9632 14084 9688 14140
rect 9736 14084 9792 14140
rect 17844 14084 17900 14140
rect 17948 14084 18004 14140
rect 18052 14084 18108 14140
rect 26160 14084 26216 14140
rect 26264 14084 26320 14140
rect 26368 14084 26424 14140
rect 34476 14084 34532 14140
rect 34580 14084 34636 14140
rect 34684 14084 34740 14140
rect 5370 13300 5426 13356
rect 5474 13300 5530 13356
rect 5578 13300 5634 13356
rect 13686 13300 13742 13356
rect 13790 13300 13846 13356
rect 13894 13300 13950 13356
rect 22002 13300 22058 13356
rect 22106 13300 22162 13356
rect 22210 13300 22266 13356
rect 30318 13300 30374 13356
rect 30422 13300 30478 13356
rect 30526 13300 30582 13356
rect 9528 12516 9584 12572
rect 9632 12516 9688 12572
rect 9736 12516 9792 12572
rect 17844 12516 17900 12572
rect 17948 12516 18004 12572
rect 18052 12516 18108 12572
rect 26160 12516 26216 12572
rect 26264 12516 26320 12572
rect 26368 12516 26424 12572
rect 34476 12516 34532 12572
rect 34580 12516 34636 12572
rect 34684 12516 34740 12572
rect 4620 11788 4676 11844
rect 5370 11732 5426 11788
rect 5474 11732 5530 11788
rect 5578 11732 5634 11788
rect 13686 11732 13742 11788
rect 13790 11732 13846 11788
rect 13894 11732 13950 11788
rect 22002 11732 22058 11788
rect 22106 11732 22162 11788
rect 22210 11732 22266 11788
rect 30318 11732 30374 11788
rect 30422 11732 30478 11788
rect 30526 11732 30582 11788
rect 4732 11564 4788 11620
rect 9528 10948 9584 11004
rect 9632 10948 9688 11004
rect 9736 10948 9792 11004
rect 17844 10948 17900 11004
rect 17948 10948 18004 11004
rect 18052 10948 18108 11004
rect 26160 10948 26216 11004
rect 26264 10948 26320 11004
rect 26368 10948 26424 11004
rect 34476 10948 34532 11004
rect 34580 10948 34636 11004
rect 34684 10948 34740 11004
rect 9324 10332 9380 10388
rect 5370 10164 5426 10220
rect 5474 10164 5530 10220
rect 5578 10164 5634 10220
rect 13686 10164 13742 10220
rect 13790 10164 13846 10220
rect 13894 10164 13950 10220
rect 22002 10164 22058 10220
rect 22106 10164 22162 10220
rect 22210 10164 22266 10220
rect 30318 10164 30374 10220
rect 30422 10164 30478 10220
rect 30526 10164 30582 10220
rect 9884 10108 9940 10164
rect 4620 9996 4676 10052
rect 6300 9884 6356 9940
rect 4732 9548 4788 9604
rect 9528 9380 9584 9436
rect 9632 9380 9688 9436
rect 9736 9380 9792 9436
rect 17844 9380 17900 9436
rect 17948 9380 18004 9436
rect 18052 9380 18108 9436
rect 26160 9380 26216 9436
rect 26264 9380 26320 9436
rect 26368 9380 26424 9436
rect 8428 8988 8484 9044
rect 34476 9380 34532 9436
rect 34580 9380 34636 9436
rect 34684 9380 34740 9436
rect 7084 8764 7140 8820
rect 5370 8596 5426 8652
rect 5474 8596 5530 8652
rect 5578 8596 5634 8652
rect 13686 8596 13742 8652
rect 13790 8596 13846 8652
rect 13894 8596 13950 8652
rect 22002 8596 22058 8652
rect 22106 8596 22162 8652
rect 22210 8596 22266 8652
rect 30318 8596 30374 8652
rect 30422 8596 30478 8652
rect 30526 8596 30582 8652
rect 7308 8428 7364 8484
rect 6972 8204 7028 8260
rect 9996 8092 10052 8148
rect 5740 7980 5796 8036
rect 9324 7868 9380 7924
rect 9528 7812 9584 7868
rect 9632 7812 9688 7868
rect 9736 7812 9792 7868
rect 17844 7812 17900 7868
rect 17948 7812 18004 7868
rect 18052 7812 18108 7868
rect 26160 7812 26216 7868
rect 26264 7812 26320 7868
rect 26368 7812 26424 7868
rect 34476 7812 34532 7868
rect 34580 7812 34636 7868
rect 34684 7812 34740 7868
rect 9996 7308 10052 7364
rect 5370 7028 5426 7084
rect 5474 7028 5530 7084
rect 5578 7028 5634 7084
rect 13686 7028 13742 7084
rect 13790 7028 13846 7084
rect 13894 7028 13950 7084
rect 9884 6972 9940 7028
rect 22002 7028 22058 7084
rect 22106 7028 22162 7084
rect 22210 7028 22266 7084
rect 30318 7028 30374 7084
rect 30422 7028 30478 7084
rect 30526 7028 30582 7084
rect 7420 6636 7476 6692
rect 7308 6300 7364 6356
rect 7532 6300 7588 6356
rect 9528 6244 9584 6300
rect 9632 6244 9688 6300
rect 9736 6244 9792 6300
rect 17844 6244 17900 6300
rect 17948 6244 18004 6300
rect 18052 6244 18108 6300
rect 26160 6244 26216 6300
rect 26264 6244 26320 6300
rect 26368 6244 26424 6300
rect 34476 6244 34532 6300
rect 34580 6244 34636 6300
rect 34684 6244 34740 6300
rect 9324 5852 9380 5908
rect 6300 5740 6356 5796
rect 6972 5740 7028 5796
rect 7420 5516 7476 5572
rect 5370 5460 5426 5516
rect 5474 5460 5530 5516
rect 5578 5460 5634 5516
rect 13686 5460 13742 5516
rect 13790 5460 13846 5516
rect 13894 5460 13950 5516
rect 22002 5460 22058 5516
rect 22106 5460 22162 5516
rect 22210 5460 22266 5516
rect 30318 5460 30374 5516
rect 30422 5460 30478 5516
rect 30526 5460 30582 5516
rect 8428 4956 8484 5012
rect 7532 4732 7588 4788
rect 9528 4676 9584 4732
rect 9632 4676 9688 4732
rect 9736 4676 9792 4732
rect 17844 4676 17900 4732
rect 17948 4676 18004 4732
rect 18052 4676 18108 4732
rect 26160 4676 26216 4732
rect 26264 4676 26320 4732
rect 26368 4676 26424 4732
rect 34476 4676 34532 4732
rect 34580 4676 34636 4732
rect 34684 4676 34740 4732
rect 4732 4508 4788 4564
rect 5740 4508 5796 4564
rect 7084 4508 7140 4564
rect 5370 3892 5426 3948
rect 5474 3892 5530 3948
rect 5578 3892 5634 3948
rect 13686 3892 13742 3948
rect 13790 3892 13846 3948
rect 13894 3892 13950 3948
rect 22002 3892 22058 3948
rect 22106 3892 22162 3948
rect 22210 3892 22266 3948
rect 30318 3892 30374 3948
rect 30422 3892 30478 3948
rect 30526 3892 30582 3948
rect 9528 3108 9584 3164
rect 9632 3108 9688 3164
rect 9736 3108 9792 3164
rect 17844 3108 17900 3164
rect 17948 3108 18004 3164
rect 18052 3108 18108 3164
rect 26160 3108 26216 3164
rect 26264 3108 26320 3164
rect 26368 3108 26424 3164
rect 34476 3108 34532 3164
rect 34580 3108 34636 3164
rect 34684 3108 34740 3164
<< metal4 >>
rect 5342 32172 5662 32204
rect 5342 32116 5370 32172
rect 5426 32116 5474 32172
rect 5530 32116 5578 32172
rect 5634 32116 5662 32172
rect 5342 30604 5662 32116
rect 5342 30548 5370 30604
rect 5426 30548 5474 30604
rect 5530 30548 5578 30604
rect 5634 30548 5662 30604
rect 5342 29036 5662 30548
rect 5342 28980 5370 29036
rect 5426 28980 5474 29036
rect 5530 28980 5578 29036
rect 5634 28980 5662 29036
rect 5342 27468 5662 28980
rect 5342 27412 5370 27468
rect 5426 27412 5474 27468
rect 5530 27412 5578 27468
rect 5634 27412 5662 27468
rect 5342 25900 5662 27412
rect 5342 25844 5370 25900
rect 5426 25844 5474 25900
rect 5530 25844 5578 25900
rect 5634 25844 5662 25900
rect 5342 24332 5662 25844
rect 5342 24276 5370 24332
rect 5426 24276 5474 24332
rect 5530 24276 5578 24332
rect 5634 24276 5662 24332
rect 5342 22764 5662 24276
rect 5342 22708 5370 22764
rect 5426 22708 5474 22764
rect 5530 22708 5578 22764
rect 5634 22708 5662 22764
rect 5342 21196 5662 22708
rect 5342 21140 5370 21196
rect 5426 21140 5474 21196
rect 5530 21140 5578 21196
rect 5634 21140 5662 21196
rect 5342 19628 5662 21140
rect 5342 19572 5370 19628
rect 5426 19572 5474 19628
rect 5530 19572 5578 19628
rect 5634 19572 5662 19628
rect 5342 18060 5662 19572
rect 5342 18004 5370 18060
rect 5426 18004 5474 18060
rect 5530 18004 5578 18060
rect 5634 18004 5662 18060
rect 5342 16492 5662 18004
rect 5342 16436 5370 16492
rect 5426 16436 5474 16492
rect 5530 16436 5578 16492
rect 5634 16436 5662 16492
rect 5342 14924 5662 16436
rect 5342 14868 5370 14924
rect 5426 14868 5474 14924
rect 5530 14868 5578 14924
rect 5634 14868 5662 14924
rect 5342 13356 5662 14868
rect 5342 13300 5370 13356
rect 5426 13300 5474 13356
rect 5530 13300 5578 13356
rect 5634 13300 5662 13356
rect 4620 11844 4676 11854
rect 4620 10052 4676 11788
rect 5342 11788 5662 13300
rect 5342 11732 5370 11788
rect 5426 11732 5474 11788
rect 5530 11732 5578 11788
rect 5634 11732 5662 11788
rect 4620 9986 4676 9996
rect 4732 11620 4788 11630
rect 4732 9604 4788 11564
rect 4732 4564 4788 9548
rect 4732 4498 4788 4508
rect 5342 10220 5662 11732
rect 9500 31388 9820 32204
rect 9500 31332 9528 31388
rect 9584 31332 9632 31388
rect 9688 31332 9736 31388
rect 9792 31332 9820 31388
rect 9500 29820 9820 31332
rect 9500 29764 9528 29820
rect 9584 29764 9632 29820
rect 9688 29764 9736 29820
rect 9792 29764 9820 29820
rect 9500 28252 9820 29764
rect 9500 28196 9528 28252
rect 9584 28196 9632 28252
rect 9688 28196 9736 28252
rect 9792 28196 9820 28252
rect 9500 26684 9820 28196
rect 9500 26628 9528 26684
rect 9584 26628 9632 26684
rect 9688 26628 9736 26684
rect 9792 26628 9820 26684
rect 9500 25116 9820 26628
rect 9500 25060 9528 25116
rect 9584 25060 9632 25116
rect 9688 25060 9736 25116
rect 9792 25060 9820 25116
rect 9500 23548 9820 25060
rect 13658 32172 13978 32204
rect 13658 32116 13686 32172
rect 13742 32116 13790 32172
rect 13846 32116 13894 32172
rect 13950 32116 13978 32172
rect 13658 30604 13978 32116
rect 13658 30548 13686 30604
rect 13742 30548 13790 30604
rect 13846 30548 13894 30604
rect 13950 30548 13978 30604
rect 13658 29036 13978 30548
rect 13658 28980 13686 29036
rect 13742 28980 13790 29036
rect 13846 28980 13894 29036
rect 13950 28980 13978 29036
rect 13658 27468 13978 28980
rect 13658 27412 13686 27468
rect 13742 27412 13790 27468
rect 13846 27412 13894 27468
rect 13950 27412 13978 27468
rect 13658 25900 13978 27412
rect 13658 25844 13686 25900
rect 13742 25844 13790 25900
rect 13846 25844 13894 25900
rect 13950 25844 13978 25900
rect 12796 24836 12852 24846
rect 12236 24724 12292 24734
rect 12236 23940 12292 24668
rect 12236 23874 12292 23884
rect 12348 24500 12404 24510
rect 12348 23828 12404 24444
rect 12796 23940 12852 24780
rect 12796 23874 12852 23884
rect 13468 24724 13524 24734
rect 12348 23762 12404 23772
rect 9500 23492 9528 23548
rect 9584 23492 9632 23548
rect 9688 23492 9736 23548
rect 9792 23492 9820 23548
rect 9500 21980 9820 23492
rect 9500 21924 9528 21980
rect 9584 21924 9632 21980
rect 9688 21924 9736 21980
rect 9792 21924 9820 21980
rect 9500 20412 9820 21924
rect 9500 20356 9528 20412
rect 9584 20356 9632 20412
rect 9688 20356 9736 20412
rect 9792 20356 9820 20412
rect 9500 18844 9820 20356
rect 13468 19684 13524 24668
rect 13468 19618 13524 19628
rect 13658 24332 13978 25844
rect 13658 24276 13686 24332
rect 13742 24276 13790 24332
rect 13846 24276 13894 24332
rect 13950 24276 13978 24332
rect 13658 22764 13978 24276
rect 17816 31388 18136 32204
rect 17816 31332 17844 31388
rect 17900 31332 17948 31388
rect 18004 31332 18052 31388
rect 18108 31332 18136 31388
rect 17816 29820 18136 31332
rect 17816 29764 17844 29820
rect 17900 29764 17948 29820
rect 18004 29764 18052 29820
rect 18108 29764 18136 29820
rect 17816 28252 18136 29764
rect 17816 28196 17844 28252
rect 17900 28196 17948 28252
rect 18004 28196 18052 28252
rect 18108 28196 18136 28252
rect 17816 26684 18136 28196
rect 17816 26628 17844 26684
rect 17900 26628 17948 26684
rect 18004 26628 18052 26684
rect 18108 26628 18136 26684
rect 17816 25116 18136 26628
rect 17816 25060 17844 25116
rect 17900 25060 17948 25116
rect 18004 25060 18052 25116
rect 18108 25060 18136 25116
rect 17816 23548 18136 25060
rect 17816 23492 17844 23548
rect 17900 23492 17948 23548
rect 18004 23492 18052 23548
rect 18108 23492 18136 23548
rect 14588 23380 14644 23390
rect 14588 23156 14644 23324
rect 14588 23090 14644 23100
rect 13658 22708 13686 22764
rect 13742 22708 13790 22764
rect 13846 22708 13894 22764
rect 13950 22708 13978 22764
rect 13658 21196 13978 22708
rect 17816 21980 18136 23492
rect 13658 21140 13686 21196
rect 13742 21140 13790 21196
rect 13846 21140 13894 21196
rect 13950 21140 13978 21196
rect 13658 19628 13978 21140
rect 9500 18788 9528 18844
rect 9584 18788 9632 18844
rect 9688 18788 9736 18844
rect 9792 18788 9820 18844
rect 9500 17276 9820 18788
rect 9500 17220 9528 17276
rect 9584 17220 9632 17276
rect 9688 17220 9736 17276
rect 9792 17220 9820 17276
rect 9500 15708 9820 17220
rect 9500 15652 9528 15708
rect 9584 15652 9632 15708
rect 9688 15652 9736 15708
rect 9792 15652 9820 15708
rect 9500 14140 9820 15652
rect 9500 14084 9528 14140
rect 9584 14084 9632 14140
rect 9688 14084 9736 14140
rect 9792 14084 9820 14140
rect 9500 12572 9820 14084
rect 9500 12516 9528 12572
rect 9584 12516 9632 12572
rect 9688 12516 9736 12572
rect 9792 12516 9820 12572
rect 9500 11004 9820 12516
rect 9500 10948 9528 11004
rect 9584 10948 9632 11004
rect 9688 10948 9736 11004
rect 9792 10948 9820 11004
rect 5342 10164 5370 10220
rect 5426 10164 5474 10220
rect 5530 10164 5578 10220
rect 5634 10164 5662 10220
rect 5342 8652 5662 10164
rect 9324 10388 9380 10398
rect 5342 8596 5370 8652
rect 5426 8596 5474 8652
rect 5530 8596 5578 8652
rect 5634 8596 5662 8652
rect 5342 7084 5662 8596
rect 6300 9940 6356 9950
rect 5342 7028 5370 7084
rect 5426 7028 5474 7084
rect 5530 7028 5578 7084
rect 5634 7028 5662 7084
rect 5342 5516 5662 7028
rect 5342 5460 5370 5516
rect 5426 5460 5474 5516
rect 5530 5460 5578 5516
rect 5634 5460 5662 5516
rect 5342 3948 5662 5460
rect 5740 8036 5796 8046
rect 5740 4564 5796 7980
rect 6300 5796 6356 9884
rect 8428 9044 8484 9054
rect 7084 8820 7140 8830
rect 6300 5730 6356 5740
rect 6972 8260 7028 8270
rect 6972 5796 7028 8204
rect 6972 5730 7028 5740
rect 5740 4498 5796 4508
rect 7084 4564 7140 8764
rect 7308 8484 7364 8494
rect 7308 6356 7364 8428
rect 7308 6290 7364 6300
rect 7420 6692 7476 6702
rect 7420 5572 7476 6636
rect 7420 5506 7476 5516
rect 7532 6356 7588 6366
rect 7532 4788 7588 6300
rect 8428 5012 8484 8988
rect 9324 7924 9380 10332
rect 9324 5908 9380 7868
rect 9324 5842 9380 5852
rect 9500 9436 9820 10948
rect 13658 19572 13686 19628
rect 13742 19572 13790 19628
rect 13846 19572 13894 19628
rect 13950 19572 13978 19628
rect 13658 18060 13978 19572
rect 13658 18004 13686 18060
rect 13742 18004 13790 18060
rect 13846 18004 13894 18060
rect 13950 18004 13978 18060
rect 13658 16492 13978 18004
rect 13658 16436 13686 16492
rect 13742 16436 13790 16492
rect 13846 16436 13894 16492
rect 13950 16436 13978 16492
rect 13658 14924 13978 16436
rect 15932 21924 15988 21934
rect 15932 16436 15988 21868
rect 15932 16370 15988 16380
rect 17816 21924 17844 21980
rect 17900 21924 17948 21980
rect 18004 21924 18052 21980
rect 18108 21924 18136 21980
rect 17816 20412 18136 21924
rect 17816 20356 17844 20412
rect 17900 20356 17948 20412
rect 18004 20356 18052 20412
rect 18108 20356 18136 20412
rect 17816 18844 18136 20356
rect 17816 18788 17844 18844
rect 17900 18788 17948 18844
rect 18004 18788 18052 18844
rect 18108 18788 18136 18844
rect 17816 17276 18136 18788
rect 17816 17220 17844 17276
rect 17900 17220 17948 17276
rect 18004 17220 18052 17276
rect 18108 17220 18136 17276
rect 13658 14868 13686 14924
rect 13742 14868 13790 14924
rect 13846 14868 13894 14924
rect 13950 14868 13978 14924
rect 13658 13356 13978 14868
rect 13658 13300 13686 13356
rect 13742 13300 13790 13356
rect 13846 13300 13894 13356
rect 13950 13300 13978 13356
rect 13658 11788 13978 13300
rect 13658 11732 13686 11788
rect 13742 11732 13790 11788
rect 13846 11732 13894 11788
rect 13950 11732 13978 11788
rect 13658 10220 13978 11732
rect 9500 9380 9528 9436
rect 9584 9380 9632 9436
rect 9688 9380 9736 9436
rect 9792 9380 9820 9436
rect 9500 7868 9820 9380
rect 9500 7812 9528 7868
rect 9584 7812 9632 7868
rect 9688 7812 9736 7868
rect 9792 7812 9820 7868
rect 9500 6300 9820 7812
rect 9884 10164 9940 10174
rect 9884 7028 9940 10108
rect 13658 10164 13686 10220
rect 13742 10164 13790 10220
rect 13846 10164 13894 10220
rect 13950 10164 13978 10220
rect 13658 8652 13978 10164
rect 13658 8596 13686 8652
rect 13742 8596 13790 8652
rect 13846 8596 13894 8652
rect 13950 8596 13978 8652
rect 9996 8148 10052 8158
rect 9996 7364 10052 8092
rect 9996 7298 10052 7308
rect 9884 6962 9940 6972
rect 13658 7084 13978 8596
rect 13658 7028 13686 7084
rect 13742 7028 13790 7084
rect 13846 7028 13894 7084
rect 13950 7028 13978 7084
rect 9500 6244 9528 6300
rect 9584 6244 9632 6300
rect 9688 6244 9736 6300
rect 9792 6244 9820 6300
rect 8428 4946 8484 4956
rect 7532 4722 7588 4732
rect 9500 4732 9820 6244
rect 7084 4498 7140 4508
rect 9500 4676 9528 4732
rect 9584 4676 9632 4732
rect 9688 4676 9736 4732
rect 9792 4676 9820 4732
rect 5342 3892 5370 3948
rect 5426 3892 5474 3948
rect 5530 3892 5578 3948
rect 5634 3892 5662 3948
rect 5342 3076 5662 3892
rect 9500 3164 9820 4676
rect 9500 3108 9528 3164
rect 9584 3108 9632 3164
rect 9688 3108 9736 3164
rect 9792 3108 9820 3164
rect 9500 3076 9820 3108
rect 13658 5516 13978 7028
rect 13658 5460 13686 5516
rect 13742 5460 13790 5516
rect 13846 5460 13894 5516
rect 13950 5460 13978 5516
rect 13658 3948 13978 5460
rect 13658 3892 13686 3948
rect 13742 3892 13790 3948
rect 13846 3892 13894 3948
rect 13950 3892 13978 3948
rect 13658 3076 13978 3892
rect 17816 15708 18136 17220
rect 17816 15652 17844 15708
rect 17900 15652 17948 15708
rect 18004 15652 18052 15708
rect 18108 15652 18136 15708
rect 17816 14140 18136 15652
rect 17816 14084 17844 14140
rect 17900 14084 17948 14140
rect 18004 14084 18052 14140
rect 18108 14084 18136 14140
rect 17816 12572 18136 14084
rect 17816 12516 17844 12572
rect 17900 12516 17948 12572
rect 18004 12516 18052 12572
rect 18108 12516 18136 12572
rect 17816 11004 18136 12516
rect 17816 10948 17844 11004
rect 17900 10948 17948 11004
rect 18004 10948 18052 11004
rect 18108 10948 18136 11004
rect 17816 9436 18136 10948
rect 17816 9380 17844 9436
rect 17900 9380 17948 9436
rect 18004 9380 18052 9436
rect 18108 9380 18136 9436
rect 17816 7868 18136 9380
rect 17816 7812 17844 7868
rect 17900 7812 17948 7868
rect 18004 7812 18052 7868
rect 18108 7812 18136 7868
rect 17816 6300 18136 7812
rect 17816 6244 17844 6300
rect 17900 6244 17948 6300
rect 18004 6244 18052 6300
rect 18108 6244 18136 6300
rect 17816 4732 18136 6244
rect 17816 4676 17844 4732
rect 17900 4676 17948 4732
rect 18004 4676 18052 4732
rect 18108 4676 18136 4732
rect 17816 3164 18136 4676
rect 17816 3108 17844 3164
rect 17900 3108 17948 3164
rect 18004 3108 18052 3164
rect 18108 3108 18136 3164
rect 17816 3076 18136 3108
rect 21974 32172 22294 32204
rect 21974 32116 22002 32172
rect 22058 32116 22106 32172
rect 22162 32116 22210 32172
rect 22266 32116 22294 32172
rect 21974 30604 22294 32116
rect 21974 30548 22002 30604
rect 22058 30548 22106 30604
rect 22162 30548 22210 30604
rect 22266 30548 22294 30604
rect 21974 29036 22294 30548
rect 21974 28980 22002 29036
rect 22058 28980 22106 29036
rect 22162 28980 22210 29036
rect 22266 28980 22294 29036
rect 21974 27468 22294 28980
rect 21974 27412 22002 27468
rect 22058 27412 22106 27468
rect 22162 27412 22210 27468
rect 22266 27412 22294 27468
rect 21974 25900 22294 27412
rect 21974 25844 22002 25900
rect 22058 25844 22106 25900
rect 22162 25844 22210 25900
rect 22266 25844 22294 25900
rect 21974 24332 22294 25844
rect 21974 24276 22002 24332
rect 22058 24276 22106 24332
rect 22162 24276 22210 24332
rect 22266 24276 22294 24332
rect 21974 22764 22294 24276
rect 21974 22708 22002 22764
rect 22058 22708 22106 22764
rect 22162 22708 22210 22764
rect 22266 22708 22294 22764
rect 21974 21196 22294 22708
rect 21974 21140 22002 21196
rect 22058 21140 22106 21196
rect 22162 21140 22210 21196
rect 22266 21140 22294 21196
rect 21974 19628 22294 21140
rect 21974 19572 22002 19628
rect 22058 19572 22106 19628
rect 22162 19572 22210 19628
rect 22266 19572 22294 19628
rect 21974 18060 22294 19572
rect 21974 18004 22002 18060
rect 22058 18004 22106 18060
rect 22162 18004 22210 18060
rect 22266 18004 22294 18060
rect 21974 16492 22294 18004
rect 21974 16436 22002 16492
rect 22058 16436 22106 16492
rect 22162 16436 22210 16492
rect 22266 16436 22294 16492
rect 21974 14924 22294 16436
rect 21974 14868 22002 14924
rect 22058 14868 22106 14924
rect 22162 14868 22210 14924
rect 22266 14868 22294 14924
rect 21974 13356 22294 14868
rect 21974 13300 22002 13356
rect 22058 13300 22106 13356
rect 22162 13300 22210 13356
rect 22266 13300 22294 13356
rect 21974 11788 22294 13300
rect 21974 11732 22002 11788
rect 22058 11732 22106 11788
rect 22162 11732 22210 11788
rect 22266 11732 22294 11788
rect 21974 10220 22294 11732
rect 21974 10164 22002 10220
rect 22058 10164 22106 10220
rect 22162 10164 22210 10220
rect 22266 10164 22294 10220
rect 21974 8652 22294 10164
rect 21974 8596 22002 8652
rect 22058 8596 22106 8652
rect 22162 8596 22210 8652
rect 22266 8596 22294 8652
rect 21974 7084 22294 8596
rect 21974 7028 22002 7084
rect 22058 7028 22106 7084
rect 22162 7028 22210 7084
rect 22266 7028 22294 7084
rect 21974 5516 22294 7028
rect 21974 5460 22002 5516
rect 22058 5460 22106 5516
rect 22162 5460 22210 5516
rect 22266 5460 22294 5516
rect 21974 3948 22294 5460
rect 21974 3892 22002 3948
rect 22058 3892 22106 3948
rect 22162 3892 22210 3948
rect 22266 3892 22294 3948
rect 21974 3076 22294 3892
rect 26132 31388 26452 32204
rect 26132 31332 26160 31388
rect 26216 31332 26264 31388
rect 26320 31332 26368 31388
rect 26424 31332 26452 31388
rect 26132 29820 26452 31332
rect 26132 29764 26160 29820
rect 26216 29764 26264 29820
rect 26320 29764 26368 29820
rect 26424 29764 26452 29820
rect 26132 28252 26452 29764
rect 26132 28196 26160 28252
rect 26216 28196 26264 28252
rect 26320 28196 26368 28252
rect 26424 28196 26452 28252
rect 26132 26684 26452 28196
rect 26132 26628 26160 26684
rect 26216 26628 26264 26684
rect 26320 26628 26368 26684
rect 26424 26628 26452 26684
rect 26132 25116 26452 26628
rect 30290 32172 30610 32204
rect 30290 32116 30318 32172
rect 30374 32116 30422 32172
rect 30478 32116 30526 32172
rect 30582 32116 30610 32172
rect 30290 30604 30610 32116
rect 30290 30548 30318 30604
rect 30374 30548 30422 30604
rect 30478 30548 30526 30604
rect 30582 30548 30610 30604
rect 30290 29036 30610 30548
rect 30290 28980 30318 29036
rect 30374 28980 30422 29036
rect 30478 28980 30526 29036
rect 30582 28980 30610 29036
rect 30290 27468 30610 28980
rect 30290 27412 30318 27468
rect 30374 27412 30422 27468
rect 30478 27412 30526 27468
rect 30582 27412 30610 27468
rect 30290 25900 30610 27412
rect 30290 25844 30318 25900
rect 30374 25844 30422 25900
rect 30478 25844 30526 25900
rect 30582 25844 30610 25900
rect 26132 25060 26160 25116
rect 26216 25060 26264 25116
rect 26320 25060 26368 25116
rect 26424 25060 26452 25116
rect 26132 23548 26452 25060
rect 26132 23492 26160 23548
rect 26216 23492 26264 23548
rect 26320 23492 26368 23548
rect 26424 23492 26452 23548
rect 26132 21980 26452 23492
rect 26796 25284 26852 25294
rect 26796 22820 26852 25228
rect 26796 22754 26852 22764
rect 30290 24332 30610 25844
rect 30290 24276 30318 24332
rect 30374 24276 30422 24332
rect 30478 24276 30526 24332
rect 30582 24276 30610 24332
rect 30290 22764 30610 24276
rect 26132 21924 26160 21980
rect 26216 21924 26264 21980
rect 26320 21924 26368 21980
rect 26424 21924 26452 21980
rect 26132 20412 26452 21924
rect 26132 20356 26160 20412
rect 26216 20356 26264 20412
rect 26320 20356 26368 20412
rect 26424 20356 26452 20412
rect 26132 18844 26452 20356
rect 26132 18788 26160 18844
rect 26216 18788 26264 18844
rect 26320 18788 26368 18844
rect 26424 18788 26452 18844
rect 26132 17276 26452 18788
rect 26132 17220 26160 17276
rect 26216 17220 26264 17276
rect 26320 17220 26368 17276
rect 26424 17220 26452 17276
rect 26132 15708 26452 17220
rect 26132 15652 26160 15708
rect 26216 15652 26264 15708
rect 26320 15652 26368 15708
rect 26424 15652 26452 15708
rect 26132 14140 26452 15652
rect 26132 14084 26160 14140
rect 26216 14084 26264 14140
rect 26320 14084 26368 14140
rect 26424 14084 26452 14140
rect 26132 12572 26452 14084
rect 26132 12516 26160 12572
rect 26216 12516 26264 12572
rect 26320 12516 26368 12572
rect 26424 12516 26452 12572
rect 26132 11004 26452 12516
rect 26132 10948 26160 11004
rect 26216 10948 26264 11004
rect 26320 10948 26368 11004
rect 26424 10948 26452 11004
rect 26132 9436 26452 10948
rect 26132 9380 26160 9436
rect 26216 9380 26264 9436
rect 26320 9380 26368 9436
rect 26424 9380 26452 9436
rect 26132 7868 26452 9380
rect 26132 7812 26160 7868
rect 26216 7812 26264 7868
rect 26320 7812 26368 7868
rect 26424 7812 26452 7868
rect 26132 6300 26452 7812
rect 26132 6244 26160 6300
rect 26216 6244 26264 6300
rect 26320 6244 26368 6300
rect 26424 6244 26452 6300
rect 26132 4732 26452 6244
rect 26132 4676 26160 4732
rect 26216 4676 26264 4732
rect 26320 4676 26368 4732
rect 26424 4676 26452 4732
rect 26132 3164 26452 4676
rect 26132 3108 26160 3164
rect 26216 3108 26264 3164
rect 26320 3108 26368 3164
rect 26424 3108 26452 3164
rect 26132 3076 26452 3108
rect 30290 22708 30318 22764
rect 30374 22708 30422 22764
rect 30478 22708 30526 22764
rect 30582 22708 30610 22764
rect 30290 21196 30610 22708
rect 30290 21140 30318 21196
rect 30374 21140 30422 21196
rect 30478 21140 30526 21196
rect 30582 21140 30610 21196
rect 30290 19628 30610 21140
rect 30290 19572 30318 19628
rect 30374 19572 30422 19628
rect 30478 19572 30526 19628
rect 30582 19572 30610 19628
rect 30290 18060 30610 19572
rect 30290 18004 30318 18060
rect 30374 18004 30422 18060
rect 30478 18004 30526 18060
rect 30582 18004 30610 18060
rect 30290 16492 30610 18004
rect 30290 16436 30318 16492
rect 30374 16436 30422 16492
rect 30478 16436 30526 16492
rect 30582 16436 30610 16492
rect 30290 14924 30610 16436
rect 30290 14868 30318 14924
rect 30374 14868 30422 14924
rect 30478 14868 30526 14924
rect 30582 14868 30610 14924
rect 30290 13356 30610 14868
rect 30290 13300 30318 13356
rect 30374 13300 30422 13356
rect 30478 13300 30526 13356
rect 30582 13300 30610 13356
rect 30290 11788 30610 13300
rect 30290 11732 30318 11788
rect 30374 11732 30422 11788
rect 30478 11732 30526 11788
rect 30582 11732 30610 11788
rect 30290 10220 30610 11732
rect 30290 10164 30318 10220
rect 30374 10164 30422 10220
rect 30478 10164 30526 10220
rect 30582 10164 30610 10220
rect 30290 8652 30610 10164
rect 30290 8596 30318 8652
rect 30374 8596 30422 8652
rect 30478 8596 30526 8652
rect 30582 8596 30610 8652
rect 30290 7084 30610 8596
rect 30290 7028 30318 7084
rect 30374 7028 30422 7084
rect 30478 7028 30526 7084
rect 30582 7028 30610 7084
rect 30290 5516 30610 7028
rect 30290 5460 30318 5516
rect 30374 5460 30422 5516
rect 30478 5460 30526 5516
rect 30582 5460 30610 5516
rect 30290 3948 30610 5460
rect 30290 3892 30318 3948
rect 30374 3892 30422 3948
rect 30478 3892 30526 3948
rect 30582 3892 30610 3948
rect 30290 3076 30610 3892
rect 34448 31388 34768 32204
rect 34448 31332 34476 31388
rect 34532 31332 34580 31388
rect 34636 31332 34684 31388
rect 34740 31332 34768 31388
rect 34448 29820 34768 31332
rect 34448 29764 34476 29820
rect 34532 29764 34580 29820
rect 34636 29764 34684 29820
rect 34740 29764 34768 29820
rect 34448 28252 34768 29764
rect 34448 28196 34476 28252
rect 34532 28196 34580 28252
rect 34636 28196 34684 28252
rect 34740 28196 34768 28252
rect 34448 26684 34768 28196
rect 34448 26628 34476 26684
rect 34532 26628 34580 26684
rect 34636 26628 34684 26684
rect 34740 26628 34768 26684
rect 34448 25116 34768 26628
rect 34448 25060 34476 25116
rect 34532 25060 34580 25116
rect 34636 25060 34684 25116
rect 34740 25060 34768 25116
rect 34448 23548 34768 25060
rect 34448 23492 34476 23548
rect 34532 23492 34580 23548
rect 34636 23492 34684 23548
rect 34740 23492 34768 23548
rect 34448 21980 34768 23492
rect 34448 21924 34476 21980
rect 34532 21924 34580 21980
rect 34636 21924 34684 21980
rect 34740 21924 34768 21980
rect 34448 20412 34768 21924
rect 34448 20356 34476 20412
rect 34532 20356 34580 20412
rect 34636 20356 34684 20412
rect 34740 20356 34768 20412
rect 34448 18844 34768 20356
rect 34448 18788 34476 18844
rect 34532 18788 34580 18844
rect 34636 18788 34684 18844
rect 34740 18788 34768 18844
rect 34448 17276 34768 18788
rect 34448 17220 34476 17276
rect 34532 17220 34580 17276
rect 34636 17220 34684 17276
rect 34740 17220 34768 17276
rect 34448 15708 34768 17220
rect 34448 15652 34476 15708
rect 34532 15652 34580 15708
rect 34636 15652 34684 15708
rect 34740 15652 34768 15708
rect 34448 14140 34768 15652
rect 34448 14084 34476 14140
rect 34532 14084 34580 14140
rect 34636 14084 34684 14140
rect 34740 14084 34768 14140
rect 34448 12572 34768 14084
rect 34448 12516 34476 12572
rect 34532 12516 34580 12572
rect 34636 12516 34684 12572
rect 34740 12516 34768 12572
rect 34448 11004 34768 12516
rect 34448 10948 34476 11004
rect 34532 10948 34580 11004
rect 34636 10948 34684 11004
rect 34740 10948 34768 11004
rect 34448 9436 34768 10948
rect 34448 9380 34476 9436
rect 34532 9380 34580 9436
rect 34636 9380 34684 9436
rect 34740 9380 34768 9436
rect 34448 7868 34768 9380
rect 34448 7812 34476 7868
rect 34532 7812 34580 7868
rect 34636 7812 34684 7868
rect 34740 7812 34768 7868
rect 34448 6300 34768 7812
rect 34448 6244 34476 6300
rect 34532 6244 34580 6300
rect 34636 6244 34684 6300
rect 34740 6244 34768 6300
rect 34448 4732 34768 6244
rect 34448 4676 34476 4732
rect 34532 4676 34580 4732
rect 34636 4676 34684 4732
rect 34740 4676 34768 4732
rect 34448 3164 34768 4676
rect 34448 3108 34476 3164
rect 34532 3108 34580 3164
rect 34636 3108 34684 3164
rect 34740 3108 34768 3164
rect 34448 3076 34768 3108
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _428_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12432 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _429_
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _430_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13888 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _431_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18816 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _432_
timestamp 1698175906
transform 1 0 16576 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _433_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 24864 0 -1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _434_
timestamp 1698175906
transform -1 0 24864 0 -1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _435_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21504 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _436_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22848 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _437_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _438_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17248 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _439_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 23632 0 -1 25088
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _440_
timestamp 1698175906
transform 1 0 4816 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _441_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 6944 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _442_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5264 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _443_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _444_
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _445_
timestamp 1698175906
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _446_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17584 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _447_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _448_
timestamp 1698175906
transform -1 0 20720 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _449_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22400 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _450_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19712 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _451_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18032 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _452_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20832 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _453_
timestamp 1698175906
transform -1 0 18032 0 1 9408
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _454_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9968 0 -1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _455_
timestamp 1698175906
transform -1 0 12320 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _456_
timestamp 1698175906
transform -1 0 18144 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _457_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17024 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _458_
timestamp 1698175906
transform -1 0 16912 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _459_
timestamp 1698175906
transform -1 0 11984 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _460_
timestamp 1698175906
transform 1 0 10976 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _461_
timestamp 1698175906
transform -1 0 11536 0 -1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _462_
timestamp 1698175906
transform -1 0 7728 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _463_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _464_
timestamp 1698175906
transform -1 0 13104 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _465_
timestamp 1698175906
transform 1 0 11872 0 1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _466_
timestamp 1698175906
transform 1 0 10416 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _467_
timestamp 1698175906
transform -1 0 11088 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _468_
timestamp 1698175906
transform 1 0 11088 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _469_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14112 0 -1 9408
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _470_
timestamp 1698175906
transform 1 0 18032 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _471_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18816 0 1 7840
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _472_
timestamp 1698175906
transform 1 0 11984 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _473_
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _474_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17024 0 -1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _475_
timestamp 1698175906
transform -1 0 15456 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _476_
timestamp 1698175906
transform -1 0 14784 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _477_
timestamp 1698175906
transform -1 0 8512 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _478_
timestamp 1698175906
transform 1 0 7840 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _479_
timestamp 1698175906
transform 1 0 18592 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _480_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15456 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _481_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15456 0 -1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _482_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11312 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _483_
timestamp 1698175906
transform -1 0 13552 0 -1 7840
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _484_
timestamp 1698175906
transform -1 0 11088 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _485_
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _486_
timestamp 1698175906
transform 1 0 6608 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _487_
timestamp 1698175906
transform 1 0 7616 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _488_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11760 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _489_
timestamp 1698175906
transform -1 0 18592 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _490_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16800 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _491_
timestamp 1698175906
transform -1 0 11760 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _492_
timestamp 1698175906
transform -1 0 3696 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _493_
timestamp 1698175906
transform 1 0 1904 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _494_
timestamp 1698175906
transform -1 0 15680 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _495_
timestamp 1698175906
transform 1 0 6608 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _496_
timestamp 1698175906
transform -1 0 13104 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _497_
timestamp 1698175906
transform -1 0 7056 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _498_
timestamp 1698175906
transform -1 0 6608 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _499_
timestamp 1698175906
transform 1 0 5040 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _500_
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _501_
timestamp 1698175906
transform 1 0 6272 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _502_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _503_
timestamp 1698175906
transform 1 0 9856 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _504_
timestamp 1698175906
transform -1 0 8512 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _505_
timestamp 1698175906
transform 1 0 2576 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _506_
timestamp 1698175906
transform 1 0 4144 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _507_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12992 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _508_
timestamp 1698175906
transform 1 0 8064 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _509_
timestamp 1698175906
transform -1 0 8400 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _510_
timestamp 1698175906
transform 1 0 13776 0 1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _511_
timestamp 1698175906
transform 1 0 5712 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _512_
timestamp 1698175906
transform 1 0 6384 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _513_
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _514_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7616 0 -1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _515_
timestamp 1698175906
transform 1 0 7280 0 -1 6272
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _516_
timestamp 1698175906
transform 1 0 8288 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _517_
timestamp 1698175906
transform 1 0 2688 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _518_
timestamp 1698175906
transform -1 0 10192 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _519_
timestamp 1698175906
transform -1 0 11088 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _520_
timestamp 1698175906
transform -1 0 10080 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _521_
timestamp 1698175906
transform 1 0 3248 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _522_
timestamp 1698175906
transform 1 0 10640 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _523_
timestamp 1698175906
transform 1 0 7728 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _524_
timestamp 1698175906
transform -1 0 12096 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _525_
timestamp 1698175906
transform -1 0 9184 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _526_
timestamp 1698175906
transform -1 0 5936 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _527_
timestamp 1698175906
transform 1 0 9408 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _528_
timestamp 1698175906
transform -1 0 10080 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _529_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _530_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _531_
timestamp 1698175906
transform -1 0 9296 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _532_
timestamp 1698175906
transform 1 0 8288 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _533_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10304 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _534_
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _535_
timestamp 1698175906
transform -1 0 5264 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _536_
timestamp 1698175906
transform -1 0 6944 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _537_
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _538_
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _539_
timestamp 1698175906
transform 1 0 2352 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _540_
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _541_
timestamp 1698175906
transform 1 0 7280 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _542_
timestamp 1698175906
transform 1 0 10640 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _543_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7616 0 1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _544_
timestamp 1698175906
transform 1 0 7504 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _545_
timestamp 1698175906
transform -1 0 7616 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _546_
timestamp 1698175906
transform 1 0 6272 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _547_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9296 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _548_
timestamp 1698175906
transform 1 0 4480 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _549_
timestamp 1698175906
transform 1 0 6496 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _550_
timestamp 1698175906
transform -1 0 2688 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _551_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 3584 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _552_
timestamp 1698175906
transform -1 0 6720 0 1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _553_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _554_
timestamp 1698175906
transform -1 0 10416 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _555_
timestamp 1698175906
transform 1 0 3360 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _556_
timestamp 1698175906
transform -1 0 3360 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _557_
timestamp 1698175906
transform 1 0 2688 0 -1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _558_
timestamp 1698175906
transform -1 0 5824 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _559_
timestamp 1698175906
transform -1 0 3024 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _560_
timestamp 1698175906
transform -1 0 5264 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _561_
timestamp 1698175906
transform 1 0 3024 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _562_
timestamp 1698175906
transform 1 0 3472 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _563_
timestamp 1698175906
transform 1 0 2688 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _564_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 3024 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _565_
timestamp 1698175906
transform 1 0 1904 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _566_
timestamp 1698175906
transform -1 0 6384 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _567_
timestamp 1698175906
transform 1 0 3360 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _568_
timestamp 1698175906
transform -1 0 5152 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _569_
timestamp 1698175906
transform -1 0 7728 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _570_
timestamp 1698175906
transform 1 0 4368 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _571_
timestamp 1698175906
transform 1 0 5824 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _572_
timestamp 1698175906
transform 1 0 2912 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _573_
timestamp 1698175906
transform -1 0 5264 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _574_
timestamp 1698175906
transform 1 0 4032 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _575_
timestamp 1698175906
transform 1 0 3472 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _576_
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _577_
timestamp 1698175906
transform 1 0 6720 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _578_
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _579_
timestamp 1698175906
transform -1 0 6944 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _580_
timestamp 1698175906
transform 1 0 23296 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _581_
timestamp 1698175906
transform -1 0 32704 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _582_
timestamp 1698175906
transform 1 0 13664 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _583_
timestamp 1698175906
transform -1 0 27664 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _584_
timestamp 1698175906
transform -1 0 23072 0 1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _585_
timestamp 1698175906
transform -1 0 33824 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _586_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22064 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _587_
timestamp 1698175906
transform 1 0 29792 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _588_
timestamp 1698175906
transform -1 0 30576 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _589_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 32144 0 -1 9408
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _590_
timestamp 1698175906
transform 1 0 26096 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _591_
timestamp 1698175906
transform -1 0 27776 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _592_
timestamp 1698175906
transform 1 0 27664 0 1 7840
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _593_
timestamp 1698175906
transform 1 0 30576 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _594_
timestamp 1698175906
transform -1 0 31920 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _595_
timestamp 1698175906
transform -1 0 26432 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _596_
timestamp 1698175906
transform 1 0 26992 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _597_
timestamp 1698175906
transform 1 0 27776 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _598_
timestamp 1698175906
transform 1 0 23072 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _599_
timestamp 1698175906
transform 1 0 23408 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _600_
timestamp 1698175906
transform 1 0 25200 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _601_
timestamp 1698175906
transform -1 0 26768 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _602_
timestamp 1698175906
transform -1 0 22288 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _603_
timestamp 1698175906
transform 1 0 17920 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _604_
timestamp 1698175906
transform -1 0 19936 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _605_
timestamp 1698175906
transform -1 0 22512 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _606_
timestamp 1698175906
transform -1 0 22064 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _607_
timestamp 1698175906
transform -1 0 27440 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _608_
timestamp 1698175906
transform -1 0 23520 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _609_
timestamp 1698175906
transform 1 0 23184 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _610_
timestamp 1698175906
transform -1 0 22288 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _611_
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _612_
timestamp 1698175906
transform 1 0 21840 0 -1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _613_
timestamp 1698175906
transform -1 0 28448 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _614_
timestamp 1698175906
transform -1 0 24416 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _615_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 24864 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _616_
timestamp 1698175906
transform 1 0 24080 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _617_
timestamp 1698175906
transform 1 0 25200 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _618_
timestamp 1698175906
transform -1 0 27216 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _619_
timestamp 1698175906
transform -1 0 28112 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _620_
timestamp 1698175906
transform -1 0 27888 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _621_
timestamp 1698175906
transform 1 0 25536 0 -1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _622_
timestamp 1698175906
transform 1 0 26880 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _623_
timestamp 1698175906
transform 1 0 28112 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _624_
timestamp 1698175906
transform 1 0 28560 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _625_
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _626_
timestamp 1698175906
transform -1 0 30352 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _627_
timestamp 1698175906
transform -1 0 29904 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _628_
timestamp 1698175906
transform 1 0 29680 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _629_
timestamp 1698175906
transform 1 0 29904 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _630_
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _631_
timestamp 1698175906
transform 1 0 30240 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _632_
timestamp 1698175906
transform 1 0 30464 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _633_
timestamp 1698175906
transform 1 0 30016 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _634_
timestamp 1698175906
transform 1 0 31360 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _635_
timestamp 1698175906
transform 1 0 29120 0 -1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _636_
timestamp 1698175906
transform 1 0 32032 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _637_
timestamp 1698175906
transform -1 0 32032 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _638_
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _639_
timestamp 1698175906
transform 1 0 30240 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _640_
timestamp 1698175906
transform -1 0 33824 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _641_
timestamp 1698175906
transform -1 0 29904 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _642_
timestamp 1698175906
transform -1 0 29904 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _643_
timestamp 1698175906
transform 1 0 28336 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _644_
timestamp 1698175906
transform 1 0 29904 0 1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _645_
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _646_
timestamp 1698175906
transform -1 0 32144 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _647_
timestamp 1698175906
transform 1 0 30912 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _648_
timestamp 1698175906
transform 1 0 31584 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _649_
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _650_
timestamp 1698175906
transform -1 0 33824 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _651_
timestamp 1698175906
transform -1 0 30800 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _652_
timestamp 1698175906
transform 1 0 32256 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _653_
timestamp 1698175906
transform 1 0 31024 0 1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _654_
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _655_
timestamp 1698175906
transform -1 0 32592 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _656_
timestamp 1698175906
transform -1 0 29904 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _657_
timestamp 1698175906
transform -1 0 29680 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _658_
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _659_
timestamp 1698175906
transform -1 0 27328 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _660_
timestamp 1698175906
transform -1 0 26208 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _661_
timestamp 1698175906
transform -1 0 26768 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _662_
timestamp 1698175906
transform 1 0 27104 0 1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _663_
timestamp 1698175906
transform -1 0 27664 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _664_
timestamp 1698175906
transform 1 0 27776 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _665_
timestamp 1698175906
transform 1 0 27776 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _666_
timestamp 1698175906
transform -1 0 27104 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _667_
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _668_
timestamp 1698175906
transform 1 0 28560 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _669_
timestamp 1698175906
transform -1 0 27888 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _670_
timestamp 1698175906
transform -1 0 27776 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _671_
timestamp 1698175906
transform -1 0 26544 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _672_
timestamp 1698175906
transform 1 0 22400 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _673_
timestamp 1698175906
transform -1 0 17920 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _674_
timestamp 1698175906
transform 1 0 17248 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _675_
timestamp 1698175906
transform 1 0 18592 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _676_
timestamp 1698175906
transform 1 0 19936 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _677_
timestamp 1698175906
transform -1 0 18816 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _678_
timestamp 1698175906
transform 1 0 20496 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _679_
timestamp 1698175906
transform -1 0 22960 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _680_
timestamp 1698175906
transform 1 0 24192 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _681_
timestamp 1698175906
transform -1 0 17248 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _682_
timestamp 1698175906
transform -1 0 15904 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _683_
timestamp 1698175906
transform 1 0 11088 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _684_
timestamp 1698175906
transform -1 0 13664 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _685_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _686_
timestamp 1698175906
transform -1 0 14000 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _687_
timestamp 1698175906
transform 1 0 13888 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _688_
timestamp 1698175906
transform 1 0 15680 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _689_
timestamp 1698175906
transform -1 0 15792 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _690_
timestamp 1698175906
transform -1 0 18592 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _691_
timestamp 1698175906
transform -1 0 18368 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _692_
timestamp 1698175906
transform -1 0 19264 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _693_
timestamp 1698175906
transform -1 0 17024 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _694_
timestamp 1698175906
transform -1 0 20048 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _695_
timestamp 1698175906
transform 1 0 14448 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _696_
timestamp 1698175906
transform -1 0 15344 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _697_
timestamp 1698175906
transform -1 0 12880 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _698_
timestamp 1698175906
transform 1 0 5376 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _699_
timestamp 1698175906
transform 1 0 6720 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _700_
timestamp 1698175906
transform -1 0 7728 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _701_
timestamp 1698175906
transform 1 0 6944 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _702_
timestamp 1698175906
transform 1 0 6608 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _703_
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _704_
timestamp 1698175906
transform -1 0 11424 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _705_
timestamp 1698175906
transform 1 0 6048 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _706_
timestamp 1698175906
transform 1 0 7504 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _707_
timestamp 1698175906
transform 1 0 8512 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _708_
timestamp 1698175906
transform 1 0 10416 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _709_
timestamp 1698175906
transform 1 0 11984 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _710_
timestamp 1698175906
transform 1 0 18144 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _711_
timestamp 1698175906
transform -1 0 18704 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _712_
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _713_
timestamp 1698175906
transform 1 0 11984 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _714_
timestamp 1698175906
transform -1 0 14672 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _715_
timestamp 1698175906
transform 1 0 9408 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _716_
timestamp 1698175906
transform -1 0 9184 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _717_
timestamp 1698175906
transform 1 0 6048 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _718_
timestamp 1698175906
transform 1 0 7952 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _719_
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _720_
timestamp 1698175906
transform 1 0 9968 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _721_
timestamp 1698175906
transform 1 0 11200 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _722_
timestamp 1698175906
transform 1 0 11872 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _723_
timestamp 1698175906
transform -1 0 11984 0 -1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _724_
timestamp 1698175906
transform -1 0 18480 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _725_
timestamp 1698175906
transform 1 0 10864 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _726_
timestamp 1698175906
transform -1 0 10192 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _727_
timestamp 1698175906
transform -1 0 11984 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _728_
timestamp 1698175906
transform 1 0 7616 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _729_
timestamp 1698175906
transform -1 0 12992 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _730_
timestamp 1698175906
transform -1 0 12320 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _731_
timestamp 1698175906
transform 1 0 9744 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _732_
timestamp 1698175906
transform 1 0 10304 0 -1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _733_
timestamp 1698175906
transform 1 0 10752 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _734_
timestamp 1698175906
transform -1 0 9184 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _735_
timestamp 1698175906
transform 1 0 7056 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _736_
timestamp 1698175906
transform 1 0 10528 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _737_
timestamp 1698175906
transform 1 0 12432 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _738_
timestamp 1698175906
transform 1 0 14336 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _739_
timestamp 1698175906
transform 1 0 15120 0 -1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _740_
timestamp 1698175906
transform 1 0 13776 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _741_
timestamp 1698175906
transform -1 0 13104 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _742_
timestamp 1698175906
transform -1 0 9184 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _743_
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _744_
timestamp 1698175906
transform 1 0 11984 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _745_
timestamp 1698175906
transform 1 0 10080 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _746_
timestamp 1698175906
transform -1 0 12544 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _747_
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _748_
timestamp 1698175906
transform -1 0 15120 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _749_
timestamp 1698175906
transform -1 0 14000 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _750_
timestamp 1698175906
transform -1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _751_
timestamp 1698175906
transform -1 0 9408 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _752_
timestamp 1698175906
transform 1 0 6832 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _753_
timestamp 1698175906
transform -1 0 10192 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _754_
timestamp 1698175906
transform -1 0 9296 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _755_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _756_
timestamp 1698175906
transform -1 0 15456 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _757_
timestamp 1698175906
transform -1 0 19376 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _758_
timestamp 1698175906
transform 1 0 16128 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _759_
timestamp 1698175906
transform 1 0 15120 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _760_
timestamp 1698175906
transform 1 0 11312 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _761_
timestamp 1698175906
transform -1 0 12880 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _762_
timestamp 1698175906
transform 1 0 10080 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _763_
timestamp 1698175906
transform -1 0 12768 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _764_
timestamp 1698175906
transform 1 0 16016 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _765_
timestamp 1698175906
transform 1 0 14224 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _766_
timestamp 1698175906
transform -1 0 20944 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _767_
timestamp 1698175906
transform -1 0 23520 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _768_
timestamp 1698175906
transform 1 0 18704 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _769_
timestamp 1698175906
transform 1 0 17808 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _770_
timestamp 1698175906
transform -1 0 23296 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _771_
timestamp 1698175906
transform 1 0 19152 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _772_
timestamp 1698175906
transform 1 0 19152 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _773_
timestamp 1698175906
transform -1 0 19376 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _774_
timestamp 1698175906
transform 1 0 18704 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _775_
timestamp 1698175906
transform 1 0 20048 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _776_
timestamp 1698175906
transform 1 0 21728 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _777_
timestamp 1698175906
transform -1 0 22736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _778_
timestamp 1698175906
transform 1 0 20272 0 -1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _779_
timestamp 1698175906
transform -1 0 22288 0 -1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _780_
timestamp 1698175906
transform -1 0 20944 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _781_
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _782_
timestamp 1698175906
transform 1 0 16352 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _783_
timestamp 1698175906
transform 1 0 25088 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _784_
timestamp 1698175906
transform 1 0 26544 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _785_
timestamp 1698175906
transform -1 0 26880 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _786_
timestamp 1698175906
transform 1 0 24192 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _787_
timestamp 1698175906
transform -1 0 26544 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _788_
timestamp 1698175906
transform 1 0 26880 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _789_
timestamp 1698175906
transform 1 0 26208 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _790_
timestamp 1698175906
transform -1 0 25984 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _791_
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _792_
timestamp 1698175906
transform 1 0 27328 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _793_
timestamp 1698175906
transform 1 0 26768 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _794_
timestamp 1698175906
transform 1 0 25984 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _795_
timestamp 1698175906
transform -1 0 26432 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _796_
timestamp 1698175906
transform -1 0 28336 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _797_
timestamp 1698175906
transform -1 0 27440 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _798_
timestamp 1698175906
transform -1 0 24192 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _799_
timestamp 1698175906
transform -1 0 19712 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _800_
timestamp 1698175906
transform 1 0 19712 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _801_
timestamp 1698175906
transform -1 0 20832 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _802_
timestamp 1698175906
transform -1 0 18592 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _803_
timestamp 1698175906
transform -1 0 17920 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _804_
timestamp 1698175906
transform 1 0 15680 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _805_
timestamp 1698175906
transform 1 0 15568 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _806_
timestamp 1698175906
transform -1 0 17920 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _807_
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _808_
timestamp 1698175906
transform 1 0 15792 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _809_
timestamp 1698175906
transform 1 0 14784 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _810_
timestamp 1698175906
transform -1 0 16016 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _811_
timestamp 1698175906
transform -1 0 15568 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _812_
timestamp 1698175906
transform -1 0 14560 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _813_
timestamp 1698175906
transform -1 0 12432 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _814_
timestamp 1698175906
transform 1 0 14560 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _815_
timestamp 1698175906
transform 1 0 15344 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _816_
timestamp 1698175906
transform -1 0 15344 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _817_
timestamp 1698175906
transform -1 0 14672 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _818_
timestamp 1698175906
transform -1 0 12992 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _819_
timestamp 1698175906
transform -1 0 17024 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _820_
timestamp 1698175906
transform -1 0 19264 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _821_
timestamp 1698175906
transform 1 0 16464 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _822_
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _823_
timestamp 1698175906
transform 1 0 18816 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _824_
timestamp 1698175906
transform -1 0 23072 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _825_
timestamp 1698175906
transform -1 0 23184 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _826_
timestamp 1698175906
transform 1 0 21504 0 1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _827_
timestamp 1698175906
transform 1 0 19936 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _828_
timestamp 1698175906
transform 1 0 21280 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _829_
timestamp 1698175906
transform -1 0 20272 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _830_
timestamp 1698175906
transform 1 0 19488 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _831_
timestamp 1698175906
transform -1 0 22624 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _832_
timestamp 1698175906
transform -1 0 20944 0 1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _833_
timestamp 1698175906
transform -1 0 16240 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _834_
timestamp 1698175906
transform -1 0 19600 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _835_
timestamp 1698175906
transform 1 0 18704 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _836_
timestamp 1698175906
transform -1 0 3472 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _837_
timestamp 1698175906
transform -1 0 18144 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _838_
timestamp 1698175906
transform -1 0 4592 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _839_
timestamp 1698175906
transform -1 0 2800 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _840_
timestamp 1698175906
transform -1 0 4144 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _841_
timestamp 1698175906
transform 1 0 4144 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _842_
timestamp 1698175906
transform 1 0 4928 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _843_
timestamp 1698175906
transform 1 0 4144 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _844_
timestamp 1698175906
transform 1 0 3248 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _845_
timestamp 1698175906
transform -1 0 6384 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _846_
timestamp 1698175906
transform 1 0 5152 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _847_
timestamp 1698175906
transform -1 0 5264 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _848_
timestamp 1698175906
transform 1 0 6048 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _849_
timestamp 1698175906
transform 1 0 6496 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _850_
timestamp 1698175906
transform -1 0 5488 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _851_
timestamp 1698175906
transform 1 0 5600 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _852_
timestamp 1698175906
transform -1 0 5264 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _853_
timestamp 1698175906
transform -1 0 3808 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _854_
timestamp 1698175906
transform -1 0 5376 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _855_
timestamp 1698175906
transform -1 0 4816 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _856_
timestamp 1698175906
transform -1 0 3136 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _857_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12096 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _858_
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _859_
timestamp 1698175906
transform 1 0 3024 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _860_
timestamp 1698175906
transform 1 0 1568 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _861_
timestamp 1698175906
transform 1 0 2016 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _862_
timestamp 1698175906
transform 1 0 5488 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _863_
timestamp 1698175906
transform 1 0 20832 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _864_
timestamp 1698175906
transform 1 0 18592 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _865_
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _866_
timestamp 1698175906
transform 1 0 19376 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _867_
timestamp 1698175906
transform 1 0 22848 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _868_
timestamp 1698175906
transform -1 0 27216 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _869_
timestamp 1698175906
transform -1 0 28896 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _870_
timestamp 1698175906
transform -1 0 32144 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _871_
timestamp 1698175906
transform 1 0 30912 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _872_
timestamp 1698175906
transform 1 0 31136 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _873_
timestamp 1698175906
transform 1 0 31136 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _874_
timestamp 1698175906
transform 1 0 31136 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _875_
timestamp 1698175906
transform 1 0 26880 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _876_
timestamp 1698175906
transform 1 0 31136 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _877_
timestamp 1698175906
transform -1 0 34384 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _878_
timestamp 1698175906
transform 1 0 31136 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _879_
timestamp 1698175906
transform 1 0 29456 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _880_
timestamp 1698175906
transform -1 0 30912 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _881_
timestamp 1698175906
transform 1 0 24304 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _882_
timestamp 1698175906
transform 1 0 23856 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _883_
timestamp 1698175906
transform 1 0 25536 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _884_
timestamp 1698175906
transform -1 0 32256 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _885_
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _886_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15120 0 1 6272
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _887_
timestamp 1698175906
transform 1 0 9296 0 1 3136
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _888_
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _889_
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _890_
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _891_
timestamp 1698175906
transform 1 0 7728 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _892_
timestamp 1698175906
transform -1 0 24864 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _893_
timestamp 1698175906
transform 1 0 18592 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _894_
timestamp 1698175906
transform 1 0 10080 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _895_
timestamp 1698175906
transform 1 0 8176 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _896_
timestamp 1698175906
transform 1 0 7168 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _897_
timestamp 1698175906
transform 1 0 6832 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _898_
timestamp 1698175906
transform 1 0 6944 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _899_
timestamp 1698175906
transform 1 0 14000 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _900_
timestamp 1698175906
transform 1 0 12880 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _901_
timestamp 1698175906
transform 1 0 17248 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _902_
timestamp 1698175906
transform 1 0 19376 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _903_
timestamp 1698175906
transform 1 0 21392 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _904_
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _905_
timestamp 1698175906
transform -1 0 30128 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _906_
timestamp 1698175906
transform -1 0 29456 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _907_
timestamp 1698175906
transform -1 0 26208 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _908_
timestamp 1698175906
transform -1 0 29680 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _909_
timestamp 1698175906
transform 1 0 22848 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _910_
timestamp 1698175906
transform 1 0 19600 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _911_
timestamp 1698175906
transform 1 0 13776 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _912_
timestamp 1698175906
transform 1 0 9856 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _913_
timestamp 1698175906
transform 1 0 10976 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _914_
timestamp 1698175906
transform -1 0 21616 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _915_
timestamp 1698175906
transform -1 0 24640 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _916_
timestamp 1698175906
transform -1 0 24416 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _917_
timestamp 1698175906
transform 1 0 18256 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _918_
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _919_
timestamp 1698175906
transform -1 0 18144 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _920_
timestamp 1698175906
transform -1 0 20048 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _921_
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _922_
timestamp 1698175906
transform 1 0 1680 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _923_
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _924_
timestamp 1698175906
transform 1 0 1904 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _925_
timestamp 1698175906
transform -1 0 8288 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _926_
timestamp 1698175906
transform 1 0 1568 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _927_
timestamp 1698175906
transform 1 0 1568 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__430__I $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__439__B
timestamp 1698175906
transform 1 0 20272 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__444__I
timestamp 1698175906
transform 1 0 18256 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__450__B
timestamp 1698175906
transform 1 0 17920 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__452__A2
timestamp 1698175906
transform -1 0 21616 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__457__A2
timestamp 1698175906
transform 1 0 18704 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__457__A3
timestamp 1698175906
transform 1 0 15344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__458__A1
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__470__A1
timestamp 1698175906
transform 1 0 21392 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__481__A2
timestamp 1698175906
transform -1 0 14000 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__490__A1
timestamp 1698175906
transform 1 0 17472 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__567__A1
timestamp 1698175906
transform 1 0 6048 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__581__I
timestamp 1698175906
transform 1 0 32928 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__599__A1
timestamp 1698175906
transform 1 0 24192 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__603__I
timestamp 1698175906
transform 1 0 19376 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__606__A1
timestamp 1698175906
transform 1 0 20944 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__674__A1
timestamp 1698175906
transform 1 0 18368 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__686__A1
timestamp 1698175906
transform -1 0 14224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__689__I
timestamp 1698175906
transform 1 0 14896 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__695__I
timestamp 1698175906
transform 1 0 16016 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__724__I
timestamp 1698175906
transform 1 0 17584 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__767__I
timestamp 1698175906
transform 1 0 22624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__780__C
timestamp 1698175906
transform 1 0 18928 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__830__A1
timestamp 1698175906
transform 1 0 20384 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__835__A1
timestamp 1698175906
transform -1 0 18704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__837__A1
timestamp 1698175906
transform -1 0 18592 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__859__CLK
timestamp 1698175906
transform 1 0 6272 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__860__CLK
timestamp 1698175906
transform 1 0 5040 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__861__CLK
timestamp 1698175906
transform 1 0 5712 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__862__CLK
timestamp 1698175906
transform 1 0 8960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__889__CLK
timestamp 1698175906
transform -1 0 5824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__890__CLK
timestamp 1698175906
transform 1 0 5040 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__891__CLK
timestamp 1698175906
transform 1 0 12544 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__912__CLK
timestamp 1698175906
transform 1 0 9632 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1698175906
transform -1 0 18032 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_0__f_wb_clk_i_I
timestamp 1698175906
transform 1 0 13552 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_1__f_wb_clk_i_I
timestamp 1698175906
transform 1 0 17024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_2__f_wb_clk_i_I
timestamp 1698175906
transform -1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_3__f_wb_clk_i_I
timestamp 1698175906
transform 1 0 19936 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_4__f_wb_clk_i_I
timestamp 1698175906
transform 1 0 22288 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_5__f_wb_clk_i_I
timestamp 1698175906
transform 1 0 26880 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_6__f_wb_clk_i_I
timestamp 1698175906
transform 1 0 22848 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_7__f_wb_clk_i_I
timestamp 1698175906
transform 1 0 26208 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698175906
transform -1 0 10864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18032 0 -1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_0__f_wb_clk_i
timestamp 1698175906
transform -1 0 12880 0 1 14112
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_1__f_wb_clk_i
timestamp 1698175906
transform 1 0 11424 0 -1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_2__f_wb_clk_i
timestamp 1698175906
transform -1 0 13104 0 1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_3__f_wb_clk_i
timestamp 1698175906
transform 1 0 13552 0 1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_4__f_wb_clk_i
timestamp 1698175906
transform -1 0 28112 0 1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_5__f_wb_clk_i
timestamp 1698175906
transform 1 0 27104 0 -1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_6__f_wb_clk_i
timestamp 1698175906
transform -1 0 28672 0 1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_7__f_wb_clk_i
timestamp 1698175906
transform 1 0 27104 0 -1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout5
timestamp 1698175906
transform 1 0 22624 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_36 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_40 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_44 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_49 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6832 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_57
timestamp 1698175906
transform 1 0 7728 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_59
timestamp 1698175906
transform 1 0 7952 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_64
timestamp 1698175906
transform 1 0 8512 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_104 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_128
timestamp 1698175906
transform 1 0 15680 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_167
timestamp 1698175906
transform 1 0 20048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698175906
transform 1 0 20272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698175906
transform 1 0 23856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698175906
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_244
timestamp 1698175906
transform 1 0 28672 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_280
timestamp 1698175906
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_284
timestamp 1698175906
transform 1 0 33152 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_292
timestamp 1698175906
transform 1 0 34048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_294
timestamp 1698175906
transform 1 0 34272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_52
timestamp 1698175906
transform 1 0 7168 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_78
timestamp 1698175906
transform 1 0 10080 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_82
timestamp 1698175906
transform 1 0 10528 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_91
timestamp 1698175906
transform 1 0 11536 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_128
timestamp 1698175906
transform 1 0 15680 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_138
timestamp 1698175906
transform 1 0 16800 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_142
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_146
timestamp 1698175906
transform 1 0 17696 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_150
timestamp 1698175906
transform 1 0 18144 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_152
timestamp 1698175906
transform 1 0 18368 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698175906
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_212
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_216
timestamp 1698175906
transform 1 0 25536 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_275
timestamp 1698175906
transform 1 0 32144 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698175906
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_290
timestamp 1698175906
transform 1 0 33824 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_294
timestamp 1698175906
transform 1 0 34272 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_4
timestamp 1698175906
transform 1 0 1792 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_39
timestamp 1698175906
transform 1 0 5712 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_81
timestamp 1698175906
transform 1 0 10416 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_104
timestamp 1698175906
transform 1 0 12992 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_148
timestamp 1698175906
transform 1 0 17920 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_187
timestamp 1698175906
transform 1 0 22288 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_189
timestamp 1698175906
transform 1 0 22512 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_198
timestamp 1698175906
transform 1 0 23520 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_237
timestamp 1698175906
transform 1 0 27888 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_255
timestamp 1698175906
transform 1 0 29904 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_257
timestamp 1698175906
transform 1 0 30128 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_10
timestamp 1698175906
transform 1 0 2464 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_21
timestamp 1698175906
transform 1 0 3696 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_31
timestamp 1698175906
transform 1 0 4816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_45
timestamp 1698175906
transform 1 0 6384 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_51
timestamp 1698175906
transform 1 0 7056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_88
timestamp 1698175906
transform 1 0 11200 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_92
timestamp 1698175906
transform 1 0 11648 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_94
timestamp 1698175906
transform 1 0 11872 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_108
timestamp 1698175906
transform 1 0 13440 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_120
timestamp 1698175906
transform 1 0 14784 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_124
timestamp 1698175906
transform 1 0 15232 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_138
timestamp 1698175906
transform 1 0 16800 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_150
timestamp 1698175906
transform 1 0 18144 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_163
timestamp 1698175906
transform 1 0 19600 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_171
timestamp 1698175906
transform 1 0 20496 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_195
timestamp 1698175906
transform 1 0 23184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_239
timestamp 1698175906
transform 1 0 28112 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_249
timestamp 1698175906
transform 1 0 29232 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_259
timestamp 1698175906
transform 1 0 30352 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_290
timestamp 1698175906
transform 1 0 33824 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_294
timestamp 1698175906
transform 1 0 34272 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_18
timestamp 1698175906
transform 1 0 3360 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_26
timestamp 1698175906
transform 1 0 4256 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_30
timestamp 1698175906
transform 1 0 4704 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_50
timestamp 1698175906
transform 1 0 6944 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_54
timestamp 1698175906
transform 1 0 7392 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_71
timestamp 1698175906
transform 1 0 9296 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_93
timestamp 1698175906
transform 1 0 11760 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_97
timestamp 1698175906
transform 1 0 12208 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_120
timestamp 1698175906
transform 1 0 14784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_122
timestamp 1698175906
transform 1 0 15008 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_160
timestamp 1698175906
transform 1 0 19264 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_168
timestamp 1698175906
transform 1 0 20160 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_172
timestamp 1698175906
transform 1 0 20608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_174
timestamp 1698175906
transform 1 0 20832 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_179
timestamp 1698175906
transform 1 0 21392 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_226
timestamp 1698175906
transform 1 0 26656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_242
timestamp 1698175906
transform 1 0 28448 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_244
timestamp 1698175906
transform 1 0 28672 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_255
timestamp 1698175906
transform 1 0 29904 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_293
timestamp 1698175906
transform 1 0 34160 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_41
timestamp 1698175906
transform 1 0 5936 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_45
timestamp 1698175906
transform 1 0 6384 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_54
timestamp 1698175906
transform 1 0 7392 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_80
timestamp 1698175906
transform 1 0 10304 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_87
timestamp 1698175906
transform 1 0 11088 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_97
timestamp 1698175906
transform 1 0 12208 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_99
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_109
timestamp 1698175906
transform 1 0 13552 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_194
timestamp 1698175906
transform 1 0 23072 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_201
timestamp 1698175906
transform 1 0 23856 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_209
timestamp 1698175906
transform 1 0 24752 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_227
timestamp 1698175906
transform 1 0 26768 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_242
timestamp 1698175906
transform 1 0 28448 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_246
timestamp 1698175906
transform 1 0 28896 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_259
timestamp 1698175906
transform 1 0 30352 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_263
timestamp 1698175906
transform 1 0 30800 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_265
timestamp 1698175906
transform 1 0 31024 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_290
timestamp 1698175906
transform 1 0 33824 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_294
timestamp 1698175906
transform 1 0 34272 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_6
timestamp 1698175906
transform 1 0 2016 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_8
timestamp 1698175906
transform 1 0 2240 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_27
timestamp 1698175906
transform 1 0 4368 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_33
timestamp 1698175906
transform 1 0 5040 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_57
timestamp 1698175906
transform 1 0 7728 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_61
timestamp 1698175906
transform 1 0 8176 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_80
timestamp 1698175906
transform 1 0 10304 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_162
timestamp 1698175906
transform 1 0 19488 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_170
timestamp 1698175906
transform 1 0 20384 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_174
timestamp 1698175906
transform 1 0 20832 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_189
timestamp 1698175906
transform 1 0 22512 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_191
timestamp 1698175906
transform 1 0 22736 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_233
timestamp 1698175906
transform 1 0 27440 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_242
timestamp 1698175906
transform 1 0 28448 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_244
timestamp 1698175906
transform 1 0 28672 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_251
timestamp 1698175906
transform 1 0 29456 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_253
timestamp 1698175906
transform 1 0 29680 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_6
timestamp 1698175906
transform 1 0 2016 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_8
timestamp 1698175906
transform 1 0 2240 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_25
timestamp 1698175906
transform 1 0 4144 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_29
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_40
timestamp 1698175906
transform 1 0 5824 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_52
timestamp 1698175906
transform 1 0 7168 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_54
timestamp 1698175906
transform 1 0 7392 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_63
timestamp 1698175906
transform 1 0 8400 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_67
timestamp 1698175906
transform 1 0 8848 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_69
timestamp 1698175906
transform 1 0 9072 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_82
timestamp 1698175906
transform 1 0 10528 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_86
timestamp 1698175906
transform 1 0 10976 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_209
timestamp 1698175906
transform 1 0 24752 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_220
timestamp 1698175906
transform 1 0 25984 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_227
timestamp 1698175906
transform 1 0 26768 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_275
timestamp 1698175906
transform 1 0 32144 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_279
timestamp 1698175906
transform 1 0 32592 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_290
timestamp 1698175906
transform 1 0 33824 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_294
timestamp 1698175906
transform 1 0 34272 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_6
timestamp 1698175906
transform 1 0 2016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_26
timestamp 1698175906
transform 1 0 4256 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_45
timestamp 1698175906
transform 1 0 6384 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_61
timestamp 1698175906
transform 1 0 8176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_75
timestamp 1698175906
transform 1 0 9744 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_93
timestamp 1698175906
transform 1 0 11760 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_168
timestamp 1698175906
transform 1 0 20160 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_172
timestamp 1698175906
transform 1 0 20608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_174
timestamp 1698175906
transform 1 0 20832 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_187
timestamp 1698175906
transform 1 0 22288 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_10
timestamp 1698175906
transform 1 0 2464 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_25
timestamp 1698175906
transform 1 0 4144 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_29
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_35
timestamp 1698175906
transform 1 0 5264 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_51
timestamp 1698175906
transform 1 0 7056 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_55
timestamp 1698175906
transform 1 0 7504 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_91
timestamp 1698175906
transform 1 0 11536 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_95
timestamp 1698175906
transform 1 0 11984 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_125
timestamp 1698175906
transform 1 0 15344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_150
timestamp 1698175906
transform 1 0 18144 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_180
timestamp 1698175906
transform 1 0 21504 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_184
timestamp 1698175906
transform 1 0 21952 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_186
timestamp 1698175906
transform 1 0 22176 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_189
timestamp 1698175906
transform 1 0 22512 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_205
timestamp 1698175906
transform 1 0 24304 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_209
timestamp 1698175906
transform 1 0 24752 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_222
timestamp 1698175906
transform 1 0 26208 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_226
timestamp 1698175906
transform 1 0 26656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_288
timestamp 1698175906
transform 1 0 33600 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_292
timestamp 1698175906
transform 1 0 34048 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_294
timestamp 1698175906
transform 1 0 34272 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_4
timestamp 1698175906
transform 1 0 1792 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_79
timestamp 1698175906
transform 1 0 10192 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_86
timestamp 1698175906
transform 1 0 10976 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_102
timestamp 1698175906
transform 1 0 12768 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_104
timestamp 1698175906
transform 1 0 12992 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_140
timestamp 1698175906
transform 1 0 17024 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_149
timestamp 1698175906
transform 1 0 18032 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_153
timestamp 1698175906
transform 1 0 18480 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_157
timestamp 1698175906
transform 1 0 18928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_159
timestamp 1698175906
transform 1 0 19152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_173
timestamp 1698175906
transform 1 0 20720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_194
timestamp 1698175906
transform 1 0 23072 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_202
timestamp 1698175906
transform 1 0 23968 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_204
timestamp 1698175906
transform 1 0 24192 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_234
timestamp 1698175906
transform 1 0 27552 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_242
timestamp 1698175906
transform 1 0 28448 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_244
timestamp 1698175906
transform 1 0 28672 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_261
timestamp 1698175906
transform 1 0 30576 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_265
timestamp 1698175906
transform 1 0 31024 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_10
timestamp 1698175906
transform 1 0 2464 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_40
timestamp 1698175906
transform 1 0 5824 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_56
timestamp 1698175906
transform 1 0 7616 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_78
timestamp 1698175906
transform 1 0 10080 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_87
timestamp 1698175906
transform 1 0 11088 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_89
timestamp 1698175906
transform 1 0 11312 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_177
timestamp 1698175906
transform 1 0 21168 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_208
timestamp 1698175906
transform 1 0 24640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_216
timestamp 1698175906
transform 1 0 25536 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_218
timestamp 1698175906
transform 1 0 25760 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_232
timestamp 1698175906
transform 1 0 27328 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_264
timestamp 1698175906
transform 1 0 30912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_266
timestamp 1698175906
transform 1 0 31136 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_275
timestamp 1698175906
transform 1 0 32144 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_279
timestamp 1698175906
transform 1 0 32592 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_290
timestamp 1698175906
transform 1 0 33824 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_294
timestamp 1698175906
transform 1 0 34272 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_18
timestamp 1698175906
transform 1 0 3360 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_52
timestamp 1698175906
transform 1 0 7168 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_98
timestamp 1698175906
transform 1 0 12320 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_102
timestamp 1698175906
transform 1 0 12768 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_104
timestamp 1698175906
transform 1 0 12992 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_109
timestamp 1698175906
transform 1 0 13552 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_116
timestamp 1698175906
transform 1 0 14336 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_124
timestamp 1698175906
transform 1 0 15232 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_127
timestamp 1698175906
transform 1 0 15568 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_135
timestamp 1698175906
transform 1 0 16464 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_139
timestamp 1698175906
transform 1 0 16912 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_142
timestamp 1698175906
transform 1 0 17248 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_146
timestamp 1698175906
transform 1 0 17696 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_179
timestamp 1698175906
transform 1 0 21392 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_195
timestamp 1698175906
transform 1 0 23184 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_199
timestamp 1698175906
transform 1 0 23632 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_235
timestamp 1698175906
transform 1 0 27664 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_243
timestamp 1698175906
transform 1 0 28560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_255
timestamp 1698175906
transform 1 0 29904 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_263
timestamp 1698175906
transform 1 0 30800 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_265
timestamp 1698175906
transform 1 0 31024 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_18
timestamp 1698175906
transform 1 0 3360 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_26
timestamp 1698175906
transform 1 0 4256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_50
timestamp 1698175906
transform 1 0 6944 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_54
timestamp 1698175906
transform 1 0 7392 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_60
timestamp 1698175906
transform 1 0 8064 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_68
timestamp 1698175906
transform 1 0 8960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_76
timestamp 1698175906
transform 1 0 9856 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_95
timestamp 1698175906
transform 1 0 11984 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_111
timestamp 1698175906
transform 1 0 13776 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_119
timestamp 1698175906
transform 1 0 14672 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_132
timestamp 1698175906
transform 1 0 16128 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_159
timestamp 1698175906
transform 1 0 19152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_163
timestamp 1698175906
transform 1 0 19600 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_165
timestamp 1698175906
transform 1 0 19824 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_172
timestamp 1698175906
transform 1 0 20608 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_176
timestamp 1698175906
transform 1 0 21056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_194
timestamp 1698175906
transform 1 0 23072 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_196
timestamp 1698175906
transform 1 0 23296 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_202
timestamp 1698175906
transform 1 0 23968 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698175906
transform 1 0 24416 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_278
timestamp 1698175906
transform 1 0 32480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_290
timestamp 1698175906
transform 1 0 33824 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_294
timestamp 1698175906
transform 1 0 34272 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_31
timestamp 1698175906
transform 1 0 4816 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_43
timestamp 1698175906
transform 1 0 6160 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_51
timestamp 1698175906
transform 1 0 7056 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_103
timestamp 1698175906
transform 1 0 12880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_111
timestamp 1698175906
transform 1 0 13776 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_127
timestamp 1698175906
transform 1 0 15568 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_133
timestamp 1698175906
transform 1 0 16240 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_153
timestamp 1698175906
transform 1 0 18480 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_157
timestamp 1698175906
transform 1 0 18928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_159
timestamp 1698175906
transform 1 0 19152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_206
timestamp 1698175906
transform 1 0 24416 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_222
timestamp 1698175906
transform 1 0 26208 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_241
timestamp 1698175906
transform 1 0 28336 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_255
timestamp 1698175906
transform 1 0 29904 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_259
timestamp 1698175906
transform 1 0 30352 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_284
timestamp 1698175906
transform 1 0 33152 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_292
timestamp 1698175906
transform 1 0 34048 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_294
timestamp 1698175906
transform 1 0 34272 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_34
timestamp 1698175906
transform 1 0 5152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_36
timestamp 1698175906
transform 1 0 5376 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_80
timestamp 1698175906
transform 1 0 10304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_84
timestamp 1698175906
transform 1 0 10752 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_115
timestamp 1698175906
transform 1 0 14224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_117
timestamp 1698175906
transform 1 0 14448 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_131
timestamp 1698175906
transform 1 0 16016 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_142
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_146
timestamp 1698175906
transform 1 0 17696 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_199
timestamp 1698175906
transform 1 0 23632 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_207
timestamp 1698175906
transform 1 0 24528 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698175906
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_212
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_216
timestamp 1698175906
transform 1 0 25536 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_218
timestamp 1698175906
transform 1 0 25760 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_225
timestamp 1698175906
transform 1 0 26544 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_229
timestamp 1698175906
transform 1 0 26992 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_231
timestamp 1698175906
transform 1 0 27216 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_237
timestamp 1698175906
transform 1 0 27888 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698175906
transform 1 0 32592 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_290
timestamp 1698175906
transform 1 0 33824 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_294
timestamp 1698175906
transform 1 0 34272 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_41
timestamp 1698175906
transform 1 0 5936 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_43
timestamp 1698175906
transform 1 0 6160 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_46
timestamp 1698175906
transform 1 0 6496 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_62
timestamp 1698175906
transform 1 0 8288 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_70
timestamp 1698175906
transform 1 0 9184 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_119
timestamp 1698175906
transform 1 0 14672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_160
timestamp 1698175906
transform 1 0 19264 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_168
timestamp 1698175906
transform 1 0 20160 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1698175906
transform 1 0 20608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698175906
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_184
timestamp 1698175906
transform 1 0 21952 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_193
timestamp 1698175906
transform 1 0 22960 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_195
timestamp 1698175906
transform 1 0 23184 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_210
timestamp 1698175906
transform 1 0 24864 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_226
timestamp 1698175906
transform 1 0 26656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_228
timestamp 1698175906
transform 1 0 26880 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698175906
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_261
timestamp 1698175906
transform 1 0 30576 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_265
timestamp 1698175906
transform 1 0 31024 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_2
timestamp 1698175906
transform 1 0 1568 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_10
timestamp 1698175906
transform 1 0 2464 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_14
timestamp 1698175906
transform 1 0 2912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_44
timestamp 1698175906
transform 1 0 6272 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_46
timestamp 1698175906
transform 1 0 6496 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_57
timestamp 1698175906
transform 1 0 7728 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_78
timestamp 1698175906
transform 1 0 10080 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_94
timestamp 1698175906
transform 1 0 11872 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_99
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_104
timestamp 1698175906
transform 1 0 12992 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_118
timestamp 1698175906
transform 1 0 14560 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_241
timestamp 1698175906
transform 1 0 28336 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_290
timestamp 1698175906
transform 1 0 33824 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_294
timestamp 1698175906
transform 1 0 34272 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_31
timestamp 1698175906
transform 1 0 4816 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_41
timestamp 1698175906
transform 1 0 5936 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_65
timestamp 1698175906
transform 1 0 8624 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_90
timestamp 1698175906
transform 1 0 11424 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_98
timestamp 1698175906
transform 1 0 12320 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_102
timestamp 1698175906
transform 1 0 12768 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_104
timestamp 1698175906
transform 1 0 12992 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_123
timestamp 1698175906
transform 1 0 15120 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_127
timestamp 1698175906
transform 1 0 15568 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_137
timestamp 1698175906
transform 1 0 16688 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_141
timestamp 1698175906
transform 1 0 17136 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_154
timestamp 1698175906
transform 1 0 18592 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_160
timestamp 1698175906
transform 1 0 19264 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_168
timestamp 1698175906
transform 1 0 20160 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_172
timestamp 1698175906
transform 1 0 20608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698175906
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_177
timestamp 1698175906
transform 1 0 21168 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_209
timestamp 1698175906
transform 1 0 24752 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_217
timestamp 1698175906
transform 1 0 25648 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_276
timestamp 1698175906
transform 1 0 32256 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_292
timestamp 1698175906
transform 1 0 34048 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_294
timestamp 1698175906
transform 1 0 34272 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_2
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_34
timestamp 1698175906
transform 1 0 5152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_103
timestamp 1698175906
transform 1 0 12880 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_150
timestamp 1698175906
transform 1 0 18144 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_183
timestamp 1698175906
transform 1 0 21840 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_187
timestamp 1698175906
transform 1 0 22288 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_189
timestamp 1698175906
transform 1 0 22512 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_204
timestamp 1698175906
transform 1 0 24192 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_208
timestamp 1698175906
transform 1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_212
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_220
timestamp 1698175906
transform 1 0 25984 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_290
timestamp 1698175906
transform 1 0 33824 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_294
timestamp 1698175906
transform 1 0 34272 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_31
timestamp 1698175906
transform 1 0 4816 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_45
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_61
timestamp 1698175906
transform 1 0 8176 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_79
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_90
timestamp 1698175906
transform 1 0 11424 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_104
timestamp 1698175906
transform 1 0 12992 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_115
timestamp 1698175906
transform 1 0 14224 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_119
timestamp 1698175906
transform 1 0 14672 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_123
timestamp 1698175906
transform 1 0 15120 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_139
timestamp 1698175906
transform 1 0 16912 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_141
timestamp 1698175906
transform 1 0 17136 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_150
timestamp 1698175906
transform 1 0 18144 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_154
timestamp 1698175906
transform 1 0 18592 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_170
timestamp 1698175906
transform 1 0 20384 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698175906
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_177
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_181
timestamp 1698175906
transform 1 0 21616 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_188
timestamp 1698175906
transform 1 0 22400 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698175906
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_247
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_279
timestamp 1698175906
transform 1 0 32592 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_40
timestamp 1698175906
transform 1 0 5824 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_48
timestamp 1698175906
transform 1 0 6720 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_50
timestamp 1698175906
transform 1 0 6944 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_63
timestamp 1698175906
transform 1 0 8400 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_103
timestamp 1698175906
transform 1 0 12880 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_129
timestamp 1698175906
transform 1 0 15792 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_133
timestamp 1698175906
transform 1 0 16240 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_160
timestamp 1698175906
transform 1 0 19264 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_164
timestamp 1698175906
transform 1 0 19712 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_166
timestamp 1698175906
transform 1 0 19936 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_208
timestamp 1698175906
transform 1 0 24640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_245
timestamp 1698175906
transform 1 0 28784 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_277
timestamp 1698175906
transform 1 0 32368 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698175906
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_290
timestamp 1698175906
transform 1 0 33824 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_294
timestamp 1698175906
transform 1 0 34272 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_6
timestamp 1698175906
transform 1 0 2016 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_33
timestamp 1698175906
transform 1 0 5040 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_74
timestamp 1698175906
transform 1 0 9632 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_93
timestamp 1698175906
transform 1 0 11760 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_97
timestamp 1698175906
transform 1 0 12208 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_104
timestamp 1698175906
transform 1 0 12992 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_118
timestamp 1698175906
transform 1 0 14560 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_126
timestamp 1698175906
transform 1 0 15456 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_154
timestamp 1698175906
transform 1 0 18592 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_170
timestamp 1698175906
transform 1 0 20384 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698175906
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_177
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_185
timestamp 1698175906
transform 1 0 22064 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_189
timestamp 1698175906
transform 1 0 22512 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_191
timestamp 1698175906
transform 1 0 22736 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_241
timestamp 1698175906
transform 1 0 28336 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_247
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_279
timestamp 1698175906
transform 1 0 32592 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_2
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_10
timestamp 1698175906
transform 1 0 2464 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_14
timestamp 1698175906
transform 1 0 2912 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_16
timestamp 1698175906
transform 1 0 3136 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_40
timestamp 1698175906
transform 1 0 5824 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_56
timestamp 1698175906
transform 1 0 7616 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_64
timestamp 1698175906
transform 1 0 8512 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698175906
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_80
timestamp 1698175906
transform 1 0 10304 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_87
timestamp 1698175906
transform 1 0 11088 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_95
timestamp 1698175906
transform 1 0 11984 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_130
timestamp 1698175906
transform 1 0 15904 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_144
timestamp 1698175906
transform 1 0 17472 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_153
timestamp 1698175906
transform 1 0 18480 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_164
timestamp 1698175906
transform 1 0 19712 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_168
timestamp 1698175906
transform 1 0 20160 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_191
timestamp 1698175906
transform 1 0 22736 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_212
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_216
timestamp 1698175906
transform 1 0 25536 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_218
timestamp 1698175906
transform 1 0 25760 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_253
timestamp 1698175906
transform 1 0 29680 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_269
timestamp 1698175906
transform 1 0 31472 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_277
timestamp 1698175906
transform 1 0 32368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698175906
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_290
timestamp 1698175906
transform 1 0 33824 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_294
timestamp 1698175906
transform 1 0 34272 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_31
timestamp 1698175906
transform 1 0 4816 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_45
timestamp 1698175906
transform 1 0 6384 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_53
timestamp 1698175906
transform 1 0 7280 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_206
timestamp 1698175906
transform 1 0 24416 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_210
timestamp 1698175906
transform 1 0 24864 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_236
timestamp 1698175906
transform 1 0 27776 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698175906
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_279
timestamp 1698175906
transform 1 0 32592 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_2
timestamp 1698175906
transform 1 0 1568 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_4
timestamp 1698175906
transform 1 0 1792 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_50
timestamp 1698175906
transform 1 0 6944 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_58
timestamp 1698175906
transform 1 0 7840 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_74
timestamp 1698175906
transform 1 0 9632 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_105
timestamp 1698175906
transform 1 0 13104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_107
timestamp 1698175906
transform 1 0 13328 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_133
timestamp 1698175906
transform 1 0 16240 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_137
timestamp 1698175906
transform 1 0 16688 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698175906
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_196
timestamp 1698175906
transform 1 0 23296 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_257
timestamp 1698175906
transform 1 0 30128 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_273
timestamp 1698175906
transform 1 0 31920 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698175906
transform 1 0 32368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_290
timestamp 1698175906
transform 1 0 33824 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_294
timestamp 1698175906
transform 1 0 34272 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_2
timestamp 1698175906
transform 1 0 1568 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_18
timestamp 1698175906
transform 1 0 3360 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_26
timestamp 1698175906
transform 1 0 4256 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_28
timestamp 1698175906
transform 1 0 4480 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_45
timestamp 1698175906
transform 1 0 6384 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_49
timestamp 1698175906
transform 1 0 6832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_79
timestamp 1698175906
transform 1 0 10192 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_83
timestamp 1698175906
transform 1 0 10640 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_99
timestamp 1698175906
transform 1 0 12432 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_150
timestamp 1698175906
transform 1 0 18144 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_154
timestamp 1698175906
transform 1 0 18592 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_167
timestamp 1698175906
transform 1 0 20048 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_171
timestamp 1698175906
transform 1 0 20496 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_177
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_209
timestamp 1698175906
transform 1 0 24752 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_231
timestamp 1698175906
transform 1 0 27216 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_239
timestamp 1698175906
transform 1 0 28112 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_243
timestamp 1698175906
transform 1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_279
timestamp 1698175906
transform 1 0 32592 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_2
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_18
timestamp 1698175906
transform 1 0 3360 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_22
timestamp 1698175906
transform 1 0 3808 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_50
timestamp 1698175906
transform 1 0 6944 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_80
timestamp 1698175906
transform 1 0 10304 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_84
timestamp 1698175906
transform 1 0 10752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_110
timestamp 1698175906
transform 1 0 13664 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_112
timestamp 1698175906
transform 1 0 13888 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_115
timestamp 1698175906
transform 1 0 14224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_117
timestamp 1698175906
transform 1 0 14448 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_130
timestamp 1698175906
transform 1 0 15904 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_138
timestamp 1698175906
transform 1 0 16800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_146
timestamp 1698175906
transform 1 0 17696 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_148
timestamp 1698175906
transform 1 0 17920 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_161
timestamp 1698175906
transform 1 0 19376 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_163
timestamp 1698175906
transform 1 0 19600 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_220
timestamp 1698175906
transform 1 0 25984 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_251
timestamp 1698175906
transform 1 0 29456 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_267
timestamp 1698175906
transform 1 0 31248 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_275
timestamp 1698175906
transform 1 0 32144 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698175906
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_290
timestamp 1698175906
transform 1 0 33824 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_294
timestamp 1698175906
transform 1 0 34272 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_2
timestamp 1698175906
transform 1 0 1568 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_22
timestamp 1698175906
transform 1 0 3808 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_45
timestamp 1698175906
transform 1 0 6384 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_78
timestamp 1698175906
transform 1 0 10080 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_102
timestamp 1698175906
transform 1 0 12768 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_104
timestamp 1698175906
transform 1 0 12992 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_139
timestamp 1698175906
transform 1 0 16912 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_155
timestamp 1698175906
transform 1 0 18704 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_172
timestamp 1698175906
transform 1 0 20608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_177
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_179
timestamp 1698175906
transform 1 0 21392 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_234
timestamp 1698175906
transform 1 0 27552 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_242
timestamp 1698175906
transform 1 0 28448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_279
timestamp 1698175906
transform 1 0 32592 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_31
timestamp 1698175906
transform 1 0 4816 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_62
timestamp 1698175906
transform 1 0 8288 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_74
timestamp 1698175906
transform 1 0 9632 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_79
timestamp 1698175906
transform 1 0 10192 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_87
timestamp 1698175906
transform 1 0 11088 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_101
timestamp 1698175906
transform 1 0 12656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_142
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_146
timestamp 1698175906
transform 1 0 17696 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_202
timestamp 1698175906
transform 1 0 23968 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_220
timestamp 1698175906
transform 1 0 25984 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_252
timestamp 1698175906
transform 1 0 29568 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_268
timestamp 1698175906
transform 1 0 31360 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698175906
transform 1 0 32256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_290
timestamp 1698175906
transform 1 0 33824 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_294
timestamp 1698175906
transform 1 0 34272 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_81
timestamp 1698175906
transform 1 0 10416 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_89
timestamp 1698175906
transform 1 0 11312 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_93
timestamp 1698175906
transform 1 0 11760 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_103
timestamp 1698175906
transform 1 0 12880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_111
timestamp 1698175906
transform 1 0 13776 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_177 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_241
timestamp 1698175906
transform 1 0 28336 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_279
timestamp 1698175906
transform 1 0 32592 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_18
timestamp 1698175906
transform 1 0 3360 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_36
timestamp 1698175906
transform 1 0 5376 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_68
timestamp 1698175906
transform 1 0 8960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_76
timestamp 1698175906
transform 1 0 9856 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_107
timestamp 1698175906
transform 1 0 13328 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_139
timestamp 1698175906
transform 1 0 16912 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_142
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_158
timestamp 1698175906
transform 1 0 19040 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_174
timestamp 1698175906
transform 1 0 20832 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698175906
transform 1 0 24416 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_290
timestamp 1698175906
transform 1 0 33824 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_294
timestamp 1698175906
transform 1 0 34272 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_53
timestamp 1698175906
transform 1 0 7280 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_90
timestamp 1698175906
transform 1 0 11424 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_98
timestamp 1698175906
transform 1 0 12320 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_102
timestamp 1698175906
transform 1 0 12768 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_104
timestamp 1698175906
transform 1 0 12992 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_279
timestamp 1698175906
transform 1 0 32592 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_290
timestamp 1698175906
transform 1 0 33824 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_294
timestamp 1698175906
transform 1 0 34272 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_279
timestamp 1698175906
transform 1 0 32592 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_290
timestamp 1698175906
transform 1 0 33824 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_294
timestamp 1698175906
transform 1 0 34272 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_36
timestamp 1698175906
transform 1 0 5376 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_70
timestamp 1698175906
transform 1 0 9184 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_104
timestamp 1698175906
transform 1 0 12992 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_138
timestamp 1698175906
transform 1 0 16800 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_172
timestamp 1698175906
transform 1 0 20608 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_206
timestamp 1698175906
transform 1 0 24416 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_240
timestamp 1698175906
transform 1 0 28224 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_274
timestamp 1698175906
transform 1 0 32032 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_290
timestamp 1698175906
transform 1 0 33824 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_294
timestamp 1698175906
transform 1 0 34272 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input1
timestamp 1698175906
transform 1 0 10864 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18032 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 25088 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform -1 0 31808 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_37 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 34608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_38
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 34608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_39
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 34608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_40
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 34608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_41
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 34608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_42
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 34608 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_43
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 34608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_44
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 34608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_45
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 34608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 34608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 34608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 34608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 34608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 34608 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 34608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 34608 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 34608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 34608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 34608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 34608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 34608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 34608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 34608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 34608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 34608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 34608 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 34608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 34608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 34608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 34608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 34608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 34608 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 34608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 34608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 34608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 34608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 34608 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_74 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_75
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_76
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_77
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_78
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_79
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_80
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_81
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_82
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_83
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_84
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_85
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_86
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_87
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_88
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_89
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_90
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_91
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_92
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_93
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_94
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_95
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_96
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_97
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_98
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_99
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_100
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_101
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_102
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_103
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_104
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_105
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_106
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_107
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_108
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_109
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_110
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_111
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_112
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_113
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_114
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_115
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_116
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_117
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_118
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_119
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_120
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_121
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_122
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_123
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_124
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_125
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_126
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_127
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_128
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_129
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_130
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_131
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_132
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_133
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_134
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_135
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_136
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_137
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_138
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_139
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_140
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_141
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_142
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_143
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_144
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_145
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_146
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_147
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_148
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_149
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_150
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_151
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_152
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_153
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_154
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_155
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_156
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_157
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_158
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_159
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_160
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_161
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_162
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_163
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_164
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_165
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_166
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_167
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_168
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_169
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_170
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_171
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_172
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_173
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_174
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_175
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_176
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_177
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_178
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_179
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_180
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_181
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_182
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_183
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_184
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_185
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_186
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_187
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_188
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_189
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_190
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_191
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_192
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_193
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_194
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_195
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_196
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_197
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_198
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_199
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_200
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_201
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_202
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_203
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_204
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_205
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_206
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_207
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_208
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_209
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_210
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_211
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_212
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_213
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_214
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_215
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_216
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_217
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_218
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_219
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_220
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_221
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_222
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_223
timestamp 1698175906
transform 1 0 8960 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_224
timestamp 1698175906
transform 1 0 12768 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_225
timestamp 1698175906
transform 1 0 16576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_226
timestamp 1698175906
transform 1 0 20384 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_227
timestamp 1698175906
transform 1 0 24192 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_228
timestamp 1698175906
transform 1 0 28000 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_229
timestamp 1698175906
transform 1 0 31808 0 1 31360
box -86 -86 310 870
<< labels >>
flabel metal2 s 17920 0 18032 800 0 FreeSans 448 90 0 0 io_out[0]
port 0 nsew signal tristate
flabel metal2 s 25088 0 25200 800 0 FreeSans 448 90 0 0 io_out[1]
port 1 nsew signal tristate
flabel metal2 s 32256 0 32368 800 0 FreeSans 448 90 0 0 io_out[2]
port 2 nsew signal tristate
flabel metal2 s 10752 0 10864 800 0 FreeSans 448 90 0 0 rst_n
port 3 nsew signal input
flabel metal4 s 5342 3076 5662 32204 0 FreeSans 1280 90 0 0 vdd
port 4 nsew power bidirectional
flabel metal4 s 13658 3076 13978 32204 0 FreeSans 1280 90 0 0 vdd
port 4 nsew power bidirectional
flabel metal4 s 21974 3076 22294 32204 0 FreeSans 1280 90 0 0 vdd
port 4 nsew power bidirectional
flabel metal4 s 30290 3076 30610 32204 0 FreeSans 1280 90 0 0 vdd
port 4 nsew power bidirectional
flabel metal4 s 9500 3076 9820 32204 0 FreeSans 1280 90 0 0 vss
port 5 nsew ground bidirectional
flabel metal4 s 17816 3076 18136 32204 0 FreeSans 1280 90 0 0 vss
port 5 nsew ground bidirectional
flabel metal4 s 26132 3076 26452 32204 0 FreeSans 1280 90 0 0 vss
port 5 nsew ground bidirectional
flabel metal4 s 34448 3076 34768 32204 0 FreeSans 1280 90 0 0 vss
port 5 nsew ground bidirectional
flabel metal2 s 3584 0 3696 800 0 FreeSans 448 90 0 0 wb_clk_i
port 6 nsew signal input
rlabel metal1 17976 32144 17976 32144 0 vdd
rlabel via1 18056 31360 18056 31360 0 vss
rlabel metal2 13104 27720 13104 27720 0 LFSR\[0\]
rlabel metal2 11760 26936 11760 26936 0 LFSR\[1\]
rlabel metal2 11144 24080 11144 24080 0 LFSR\[2\]
rlabel metal2 9912 24416 9912 24416 0 LFSR\[3\]
rlabel metal2 11704 23352 11704 23352 0 LFSR\[4\]
rlabel metal2 16912 27160 16912 27160 0 LFSR\[5\]
rlabel metal2 15288 24528 15288 24528 0 LFSR\[6\]
rlabel metal2 21672 17248 21672 17248 0 OP_reg
rlabel metal2 17472 8232 17472 8232 0 PC\[0\]
rlabel metal2 16744 9744 16744 9744 0 PC\[1\]
rlabel metal2 17864 5712 17864 5712 0 PC\[2\]
rlabel metal2 3920 12152 3920 12152 0 PC\[3\]
rlabel metal2 5656 14560 5656 14560 0 PC\[4\]
rlabel metal3 11200 13832 11200 13832 0 PC\[5\]
rlabel metal2 13048 10976 13048 10976 0 _000_
rlabel metal3 12488 11480 12488 11480 0 _001_
rlabel metal2 5152 16856 5152 16856 0 _002_
rlabel metal2 2408 14504 2408 14504 0 _003_
rlabel metal2 2968 15120 2968 15120 0 _004_
rlabel metal2 6496 13944 6496 13944 0 _005_
rlabel metal2 21784 9520 21784 9520 0 _006_
rlabel metal2 21336 6048 21336 6048 0 _007_
rlabel metal2 21560 4312 21560 4312 0 _008_
rlabel metal3 22008 4200 22008 4200 0 _009_
rlabel metal2 23912 8344 23912 8344 0 _010_
rlabel metal2 26264 5432 26264 5432 0 _011_
rlabel metal2 27944 4760 27944 4760 0 _012_
rlabel metal2 31192 4648 31192 4648 0 _013_
rlabel metal2 30520 5264 30520 5264 0 _014_
rlabel metal2 32088 5432 32088 5432 0 _015_
rlabel metal2 31752 7896 31752 7896 0 _016_
rlabel metal2 33040 7560 33040 7560 0 _017_
rlabel metal2 27832 9352 27832 9352 0 _018_
rlabel metal2 31416 11704 31416 11704 0 _019_
rlabel metal2 33432 13384 33432 13384 0 _020_
rlabel metal2 32088 15904 32088 15904 0 _021_
rlabel metal2 31976 15904 31976 15904 0 _022_
rlabel metal2 29960 14112 29960 14112 0 _023_
rlabel metal2 25704 10864 25704 10864 0 _024_
rlabel metal2 24808 13272 24808 13272 0 _025_
rlabel metal2 26600 19096 26600 19096 0 _026_
rlabel metal2 28952 17304 28952 17304 0 _027_
rlabel metal2 26040 15960 26040 15960 0 _028_
rlabel metal2 16072 5936 16072 5936 0 _029_
rlabel metal2 9016 4032 9016 4032 0 _030_
rlabel metal2 11480 5936 11480 5936 0 _031_
rlabel metal2 3136 4984 3136 4984 0 _032_
rlabel metal2 2520 13944 2520 13944 0 _033_
rlabel metal3 9800 12264 9800 12264 0 _034_
rlabel metal2 24472 16464 24472 16464 0 _035_
rlabel metal2 19544 18816 19544 18816 0 _036_
rlabel metal2 12264 27440 12264 27440 0 _037_
rlabel metal2 9520 28504 9520 28504 0 _038_
rlabel metal2 8904 25704 8904 25704 0 _039_
rlabel metal2 8904 23744 8904 23744 0 _040_
rlabel metal2 8400 23352 8400 23352 0 _041_
rlabel metal2 15008 26936 15008 26936 0 _042_
rlabel metal2 14504 25872 14504 25872 0 _043_
rlabel metal2 18200 26712 18200 26712 0 _044_
rlabel metal3 19656 23240 19656 23240 0 _045_
rlabel metal2 22344 19432 22344 19432 0 _046_
rlabel metal3 21392 22232 21392 22232 0 _047_
rlabel metal3 28112 23240 28112 23240 0 _048_
rlabel metal2 28504 25200 28504 25200 0 _049_
rlabel metal2 25312 25592 25312 25592 0 _050_
rlabel metal3 28392 20888 28392 20888 0 _051_
rlabel metal2 23912 19544 23912 19544 0 _052_
rlabel metal2 20552 27048 20552 27048 0 _053_
rlabel metal2 16072 18032 16072 18032 0 _054_
rlabel metal2 10808 16520 10808 16520 0 _055_
rlabel metal2 11928 15624 11928 15624 0 _056_
rlabel metal2 20664 17192 20664 17192 0 _057_
rlabel metal2 23688 12488 23688 12488 0 _058_
rlabel metal3 22512 14616 22512 14616 0 _059_
rlabel metal2 19656 9800 19656 9800 0 _060_
rlabel metal2 18200 12488 18200 12488 0 _061_
rlabel metal2 15960 23576 15960 23576 0 _062_
rlabel metal2 19096 3920 19096 3920 0 _063_
rlabel metal2 2520 19936 2520 19936 0 _064_
rlabel metal3 3920 19880 3920 19880 0 _065_
rlabel metal3 4088 22232 4088 22232 0 _066_
rlabel metal3 4816 23016 4816 23016 0 _067_
rlabel metal3 6832 26376 6832 26376 0 _068_
rlabel metal2 3304 26040 3304 26040 0 _069_
rlabel metal2 2632 25928 2632 25928 0 _070_
rlabel metal2 6776 5880 6776 5880 0 _071_
rlabel metal2 6944 11592 6944 11592 0 _072_
rlabel metal3 12992 9576 12992 9576 0 _073_
rlabel metal2 19096 8680 19096 8680 0 _074_
rlabel metal2 16912 11144 16912 11144 0 _075_
rlabel metal2 22792 25144 22792 25144 0 _076_
rlabel metal2 22568 25424 22568 25424 0 _077_
rlabel metal2 20888 25032 20888 25032 0 _078_
rlabel metal2 23016 24976 23016 24976 0 _079_
rlabel metal3 16744 14504 16744 14504 0 _080_
rlabel metal2 20216 24640 20216 24640 0 _081_
rlabel metal3 19432 19320 19432 19320 0 _082_
rlabel metal2 4648 25424 4648 25424 0 _083_
rlabel metal2 6328 22680 6328 22680 0 _084_
rlabel metal2 5768 21112 5768 21112 0 _085_
rlabel metal2 16520 11816 16520 11816 0 _086_
rlabel metal2 17752 19320 17752 19320 0 _087_
rlabel metal2 17192 15400 17192 15400 0 _088_
rlabel metal3 18592 15848 18592 15848 0 _089_
rlabel metal2 17752 12600 17752 12600 0 _090_
rlabel metal3 20160 11592 20160 11592 0 _091_
rlabel metal2 19544 13216 19544 13216 0 _092_
rlabel metal2 18424 12488 18424 12488 0 _093_
rlabel metal2 19376 9800 19376 9800 0 _094_
rlabel metal2 17304 9408 17304 9408 0 _095_
rlabel metal2 10136 13608 10136 13608 0 _096_
rlabel metal2 10696 14000 10696 14000 0 _097_
rlabel metal3 11704 12712 11704 12712 0 _098_
rlabel metal2 16296 7280 16296 7280 0 _099_
rlabel metal2 15848 9240 15848 9240 0 _100_
rlabel metal2 11928 9464 11928 9464 0 _101_
rlabel metal2 11704 13216 11704 13216 0 _102_
rlabel metal2 11256 13384 11256 13384 0 _103_
rlabel metal3 10416 12376 10416 12376 0 _104_
rlabel metal3 2464 12152 2464 12152 0 _105_
rlabel metal2 15400 8400 15400 8400 0 _106_
rlabel metal2 11704 8288 11704 8288 0 _107_
rlabel metal2 2520 7672 2520 7672 0 _108_
rlabel metal2 5656 8288 5656 8288 0 _109_
rlabel metal3 13496 6552 13496 6552 0 _110_
rlabel metal2 6888 6160 6888 6160 0 _111_
rlabel metal2 18312 8960 18312 8960 0 _112_
rlabel metal2 17192 7224 17192 7224 0 _113_
rlabel metal2 12040 6104 12040 6104 0 _114_
rlabel metal2 17752 5712 17752 5712 0 _115_
rlabel metal2 15568 3640 15568 3640 0 _116_
rlabel metal2 15288 4368 15288 4368 0 _117_
rlabel metal2 8904 6328 8904 6328 0 _118_
rlabel metal2 8176 4312 8176 4312 0 _119_
rlabel metal2 17976 22568 17976 22568 0 _120_
rlabel metal2 16632 6664 16632 6664 0 _121_
rlabel metal3 3108 8120 3108 8120 0 _122_
rlabel metal2 11592 8344 11592 8344 0 _123_
rlabel metal2 10920 6944 10920 6944 0 _124_
rlabel metal2 11480 9520 11480 9520 0 _125_
rlabel metal3 6216 12936 6216 12936 0 _126_
rlabel metal2 7112 13048 7112 13048 0 _127_
rlabel metal2 11368 10136 11368 10136 0 _128_
rlabel metal2 10136 9800 10136 9800 0 _129_
rlabel metal2 16632 4984 16632 4984 0 _130_
rlabel metal2 16072 4648 16072 4648 0 _131_
rlabel metal2 8232 7392 8232 7392 0 _132_
rlabel metal2 2856 5488 2856 5488 0 _133_
rlabel metal2 2744 5152 2744 5152 0 _134_
rlabel metal2 6776 4032 6776 4032 0 _135_
rlabel metal2 7672 8904 7672 8904 0 _136_
rlabel metal2 8008 6440 8008 6440 0 _137_
rlabel metal2 6496 4536 6496 4536 0 _138_
rlabel metal2 4872 5488 4872 5488 0 _139_
rlabel metal3 6608 6104 6608 6104 0 _140_
rlabel metal2 9800 7672 9800 7672 0 _141_
rlabel metal3 7056 12264 7056 12264 0 _142_
rlabel metal2 10024 9520 10024 9520 0 _143_
rlabel metal2 10360 9632 10360 9632 0 _144_
rlabel metal2 8008 12152 8008 12152 0 _145_
rlabel metal2 3080 6776 3080 6776 0 _146_
rlabel metal2 8232 6160 8232 6160 0 _147_
rlabel metal2 10808 5264 10808 5264 0 _148_
rlabel metal2 8288 11256 8288 11256 0 _149_
rlabel metal3 8792 11256 8792 11256 0 _150_
rlabel metal2 5768 4256 5768 4256 0 _151_
rlabel metal2 6216 6272 6216 6272 0 _152_
rlabel metal2 6664 6608 6664 6608 0 _153_
rlabel metal2 8120 7840 8120 7840 0 _154_
rlabel metal3 8400 6104 8400 6104 0 _155_
rlabel metal2 9240 8960 9240 8960 0 _156_
rlabel metal2 3304 10920 3304 10920 0 _157_
rlabel metal2 9968 11480 9968 11480 0 _158_
rlabel metal3 10024 11592 10024 11592 0 _159_
rlabel metal2 3976 5880 3976 5880 0 _160_
rlabel metal2 10472 10752 10472 10752 0 _161_
rlabel metal2 8232 10528 8232 10528 0 _162_
rlabel metal2 9912 8288 9912 8288 0 _163_
rlabel metal3 6216 7224 6216 7224 0 _164_
rlabel metal2 5600 7448 5600 7448 0 _165_
rlabel metal2 9688 8792 9688 8792 0 _166_
rlabel metal2 9576 12012 9576 12012 0 _167_
rlabel metal2 10360 10920 10360 10920 0 _168_
rlabel metal2 8680 10136 8680 10136 0 _169_
rlabel metal2 8568 10920 8568 10920 0 _170_
rlabel metal2 9072 10696 9072 10696 0 _171_
rlabel metal2 8680 6496 8680 6496 0 _172_
rlabel metal3 4536 6664 4536 6664 0 _173_
rlabel metal3 4144 12152 4144 12152 0 _174_
rlabel metal2 5768 6832 5768 6832 0 _175_
rlabel metal3 3108 9128 3108 9128 0 _176_
rlabel metal2 5152 7672 5152 7672 0 _177_
rlabel metal3 8456 4536 8456 4536 0 _178_
rlabel metal3 7560 9016 7560 9016 0 _179_
rlabel metal3 5208 9016 5208 9016 0 _180_
rlabel metal3 6048 8904 6048 8904 0 _181_
rlabel metal2 2968 9520 2968 9520 0 _182_
rlabel metal3 5432 8232 5432 8232 0 _183_
rlabel metal2 6776 7728 6776 7728 0 _184_
rlabel metal2 2184 7448 2184 7448 0 _185_
rlabel metal2 4536 7616 4536 7616 0 _186_
rlabel metal2 5208 8512 5208 8512 0 _187_
rlabel metal2 2912 7448 2912 7448 0 _188_
rlabel metal2 3080 10080 3080 10080 0 _189_
rlabel metal2 2296 10304 2296 10304 0 _190_
rlabel metal2 2520 10976 2520 10976 0 _191_
rlabel metal2 5320 12544 5320 12544 0 _192_
rlabel metal2 2744 8372 2744 8372 0 _193_
rlabel metal2 3752 6832 3752 6832 0 _194_
rlabel metal2 3416 9800 3416 9800 0 _195_
rlabel metal2 3696 10808 3696 10808 0 _196_
rlabel metal2 2968 7952 2968 7952 0 _197_
rlabel metal2 2184 9912 2184 9912 0 _198_
rlabel metal2 5880 12432 5880 12432 0 _199_
rlabel metal2 4536 12208 4536 12208 0 _200_
rlabel metal2 3864 12544 3864 12544 0 _201_
rlabel metal2 7224 9184 7224 9184 0 _202_
rlabel metal2 3640 13048 3640 13048 0 _203_
rlabel metal2 6328 10640 6328 10640 0 _204_
rlabel metal2 3920 11368 3920 11368 0 _205_
rlabel metal2 4760 10920 4760 10920 0 _206_
rlabel metal2 4312 12348 4312 12348 0 _207_
rlabel metal2 6552 13440 6552 13440 0 _208_
rlabel metal3 6664 11256 6664 11256 0 _209_
rlabel metal2 6328 12824 6328 12824 0 _210_
rlabel metal3 26936 9184 26936 9184 0 _211_
rlabel metal2 23632 13944 23632 13944 0 _212_
rlabel metal2 27160 11760 27160 11760 0 _213_
rlabel metal3 23912 6552 23912 6552 0 _214_
rlabel metal2 29624 7056 29624 7056 0 _215_
rlabel metal2 23072 5992 23072 5992 0 _216_
rlabel metal2 30184 9016 30184 9016 0 _217_
rlabel metal2 31864 9072 31864 9072 0 _218_
rlabel metal3 29344 8904 29344 8904 0 _219_
rlabel metal2 27384 7000 27384 7000 0 _220_
rlabel metal2 27496 7952 27496 7952 0 _221_
rlabel metal2 28168 8008 28168 8008 0 _222_
rlabel metal2 30856 14784 30856 14784 0 _223_
rlabel metal3 29176 15848 29176 15848 0 _224_
rlabel metal2 25928 16912 25928 16912 0 _225_
rlabel metal2 28000 14728 28000 14728 0 _226_
rlabel metal2 24136 6944 24136 6944 0 _227_
rlabel metal2 23800 6328 23800 6328 0 _228_
rlabel metal2 28616 14560 28616 14560 0 _229_
rlabel metal2 27048 13832 27048 13832 0 _230_
rlabel metal2 25816 12544 25816 12544 0 _231_
rlabel metal2 19656 14224 19656 14224 0 _232_
rlabel metal2 18984 20832 18984 20832 0 _233_
rlabel metal2 23352 7784 23352 7784 0 _234_
rlabel metal2 27496 5432 27496 5432 0 _235_
rlabel metal3 22344 4536 22344 4536 0 _236_
rlabel metal2 21952 5320 21952 5320 0 _237_
rlabel metal2 24696 3752 24696 3752 0 _238_
rlabel metal2 28168 6832 28168 6832 0 _239_
rlabel metal2 27048 5936 27048 5936 0 _240_
rlabel metal2 24192 5656 24192 5656 0 _241_
rlabel metal2 27720 5600 27720 5600 0 _242_
rlabel metal3 27384 5768 27384 5768 0 _243_
rlabel metal2 27328 5320 27328 5320 0 _244_
rlabel metal2 27104 6888 27104 6888 0 _245_
rlabel metal2 29288 6104 29288 6104 0 _246_
rlabel metal2 29288 5096 29288 5096 0 _247_
rlabel via2 30072 6776 30072 6776 0 _248_
rlabel metal2 29848 5936 29848 5936 0 _249_
rlabel metal2 29960 16072 29960 16072 0 _250_
rlabel metal2 29176 10864 29176 10864 0 _251_
rlabel metal2 30968 5208 30968 5208 0 _252_
rlabel metal3 31248 5768 31248 5768 0 _253_
rlabel metal2 30744 6944 30744 6944 0 _254_
rlabel metal2 30632 7952 30632 7952 0 _255_
rlabel metal2 32088 7448 32088 7448 0 _256_
rlabel metal2 33376 7448 33376 7448 0 _257_
rlabel metal2 31024 8008 31024 8008 0 _258_
rlabel metal2 29288 10080 29288 10080 0 _259_
rlabel metal2 31528 12880 31528 12880 0 _260_
rlabel metal2 31752 11536 31752 11536 0 _261_
rlabel metal2 31864 11144 31864 11144 0 _262_
rlabel metal3 32368 13496 32368 13496 0 _263_
rlabel metal2 33208 14448 33208 14448 0 _264_
rlabel metal2 33152 15512 33152 15512 0 _265_
rlabel metal2 30520 15120 30520 15120 0 _266_
rlabel metal2 29512 15456 29512 15456 0 _267_
rlabel metal2 32424 15680 32424 15680 0 _268_
rlabel metal2 29176 13832 29176 13832 0 _269_
rlabel metal2 29288 14952 29288 14952 0 _270_
rlabel metal2 26040 11424 26040 11424 0 _271_
rlabel metal3 26880 13608 26880 13608 0 _272_
rlabel metal2 27944 16240 27944 16240 0 _273_
rlabel metal2 28504 17920 28504 17920 0 _274_
rlabel metal3 27496 16184 27496 16184 0 _275_
rlabel metal2 29288 16520 29288 16520 0 _276_
rlabel metal2 27440 15512 27440 15512 0 _277_
rlabel metal2 26488 15400 26488 15400 0 _278_
rlabel metal2 23688 18368 23688 18368 0 _279_
rlabel metal3 17640 21784 17640 21784 0 _280_
rlabel metal2 18424 16968 18424 16968 0 _281_
rlabel metal3 19600 13720 19600 13720 0 _282_
rlabel metal2 22792 15540 22792 15540 0 _283_
rlabel metal3 19600 12376 19600 12376 0 _284_
rlabel metal2 22232 15540 22232 15540 0 _285_
rlabel metal3 23520 15960 23520 15960 0 _286_
rlabel metal2 15848 21336 15848 21336 0 _287_
rlabel metal2 15624 24192 15624 24192 0 _288_
rlabel metal2 11816 23464 11816 23464 0 _289_
rlabel metal2 13440 23912 13440 23912 0 _290_
rlabel metal2 13832 23688 13832 23688 0 _291_
rlabel metal2 12712 22064 12712 22064 0 _292_
rlabel metal2 14392 20720 14392 20720 0 _293_
rlabel metal3 17304 19992 17304 19992 0 _294_
rlabel metal2 16632 19936 16632 19936 0 _295_
rlabel metal2 17976 20552 17976 20552 0 _296_
rlabel metal2 18536 19824 18536 19824 0 _297_
rlabel metal2 16520 21504 16520 21504 0 _298_
rlabel metal2 20664 27496 20664 27496 0 _299_
rlabel metal2 18648 16016 18648 16016 0 _300_
rlabel metal3 11088 23352 11088 23352 0 _301_
rlabel metal2 12376 21616 12376 21616 0 _302_
rlabel metal3 6496 18312 6496 18312 0 _303_
rlabel metal2 11480 18648 11480 18648 0 _304_
rlabel metal2 7392 17080 7392 17080 0 _305_
rlabel metal2 10472 17248 10472 17248 0 _306_
rlabel metal2 8232 18704 8232 18704 0 _307_
rlabel metal2 11368 18480 11368 18480 0 _308_
rlabel metal2 10808 19376 10808 19376 0 _309_
rlabel metal3 7112 19880 7112 19880 0 _310_
rlabel metal2 8680 19488 8680 19488 0 _311_
rlabel metal2 9464 18536 9464 18536 0 _312_
rlabel metal2 12208 20216 12208 20216 0 _313_
rlabel metal3 12264 24584 12264 24584 0 _314_
rlabel metal2 18704 23240 18704 23240 0 _315_
rlabel metal2 18256 24808 18256 24808 0 _316_
rlabel metal3 13160 25592 13160 25592 0 _317_
rlabel metal2 14224 23352 14224 23352 0 _318_
rlabel metal2 9912 17920 9912 17920 0 _319_
rlabel metal3 8456 18536 8456 18536 0 _320_
rlabel metal2 7336 18480 7336 18480 0 _321_
rlabel metal2 8680 18536 8680 18536 0 _322_
rlabel metal3 9520 18200 9520 18200 0 _323_
rlabel metal2 10696 18816 10696 18816 0 _324_
rlabel metal2 11480 21280 11480 21280 0 _325_
rlabel metal2 12040 24136 12040 24136 0 _326_
rlabel metal2 11536 24696 11536 24696 0 _327_
rlabel metal2 15400 23576 15400 23576 0 _328_
rlabel metal2 10024 25536 10024 25536 0 _329_
rlabel metal2 11704 19208 11704 19208 0 _330_
rlabel metal2 8120 18200 8120 18200 0 _331_
rlabel metal2 12600 19432 12600 19432 0 _332_
rlabel metal2 12040 20944 12040 20944 0 _333_
rlabel metal2 10248 23184 10248 23184 0 _334_
rlabel metal2 11032 23408 11032 23408 0 _335_
rlabel metal2 9016 24304 9016 24304 0 _336_
rlabel metal2 10248 20384 10248 20384 0 _337_
rlabel metal2 12600 21056 12600 21056 0 _338_
rlabel metal2 15512 21280 15512 21280 0 _339_
rlabel metal2 15176 22456 15176 22456 0 _340_
rlabel metal2 12488 22288 12488 22288 0 _341_
rlabel metal2 13048 21784 13048 21784 0 _342_
rlabel metal3 10808 23016 10808 23016 0 _343_
rlabel metal2 9912 18368 9912 18368 0 _344_
rlabel metal2 12656 18648 12656 18648 0 _345_
rlabel metal2 10472 18200 10472 18200 0 _346_
rlabel metal3 12824 19320 12824 19320 0 _347_
rlabel metal2 13832 20832 13832 20832 0 _348_
rlabel metal3 14168 21672 14168 21672 0 _349_
rlabel metal2 13720 22008 13720 22008 0 _350_
rlabel metal2 10472 20272 10472 20272 0 _351_
rlabel metal2 8008 19600 8008 19600 0 _352_
rlabel metal2 9240 19264 9240 19264 0 _353_
rlabel metal3 9800 19320 9800 19320 0 _354_
rlabel metal2 10248 19656 10248 19656 0 _355_
rlabel metal2 15176 25200 15176 25200 0 _356_
rlabel metal2 16184 25536 16184 25536 0 _357_
rlabel metal2 15960 25480 15960 25480 0 _358_
rlabel metal2 12600 25816 12600 25816 0 _359_
rlabel metal2 12600 19712 12600 19712 0 _360_
rlabel metal2 11032 21280 11032 21280 0 _361_
rlabel metal2 14280 25592 14280 25592 0 _362_
rlabel metal3 15624 25368 15624 25368 0 _363_
rlabel metal3 19488 26936 19488 26936 0 _364_
rlabel metal2 23016 18368 23016 18368 0 _365_
rlabel metal2 18536 26432 18536 26432 0 _366_
rlabel metal2 21784 21728 21784 21728 0 _367_
rlabel metal2 19432 23184 19432 23184 0 _368_
rlabel metal2 19432 20664 19432 20664 0 _369_
rlabel metal2 18872 23576 18872 23576 0 _370_
rlabel metal2 21896 19656 21896 19656 0 _371_
rlabel metal3 21504 21560 21504 21560 0 _372_
rlabel metal2 20776 21840 20776 21840 0 _373_
rlabel metal2 25256 22624 25256 22624 0 _374_
rlabel metal2 26544 23128 26544 23128 0 _375_
rlabel metal2 16912 20104 16912 20104 0 _376_
rlabel metal2 25480 22456 25480 22456 0 _377_
rlabel metal3 25312 23128 25312 23128 0 _378_
rlabel metal2 26936 22568 26936 22568 0 _379_
rlabel metal2 26264 24192 26264 24192 0 _380_
rlabel metal2 27048 22288 27048 22288 0 _381_
rlabel metal2 25704 25592 25704 25592 0 _382_
rlabel metal2 27832 21448 27832 21448 0 _383_
rlabel metal2 28168 20608 28168 20608 0 _384_
rlabel metal2 26264 21728 26264 21728 0 _385_
rlabel metal2 27608 21056 27608 21056 0 _386_
rlabel metal2 24024 19264 24024 19264 0 _387_
rlabel metal2 19264 27832 19264 27832 0 _388_
rlabel metal2 20104 27356 20104 27356 0 _389_
rlabel metal2 16184 17584 16184 17584 0 _390_
rlabel metal2 15624 15960 15624 15960 0 _391_
rlabel metal2 16632 16464 16632 16464 0 _392_
rlabel metal2 15848 17360 15848 17360 0 _393_
rlabel metal2 17416 17976 17416 17976 0 _394_
rlabel metal2 16520 17976 16520 17976 0 _395_
rlabel metal2 15960 13888 15960 13888 0 _396_
rlabel metal2 15512 15568 15512 15568 0 _397_
rlabel metal2 13944 16744 13944 16744 0 _398_
rlabel metal2 12264 16800 12264 16800 0 _399_
rlabel metal2 15512 15960 15512 15960 0 _400_
rlabel metal3 15624 15960 15624 15960 0 _401_
rlabel metal3 14448 15960 14448 15960 0 _402_
rlabel metal3 13272 16184 13272 16184 0 _403_
rlabel metal2 19096 16352 19096 16352 0 _404_
rlabel metal3 17752 15960 17752 15960 0 _405_
rlabel metal2 17416 16296 17416 16296 0 _406_
rlabel metal2 18200 17136 18200 17136 0 _407_
rlabel metal2 22792 12208 22792 12208 0 _408_
rlabel metal3 22288 12824 22288 12824 0 _409_
rlabel metal2 21448 15540 21448 15540 0 _410_
rlabel metal2 19656 10304 19656 10304 0 _411_
rlabel metal2 21448 12208 21448 12208 0 _412_
rlabel metal2 18816 4424 18816 4424 0 _413_
rlabel metal3 2688 20552 2688 20552 0 _414_
rlabel metal3 10640 23128 10640 23128 0 _415_
rlabel metal2 2632 23240 2632 23240 0 _416_
rlabel metal2 4536 20272 4536 20272 0 _417_
rlabel metal2 5544 20048 5544 20048 0 _418_
rlabel metal2 5544 23464 5544 23464 0 _419_
rlabel metal2 3640 22064 3640 22064 0 _420_
rlabel metal2 5096 24752 5096 24752 0 _421_
rlabel metal2 6216 23184 6216 23184 0 _422_
rlabel metal3 6384 27048 6384 27048 0 _423_
rlabel metal3 5544 27272 5544 27272 0 _424_
rlabel metal2 3864 25368 3864 25368 0 _425_
rlabel metal2 4704 27832 4704 27832 0 _426_
rlabel metal2 2968 26712 2968 26712 0 _427_
rlabel metal2 27104 10584 27104 10584 0 clknet_0_wb_clk_i
rlabel metal2 3304 15456 3304 15456 0 clknet_3_0__leaf_wb_clk_i
rlabel metal3 12376 15288 12376 15288 0 clknet_3_1__leaf_wb_clk_i
rlabel metal2 2072 22736 2072 22736 0 clknet_3_2__leaf_wb_clk_i
rlabel metal3 15904 27048 15904 27048 0 clknet_3_3__leaf_wb_clk_i
rlabel metal2 18480 10584 18480 10584 0 clknet_3_4__leaf_wb_clk_i
rlabel metal2 27104 5096 27104 5096 0 clknet_3_5__leaf_wb_clk_i
rlabel metal2 26040 22400 26040 22400 0 clknet_3_6__leaf_wb_clk_i
rlabel metal2 29848 23912 29848 23912 0 clknet_3_7__leaf_wb_clk_i
rlabel metal2 23128 23968 23128 23968 0 clock_div\[0\]
rlabel metal2 24136 20720 24136 20720 0 clock_div\[1\]
rlabel metal2 24248 22064 24248 22064 0 clock_div\[2\]
rlabel metal2 26992 23016 26992 23016 0 clock_div\[3\]
rlabel metal2 26376 24640 26376 24640 0 clock_div\[4\]
rlabel metal2 24584 25144 24584 25144 0 clock_div\[5\]
rlabel metal2 27496 22176 27496 22176 0 clock_div\[6\]
rlabel metal2 25928 21168 25928 21168 0 clock_div\[7\]
rlabel metal3 20888 25480 20888 25480 0 clock_div\[8\]
rlabel metal2 22344 8400 22344 8400 0 counter\[0\]
rlabel metal3 30016 8120 30016 8120 0 counter\[10\]
rlabel metal3 30184 8344 30184 8344 0 counter\[11\]
rlabel metal2 30408 9856 30408 9856 0 counter\[12\]
rlabel metal2 31248 9016 31248 9016 0 counter\[13\]
rlabel metal2 31024 14392 31024 14392 0 counter\[14\]
rlabel metal2 31248 14616 31248 14616 0 counter\[15\]
rlabel metal2 31752 15960 31752 15960 0 counter\[16\]
rlabel metal3 30408 15400 30408 15400 0 counter\[17\]
rlabel metal2 27552 12936 27552 12936 0 counter\[18\]
rlabel metal2 27384 13048 27384 13048 0 counter\[19\]
rlabel metal3 22400 7448 22400 7448 0 counter\[1\]
rlabel metal2 27944 17808 27944 17808 0 counter\[20\]
rlabel metal2 29176 17696 29176 17696 0 counter\[21\]
rlabel metal3 27720 16744 27720 16744 0 counter\[22\]
rlabel metal2 22456 3864 22456 3864 0 counter\[3\]
rlabel metal2 25928 8288 25928 8288 0 counter\[4\]
rlabel metal2 25368 5656 25368 5656 0 counter\[5\]
rlabel metal2 28280 7784 28280 7784 0 counter\[6\]
rlabel metal3 28448 7448 28448 7448 0 counter\[7\]
rlabel metal2 30968 6048 30968 6048 0 counter\[8\]
rlabel metal2 31192 5656 31192 5656 0 counter\[9\]
rlabel metal2 17976 1582 17976 1582 0 io_out[0]
rlabel metal2 25144 2086 25144 2086 0 io_out[1]
rlabel metal2 32312 2086 32312 2086 0 io_out[2]
rlabel metal3 22120 16072 22120 16072 0 just_inc
rlabel metal2 15064 24360 15064 24360 0 just_rst
rlabel metal2 4536 21280 4536 21280 0 master_clk_div\[0\]
rlabel metal3 6104 20664 6104 20664 0 master_clk_div\[1\]
rlabel metal3 4312 21672 4312 21672 0 master_clk_div\[2\]
rlabel metal2 5320 22960 5320 22960 0 master_clk_div\[3\]
rlabel metal3 6048 26936 6048 26936 0 master_clk_div\[4\]
rlabel metal2 5040 27160 5040 27160 0 master_clk_div\[5\]
rlabel metal2 4312 27356 4312 27356 0 master_clk_div\[6\]
rlabel metal2 11200 5096 11200 5096 0 net1
rlabel metal3 17584 5096 17584 5096 0 net2
rlabel metal2 22792 6272 22792 6272 0 net3
rlabel metal2 32200 3472 32200 3472 0 net4
rlabel metal2 23352 4144 23352 4144 0 net5
rlabel metal3 21616 25704 21616 25704 0 prev_clk_div
rlabel metal2 16856 16576 16856 16576 0 rhythm_LFSR\[0\]
rlabel metal3 17304 16968 17304 16968 0 rhythm_LFSR\[1\]
rlabel metal2 17920 14728 17920 14728 0 rhythm_LFSR\[2\]
rlabel metal2 17640 16856 17640 16856 0 rhythm_LFSR\[3\]
rlabel metal2 11032 4256 11032 4256 0 rst_n
rlabel metal2 21560 12768 21560 12768 0 tempo_LFSR\[0\]
rlabel metal3 22512 13496 22512 13496 0 tempo_LFSR\[1\]
rlabel metal2 22232 14056 22232 14056 0 tempo_LFSR\[2\]
rlabel metal2 20552 11760 20552 11760 0 tempo_LFSR\[3\]
rlabel metal2 15736 15904 15736 15904 0 tune_ROM\[0\]
rlabel metal2 15848 12600 15848 12600 0 tune_ROM\[1\]
rlabel metal2 6216 17192 6216 17192 0 tune_ROM\[2\]
rlabel metal3 6048 18424 6048 18424 0 tune_ROM\[3\]
rlabel metal3 6048 16856 6048 16856 0 tune_ROM\[4\]
rlabel metal2 8904 16016 8904 16016 0 tune_ROM\[5\]
rlabel metal2 1624 9688 1624 9688 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 36000 36000
<< end >>
