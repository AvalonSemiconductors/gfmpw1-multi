VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO multiplexer
  CLASS BLOCK ;
  FOREIGN multiplexer ;
  ORIGIN 0.000 0.000 ;
  SIZE 750.000 BY 700.000 ;
  PIN ay8913_do[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 196.000 696.000 196.560 700.000 ;
    END
  END ay8913_do[0]
  PIN ay8913_do[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 229.600 696.000 230.160 700.000 ;
    END
  END ay8913_do[10]
  PIN ay8913_do[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 232.960 696.000 233.520 700.000 ;
    END
  END ay8913_do[11]
  PIN ay8913_do[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 236.320 696.000 236.880 700.000 ;
    END
  END ay8913_do[12]
  PIN ay8913_do[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 239.680 696.000 240.240 700.000 ;
    END
  END ay8913_do[13]
  PIN ay8913_do[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 243.040 696.000 243.600 700.000 ;
    END
  END ay8913_do[14]
  PIN ay8913_do[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 246.400 696.000 246.960 700.000 ;
    END
  END ay8913_do[15]
  PIN ay8913_do[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 249.760 696.000 250.320 700.000 ;
    END
  END ay8913_do[16]
  PIN ay8913_do[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 253.120 696.000 253.680 700.000 ;
    END
  END ay8913_do[17]
  PIN ay8913_do[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 256.480 696.000 257.040 700.000 ;
    END
  END ay8913_do[18]
  PIN ay8913_do[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 259.840 696.000 260.400 700.000 ;
    END
  END ay8913_do[19]
  PIN ay8913_do[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 199.360 696.000 199.920 700.000 ;
    END
  END ay8913_do[1]
  PIN ay8913_do[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 263.200 696.000 263.760 700.000 ;
    END
  END ay8913_do[20]
  PIN ay8913_do[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 266.560 696.000 267.120 700.000 ;
    END
  END ay8913_do[21]
  PIN ay8913_do[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 269.920 696.000 270.480 700.000 ;
    END
  END ay8913_do[22]
  PIN ay8913_do[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 273.280 696.000 273.840 700.000 ;
    END
  END ay8913_do[23]
  PIN ay8913_do[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 276.640 696.000 277.200 700.000 ;
    END
  END ay8913_do[24]
  PIN ay8913_do[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 280.000 696.000 280.560 700.000 ;
    END
  END ay8913_do[25]
  PIN ay8913_do[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 283.360 696.000 283.920 700.000 ;
    END
  END ay8913_do[26]
  PIN ay8913_do[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 286.720 696.000 287.280 700.000 ;
    END
  END ay8913_do[27]
  PIN ay8913_do[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 202.720 696.000 203.280 700.000 ;
    END
  END ay8913_do[2]
  PIN ay8913_do[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 206.080 696.000 206.640 700.000 ;
    END
  END ay8913_do[3]
  PIN ay8913_do[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 209.440 696.000 210.000 700.000 ;
    END
  END ay8913_do[4]
  PIN ay8913_do[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 212.800 696.000 213.360 700.000 ;
    END
  END ay8913_do[5]
  PIN ay8913_do[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 216.160 696.000 216.720 700.000 ;
    END
  END ay8913_do[6]
  PIN ay8913_do[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 219.520 696.000 220.080 700.000 ;
    END
  END ay8913_do[7]
  PIN ay8913_do[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 222.880 696.000 223.440 700.000 ;
    END
  END ay8913_do[8]
  PIN ay8913_do[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 226.240 696.000 226.800 700.000 ;
    END
  END ay8913_do[9]
  PIN blinker_do[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 631.680 4.000 632.240 ;
    END
  END blinker_do[0]
  PIN blinker_do[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 637.280 4.000 637.840 ;
    END
  END blinker_do[1]
  PIN blinker_do[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 642.880 4.000 643.440 ;
    END
  END blinker_do[2]
  PIN custom_settings[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 190.400 750.000 190.960 ;
    END
  END custom_settings[0]
  PIN custom_settings[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 235.200 750.000 235.760 ;
    END
  END custom_settings[10]
  PIN custom_settings[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 239.680 750.000 240.240 ;
    END
  END custom_settings[11]
  PIN custom_settings[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 244.160 750.000 244.720 ;
    END
  END custom_settings[12]
  PIN custom_settings[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 248.640 750.000 249.200 ;
    END
  END custom_settings[13]
  PIN custom_settings[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 253.120 750.000 253.680 ;
    END
  END custom_settings[14]
  PIN custom_settings[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 257.600 750.000 258.160 ;
    END
  END custom_settings[15]
  PIN custom_settings[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 262.080 750.000 262.640 ;
    END
  END custom_settings[16]
  PIN custom_settings[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 266.560 750.000 267.120 ;
    END
  END custom_settings[17]
  PIN custom_settings[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 271.040 750.000 271.600 ;
    END
  END custom_settings[18]
  PIN custom_settings[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 275.520 750.000 276.080 ;
    END
  END custom_settings[19]
  PIN custom_settings[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 194.880 750.000 195.440 ;
    END
  END custom_settings[1]
  PIN custom_settings[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 280.000 750.000 280.560 ;
    END
  END custom_settings[20]
  PIN custom_settings[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 284.480 750.000 285.040 ;
    END
  END custom_settings[21]
  PIN custom_settings[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 288.960 750.000 289.520 ;
    END
  END custom_settings[22]
  PIN custom_settings[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 293.440 750.000 294.000 ;
    END
  END custom_settings[23]
  PIN custom_settings[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 297.920 750.000 298.480 ;
    END
  END custom_settings[24]
  PIN custom_settings[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 302.400 750.000 302.960 ;
    END
  END custom_settings[25]
  PIN custom_settings[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 306.880 750.000 307.440 ;
    END
  END custom_settings[26]
  PIN custom_settings[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 311.360 750.000 311.920 ;
    END
  END custom_settings[27]
  PIN custom_settings[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 315.840 750.000 316.400 ;
    END
  END custom_settings[28]
  PIN custom_settings[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 320.320 750.000 320.880 ;
    END
  END custom_settings[29]
  PIN custom_settings[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 199.360 750.000 199.920 ;
    END
  END custom_settings[2]
  PIN custom_settings[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 324.800 750.000 325.360 ;
    END
  END custom_settings[30]
  PIN custom_settings[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 329.280 750.000 329.840 ;
    END
  END custom_settings[31]
  PIN custom_settings[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 203.840 750.000 204.400 ;
    END
  END custom_settings[3]
  PIN custom_settings[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 208.320 750.000 208.880 ;
    END
  END custom_settings[4]
  PIN custom_settings[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 212.800 750.000 213.360 ;
    END
  END custom_settings[5]
  PIN custom_settings[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 217.280 750.000 217.840 ;
    END
  END custom_settings[6]
  PIN custom_settings[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 221.760 750.000 222.320 ;
    END
  END custom_settings[7]
  PIN custom_settings[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 226.240 750.000 226.800 ;
    END
  END custom_settings[8]
  PIN custom_settings[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 230.720 750.000 231.280 ;
    END
  END custom_settings[9]
  PIN diceroll_do[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 629.440 696.000 630.000 700.000 ;
    END
  END diceroll_do[0]
  PIN diceroll_do[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 632.800 696.000 633.360 700.000 ;
    END
  END diceroll_do[1]
  PIN diceroll_do[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 636.160 696.000 636.720 700.000 ;
    END
  END diceroll_do[2]
  PIN diceroll_do[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 639.520 696.000 640.080 700.000 ;
    END
  END diceroll_do[3]
  PIN diceroll_do[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 642.880 696.000 643.440 700.000 ;
    END
  END diceroll_do[4]
  PIN diceroll_do[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 646.240 696.000 646.800 700.000 ;
    END
  END diceroll_do[5]
  PIN diceroll_do[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 649.600 696.000 650.160 700.000 ;
    END
  END diceroll_do[6]
  PIN diceroll_do[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 652.960 696.000 653.520 700.000 ;
    END
  END diceroll_do[7]
  PIN diceroll_do[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 656.320 696.000 656.880 700.000 ;
    END
  END diceroll_do[8]
  PIN hellorld_do
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 586.880 4.000 587.440 ;
    END
  END hellorld_do
  PIN io_in_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 51.520 696.000 52.080 700.000 ;
    END
  END io_in_0
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 54.880 4.000 55.440 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 110.880 4.000 111.440 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 116.480 4.000 117.040 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 122.080 4.000 122.640 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 127.680 4.000 128.240 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 133.280 4.000 133.840 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 138.880 4.000 139.440 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 144.480 4.000 145.040 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 150.080 4.000 150.640 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 155.680 4.000 156.240 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 161.280 4.000 161.840 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 60.480 4.000 61.040 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 166.880 4.000 167.440 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 172.480 4.000 173.040 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 178.080 4.000 178.640 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 183.680 4.000 184.240 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 189.280 4.000 189.840 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 194.880 4.000 195.440 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 200.480 4.000 201.040 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 206.080 4.000 206.640 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 211.680 4.000 212.240 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 217.280 4.000 217.840 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 66.080 4.000 66.640 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 222.880 4.000 223.440 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 228.480 4.000 229.040 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 234.080 4.000 234.640 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 239.680 4.000 240.240 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 245.280 4.000 245.840 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 250.880 4.000 251.440 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 256.480 4.000 257.040 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 262.080 4.000 262.640 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 71.680 4.000 72.240 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 77.280 4.000 77.840 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 82.880 4.000 83.440 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 88.480 4.000 89.040 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 94.080 4.000 94.640 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 99.680 4.000 100.240 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 105.280 4.000 105.840 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 54.880 696.000 55.440 700.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 88.480 696.000 89.040 700.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 91.840 696.000 92.400 700.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 696.000 95.760 700.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 98.560 696.000 99.120 700.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 101.920 696.000 102.480 700.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 105.280 696.000 105.840 700.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 108.640 696.000 109.200 700.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 112.000 696.000 112.560 700.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 115.360 696.000 115.920 700.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 118.720 696.000 119.280 700.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.240 696.000 58.800 700.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 122.080 696.000 122.640 700.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 125.440 696.000 126.000 700.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 128.800 696.000 129.360 700.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 132.160 696.000 132.720 700.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 135.520 696.000 136.080 700.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 138.880 696.000 139.440 700.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 142.240 696.000 142.800 700.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 145.600 696.000 146.160 700.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 148.960 696.000 149.520 700.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 152.320 696.000 152.880 700.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 61.600 696.000 62.160 700.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 155.680 696.000 156.240 700.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 159.040 696.000 159.600 700.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 162.400 696.000 162.960 700.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 165.760 696.000 166.320 700.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 169.120 696.000 169.680 700.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 172.480 696.000 173.040 700.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 175.840 696.000 176.400 700.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 179.200 696.000 179.760 700.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 64.960 696.000 65.520 700.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.320 696.000 68.880 700.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 71.680 696.000 72.240 700.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 75.040 696.000 75.600 700.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 78.400 696.000 78.960 700.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 81.760 696.000 82.320 700.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 85.120 696.000 85.680 700.000 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 182.560 696.000 183.120 700.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 185.920 696.000 186.480 700.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 189.280 696.000 189.840 700.000 ;
    END
  END irq[2]
  PIN mc14500_do[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 407.680 4.000 408.240 ;
    END
  END mc14500_do[0]
  PIN mc14500_do[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 463.680 4.000 464.240 ;
    END
  END mc14500_do[10]
  PIN mc14500_do[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 469.280 4.000 469.840 ;
    END
  END mc14500_do[11]
  PIN mc14500_do[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 474.880 4.000 475.440 ;
    END
  END mc14500_do[12]
  PIN mc14500_do[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 480.480 4.000 481.040 ;
    END
  END mc14500_do[13]
  PIN mc14500_do[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 486.080 4.000 486.640 ;
    END
  END mc14500_do[14]
  PIN mc14500_do[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 491.680 4.000 492.240 ;
    END
  END mc14500_do[15]
  PIN mc14500_do[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 497.280 4.000 497.840 ;
    END
  END mc14500_do[16]
  PIN mc14500_do[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 502.880 4.000 503.440 ;
    END
  END mc14500_do[17]
  PIN mc14500_do[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 508.480 4.000 509.040 ;
    END
  END mc14500_do[18]
  PIN mc14500_do[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 514.080 4.000 514.640 ;
    END
  END mc14500_do[19]
  PIN mc14500_do[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 413.280 4.000 413.840 ;
    END
  END mc14500_do[1]
  PIN mc14500_do[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 519.680 4.000 520.240 ;
    END
  END mc14500_do[20]
  PIN mc14500_do[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 525.280 4.000 525.840 ;
    END
  END mc14500_do[21]
  PIN mc14500_do[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 530.880 4.000 531.440 ;
    END
  END mc14500_do[22]
  PIN mc14500_do[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 536.480 4.000 537.040 ;
    END
  END mc14500_do[23]
  PIN mc14500_do[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 542.080 4.000 542.640 ;
    END
  END mc14500_do[24]
  PIN mc14500_do[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 547.680 4.000 548.240 ;
    END
  END mc14500_do[25]
  PIN mc14500_do[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 553.280 4.000 553.840 ;
    END
  END mc14500_do[26]
  PIN mc14500_do[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 558.880 4.000 559.440 ;
    END
  END mc14500_do[27]
  PIN mc14500_do[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 564.480 4.000 565.040 ;
    END
  END mc14500_do[28]
  PIN mc14500_do[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 570.080 4.000 570.640 ;
    END
  END mc14500_do[29]
  PIN mc14500_do[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 418.880 4.000 419.440 ;
    END
  END mc14500_do[2]
  PIN mc14500_do[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 575.680 4.000 576.240 ;
    END
  END mc14500_do[30]
  PIN mc14500_do[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 424.480 4.000 425.040 ;
    END
  END mc14500_do[3]
  PIN mc14500_do[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 430.080 4.000 430.640 ;
    END
  END mc14500_do[4]
  PIN mc14500_do[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 435.680 4.000 436.240 ;
    END
  END mc14500_do[5]
  PIN mc14500_do[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 441.280 4.000 441.840 ;
    END
  END mc14500_do[6]
  PIN mc14500_do[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 446.880 4.000 447.440 ;
    END
  END mc14500_do[7]
  PIN mc14500_do[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 452.480 4.000 453.040 ;
    END
  END mc14500_do[8]
  PIN mc14500_do[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 458.080 4.000 458.640 ;
    END
  END mc14500_do[9]
  PIN mc14500_sram_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 660.800 0.000 661.360 4.000 ;
    END
  END mc14500_sram_addr[0]
  PIN mc14500_sram_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 665.280 0.000 665.840 4.000 ;
    END
  END mc14500_sram_addr[1]
  PIN mc14500_sram_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 669.760 0.000 670.320 4.000 ;
    END
  END mc14500_sram_addr[2]
  PIN mc14500_sram_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 674.240 0.000 674.800 4.000 ;
    END
  END mc14500_sram_addr[3]
  PIN mc14500_sram_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 678.720 0.000 679.280 4.000 ;
    END
  END mc14500_sram_addr[4]
  PIN mc14500_sram_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 683.200 0.000 683.760 4.000 ;
    END
  END mc14500_sram_addr[5]
  PIN mc14500_sram_gwe
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 723.520 0.000 724.080 4.000 ;
    END
  END mc14500_sram_gwe
  PIN mc14500_sram_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 687.680 0.000 688.240 4.000 ;
    END
  END mc14500_sram_in[0]
  PIN mc14500_sram_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 692.160 0.000 692.720 4.000 ;
    END
  END mc14500_sram_in[1]
  PIN mc14500_sram_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 696.640 0.000 697.200 4.000 ;
    END
  END mc14500_sram_in[2]
  PIN mc14500_sram_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 701.120 0.000 701.680 4.000 ;
    END
  END mc14500_sram_in[3]
  PIN mc14500_sram_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 705.600 0.000 706.160 4.000 ;
    END
  END mc14500_sram_in[4]
  PIN mc14500_sram_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 710.080 0.000 710.640 4.000 ;
    END
  END mc14500_sram_in[5]
  PIN mc14500_sram_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 714.560 0.000 715.120 4.000 ;
    END
  END mc14500_sram_in[6]
  PIN mc14500_sram_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 719.040 0.000 719.600 4.000 ;
    END
  END mc14500_sram_in[7]
  PIN pdp11_do[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 290.080 696.000 290.640 700.000 ;
    END
  END pdp11_do[0]
  PIN pdp11_do[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 357.280 696.000 357.840 700.000 ;
    END
  END pdp11_do[10]
  PIN pdp11_do[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 364.000 696.000 364.560 700.000 ;
    END
  END pdp11_do[11]
  PIN pdp11_do[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 370.720 696.000 371.280 700.000 ;
    END
  END pdp11_do[12]
  PIN pdp11_do[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 377.440 696.000 378.000 700.000 ;
    END
  END pdp11_do[13]
  PIN pdp11_do[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 384.160 696.000 384.720 700.000 ;
    END
  END pdp11_do[14]
  PIN pdp11_do[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 390.880 696.000 391.440 700.000 ;
    END
  END pdp11_do[15]
  PIN pdp11_do[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 397.600 696.000 398.160 700.000 ;
    END
  END pdp11_do[16]
  PIN pdp11_do[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 404.320 696.000 404.880 700.000 ;
    END
  END pdp11_do[17]
  PIN pdp11_do[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 411.040 696.000 411.600 700.000 ;
    END
  END pdp11_do[18]
  PIN pdp11_do[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 417.760 696.000 418.320 700.000 ;
    END
  END pdp11_do[19]
  PIN pdp11_do[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 296.800 696.000 297.360 700.000 ;
    END
  END pdp11_do[1]
  PIN pdp11_do[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 424.480 696.000 425.040 700.000 ;
    END
  END pdp11_do[20]
  PIN pdp11_do[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 431.200 696.000 431.760 700.000 ;
    END
  END pdp11_do[21]
  PIN pdp11_do[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 437.920 696.000 438.480 700.000 ;
    END
  END pdp11_do[22]
  PIN pdp11_do[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 444.640 696.000 445.200 700.000 ;
    END
  END pdp11_do[23]
  PIN pdp11_do[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 451.360 696.000 451.920 700.000 ;
    END
  END pdp11_do[24]
  PIN pdp11_do[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 458.080 696.000 458.640 700.000 ;
    END
  END pdp11_do[25]
  PIN pdp11_do[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 464.800 696.000 465.360 700.000 ;
    END
  END pdp11_do[26]
  PIN pdp11_do[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 471.520 696.000 472.080 700.000 ;
    END
  END pdp11_do[27]
  PIN pdp11_do[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 478.240 696.000 478.800 700.000 ;
    END
  END pdp11_do[28]
  PIN pdp11_do[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 484.960 696.000 485.520 700.000 ;
    END
  END pdp11_do[29]
  PIN pdp11_do[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 303.520 696.000 304.080 700.000 ;
    END
  END pdp11_do[2]
  PIN pdp11_do[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 491.680 696.000 492.240 700.000 ;
    END
  END pdp11_do[30]
  PIN pdp11_do[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 498.400 696.000 498.960 700.000 ;
    END
  END pdp11_do[31]
  PIN pdp11_do[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 505.120 696.000 505.680 700.000 ;
    END
  END pdp11_do[32]
  PIN pdp11_do[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 310.240 696.000 310.800 700.000 ;
    END
  END pdp11_do[3]
  PIN pdp11_do[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 316.960 696.000 317.520 700.000 ;
    END
  END pdp11_do[4]
  PIN pdp11_do[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 323.680 696.000 324.240 700.000 ;
    END
  END pdp11_do[5]
  PIN pdp11_do[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 330.400 696.000 330.960 700.000 ;
    END
  END pdp11_do[6]
  PIN pdp11_do[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 337.120 696.000 337.680 700.000 ;
    END
  END pdp11_do[7]
  PIN pdp11_do[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 343.840 696.000 344.400 700.000 ;
    END
  END pdp11_do[8]
  PIN pdp11_do[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 350.560 696.000 351.120 700.000 ;
    END
  END pdp11_do[9]
  PIN pdp11_oeb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 293.440 696.000 294.000 700.000 ;
    END
  END pdp11_oeb[0]
  PIN pdp11_oeb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 360.640 696.000 361.200 700.000 ;
    END
  END pdp11_oeb[10]
  PIN pdp11_oeb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 367.360 696.000 367.920 700.000 ;
    END
  END pdp11_oeb[11]
  PIN pdp11_oeb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 374.080 696.000 374.640 700.000 ;
    END
  END pdp11_oeb[12]
  PIN pdp11_oeb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 380.800 696.000 381.360 700.000 ;
    END
  END pdp11_oeb[13]
  PIN pdp11_oeb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 387.520 696.000 388.080 700.000 ;
    END
  END pdp11_oeb[14]
  PIN pdp11_oeb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 394.240 696.000 394.800 700.000 ;
    END
  END pdp11_oeb[15]
  PIN pdp11_oeb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 400.960 696.000 401.520 700.000 ;
    END
  END pdp11_oeb[16]
  PIN pdp11_oeb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 407.680 696.000 408.240 700.000 ;
    END
  END pdp11_oeb[17]
  PIN pdp11_oeb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 414.400 696.000 414.960 700.000 ;
    END
  END pdp11_oeb[18]
  PIN pdp11_oeb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 421.120 696.000 421.680 700.000 ;
    END
  END pdp11_oeb[19]
  PIN pdp11_oeb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 300.160 696.000 300.720 700.000 ;
    END
  END pdp11_oeb[1]
  PIN pdp11_oeb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 427.840 696.000 428.400 700.000 ;
    END
  END pdp11_oeb[20]
  PIN pdp11_oeb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 434.560 696.000 435.120 700.000 ;
    END
  END pdp11_oeb[21]
  PIN pdp11_oeb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 441.280 696.000 441.840 700.000 ;
    END
  END pdp11_oeb[22]
  PIN pdp11_oeb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 448.000 696.000 448.560 700.000 ;
    END
  END pdp11_oeb[23]
  PIN pdp11_oeb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 454.720 696.000 455.280 700.000 ;
    END
  END pdp11_oeb[24]
  PIN pdp11_oeb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 461.440 696.000 462.000 700.000 ;
    END
  END pdp11_oeb[25]
  PIN pdp11_oeb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 468.160 696.000 468.720 700.000 ;
    END
  END pdp11_oeb[26]
  PIN pdp11_oeb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 474.880 696.000 475.440 700.000 ;
    END
  END pdp11_oeb[27]
  PIN pdp11_oeb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 481.600 696.000 482.160 700.000 ;
    END
  END pdp11_oeb[28]
  PIN pdp11_oeb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 488.320 696.000 488.880 700.000 ;
    END
  END pdp11_oeb[29]
  PIN pdp11_oeb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 306.880 696.000 307.440 700.000 ;
    END
  END pdp11_oeb[2]
  PIN pdp11_oeb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 495.040 696.000 495.600 700.000 ;
    END
  END pdp11_oeb[30]
  PIN pdp11_oeb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 501.760 696.000 502.320 700.000 ;
    END
  END pdp11_oeb[31]
  PIN pdp11_oeb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 508.480 696.000 509.040 700.000 ;
    END
  END pdp11_oeb[32]
  PIN pdp11_oeb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 313.600 696.000 314.160 700.000 ;
    END
  END pdp11_oeb[3]
  PIN pdp11_oeb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 320.320 696.000 320.880 700.000 ;
    END
  END pdp11_oeb[4]
  PIN pdp11_oeb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 327.040 696.000 327.600 700.000 ;
    END
  END pdp11_oeb[5]
  PIN pdp11_oeb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 333.760 696.000 334.320 700.000 ;
    END
  END pdp11_oeb[6]
  PIN pdp11_oeb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 340.480 696.000 341.040 700.000 ;
    END
  END pdp11_oeb[7]
  PIN pdp11_oeb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 347.200 696.000 347.760 700.000 ;
    END
  END pdp11_oeb[8]
  PIN pdp11_oeb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 353.920 696.000 354.480 700.000 ;
    END
  END pdp11_oeb[9]
  PIN qcpu_do[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 445.760 0.000 446.320 4.000 ;
    END
  END qcpu_do[0]
  PIN qcpu_do[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 490.560 0.000 491.120 4.000 ;
    END
  END qcpu_do[10]
  PIN qcpu_do[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 495.040 0.000 495.600 4.000 ;
    END
  END qcpu_do[11]
  PIN qcpu_do[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 499.520 0.000 500.080 4.000 ;
    END
  END qcpu_do[12]
  PIN qcpu_do[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 504.000 0.000 504.560 4.000 ;
    END
  END qcpu_do[13]
  PIN qcpu_do[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 508.480 0.000 509.040 4.000 ;
    END
  END qcpu_do[14]
  PIN qcpu_do[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 512.960 0.000 513.520 4.000 ;
    END
  END qcpu_do[15]
  PIN qcpu_do[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 517.440 0.000 518.000 4.000 ;
    END
  END qcpu_do[16]
  PIN qcpu_do[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 521.920 0.000 522.480 4.000 ;
    END
  END qcpu_do[17]
  PIN qcpu_do[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 526.400 0.000 526.960 4.000 ;
    END
  END qcpu_do[18]
  PIN qcpu_do[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 530.880 0.000 531.440 4.000 ;
    END
  END qcpu_do[19]
  PIN qcpu_do[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 450.240 0.000 450.800 4.000 ;
    END
  END qcpu_do[1]
  PIN qcpu_do[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 535.360 0.000 535.920 4.000 ;
    END
  END qcpu_do[20]
  PIN qcpu_do[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 539.840 0.000 540.400 4.000 ;
    END
  END qcpu_do[21]
  PIN qcpu_do[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 544.320 0.000 544.880 4.000 ;
    END
  END qcpu_do[22]
  PIN qcpu_do[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 548.800 0.000 549.360 4.000 ;
    END
  END qcpu_do[23]
  PIN qcpu_do[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 553.280 0.000 553.840 4.000 ;
    END
  END qcpu_do[24]
  PIN qcpu_do[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 557.760 0.000 558.320 4.000 ;
    END
  END qcpu_do[25]
  PIN qcpu_do[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 562.240 0.000 562.800 4.000 ;
    END
  END qcpu_do[26]
  PIN qcpu_do[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 566.720 0.000 567.280 4.000 ;
    END
  END qcpu_do[27]
  PIN qcpu_do[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 571.200 0.000 571.760 4.000 ;
    END
  END qcpu_do[28]
  PIN qcpu_do[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 575.680 0.000 576.240 4.000 ;
    END
  END qcpu_do[29]
  PIN qcpu_do[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 454.720 0.000 455.280 4.000 ;
    END
  END qcpu_do[2]
  PIN qcpu_do[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 580.160 0.000 580.720 4.000 ;
    END
  END qcpu_do[30]
  PIN qcpu_do[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 584.640 0.000 585.200 4.000 ;
    END
  END qcpu_do[31]
  PIN qcpu_do[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 589.120 0.000 589.680 4.000 ;
    END
  END qcpu_do[32]
  PIN qcpu_do[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 459.200 0.000 459.760 4.000 ;
    END
  END qcpu_do[3]
  PIN qcpu_do[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 463.680 0.000 464.240 4.000 ;
    END
  END qcpu_do[4]
  PIN qcpu_do[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 468.160 0.000 468.720 4.000 ;
    END
  END qcpu_do[5]
  PIN qcpu_do[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 472.640 0.000 473.200 4.000 ;
    END
  END qcpu_do[6]
  PIN qcpu_do[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 477.120 0.000 477.680 4.000 ;
    END
  END qcpu_do[7]
  PIN qcpu_do[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 481.600 0.000 482.160 4.000 ;
    END
  END qcpu_do[8]
  PIN qcpu_do[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 486.080 0.000 486.640 4.000 ;
    END
  END qcpu_do[9]
  PIN qcpu_oeb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 333.760 750.000 334.320 ;
    END
  END qcpu_oeb[0]
  PIN qcpu_oeb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 378.560 750.000 379.120 ;
    END
  END qcpu_oeb[10]
  PIN qcpu_oeb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 383.040 750.000 383.600 ;
    END
  END qcpu_oeb[11]
  PIN qcpu_oeb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 387.520 750.000 388.080 ;
    END
  END qcpu_oeb[12]
  PIN qcpu_oeb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 392.000 750.000 392.560 ;
    END
  END qcpu_oeb[13]
  PIN qcpu_oeb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 396.480 750.000 397.040 ;
    END
  END qcpu_oeb[14]
  PIN qcpu_oeb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 400.960 750.000 401.520 ;
    END
  END qcpu_oeb[15]
  PIN qcpu_oeb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 405.440 750.000 406.000 ;
    END
  END qcpu_oeb[16]
  PIN qcpu_oeb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 409.920 750.000 410.480 ;
    END
  END qcpu_oeb[17]
  PIN qcpu_oeb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 414.400 750.000 414.960 ;
    END
  END qcpu_oeb[18]
  PIN qcpu_oeb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 418.880 750.000 419.440 ;
    END
  END qcpu_oeb[19]
  PIN qcpu_oeb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 338.240 750.000 338.800 ;
    END
  END qcpu_oeb[1]
  PIN qcpu_oeb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 423.360 750.000 423.920 ;
    END
  END qcpu_oeb[20]
  PIN qcpu_oeb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 427.840 750.000 428.400 ;
    END
  END qcpu_oeb[21]
  PIN qcpu_oeb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 432.320 750.000 432.880 ;
    END
  END qcpu_oeb[22]
  PIN qcpu_oeb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 436.800 750.000 437.360 ;
    END
  END qcpu_oeb[23]
  PIN qcpu_oeb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 441.280 750.000 441.840 ;
    END
  END qcpu_oeb[24]
  PIN qcpu_oeb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 445.760 750.000 446.320 ;
    END
  END qcpu_oeb[25]
  PIN qcpu_oeb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 450.240 750.000 450.800 ;
    END
  END qcpu_oeb[26]
  PIN qcpu_oeb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 454.720 750.000 455.280 ;
    END
  END qcpu_oeb[27]
  PIN qcpu_oeb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 459.200 750.000 459.760 ;
    END
  END qcpu_oeb[28]
  PIN qcpu_oeb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 463.680 750.000 464.240 ;
    END
  END qcpu_oeb[29]
  PIN qcpu_oeb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 342.720 750.000 343.280 ;
    END
  END qcpu_oeb[2]
  PIN qcpu_oeb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 468.160 750.000 468.720 ;
    END
  END qcpu_oeb[30]
  PIN qcpu_oeb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 472.640 750.000 473.200 ;
    END
  END qcpu_oeb[31]
  PIN qcpu_oeb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 477.120 750.000 477.680 ;
    END
  END qcpu_oeb[32]
  PIN qcpu_oeb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 347.200 750.000 347.760 ;
    END
  END qcpu_oeb[3]
  PIN qcpu_oeb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 351.680 750.000 352.240 ;
    END
  END qcpu_oeb[4]
  PIN qcpu_oeb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 356.160 750.000 356.720 ;
    END
  END qcpu_oeb[5]
  PIN qcpu_oeb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 360.640 750.000 361.200 ;
    END
  END qcpu_oeb[6]
  PIN qcpu_oeb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 365.120 750.000 365.680 ;
    END
  END qcpu_oeb[7]
  PIN qcpu_oeb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 369.600 750.000 370.160 ;
    END
  END qcpu_oeb[8]
  PIN qcpu_oeb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 374.080 750.000 374.640 ;
    END
  END qcpu_oeb[9]
  PIN qcpu_sram_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 593.600 0.000 594.160 4.000 ;
    END
  END qcpu_sram_addr[0]
  PIN qcpu_sram_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 598.080 0.000 598.640 4.000 ;
    END
  END qcpu_sram_addr[1]
  PIN qcpu_sram_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 602.560 0.000 603.120 4.000 ;
    END
  END qcpu_sram_addr[2]
  PIN qcpu_sram_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 607.040 0.000 607.600 4.000 ;
    END
  END qcpu_sram_addr[3]
  PIN qcpu_sram_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 611.520 0.000 612.080 4.000 ;
    END
  END qcpu_sram_addr[4]
  PIN qcpu_sram_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 616.000 0.000 616.560 4.000 ;
    END
  END qcpu_sram_addr[5]
  PIN qcpu_sram_gwe
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 620.480 0.000 621.040 4.000 ;
    END
  END qcpu_sram_gwe
  PIN qcpu_sram_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 624.960 0.000 625.520 4.000 ;
    END
  END qcpu_sram_in[0]
  PIN qcpu_sram_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 629.440 0.000 630.000 4.000 ;
    END
  END qcpu_sram_in[1]
  PIN qcpu_sram_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 633.920 0.000 634.480 4.000 ;
    END
  END qcpu_sram_in[2]
  PIN qcpu_sram_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 638.400 0.000 638.960 4.000 ;
    END
  END qcpu_sram_in[3]
  PIN qcpu_sram_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 642.880 0.000 643.440 4.000 ;
    END
  END qcpu_sram_in[4]
  PIN qcpu_sram_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 647.360 0.000 647.920 4.000 ;
    END
  END qcpu_sram_in[5]
  PIN qcpu_sram_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 651.840 0.000 652.400 4.000 ;
    END
  END qcpu_sram_in[6]
  PIN qcpu_sram_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 656.320 0.000 656.880 4.000 ;
    END
  END qcpu_sram_in[7]
  PIN qcpu_sram_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 481.600 750.000 482.160 ;
    END
  END qcpu_sram_out[0]
  PIN qcpu_sram_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 486.080 750.000 486.640 ;
    END
  END qcpu_sram_out[1]
  PIN qcpu_sram_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 490.560 750.000 491.120 ;
    END
  END qcpu_sram_out[2]
  PIN qcpu_sram_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 495.040 750.000 495.600 ;
    END
  END qcpu_sram_out[3]
  PIN qcpu_sram_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 499.520 750.000 500.080 ;
    END
  END qcpu_sram_out[4]
  PIN qcpu_sram_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 504.000 750.000 504.560 ;
    END
  END qcpu_sram_out[5]
  PIN qcpu_sram_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 508.480 750.000 509.040 ;
    END
  END qcpu_sram_out[6]
  PIN qcpu_sram_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 512.960 750.000 513.520 ;
    END
  END qcpu_sram_out[7]
  PIN rst_ay8913
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 517.440 750.000 518.000 ;
    END
  END rst_ay8913
  PIN rst_blinker
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 626.080 4.000 626.640 ;
    END
  END rst_blinker
  PIN rst_diceroll
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 626.080 696.000 626.640 700.000 ;
    END
  END rst_diceroll
  PIN rst_hellorld
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 581.280 4.000 581.840 ;
    END
  END rst_hellorld
  PIN rst_mc14500
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 402.080 4.000 402.640 ;
    END
  END rst_mc14500
  PIN rst_pdp11
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 521.920 750.000 522.480 ;
    END
  END rst_pdp11
  PIN rst_qcpu
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 396.480 4.000 397.040 ;
    END
  END rst_qcpu
  PIN rst_sid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 267.680 4.000 268.240 ;
    END
  END rst_sid
  PIN rst_sn76489
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 192.640 696.000 193.200 700.000 ;
    END
  END rst_sn76489
  PIN rst_tbb1143
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 592.480 4.000 593.040 ;
    END
  END rst_tbb1143
  PIN rst_tholin_riscv
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 511.840 696.000 512.400 700.000 ;
    END
  END rst_tholin_riscv
  PIN rst_ue1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 659.680 696.000 660.240 700.000 ;
    END
  END rst_ue1
  PIN sid_do[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 273.280 4.000 273.840 ;
    END
  END sid_do[0]
  PIN sid_do[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 329.280 4.000 329.840 ;
    END
  END sid_do[10]
  PIN sid_do[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 334.880 4.000 335.440 ;
    END
  END sid_do[11]
  PIN sid_do[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 340.480 4.000 341.040 ;
    END
  END sid_do[12]
  PIN sid_do[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 346.080 4.000 346.640 ;
    END
  END sid_do[13]
  PIN sid_do[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 351.680 4.000 352.240 ;
    END
  END sid_do[14]
  PIN sid_do[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 357.280 4.000 357.840 ;
    END
  END sid_do[15]
  PIN sid_do[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 362.880 4.000 363.440 ;
    END
  END sid_do[16]
  PIN sid_do[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 368.480 4.000 369.040 ;
    END
  END sid_do[17]
  PIN sid_do[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 374.080 4.000 374.640 ;
    END
  END sid_do[18]
  PIN sid_do[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 379.680 4.000 380.240 ;
    END
  END sid_do[19]
  PIN sid_do[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 278.880 4.000 279.440 ;
    END
  END sid_do[1]
  PIN sid_do[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 385.280 4.000 385.840 ;
    END
  END sid_do[20]
  PIN sid_do[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 284.480 4.000 285.040 ;
    END
  END sid_do[2]
  PIN sid_do[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 290.080 4.000 290.640 ;
    END
  END sid_do[3]
  PIN sid_do[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 295.680 4.000 296.240 ;
    END
  END sid_do[4]
  PIN sid_do[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 301.280 4.000 301.840 ;
    END
  END sid_do[5]
  PIN sid_do[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 306.880 4.000 307.440 ;
    END
  END sid_do[6]
  PIN sid_do[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 312.480 4.000 313.040 ;
    END
  END sid_do[7]
  PIN sid_do[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 318.080 4.000 318.640 ;
    END
  END sid_do[8]
  PIN sid_do[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 323.680 4.000 324.240 ;
    END
  END sid_do[9]
  PIN sid_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 390.880 4.000 391.440 ;
    END
  END sid_oeb
  PIN sn76489_do[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 320.320 0.000 320.880 4.000 ;
    END
  END sn76489_do[0]
  PIN sn76489_do[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 365.120 0.000 365.680 4.000 ;
    END
  END sn76489_do[10]
  PIN sn76489_do[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 369.600 0.000 370.160 4.000 ;
    END
  END sn76489_do[11]
  PIN sn76489_do[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 374.080 0.000 374.640 4.000 ;
    END
  END sn76489_do[12]
  PIN sn76489_do[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 378.560 0.000 379.120 4.000 ;
    END
  END sn76489_do[13]
  PIN sn76489_do[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 383.040 0.000 383.600 4.000 ;
    END
  END sn76489_do[14]
  PIN sn76489_do[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 387.520 0.000 388.080 4.000 ;
    END
  END sn76489_do[15]
  PIN sn76489_do[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 392.000 0.000 392.560 4.000 ;
    END
  END sn76489_do[16]
  PIN sn76489_do[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 396.480 0.000 397.040 4.000 ;
    END
  END sn76489_do[17]
  PIN sn76489_do[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 400.960 0.000 401.520 4.000 ;
    END
  END sn76489_do[18]
  PIN sn76489_do[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 405.440 0.000 406.000 4.000 ;
    END
  END sn76489_do[19]
  PIN sn76489_do[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 324.800 0.000 325.360 4.000 ;
    END
  END sn76489_do[1]
  PIN sn76489_do[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 409.920 0.000 410.480 4.000 ;
    END
  END sn76489_do[20]
  PIN sn76489_do[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 414.400 0.000 414.960 4.000 ;
    END
  END sn76489_do[21]
  PIN sn76489_do[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 418.880 0.000 419.440 4.000 ;
    END
  END sn76489_do[22]
  PIN sn76489_do[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 423.360 0.000 423.920 4.000 ;
    END
  END sn76489_do[23]
  PIN sn76489_do[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 427.840 0.000 428.400 4.000 ;
    END
  END sn76489_do[24]
  PIN sn76489_do[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 432.320 0.000 432.880 4.000 ;
    END
  END sn76489_do[25]
  PIN sn76489_do[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 436.800 0.000 437.360 4.000 ;
    END
  END sn76489_do[26]
  PIN sn76489_do[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 441.280 0.000 441.840 4.000 ;
    END
  END sn76489_do[27]
  PIN sn76489_do[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 329.280 0.000 329.840 4.000 ;
    END
  END sn76489_do[2]
  PIN sn76489_do[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 333.760 0.000 334.320 4.000 ;
    END
  END sn76489_do[3]
  PIN sn76489_do[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 338.240 0.000 338.800 4.000 ;
    END
  END sn76489_do[4]
  PIN sn76489_do[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 342.720 0.000 343.280 4.000 ;
    END
  END sn76489_do[5]
  PIN sn76489_do[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 347.200 0.000 347.760 4.000 ;
    END
  END sn76489_do[6]
  PIN sn76489_do[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 351.680 0.000 352.240 4.000 ;
    END
  END sn76489_do[7]
  PIN sn76489_do[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 356.160 0.000 356.720 4.000 ;
    END
  END sn76489_do[8]
  PIN sn76489_do[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 360.640 0.000 361.200 4.000 ;
    END
  END sn76489_do[9]
  PIN tbb1143_do[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 598.080 4.000 598.640 ;
    END
  END tbb1143_do[0]
  PIN tbb1143_do[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 603.680 4.000 604.240 ;
    END
  END tbb1143_do[1]
  PIN tbb1143_do[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 609.280 4.000 609.840 ;
    END
  END tbb1143_do[2]
  PIN tbb1143_do[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 614.880 4.000 615.440 ;
    END
  END tbb1143_do[3]
  PIN tbb1143_do[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 620.480 4.000 621.040 ;
    END
  END tbb1143_do[4]
  PIN tholin_riscv_do[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 526.400 750.000 526.960 ;
    END
  END tholin_riscv_do[0]
  PIN tholin_riscv_do[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 571.200 750.000 571.760 ;
    END
  END tholin_riscv_do[10]
  PIN tholin_riscv_do[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 575.680 750.000 576.240 ;
    END
  END tholin_riscv_do[11]
  PIN tholin_riscv_do[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 580.160 750.000 580.720 ;
    END
  END tholin_riscv_do[12]
  PIN tholin_riscv_do[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 584.640 750.000 585.200 ;
    END
  END tholin_riscv_do[13]
  PIN tholin_riscv_do[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 589.120 750.000 589.680 ;
    END
  END tholin_riscv_do[14]
  PIN tholin_riscv_do[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 593.600 750.000 594.160 ;
    END
  END tholin_riscv_do[15]
  PIN tholin_riscv_do[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 598.080 750.000 598.640 ;
    END
  END tholin_riscv_do[16]
  PIN tholin_riscv_do[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 602.560 750.000 603.120 ;
    END
  END tholin_riscv_do[17]
  PIN tholin_riscv_do[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 607.040 750.000 607.600 ;
    END
  END tholin_riscv_do[18]
  PIN tholin_riscv_do[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 611.520 750.000 612.080 ;
    END
  END tholin_riscv_do[19]
  PIN tholin_riscv_do[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 530.880 750.000 531.440 ;
    END
  END tholin_riscv_do[1]
  PIN tholin_riscv_do[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 616.000 750.000 616.560 ;
    END
  END tholin_riscv_do[20]
  PIN tholin_riscv_do[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 620.480 750.000 621.040 ;
    END
  END tholin_riscv_do[21]
  PIN tholin_riscv_do[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 624.960 750.000 625.520 ;
    END
  END tholin_riscv_do[22]
  PIN tholin_riscv_do[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 629.440 750.000 630.000 ;
    END
  END tholin_riscv_do[23]
  PIN tholin_riscv_do[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 633.920 750.000 634.480 ;
    END
  END tholin_riscv_do[24]
  PIN tholin_riscv_do[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 638.400 750.000 638.960 ;
    END
  END tholin_riscv_do[25]
  PIN tholin_riscv_do[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 642.880 750.000 643.440 ;
    END
  END tholin_riscv_do[26]
  PIN tholin_riscv_do[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 647.360 750.000 647.920 ;
    END
  END tholin_riscv_do[27]
  PIN tholin_riscv_do[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 651.840 750.000 652.400 ;
    END
  END tholin_riscv_do[28]
  PIN tholin_riscv_do[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 656.320 750.000 656.880 ;
    END
  END tholin_riscv_do[29]
  PIN tholin_riscv_do[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 535.360 750.000 535.920 ;
    END
  END tholin_riscv_do[2]
  PIN tholin_riscv_do[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 660.800 750.000 661.360 ;
    END
  END tholin_riscv_do[30]
  PIN tholin_riscv_do[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 665.280 750.000 665.840 ;
    END
  END tholin_riscv_do[31]
  PIN tholin_riscv_do[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 669.760 750.000 670.320 ;
    END
  END tholin_riscv_do[32]
  PIN tholin_riscv_do[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 539.840 750.000 540.400 ;
    END
  END tholin_riscv_do[3]
  PIN tholin_riscv_do[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 544.320 750.000 544.880 ;
    END
  END tholin_riscv_do[4]
  PIN tholin_riscv_do[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 548.800 750.000 549.360 ;
    END
  END tholin_riscv_do[5]
  PIN tholin_riscv_do[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 553.280 750.000 553.840 ;
    END
  END tholin_riscv_do[6]
  PIN tholin_riscv_do[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 557.760 750.000 558.320 ;
    END
  END tholin_riscv_do[7]
  PIN tholin_riscv_do[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 562.240 750.000 562.800 ;
    END
  END tholin_riscv_do[8]
  PIN tholin_riscv_do[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 566.720 750.000 567.280 ;
    END
  END tholin_riscv_do[9]
  PIN tholin_riscv_oeb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 515.200 696.000 515.760 700.000 ;
    END
  END tholin_riscv_oeb[0]
  PIN tholin_riscv_oeb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 548.800 696.000 549.360 700.000 ;
    END
  END tholin_riscv_oeb[10]
  PIN tholin_riscv_oeb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 552.160 696.000 552.720 700.000 ;
    END
  END tholin_riscv_oeb[11]
  PIN tholin_riscv_oeb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 555.520 696.000 556.080 700.000 ;
    END
  END tholin_riscv_oeb[12]
  PIN tholin_riscv_oeb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 558.880 696.000 559.440 700.000 ;
    END
  END tholin_riscv_oeb[13]
  PIN tholin_riscv_oeb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 562.240 696.000 562.800 700.000 ;
    END
  END tholin_riscv_oeb[14]
  PIN tholin_riscv_oeb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 565.600 696.000 566.160 700.000 ;
    END
  END tholin_riscv_oeb[15]
  PIN tholin_riscv_oeb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 568.960 696.000 569.520 700.000 ;
    END
  END tholin_riscv_oeb[16]
  PIN tholin_riscv_oeb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 572.320 696.000 572.880 700.000 ;
    END
  END tholin_riscv_oeb[17]
  PIN tholin_riscv_oeb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 575.680 696.000 576.240 700.000 ;
    END
  END tholin_riscv_oeb[18]
  PIN tholin_riscv_oeb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 579.040 696.000 579.600 700.000 ;
    END
  END tholin_riscv_oeb[19]
  PIN tholin_riscv_oeb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 518.560 696.000 519.120 700.000 ;
    END
  END tholin_riscv_oeb[1]
  PIN tholin_riscv_oeb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 582.400 696.000 582.960 700.000 ;
    END
  END tholin_riscv_oeb[20]
  PIN tholin_riscv_oeb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 585.760 696.000 586.320 700.000 ;
    END
  END tholin_riscv_oeb[21]
  PIN tholin_riscv_oeb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 589.120 696.000 589.680 700.000 ;
    END
  END tholin_riscv_oeb[22]
  PIN tholin_riscv_oeb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 592.480 696.000 593.040 700.000 ;
    END
  END tholin_riscv_oeb[23]
  PIN tholin_riscv_oeb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 595.840 696.000 596.400 700.000 ;
    END
  END tholin_riscv_oeb[24]
  PIN tholin_riscv_oeb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 599.200 696.000 599.760 700.000 ;
    END
  END tholin_riscv_oeb[25]
  PIN tholin_riscv_oeb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 602.560 696.000 603.120 700.000 ;
    END
  END tholin_riscv_oeb[26]
  PIN tholin_riscv_oeb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 605.920 696.000 606.480 700.000 ;
    END
  END tholin_riscv_oeb[27]
  PIN tholin_riscv_oeb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 609.280 696.000 609.840 700.000 ;
    END
  END tholin_riscv_oeb[28]
  PIN tholin_riscv_oeb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 612.640 696.000 613.200 700.000 ;
    END
  END tholin_riscv_oeb[29]
  PIN tholin_riscv_oeb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 521.920 696.000 522.480 700.000 ;
    END
  END tholin_riscv_oeb[2]
  PIN tholin_riscv_oeb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 616.000 696.000 616.560 700.000 ;
    END
  END tholin_riscv_oeb[30]
  PIN tholin_riscv_oeb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 619.360 696.000 619.920 700.000 ;
    END
  END tholin_riscv_oeb[31]
  PIN tholin_riscv_oeb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 622.720 696.000 623.280 700.000 ;
    END
  END tholin_riscv_oeb[32]
  PIN tholin_riscv_oeb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 525.280 696.000 525.840 700.000 ;
    END
  END tholin_riscv_oeb[3]
  PIN tholin_riscv_oeb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 528.640 696.000 529.200 700.000 ;
    END
  END tholin_riscv_oeb[4]
  PIN tholin_riscv_oeb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 532.000 696.000 532.560 700.000 ;
    END
  END tholin_riscv_oeb[5]
  PIN tholin_riscv_oeb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 535.360 696.000 535.920 700.000 ;
    END
  END tholin_riscv_oeb[6]
  PIN tholin_riscv_oeb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 538.720 696.000 539.280 700.000 ;
    END
  END tholin_riscv_oeb[7]
  PIN tholin_riscv_oeb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 542.080 696.000 542.640 700.000 ;
    END
  END tholin_riscv_oeb[8]
  PIN tholin_riscv_oeb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 545.440 696.000 546.000 700.000 ;
    END
  END tholin_riscv_oeb[9]
  PIN ue1_do[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 666.400 696.000 666.960 700.000 ;
    END
  END ue1_do[0]
  PIN ue1_do[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 669.760 696.000 670.320 700.000 ;
    END
  END ue1_do[1]
  PIN ue1_do[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 673.120 696.000 673.680 700.000 ;
    END
  END ue1_do[2]
  PIN ue1_do[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 676.480 696.000 677.040 700.000 ;
    END
  END ue1_do[3]
  PIN ue1_do[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 679.840 696.000 680.400 700.000 ;
    END
  END ue1_do[4]
  PIN ue1_do[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 683.200 696.000 683.760 700.000 ;
    END
  END ue1_do[5]
  PIN ue1_do[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 686.560 696.000 687.120 700.000 ;
    END
  END ue1_do[6]
  PIN ue1_do[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 689.920 696.000 690.480 700.000 ;
    END
  END ue1_do[7]
  PIN ue1_do[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 693.280 696.000 693.840 700.000 ;
    END
  END ue1_do[8]
  PIN ue1_do[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 696.640 696.000 697.200 700.000 ;
    END
  END ue1_do[9]
  PIN ue1_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 663.040 696.000 663.600 700.000 ;
    END
  END ue1_oeb
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 682.380 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 682.380 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 24.640 0.000 25.200 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 29.120 0.000 29.680 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 185.920 750.000 186.480 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 0.000 34.160 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 78.400 0.000 78.960 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 82.880 0.000 83.440 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 0.000 87.920 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 91.840 0.000 92.400 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 96.320 0.000 96.880 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 0.000 101.360 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 105.280 0.000 105.840 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 109.760 0.000 110.320 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 0.000 114.800 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 118.720 0.000 119.280 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 38.080 0.000 38.640 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 123.200 0.000 123.760 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 0.000 128.240 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 132.160 0.000 132.720 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 136.640 0.000 137.200 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 0.000 141.680 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 145.600 0.000 146.160 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 150.080 0.000 150.640 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 0.000 155.120 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 159.040 0.000 159.600 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 163.520 0.000 164.080 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 42.560 0.000 43.120 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 0.000 168.560 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 172.480 0.000 173.040 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 0.000 47.600 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 51.520 0.000 52.080 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 56.000 0.000 56.560 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 0.000 61.040 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 64.960 0.000 65.520 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 69.440 0.000 70.000 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 0.000 74.480 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 176.960 750.000 177.520 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 176.960 0.000 177.520 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 0.000 222.320 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 226.240 0.000 226.800 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 230.720 0.000 231.280 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 235.200 0.000 235.760 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 239.680 0.000 240.240 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 244.160 0.000 244.720 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 0.000 249.200 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 253.120 0.000 253.680 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 257.600 0.000 258.160 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 0.000 262.640 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 181.440 0.000 182.000 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 266.560 0.000 267.120 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 271.040 0.000 271.600 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 0.000 276.080 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 280.000 0.000 280.560 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 284.480 0.000 285.040 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 288.960 0.000 289.520 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 293.440 0.000 294.000 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 297.920 0.000 298.480 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 302.400 0.000 302.960 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 306.880 0.000 307.440 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 185.920 0.000 186.480 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 311.360 0.000 311.920 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 315.840 0.000 316.400 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 190.400 0.000 190.960 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 0.000 195.440 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 199.360 0.000 199.920 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 203.840 0.000 204.400 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 208.320 0.000 208.880 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 212.800 0.000 213.360 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 217.280 0.000 217.840 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 29.120 750.000 29.680 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 73.920 750.000 74.480 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 78.400 750.000 78.960 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 82.880 750.000 83.440 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 87.360 750.000 87.920 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 91.840 750.000 92.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 96.320 750.000 96.880 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 100.800 750.000 101.360 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 105.280 750.000 105.840 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 109.760 750.000 110.320 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 114.240 750.000 114.800 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 33.600 750.000 34.160 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 118.720 750.000 119.280 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 123.200 750.000 123.760 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 127.680 750.000 128.240 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 132.160 750.000 132.720 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 136.640 750.000 137.200 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 141.120 750.000 141.680 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 145.600 750.000 146.160 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 150.080 750.000 150.640 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 154.560 750.000 155.120 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 159.040 750.000 159.600 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 38.080 750.000 38.640 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 163.520 750.000 164.080 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 168.000 750.000 168.560 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 42.560 750.000 43.120 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 47.040 750.000 47.600 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 51.520 750.000 52.080 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 56.000 750.000 56.560 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 60.480 750.000 61.040 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 64.960 750.000 65.520 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 69.440 750.000 70.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 181.440 750.000 182.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 172.480 750.000 173.040 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 13.590 743.120 683.050 ;
      LAYER Metal2 ;
        RECT 7.980 695.700 51.220 696.000 ;
        RECT 52.380 695.700 54.580 696.000 ;
        RECT 55.740 695.700 57.940 696.000 ;
        RECT 59.100 695.700 61.300 696.000 ;
        RECT 62.460 695.700 64.660 696.000 ;
        RECT 65.820 695.700 68.020 696.000 ;
        RECT 69.180 695.700 71.380 696.000 ;
        RECT 72.540 695.700 74.740 696.000 ;
        RECT 75.900 695.700 78.100 696.000 ;
        RECT 79.260 695.700 81.460 696.000 ;
        RECT 82.620 695.700 84.820 696.000 ;
        RECT 85.980 695.700 88.180 696.000 ;
        RECT 89.340 695.700 91.540 696.000 ;
        RECT 92.700 695.700 94.900 696.000 ;
        RECT 96.060 695.700 98.260 696.000 ;
        RECT 99.420 695.700 101.620 696.000 ;
        RECT 102.780 695.700 104.980 696.000 ;
        RECT 106.140 695.700 108.340 696.000 ;
        RECT 109.500 695.700 111.700 696.000 ;
        RECT 112.860 695.700 115.060 696.000 ;
        RECT 116.220 695.700 118.420 696.000 ;
        RECT 119.580 695.700 121.780 696.000 ;
        RECT 122.940 695.700 125.140 696.000 ;
        RECT 126.300 695.700 128.500 696.000 ;
        RECT 129.660 695.700 131.860 696.000 ;
        RECT 133.020 695.700 135.220 696.000 ;
        RECT 136.380 695.700 138.580 696.000 ;
        RECT 139.740 695.700 141.940 696.000 ;
        RECT 143.100 695.700 145.300 696.000 ;
        RECT 146.460 695.700 148.660 696.000 ;
        RECT 149.820 695.700 152.020 696.000 ;
        RECT 153.180 695.700 155.380 696.000 ;
        RECT 156.540 695.700 158.740 696.000 ;
        RECT 159.900 695.700 162.100 696.000 ;
        RECT 163.260 695.700 165.460 696.000 ;
        RECT 166.620 695.700 168.820 696.000 ;
        RECT 169.980 695.700 172.180 696.000 ;
        RECT 173.340 695.700 175.540 696.000 ;
        RECT 176.700 695.700 178.900 696.000 ;
        RECT 180.060 695.700 182.260 696.000 ;
        RECT 183.420 695.700 185.620 696.000 ;
        RECT 186.780 695.700 188.980 696.000 ;
        RECT 190.140 695.700 192.340 696.000 ;
        RECT 193.500 695.700 195.700 696.000 ;
        RECT 196.860 695.700 199.060 696.000 ;
        RECT 200.220 695.700 202.420 696.000 ;
        RECT 203.580 695.700 205.780 696.000 ;
        RECT 206.940 695.700 209.140 696.000 ;
        RECT 210.300 695.700 212.500 696.000 ;
        RECT 213.660 695.700 215.860 696.000 ;
        RECT 217.020 695.700 219.220 696.000 ;
        RECT 220.380 695.700 222.580 696.000 ;
        RECT 223.740 695.700 225.940 696.000 ;
        RECT 227.100 695.700 229.300 696.000 ;
        RECT 230.460 695.700 232.660 696.000 ;
        RECT 233.820 695.700 236.020 696.000 ;
        RECT 237.180 695.700 239.380 696.000 ;
        RECT 240.540 695.700 242.740 696.000 ;
        RECT 243.900 695.700 246.100 696.000 ;
        RECT 247.260 695.700 249.460 696.000 ;
        RECT 250.620 695.700 252.820 696.000 ;
        RECT 253.980 695.700 256.180 696.000 ;
        RECT 257.340 695.700 259.540 696.000 ;
        RECT 260.700 695.700 262.900 696.000 ;
        RECT 264.060 695.700 266.260 696.000 ;
        RECT 267.420 695.700 269.620 696.000 ;
        RECT 270.780 695.700 272.980 696.000 ;
        RECT 274.140 695.700 276.340 696.000 ;
        RECT 277.500 695.700 279.700 696.000 ;
        RECT 280.860 695.700 283.060 696.000 ;
        RECT 284.220 695.700 286.420 696.000 ;
        RECT 287.580 695.700 289.780 696.000 ;
        RECT 290.940 695.700 293.140 696.000 ;
        RECT 294.300 695.700 296.500 696.000 ;
        RECT 297.660 695.700 299.860 696.000 ;
        RECT 301.020 695.700 303.220 696.000 ;
        RECT 304.380 695.700 306.580 696.000 ;
        RECT 307.740 695.700 309.940 696.000 ;
        RECT 311.100 695.700 313.300 696.000 ;
        RECT 314.460 695.700 316.660 696.000 ;
        RECT 317.820 695.700 320.020 696.000 ;
        RECT 321.180 695.700 323.380 696.000 ;
        RECT 324.540 695.700 326.740 696.000 ;
        RECT 327.900 695.700 330.100 696.000 ;
        RECT 331.260 695.700 333.460 696.000 ;
        RECT 334.620 695.700 336.820 696.000 ;
        RECT 337.980 695.700 340.180 696.000 ;
        RECT 341.340 695.700 343.540 696.000 ;
        RECT 344.700 695.700 346.900 696.000 ;
        RECT 348.060 695.700 350.260 696.000 ;
        RECT 351.420 695.700 353.620 696.000 ;
        RECT 354.780 695.700 356.980 696.000 ;
        RECT 358.140 695.700 360.340 696.000 ;
        RECT 361.500 695.700 363.700 696.000 ;
        RECT 364.860 695.700 367.060 696.000 ;
        RECT 368.220 695.700 370.420 696.000 ;
        RECT 371.580 695.700 373.780 696.000 ;
        RECT 374.940 695.700 377.140 696.000 ;
        RECT 378.300 695.700 380.500 696.000 ;
        RECT 381.660 695.700 383.860 696.000 ;
        RECT 385.020 695.700 387.220 696.000 ;
        RECT 388.380 695.700 390.580 696.000 ;
        RECT 391.740 695.700 393.940 696.000 ;
        RECT 395.100 695.700 397.300 696.000 ;
        RECT 398.460 695.700 400.660 696.000 ;
        RECT 401.820 695.700 404.020 696.000 ;
        RECT 405.180 695.700 407.380 696.000 ;
        RECT 408.540 695.700 410.740 696.000 ;
        RECT 411.900 695.700 414.100 696.000 ;
        RECT 415.260 695.700 417.460 696.000 ;
        RECT 418.620 695.700 420.820 696.000 ;
        RECT 421.980 695.700 424.180 696.000 ;
        RECT 425.340 695.700 427.540 696.000 ;
        RECT 428.700 695.700 430.900 696.000 ;
        RECT 432.060 695.700 434.260 696.000 ;
        RECT 435.420 695.700 437.620 696.000 ;
        RECT 438.780 695.700 440.980 696.000 ;
        RECT 442.140 695.700 444.340 696.000 ;
        RECT 445.500 695.700 447.700 696.000 ;
        RECT 448.860 695.700 451.060 696.000 ;
        RECT 452.220 695.700 454.420 696.000 ;
        RECT 455.580 695.700 457.780 696.000 ;
        RECT 458.940 695.700 461.140 696.000 ;
        RECT 462.300 695.700 464.500 696.000 ;
        RECT 465.660 695.700 467.860 696.000 ;
        RECT 469.020 695.700 471.220 696.000 ;
        RECT 472.380 695.700 474.580 696.000 ;
        RECT 475.740 695.700 477.940 696.000 ;
        RECT 479.100 695.700 481.300 696.000 ;
        RECT 482.460 695.700 484.660 696.000 ;
        RECT 485.820 695.700 488.020 696.000 ;
        RECT 489.180 695.700 491.380 696.000 ;
        RECT 492.540 695.700 494.740 696.000 ;
        RECT 495.900 695.700 498.100 696.000 ;
        RECT 499.260 695.700 501.460 696.000 ;
        RECT 502.620 695.700 504.820 696.000 ;
        RECT 505.980 695.700 508.180 696.000 ;
        RECT 509.340 695.700 511.540 696.000 ;
        RECT 512.700 695.700 514.900 696.000 ;
        RECT 516.060 695.700 518.260 696.000 ;
        RECT 519.420 695.700 521.620 696.000 ;
        RECT 522.780 695.700 524.980 696.000 ;
        RECT 526.140 695.700 528.340 696.000 ;
        RECT 529.500 695.700 531.700 696.000 ;
        RECT 532.860 695.700 535.060 696.000 ;
        RECT 536.220 695.700 538.420 696.000 ;
        RECT 539.580 695.700 541.780 696.000 ;
        RECT 542.940 695.700 545.140 696.000 ;
        RECT 546.300 695.700 548.500 696.000 ;
        RECT 549.660 695.700 551.860 696.000 ;
        RECT 553.020 695.700 555.220 696.000 ;
        RECT 556.380 695.700 558.580 696.000 ;
        RECT 559.740 695.700 561.940 696.000 ;
        RECT 563.100 695.700 565.300 696.000 ;
        RECT 566.460 695.700 568.660 696.000 ;
        RECT 569.820 695.700 572.020 696.000 ;
        RECT 573.180 695.700 575.380 696.000 ;
        RECT 576.540 695.700 578.740 696.000 ;
        RECT 579.900 695.700 582.100 696.000 ;
        RECT 583.260 695.700 585.460 696.000 ;
        RECT 586.620 695.700 588.820 696.000 ;
        RECT 589.980 695.700 592.180 696.000 ;
        RECT 593.340 695.700 595.540 696.000 ;
        RECT 596.700 695.700 598.900 696.000 ;
        RECT 600.060 695.700 602.260 696.000 ;
        RECT 603.420 695.700 605.620 696.000 ;
        RECT 606.780 695.700 608.980 696.000 ;
        RECT 610.140 695.700 612.340 696.000 ;
        RECT 613.500 695.700 615.700 696.000 ;
        RECT 616.860 695.700 619.060 696.000 ;
        RECT 620.220 695.700 622.420 696.000 ;
        RECT 623.580 695.700 625.780 696.000 ;
        RECT 626.940 695.700 629.140 696.000 ;
        RECT 630.300 695.700 632.500 696.000 ;
        RECT 633.660 695.700 635.860 696.000 ;
        RECT 637.020 695.700 639.220 696.000 ;
        RECT 640.380 695.700 642.580 696.000 ;
        RECT 643.740 695.700 645.940 696.000 ;
        RECT 647.100 695.700 649.300 696.000 ;
        RECT 650.460 695.700 652.660 696.000 ;
        RECT 653.820 695.700 656.020 696.000 ;
        RECT 657.180 695.700 659.380 696.000 ;
        RECT 660.540 695.700 662.740 696.000 ;
        RECT 663.900 695.700 666.100 696.000 ;
        RECT 667.260 695.700 669.460 696.000 ;
        RECT 670.620 695.700 672.820 696.000 ;
        RECT 673.980 695.700 676.180 696.000 ;
        RECT 677.340 695.700 679.540 696.000 ;
        RECT 680.700 695.700 682.900 696.000 ;
        RECT 684.060 695.700 686.260 696.000 ;
        RECT 687.420 695.700 689.620 696.000 ;
        RECT 690.780 695.700 692.980 696.000 ;
        RECT 694.140 695.700 696.340 696.000 ;
        RECT 697.500 695.700 741.860 696.000 ;
        RECT 7.980 4.300 741.860 695.700 ;
        RECT 7.980 3.450 24.340 4.300 ;
        RECT 25.500 3.450 28.820 4.300 ;
        RECT 29.980 3.450 33.300 4.300 ;
        RECT 34.460 3.450 37.780 4.300 ;
        RECT 38.940 3.450 42.260 4.300 ;
        RECT 43.420 3.450 46.740 4.300 ;
        RECT 47.900 3.450 51.220 4.300 ;
        RECT 52.380 3.450 55.700 4.300 ;
        RECT 56.860 3.450 60.180 4.300 ;
        RECT 61.340 3.450 64.660 4.300 ;
        RECT 65.820 3.450 69.140 4.300 ;
        RECT 70.300 3.450 73.620 4.300 ;
        RECT 74.780 3.450 78.100 4.300 ;
        RECT 79.260 3.450 82.580 4.300 ;
        RECT 83.740 3.450 87.060 4.300 ;
        RECT 88.220 3.450 91.540 4.300 ;
        RECT 92.700 3.450 96.020 4.300 ;
        RECT 97.180 3.450 100.500 4.300 ;
        RECT 101.660 3.450 104.980 4.300 ;
        RECT 106.140 3.450 109.460 4.300 ;
        RECT 110.620 3.450 113.940 4.300 ;
        RECT 115.100 3.450 118.420 4.300 ;
        RECT 119.580 3.450 122.900 4.300 ;
        RECT 124.060 3.450 127.380 4.300 ;
        RECT 128.540 3.450 131.860 4.300 ;
        RECT 133.020 3.450 136.340 4.300 ;
        RECT 137.500 3.450 140.820 4.300 ;
        RECT 141.980 3.450 145.300 4.300 ;
        RECT 146.460 3.450 149.780 4.300 ;
        RECT 150.940 3.450 154.260 4.300 ;
        RECT 155.420 3.450 158.740 4.300 ;
        RECT 159.900 3.450 163.220 4.300 ;
        RECT 164.380 3.450 167.700 4.300 ;
        RECT 168.860 3.450 172.180 4.300 ;
        RECT 173.340 3.450 176.660 4.300 ;
        RECT 177.820 3.450 181.140 4.300 ;
        RECT 182.300 3.450 185.620 4.300 ;
        RECT 186.780 3.450 190.100 4.300 ;
        RECT 191.260 3.450 194.580 4.300 ;
        RECT 195.740 3.450 199.060 4.300 ;
        RECT 200.220 3.450 203.540 4.300 ;
        RECT 204.700 3.450 208.020 4.300 ;
        RECT 209.180 3.450 212.500 4.300 ;
        RECT 213.660 3.450 216.980 4.300 ;
        RECT 218.140 3.450 221.460 4.300 ;
        RECT 222.620 3.450 225.940 4.300 ;
        RECT 227.100 3.450 230.420 4.300 ;
        RECT 231.580 3.450 234.900 4.300 ;
        RECT 236.060 3.450 239.380 4.300 ;
        RECT 240.540 3.450 243.860 4.300 ;
        RECT 245.020 3.450 248.340 4.300 ;
        RECT 249.500 3.450 252.820 4.300 ;
        RECT 253.980 3.450 257.300 4.300 ;
        RECT 258.460 3.450 261.780 4.300 ;
        RECT 262.940 3.450 266.260 4.300 ;
        RECT 267.420 3.450 270.740 4.300 ;
        RECT 271.900 3.450 275.220 4.300 ;
        RECT 276.380 3.450 279.700 4.300 ;
        RECT 280.860 3.450 284.180 4.300 ;
        RECT 285.340 3.450 288.660 4.300 ;
        RECT 289.820 3.450 293.140 4.300 ;
        RECT 294.300 3.450 297.620 4.300 ;
        RECT 298.780 3.450 302.100 4.300 ;
        RECT 303.260 3.450 306.580 4.300 ;
        RECT 307.740 3.450 311.060 4.300 ;
        RECT 312.220 3.450 315.540 4.300 ;
        RECT 316.700 3.450 320.020 4.300 ;
        RECT 321.180 3.450 324.500 4.300 ;
        RECT 325.660 3.450 328.980 4.300 ;
        RECT 330.140 3.450 333.460 4.300 ;
        RECT 334.620 3.450 337.940 4.300 ;
        RECT 339.100 3.450 342.420 4.300 ;
        RECT 343.580 3.450 346.900 4.300 ;
        RECT 348.060 3.450 351.380 4.300 ;
        RECT 352.540 3.450 355.860 4.300 ;
        RECT 357.020 3.450 360.340 4.300 ;
        RECT 361.500 3.450 364.820 4.300 ;
        RECT 365.980 3.450 369.300 4.300 ;
        RECT 370.460 3.450 373.780 4.300 ;
        RECT 374.940 3.450 378.260 4.300 ;
        RECT 379.420 3.450 382.740 4.300 ;
        RECT 383.900 3.450 387.220 4.300 ;
        RECT 388.380 3.450 391.700 4.300 ;
        RECT 392.860 3.450 396.180 4.300 ;
        RECT 397.340 3.450 400.660 4.300 ;
        RECT 401.820 3.450 405.140 4.300 ;
        RECT 406.300 3.450 409.620 4.300 ;
        RECT 410.780 3.450 414.100 4.300 ;
        RECT 415.260 3.450 418.580 4.300 ;
        RECT 419.740 3.450 423.060 4.300 ;
        RECT 424.220 3.450 427.540 4.300 ;
        RECT 428.700 3.450 432.020 4.300 ;
        RECT 433.180 3.450 436.500 4.300 ;
        RECT 437.660 3.450 440.980 4.300 ;
        RECT 442.140 3.450 445.460 4.300 ;
        RECT 446.620 3.450 449.940 4.300 ;
        RECT 451.100 3.450 454.420 4.300 ;
        RECT 455.580 3.450 458.900 4.300 ;
        RECT 460.060 3.450 463.380 4.300 ;
        RECT 464.540 3.450 467.860 4.300 ;
        RECT 469.020 3.450 472.340 4.300 ;
        RECT 473.500 3.450 476.820 4.300 ;
        RECT 477.980 3.450 481.300 4.300 ;
        RECT 482.460 3.450 485.780 4.300 ;
        RECT 486.940 3.450 490.260 4.300 ;
        RECT 491.420 3.450 494.740 4.300 ;
        RECT 495.900 3.450 499.220 4.300 ;
        RECT 500.380 3.450 503.700 4.300 ;
        RECT 504.860 3.450 508.180 4.300 ;
        RECT 509.340 3.450 512.660 4.300 ;
        RECT 513.820 3.450 517.140 4.300 ;
        RECT 518.300 3.450 521.620 4.300 ;
        RECT 522.780 3.450 526.100 4.300 ;
        RECT 527.260 3.450 530.580 4.300 ;
        RECT 531.740 3.450 535.060 4.300 ;
        RECT 536.220 3.450 539.540 4.300 ;
        RECT 540.700 3.450 544.020 4.300 ;
        RECT 545.180 3.450 548.500 4.300 ;
        RECT 549.660 3.450 552.980 4.300 ;
        RECT 554.140 3.450 557.460 4.300 ;
        RECT 558.620 3.450 561.940 4.300 ;
        RECT 563.100 3.450 566.420 4.300 ;
        RECT 567.580 3.450 570.900 4.300 ;
        RECT 572.060 3.450 575.380 4.300 ;
        RECT 576.540 3.450 579.860 4.300 ;
        RECT 581.020 3.450 584.340 4.300 ;
        RECT 585.500 3.450 588.820 4.300 ;
        RECT 589.980 3.450 593.300 4.300 ;
        RECT 594.460 3.450 597.780 4.300 ;
        RECT 598.940 3.450 602.260 4.300 ;
        RECT 603.420 3.450 606.740 4.300 ;
        RECT 607.900 3.450 611.220 4.300 ;
        RECT 612.380 3.450 615.700 4.300 ;
        RECT 616.860 3.450 620.180 4.300 ;
        RECT 621.340 3.450 624.660 4.300 ;
        RECT 625.820 3.450 629.140 4.300 ;
        RECT 630.300 3.450 633.620 4.300 ;
        RECT 634.780 3.450 638.100 4.300 ;
        RECT 639.260 3.450 642.580 4.300 ;
        RECT 643.740 3.450 647.060 4.300 ;
        RECT 648.220 3.450 651.540 4.300 ;
        RECT 652.700 3.450 656.020 4.300 ;
        RECT 657.180 3.450 660.500 4.300 ;
        RECT 661.660 3.450 664.980 4.300 ;
        RECT 666.140 3.450 669.460 4.300 ;
        RECT 670.620 3.450 673.940 4.300 ;
        RECT 675.100 3.450 678.420 4.300 ;
        RECT 679.580 3.450 682.900 4.300 ;
        RECT 684.060 3.450 687.380 4.300 ;
        RECT 688.540 3.450 691.860 4.300 ;
        RECT 693.020 3.450 696.340 4.300 ;
        RECT 697.500 3.450 700.820 4.300 ;
        RECT 701.980 3.450 705.300 4.300 ;
        RECT 706.460 3.450 709.780 4.300 ;
        RECT 710.940 3.450 714.260 4.300 ;
        RECT 715.420 3.450 718.740 4.300 ;
        RECT 719.900 3.450 723.220 4.300 ;
        RECT 724.380 3.450 741.860 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 670.620 746.340 692.580 ;
        RECT 4.000 669.460 745.700 670.620 ;
        RECT 4.000 666.140 746.340 669.460 ;
        RECT 4.000 664.980 745.700 666.140 ;
        RECT 4.000 661.660 746.340 664.980 ;
        RECT 4.000 660.500 745.700 661.660 ;
        RECT 4.000 657.180 746.340 660.500 ;
        RECT 4.000 656.020 745.700 657.180 ;
        RECT 4.000 652.700 746.340 656.020 ;
        RECT 4.000 651.540 745.700 652.700 ;
        RECT 4.000 648.220 746.340 651.540 ;
        RECT 4.000 647.060 745.700 648.220 ;
        RECT 4.000 643.740 746.340 647.060 ;
        RECT 4.300 642.580 745.700 643.740 ;
        RECT 4.000 639.260 746.340 642.580 ;
        RECT 4.000 638.140 745.700 639.260 ;
        RECT 4.300 638.100 745.700 638.140 ;
        RECT 4.300 636.980 746.340 638.100 ;
        RECT 4.000 634.780 746.340 636.980 ;
        RECT 4.000 633.620 745.700 634.780 ;
        RECT 4.000 632.540 746.340 633.620 ;
        RECT 4.300 631.380 746.340 632.540 ;
        RECT 4.000 630.300 746.340 631.380 ;
        RECT 4.000 629.140 745.700 630.300 ;
        RECT 4.000 626.940 746.340 629.140 ;
        RECT 4.300 625.820 746.340 626.940 ;
        RECT 4.300 625.780 745.700 625.820 ;
        RECT 4.000 624.660 745.700 625.780 ;
        RECT 4.000 621.340 746.340 624.660 ;
        RECT 4.300 620.180 745.700 621.340 ;
        RECT 4.000 616.860 746.340 620.180 ;
        RECT 4.000 615.740 745.700 616.860 ;
        RECT 4.300 615.700 745.700 615.740 ;
        RECT 4.300 614.580 746.340 615.700 ;
        RECT 4.000 612.380 746.340 614.580 ;
        RECT 4.000 611.220 745.700 612.380 ;
        RECT 4.000 610.140 746.340 611.220 ;
        RECT 4.300 608.980 746.340 610.140 ;
        RECT 4.000 607.900 746.340 608.980 ;
        RECT 4.000 606.740 745.700 607.900 ;
        RECT 4.000 604.540 746.340 606.740 ;
        RECT 4.300 603.420 746.340 604.540 ;
        RECT 4.300 603.380 745.700 603.420 ;
        RECT 4.000 602.260 745.700 603.380 ;
        RECT 4.000 598.940 746.340 602.260 ;
        RECT 4.300 597.780 745.700 598.940 ;
        RECT 4.000 594.460 746.340 597.780 ;
        RECT 4.000 593.340 745.700 594.460 ;
        RECT 4.300 593.300 745.700 593.340 ;
        RECT 4.300 592.180 746.340 593.300 ;
        RECT 4.000 589.980 746.340 592.180 ;
        RECT 4.000 588.820 745.700 589.980 ;
        RECT 4.000 587.740 746.340 588.820 ;
        RECT 4.300 586.580 746.340 587.740 ;
        RECT 4.000 585.500 746.340 586.580 ;
        RECT 4.000 584.340 745.700 585.500 ;
        RECT 4.000 582.140 746.340 584.340 ;
        RECT 4.300 581.020 746.340 582.140 ;
        RECT 4.300 580.980 745.700 581.020 ;
        RECT 4.000 579.860 745.700 580.980 ;
        RECT 4.000 576.540 746.340 579.860 ;
        RECT 4.300 575.380 745.700 576.540 ;
        RECT 4.000 572.060 746.340 575.380 ;
        RECT 4.000 570.940 745.700 572.060 ;
        RECT 4.300 570.900 745.700 570.940 ;
        RECT 4.300 569.780 746.340 570.900 ;
        RECT 4.000 567.580 746.340 569.780 ;
        RECT 4.000 566.420 745.700 567.580 ;
        RECT 4.000 565.340 746.340 566.420 ;
        RECT 4.300 564.180 746.340 565.340 ;
        RECT 4.000 563.100 746.340 564.180 ;
        RECT 4.000 561.940 745.700 563.100 ;
        RECT 4.000 559.740 746.340 561.940 ;
        RECT 4.300 558.620 746.340 559.740 ;
        RECT 4.300 558.580 745.700 558.620 ;
        RECT 4.000 557.460 745.700 558.580 ;
        RECT 4.000 554.140 746.340 557.460 ;
        RECT 4.300 552.980 745.700 554.140 ;
        RECT 4.000 549.660 746.340 552.980 ;
        RECT 4.000 548.540 745.700 549.660 ;
        RECT 4.300 548.500 745.700 548.540 ;
        RECT 4.300 547.380 746.340 548.500 ;
        RECT 4.000 545.180 746.340 547.380 ;
        RECT 4.000 544.020 745.700 545.180 ;
        RECT 4.000 542.940 746.340 544.020 ;
        RECT 4.300 541.780 746.340 542.940 ;
        RECT 4.000 540.700 746.340 541.780 ;
        RECT 4.000 539.540 745.700 540.700 ;
        RECT 4.000 537.340 746.340 539.540 ;
        RECT 4.300 536.220 746.340 537.340 ;
        RECT 4.300 536.180 745.700 536.220 ;
        RECT 4.000 535.060 745.700 536.180 ;
        RECT 4.000 531.740 746.340 535.060 ;
        RECT 4.300 530.580 745.700 531.740 ;
        RECT 4.000 527.260 746.340 530.580 ;
        RECT 4.000 526.140 745.700 527.260 ;
        RECT 4.300 526.100 745.700 526.140 ;
        RECT 4.300 524.980 746.340 526.100 ;
        RECT 4.000 522.780 746.340 524.980 ;
        RECT 4.000 521.620 745.700 522.780 ;
        RECT 4.000 520.540 746.340 521.620 ;
        RECT 4.300 519.380 746.340 520.540 ;
        RECT 4.000 518.300 746.340 519.380 ;
        RECT 4.000 517.140 745.700 518.300 ;
        RECT 4.000 514.940 746.340 517.140 ;
        RECT 4.300 513.820 746.340 514.940 ;
        RECT 4.300 513.780 745.700 513.820 ;
        RECT 4.000 512.660 745.700 513.780 ;
        RECT 4.000 509.340 746.340 512.660 ;
        RECT 4.300 508.180 745.700 509.340 ;
        RECT 4.000 504.860 746.340 508.180 ;
        RECT 4.000 503.740 745.700 504.860 ;
        RECT 4.300 503.700 745.700 503.740 ;
        RECT 4.300 502.580 746.340 503.700 ;
        RECT 4.000 500.380 746.340 502.580 ;
        RECT 4.000 499.220 745.700 500.380 ;
        RECT 4.000 498.140 746.340 499.220 ;
        RECT 4.300 496.980 746.340 498.140 ;
        RECT 4.000 495.900 746.340 496.980 ;
        RECT 4.000 494.740 745.700 495.900 ;
        RECT 4.000 492.540 746.340 494.740 ;
        RECT 4.300 491.420 746.340 492.540 ;
        RECT 4.300 491.380 745.700 491.420 ;
        RECT 4.000 490.260 745.700 491.380 ;
        RECT 4.000 486.940 746.340 490.260 ;
        RECT 4.300 485.780 745.700 486.940 ;
        RECT 4.000 482.460 746.340 485.780 ;
        RECT 4.000 481.340 745.700 482.460 ;
        RECT 4.300 481.300 745.700 481.340 ;
        RECT 4.300 480.180 746.340 481.300 ;
        RECT 4.000 477.980 746.340 480.180 ;
        RECT 4.000 476.820 745.700 477.980 ;
        RECT 4.000 475.740 746.340 476.820 ;
        RECT 4.300 474.580 746.340 475.740 ;
        RECT 4.000 473.500 746.340 474.580 ;
        RECT 4.000 472.340 745.700 473.500 ;
        RECT 4.000 470.140 746.340 472.340 ;
        RECT 4.300 469.020 746.340 470.140 ;
        RECT 4.300 468.980 745.700 469.020 ;
        RECT 4.000 467.860 745.700 468.980 ;
        RECT 4.000 464.540 746.340 467.860 ;
        RECT 4.300 463.380 745.700 464.540 ;
        RECT 4.000 460.060 746.340 463.380 ;
        RECT 4.000 458.940 745.700 460.060 ;
        RECT 4.300 458.900 745.700 458.940 ;
        RECT 4.300 457.780 746.340 458.900 ;
        RECT 4.000 455.580 746.340 457.780 ;
        RECT 4.000 454.420 745.700 455.580 ;
        RECT 4.000 453.340 746.340 454.420 ;
        RECT 4.300 452.180 746.340 453.340 ;
        RECT 4.000 451.100 746.340 452.180 ;
        RECT 4.000 449.940 745.700 451.100 ;
        RECT 4.000 447.740 746.340 449.940 ;
        RECT 4.300 446.620 746.340 447.740 ;
        RECT 4.300 446.580 745.700 446.620 ;
        RECT 4.000 445.460 745.700 446.580 ;
        RECT 4.000 442.140 746.340 445.460 ;
        RECT 4.300 440.980 745.700 442.140 ;
        RECT 4.000 437.660 746.340 440.980 ;
        RECT 4.000 436.540 745.700 437.660 ;
        RECT 4.300 436.500 745.700 436.540 ;
        RECT 4.300 435.380 746.340 436.500 ;
        RECT 4.000 433.180 746.340 435.380 ;
        RECT 4.000 432.020 745.700 433.180 ;
        RECT 4.000 430.940 746.340 432.020 ;
        RECT 4.300 429.780 746.340 430.940 ;
        RECT 4.000 428.700 746.340 429.780 ;
        RECT 4.000 427.540 745.700 428.700 ;
        RECT 4.000 425.340 746.340 427.540 ;
        RECT 4.300 424.220 746.340 425.340 ;
        RECT 4.300 424.180 745.700 424.220 ;
        RECT 4.000 423.060 745.700 424.180 ;
        RECT 4.000 419.740 746.340 423.060 ;
        RECT 4.300 418.580 745.700 419.740 ;
        RECT 4.000 415.260 746.340 418.580 ;
        RECT 4.000 414.140 745.700 415.260 ;
        RECT 4.300 414.100 745.700 414.140 ;
        RECT 4.300 412.980 746.340 414.100 ;
        RECT 4.000 410.780 746.340 412.980 ;
        RECT 4.000 409.620 745.700 410.780 ;
        RECT 4.000 408.540 746.340 409.620 ;
        RECT 4.300 407.380 746.340 408.540 ;
        RECT 4.000 406.300 746.340 407.380 ;
        RECT 4.000 405.140 745.700 406.300 ;
        RECT 4.000 402.940 746.340 405.140 ;
        RECT 4.300 401.820 746.340 402.940 ;
        RECT 4.300 401.780 745.700 401.820 ;
        RECT 4.000 400.660 745.700 401.780 ;
        RECT 4.000 397.340 746.340 400.660 ;
        RECT 4.300 396.180 745.700 397.340 ;
        RECT 4.000 392.860 746.340 396.180 ;
        RECT 4.000 391.740 745.700 392.860 ;
        RECT 4.300 391.700 745.700 391.740 ;
        RECT 4.300 390.580 746.340 391.700 ;
        RECT 4.000 388.380 746.340 390.580 ;
        RECT 4.000 387.220 745.700 388.380 ;
        RECT 4.000 386.140 746.340 387.220 ;
        RECT 4.300 384.980 746.340 386.140 ;
        RECT 4.000 383.900 746.340 384.980 ;
        RECT 4.000 382.740 745.700 383.900 ;
        RECT 4.000 380.540 746.340 382.740 ;
        RECT 4.300 379.420 746.340 380.540 ;
        RECT 4.300 379.380 745.700 379.420 ;
        RECT 4.000 378.260 745.700 379.380 ;
        RECT 4.000 374.940 746.340 378.260 ;
        RECT 4.300 373.780 745.700 374.940 ;
        RECT 4.000 370.460 746.340 373.780 ;
        RECT 4.000 369.340 745.700 370.460 ;
        RECT 4.300 369.300 745.700 369.340 ;
        RECT 4.300 368.180 746.340 369.300 ;
        RECT 4.000 365.980 746.340 368.180 ;
        RECT 4.000 364.820 745.700 365.980 ;
        RECT 4.000 363.740 746.340 364.820 ;
        RECT 4.300 362.580 746.340 363.740 ;
        RECT 4.000 361.500 746.340 362.580 ;
        RECT 4.000 360.340 745.700 361.500 ;
        RECT 4.000 358.140 746.340 360.340 ;
        RECT 4.300 357.020 746.340 358.140 ;
        RECT 4.300 356.980 745.700 357.020 ;
        RECT 4.000 355.860 745.700 356.980 ;
        RECT 4.000 352.540 746.340 355.860 ;
        RECT 4.300 351.380 745.700 352.540 ;
        RECT 4.000 348.060 746.340 351.380 ;
        RECT 4.000 346.940 745.700 348.060 ;
        RECT 4.300 346.900 745.700 346.940 ;
        RECT 4.300 345.780 746.340 346.900 ;
        RECT 4.000 343.580 746.340 345.780 ;
        RECT 4.000 342.420 745.700 343.580 ;
        RECT 4.000 341.340 746.340 342.420 ;
        RECT 4.300 340.180 746.340 341.340 ;
        RECT 4.000 339.100 746.340 340.180 ;
        RECT 4.000 337.940 745.700 339.100 ;
        RECT 4.000 335.740 746.340 337.940 ;
        RECT 4.300 334.620 746.340 335.740 ;
        RECT 4.300 334.580 745.700 334.620 ;
        RECT 4.000 333.460 745.700 334.580 ;
        RECT 4.000 330.140 746.340 333.460 ;
        RECT 4.300 328.980 745.700 330.140 ;
        RECT 4.000 325.660 746.340 328.980 ;
        RECT 4.000 324.540 745.700 325.660 ;
        RECT 4.300 324.500 745.700 324.540 ;
        RECT 4.300 323.380 746.340 324.500 ;
        RECT 4.000 321.180 746.340 323.380 ;
        RECT 4.000 320.020 745.700 321.180 ;
        RECT 4.000 318.940 746.340 320.020 ;
        RECT 4.300 317.780 746.340 318.940 ;
        RECT 4.000 316.700 746.340 317.780 ;
        RECT 4.000 315.540 745.700 316.700 ;
        RECT 4.000 313.340 746.340 315.540 ;
        RECT 4.300 312.220 746.340 313.340 ;
        RECT 4.300 312.180 745.700 312.220 ;
        RECT 4.000 311.060 745.700 312.180 ;
        RECT 4.000 307.740 746.340 311.060 ;
        RECT 4.300 306.580 745.700 307.740 ;
        RECT 4.000 303.260 746.340 306.580 ;
        RECT 4.000 302.140 745.700 303.260 ;
        RECT 4.300 302.100 745.700 302.140 ;
        RECT 4.300 300.980 746.340 302.100 ;
        RECT 4.000 298.780 746.340 300.980 ;
        RECT 4.000 297.620 745.700 298.780 ;
        RECT 4.000 296.540 746.340 297.620 ;
        RECT 4.300 295.380 746.340 296.540 ;
        RECT 4.000 294.300 746.340 295.380 ;
        RECT 4.000 293.140 745.700 294.300 ;
        RECT 4.000 290.940 746.340 293.140 ;
        RECT 4.300 289.820 746.340 290.940 ;
        RECT 4.300 289.780 745.700 289.820 ;
        RECT 4.000 288.660 745.700 289.780 ;
        RECT 4.000 285.340 746.340 288.660 ;
        RECT 4.300 284.180 745.700 285.340 ;
        RECT 4.000 280.860 746.340 284.180 ;
        RECT 4.000 279.740 745.700 280.860 ;
        RECT 4.300 279.700 745.700 279.740 ;
        RECT 4.300 278.580 746.340 279.700 ;
        RECT 4.000 276.380 746.340 278.580 ;
        RECT 4.000 275.220 745.700 276.380 ;
        RECT 4.000 274.140 746.340 275.220 ;
        RECT 4.300 272.980 746.340 274.140 ;
        RECT 4.000 271.900 746.340 272.980 ;
        RECT 4.000 270.740 745.700 271.900 ;
        RECT 4.000 268.540 746.340 270.740 ;
        RECT 4.300 267.420 746.340 268.540 ;
        RECT 4.300 267.380 745.700 267.420 ;
        RECT 4.000 266.260 745.700 267.380 ;
        RECT 4.000 262.940 746.340 266.260 ;
        RECT 4.300 261.780 745.700 262.940 ;
        RECT 4.000 258.460 746.340 261.780 ;
        RECT 4.000 257.340 745.700 258.460 ;
        RECT 4.300 257.300 745.700 257.340 ;
        RECT 4.300 256.180 746.340 257.300 ;
        RECT 4.000 253.980 746.340 256.180 ;
        RECT 4.000 252.820 745.700 253.980 ;
        RECT 4.000 251.740 746.340 252.820 ;
        RECT 4.300 250.580 746.340 251.740 ;
        RECT 4.000 249.500 746.340 250.580 ;
        RECT 4.000 248.340 745.700 249.500 ;
        RECT 4.000 246.140 746.340 248.340 ;
        RECT 4.300 245.020 746.340 246.140 ;
        RECT 4.300 244.980 745.700 245.020 ;
        RECT 4.000 243.860 745.700 244.980 ;
        RECT 4.000 240.540 746.340 243.860 ;
        RECT 4.300 239.380 745.700 240.540 ;
        RECT 4.000 236.060 746.340 239.380 ;
        RECT 4.000 234.940 745.700 236.060 ;
        RECT 4.300 234.900 745.700 234.940 ;
        RECT 4.300 233.780 746.340 234.900 ;
        RECT 4.000 231.580 746.340 233.780 ;
        RECT 4.000 230.420 745.700 231.580 ;
        RECT 4.000 229.340 746.340 230.420 ;
        RECT 4.300 228.180 746.340 229.340 ;
        RECT 4.000 227.100 746.340 228.180 ;
        RECT 4.000 225.940 745.700 227.100 ;
        RECT 4.000 223.740 746.340 225.940 ;
        RECT 4.300 222.620 746.340 223.740 ;
        RECT 4.300 222.580 745.700 222.620 ;
        RECT 4.000 221.460 745.700 222.580 ;
        RECT 4.000 218.140 746.340 221.460 ;
        RECT 4.300 216.980 745.700 218.140 ;
        RECT 4.000 213.660 746.340 216.980 ;
        RECT 4.000 212.540 745.700 213.660 ;
        RECT 4.300 212.500 745.700 212.540 ;
        RECT 4.300 211.380 746.340 212.500 ;
        RECT 4.000 209.180 746.340 211.380 ;
        RECT 4.000 208.020 745.700 209.180 ;
        RECT 4.000 206.940 746.340 208.020 ;
        RECT 4.300 205.780 746.340 206.940 ;
        RECT 4.000 204.700 746.340 205.780 ;
        RECT 4.000 203.540 745.700 204.700 ;
        RECT 4.000 201.340 746.340 203.540 ;
        RECT 4.300 200.220 746.340 201.340 ;
        RECT 4.300 200.180 745.700 200.220 ;
        RECT 4.000 199.060 745.700 200.180 ;
        RECT 4.000 195.740 746.340 199.060 ;
        RECT 4.300 194.580 745.700 195.740 ;
        RECT 4.000 191.260 746.340 194.580 ;
        RECT 4.000 190.140 745.700 191.260 ;
        RECT 4.300 190.100 745.700 190.140 ;
        RECT 4.300 188.980 746.340 190.100 ;
        RECT 4.000 186.780 746.340 188.980 ;
        RECT 4.000 185.620 745.700 186.780 ;
        RECT 4.000 184.540 746.340 185.620 ;
        RECT 4.300 183.380 746.340 184.540 ;
        RECT 4.000 182.300 746.340 183.380 ;
        RECT 4.000 181.140 745.700 182.300 ;
        RECT 4.000 178.940 746.340 181.140 ;
        RECT 4.300 177.820 746.340 178.940 ;
        RECT 4.300 177.780 745.700 177.820 ;
        RECT 4.000 176.660 745.700 177.780 ;
        RECT 4.000 173.340 746.340 176.660 ;
        RECT 4.300 172.180 745.700 173.340 ;
        RECT 4.000 168.860 746.340 172.180 ;
        RECT 4.000 167.740 745.700 168.860 ;
        RECT 4.300 167.700 745.700 167.740 ;
        RECT 4.300 166.580 746.340 167.700 ;
        RECT 4.000 164.380 746.340 166.580 ;
        RECT 4.000 163.220 745.700 164.380 ;
        RECT 4.000 162.140 746.340 163.220 ;
        RECT 4.300 160.980 746.340 162.140 ;
        RECT 4.000 159.900 746.340 160.980 ;
        RECT 4.000 158.740 745.700 159.900 ;
        RECT 4.000 156.540 746.340 158.740 ;
        RECT 4.300 155.420 746.340 156.540 ;
        RECT 4.300 155.380 745.700 155.420 ;
        RECT 4.000 154.260 745.700 155.380 ;
        RECT 4.000 150.940 746.340 154.260 ;
        RECT 4.300 149.780 745.700 150.940 ;
        RECT 4.000 146.460 746.340 149.780 ;
        RECT 4.000 145.340 745.700 146.460 ;
        RECT 4.300 145.300 745.700 145.340 ;
        RECT 4.300 144.180 746.340 145.300 ;
        RECT 4.000 141.980 746.340 144.180 ;
        RECT 4.000 140.820 745.700 141.980 ;
        RECT 4.000 139.740 746.340 140.820 ;
        RECT 4.300 138.580 746.340 139.740 ;
        RECT 4.000 137.500 746.340 138.580 ;
        RECT 4.000 136.340 745.700 137.500 ;
        RECT 4.000 134.140 746.340 136.340 ;
        RECT 4.300 133.020 746.340 134.140 ;
        RECT 4.300 132.980 745.700 133.020 ;
        RECT 4.000 131.860 745.700 132.980 ;
        RECT 4.000 128.540 746.340 131.860 ;
        RECT 4.300 127.380 745.700 128.540 ;
        RECT 4.000 124.060 746.340 127.380 ;
        RECT 4.000 122.940 745.700 124.060 ;
        RECT 4.300 122.900 745.700 122.940 ;
        RECT 4.300 121.780 746.340 122.900 ;
        RECT 4.000 119.580 746.340 121.780 ;
        RECT 4.000 118.420 745.700 119.580 ;
        RECT 4.000 117.340 746.340 118.420 ;
        RECT 4.300 116.180 746.340 117.340 ;
        RECT 4.000 115.100 746.340 116.180 ;
        RECT 4.000 113.940 745.700 115.100 ;
        RECT 4.000 111.740 746.340 113.940 ;
        RECT 4.300 110.620 746.340 111.740 ;
        RECT 4.300 110.580 745.700 110.620 ;
        RECT 4.000 109.460 745.700 110.580 ;
        RECT 4.000 106.140 746.340 109.460 ;
        RECT 4.300 104.980 745.700 106.140 ;
        RECT 4.000 101.660 746.340 104.980 ;
        RECT 4.000 100.540 745.700 101.660 ;
        RECT 4.300 100.500 745.700 100.540 ;
        RECT 4.300 99.380 746.340 100.500 ;
        RECT 4.000 97.180 746.340 99.380 ;
        RECT 4.000 96.020 745.700 97.180 ;
        RECT 4.000 94.940 746.340 96.020 ;
        RECT 4.300 93.780 746.340 94.940 ;
        RECT 4.000 92.700 746.340 93.780 ;
        RECT 4.000 91.540 745.700 92.700 ;
        RECT 4.000 89.340 746.340 91.540 ;
        RECT 4.300 88.220 746.340 89.340 ;
        RECT 4.300 88.180 745.700 88.220 ;
        RECT 4.000 87.060 745.700 88.180 ;
        RECT 4.000 83.740 746.340 87.060 ;
        RECT 4.300 82.580 745.700 83.740 ;
        RECT 4.000 79.260 746.340 82.580 ;
        RECT 4.000 78.140 745.700 79.260 ;
        RECT 4.300 78.100 745.700 78.140 ;
        RECT 4.300 76.980 746.340 78.100 ;
        RECT 4.000 74.780 746.340 76.980 ;
        RECT 4.000 73.620 745.700 74.780 ;
        RECT 4.000 72.540 746.340 73.620 ;
        RECT 4.300 71.380 746.340 72.540 ;
        RECT 4.000 70.300 746.340 71.380 ;
        RECT 4.000 69.140 745.700 70.300 ;
        RECT 4.000 66.940 746.340 69.140 ;
        RECT 4.300 65.820 746.340 66.940 ;
        RECT 4.300 65.780 745.700 65.820 ;
        RECT 4.000 64.660 745.700 65.780 ;
        RECT 4.000 61.340 746.340 64.660 ;
        RECT 4.300 60.180 745.700 61.340 ;
        RECT 4.000 56.860 746.340 60.180 ;
        RECT 4.000 55.740 745.700 56.860 ;
        RECT 4.300 55.700 745.700 55.740 ;
        RECT 4.300 54.580 746.340 55.700 ;
        RECT 4.000 52.380 746.340 54.580 ;
        RECT 4.000 51.220 745.700 52.380 ;
        RECT 4.000 47.900 746.340 51.220 ;
        RECT 4.000 46.740 745.700 47.900 ;
        RECT 4.000 43.420 746.340 46.740 ;
        RECT 4.000 42.260 745.700 43.420 ;
        RECT 4.000 38.940 746.340 42.260 ;
        RECT 4.000 37.780 745.700 38.940 ;
        RECT 4.000 34.460 746.340 37.780 ;
        RECT 4.000 33.300 745.700 34.460 ;
        RECT 4.000 29.980 746.340 33.300 ;
        RECT 4.000 28.820 745.700 29.980 ;
        RECT 4.000 3.500 746.340 28.820 ;
      LAYER Metal4 ;
        RECT 262.780 682.680 738.500 692.630 ;
        RECT 262.780 15.080 329.140 682.680 ;
        RECT 331.340 15.080 405.940 682.680 ;
        RECT 408.140 15.080 482.740 682.680 ;
        RECT 484.940 15.080 559.540 682.680 ;
        RECT 561.740 15.080 636.340 682.680 ;
        RECT 638.540 15.080 713.140 682.680 ;
        RECT 715.340 15.080 738.500 682.680 ;
        RECT 262.780 10.730 738.500 15.080 ;
  END
END multiplexer
END LIBRARY

